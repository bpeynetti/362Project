
module PipeCtlRegN_WIDTH108 ( out, in, ctl, clk, reset );
  output [0:107] out;
  input [0:107] in;
  input ctl, clk, reset;
  wire   n217, n218, n219, n220, n221, n222;

  SDFFR_X2 \out_reg[0]  ( .D(1'b0), .SI(n219), .SE(in[0]), .CK(clk), .RN(reset), .Q(out[0]) );
  SDFFR_X2 \out_reg[1]  ( .D(1'b0), .SI(n220), .SE(in[1]), .CK(clk), .RN(reset), .Q(out[1]) );
  SDFFR_X2 \out_reg[2]  ( .D(1'b0), .SI(n221), .SE(in[2]), .CK(clk), .RN(reset), .Q(out[2]) );
  SDFFR_X2 \out_reg[3]  ( .D(1'b0), .SI(n222), .SE(in[3]), .CK(clk), .RN(reset), .Q(out[3]) );
  SDFFR_X2 \out_reg[4]  ( .D(1'b0), .SI(n219), .SE(in[4]), .CK(clk), .RN(reset), .Q(out[4]) );
  SDFFR_X2 \out_reg[5]  ( .D(1'b0), .SI(n220), .SE(in[5]), .CK(clk), .RN(reset), .Q(out[5]) );
  SDFFR_X2 \out_reg[6]  ( .D(1'b0), .SI(n221), .SE(in[6]), .CK(clk), .RN(reset), .Q(out[6]) );
  SDFFR_X2 \out_reg[7]  ( .D(1'b0), .SI(n222), .SE(in[7]), .CK(clk), .RN(reset), .Q(out[7]) );
  SDFFR_X2 \out_reg[8]  ( .D(1'b0), .SI(n219), .SE(in[8]), .CK(clk), .RN(reset), .Q(out[8]) );
  SDFFR_X2 \out_reg[9]  ( .D(1'b0), .SI(n220), .SE(in[9]), .CK(clk), .RN(reset), .Q(out[9]) );
  SDFFR_X2 \out_reg[10]  ( .D(1'b0), .SI(n221), .SE(in[10]), .CK(clk), .RN(
        reset), .Q(out[10]) );
  SDFFR_X2 \out_reg[11]  ( .D(1'b0), .SI(n222), .SE(in[11]), .CK(clk), .RN(
        reset), .Q(out[11]) );
  SDFFR_X2 \out_reg[12]  ( .D(1'b0), .SI(n219), .SE(in[12]), .CK(clk), .RN(
        reset), .Q(out[12]) );
  SDFFR_X2 \out_reg[13]  ( .D(1'b0), .SI(n220), .SE(in[13]), .CK(clk), .RN(
        reset), .Q(out[13]) );
  SDFFR_X2 \out_reg[14]  ( .D(1'b0), .SI(n221), .SE(in[14]), .CK(clk), .RN(
        reset), .Q(out[14]) );
  SDFFR_X2 \out_reg[15]  ( .D(1'b0), .SI(n222), .SE(in[15]), .CK(clk), .RN(
        reset), .Q(out[15]) );
  SDFFR_X2 \out_reg[16]  ( .D(1'b0), .SI(n219), .SE(in[16]), .CK(clk), .RN(
        reset), .Q(out[16]) );
  SDFFR_X2 \out_reg[17]  ( .D(1'b0), .SI(n220), .SE(in[17]), .CK(clk), .RN(
        reset), .Q(out[17]) );
  SDFFR_X2 \out_reg[18]  ( .D(1'b0), .SI(n221), .SE(in[18]), .CK(clk), .RN(
        reset), .Q(out[18]) );
  SDFFR_X2 \out_reg[19]  ( .D(1'b0), .SI(n222), .SE(in[19]), .CK(clk), .RN(
        reset), .Q(out[19]) );
  SDFFR_X2 \out_reg[20]  ( .D(1'b0), .SI(n219), .SE(in[20]), .CK(clk), .RN(
        reset), .Q(out[20]) );
  SDFFR_X2 \out_reg[21]  ( .D(1'b0), .SI(n220), .SE(in[21]), .CK(clk), .RN(
        reset), .Q(out[21]) );
  SDFFR_X2 \out_reg[22]  ( .D(1'b0), .SI(n221), .SE(in[22]), .CK(clk), .RN(
        reset), .Q(out[22]) );
  SDFFR_X2 \out_reg[23]  ( .D(1'b0), .SI(n222), .SE(in[23]), .CK(clk), .RN(
        reset), .Q(out[23]) );
  SDFFR_X2 \out_reg[24]  ( .D(1'b0), .SI(n219), .SE(in[24]), .CK(clk), .RN(
        reset), .Q(out[24]) );
  SDFFR_X2 \out_reg[25]  ( .D(1'b0), .SI(n220), .SE(in[25]), .CK(clk), .RN(
        reset), .Q(out[25]) );
  SDFFR_X2 \out_reg[26]  ( .D(1'b0), .SI(n221), .SE(in[26]), .CK(clk), .RN(
        reset), .Q(out[26]) );
  SDFFR_X2 \out_reg[27]  ( .D(1'b0), .SI(n222), .SE(in[27]), .CK(clk), .RN(
        reset), .Q(out[27]) );
  SDFFR_X2 \out_reg[28]  ( .D(1'b0), .SI(n219), .SE(in[28]), .CK(clk), .RN(
        reset), .Q(out[28]) );
  SDFFR_X2 \out_reg[29]  ( .D(1'b0), .SI(n220), .SE(in[29]), .CK(clk), .RN(
        reset), .Q(out[29]) );
  SDFFR_X2 \out_reg[30]  ( .D(1'b0), .SI(n221), .SE(in[30]), .CK(clk), .RN(
        reset), .Q(out[30]) );
  SDFFR_X2 \out_reg[31]  ( .D(1'b0), .SI(n222), .SE(in[31]), .CK(clk), .RN(
        reset), .Q(out[31]) );
  SDFFR_X2 \out_reg[32]  ( .D(1'b0), .SI(n219), .SE(in[32]), .CK(clk), .RN(
        reset), .Q(out[32]) );
  SDFFR_X2 \out_reg[33]  ( .D(1'b0), .SI(n220), .SE(in[33]), .CK(clk), .RN(
        reset), .Q(out[33]) );
  SDFFR_X2 \out_reg[34]  ( .D(1'b0), .SI(n221), .SE(in[34]), .CK(clk), .RN(
        reset), .Q(out[34]) );
  SDFFR_X2 \out_reg[35]  ( .D(1'b0), .SI(n222), .SE(in[35]), .CK(clk), .RN(
        reset), .Q(out[35]) );
  SDFFR_X2 \out_reg[36]  ( .D(1'b0), .SI(n219), .SE(in[36]), .CK(clk), .RN(
        reset), .Q(out[36]) );
  SDFFR_X2 \out_reg[37]  ( .D(1'b0), .SI(n220), .SE(in[37]), .CK(clk), .RN(
        reset), .Q(out[37]) );
  SDFFR_X2 \out_reg[38]  ( .D(1'b0), .SI(n221), .SE(in[38]), .CK(clk), .RN(
        reset), .Q(out[38]) );
  SDFFR_X2 \out_reg[39]  ( .D(1'b0), .SI(n222), .SE(in[39]), .CK(clk), .RN(
        reset), .Q(out[39]) );
  SDFFR_X2 \out_reg[40]  ( .D(1'b0), .SI(n219), .SE(in[40]), .CK(clk), .RN(
        reset), .Q(out[40]) );
  SDFFR_X2 \out_reg[41]  ( .D(1'b0), .SI(n220), .SE(in[41]), .CK(clk), .RN(
        reset), .Q(out[41]) );
  SDFFR_X2 \out_reg[42]  ( .D(1'b0), .SI(n221), .SE(in[42]), .CK(clk), .RN(
        reset), .Q(out[42]) );
  SDFFR_X2 \out_reg[43]  ( .D(1'b0), .SI(n222), .SE(in[43]), .CK(clk), .RN(
        reset), .Q(out[43]) );
  SDFFR_X2 \out_reg[44]  ( .D(1'b0), .SI(n219), .SE(in[44]), .CK(clk), .RN(
        reset), .Q(out[44]) );
  SDFFR_X2 \out_reg[45]  ( .D(1'b0), .SI(n220), .SE(in[45]), .CK(clk), .RN(
        reset), .Q(out[45]) );
  SDFFR_X2 \out_reg[46]  ( .D(1'b0), .SI(n221), .SE(in[46]), .CK(clk), .RN(
        reset), .Q(out[46]) );
  SDFFR_X2 \out_reg[47]  ( .D(1'b0), .SI(n222), .SE(in[47]), .CK(clk), .RN(
        reset), .Q(out[47]) );
  SDFFR_X2 \out_reg[48]  ( .D(1'b0), .SI(n219), .SE(in[48]), .CK(clk), .RN(
        reset), .Q(out[48]) );
  SDFFR_X2 \out_reg[49]  ( .D(1'b0), .SI(n220), .SE(in[49]), .CK(clk), .RN(
        reset), .Q(out[49]) );
  SDFFR_X2 \out_reg[50]  ( .D(1'b0), .SI(n221), .SE(in[50]), .CK(clk), .RN(
        reset), .Q(out[50]) );
  SDFFR_X2 \out_reg[51]  ( .D(1'b0), .SI(n222), .SE(in[51]), .CK(clk), .RN(
        reset), .Q(out[51]) );
  SDFFR_X2 \out_reg[52]  ( .D(1'b0), .SI(n219), .SE(in[52]), .CK(clk), .RN(
        reset), .Q(out[52]) );
  SDFFR_X2 \out_reg[53]  ( .D(1'b0), .SI(n220), .SE(in[53]), .CK(clk), .RN(
        reset), .Q(out[53]) );
  SDFFR_X2 \out_reg[54]  ( .D(1'b0), .SI(n221), .SE(in[54]), .CK(clk), .RN(
        reset), .Q(out[54]) );
  SDFFR_X2 \out_reg[55]  ( .D(1'b0), .SI(n222), .SE(in[55]), .CK(clk), .RN(
        reset), .Q(out[55]) );
  SDFFR_X2 \out_reg[56]  ( .D(1'b0), .SI(n219), .SE(in[56]), .CK(clk), .RN(
        reset), .Q(out[56]) );
  SDFFR_X2 \out_reg[57]  ( .D(1'b0), .SI(n220), .SE(in[57]), .CK(clk), .RN(
        reset), .Q(out[57]) );
  SDFFR_X2 \out_reg[58]  ( .D(1'b0), .SI(n221), .SE(in[58]), .CK(clk), .RN(
        reset), .Q(out[58]) );
  SDFFR_X2 \out_reg[59]  ( .D(1'b0), .SI(n222), .SE(in[59]), .CK(clk), .RN(
        reset), .Q(out[59]) );
  SDFFR_X2 \out_reg[60]  ( .D(1'b0), .SI(n219), .SE(in[60]), .CK(clk), .RN(
        reset), .Q(out[60]) );
  SDFFR_X2 \out_reg[61]  ( .D(1'b0), .SI(n220), .SE(in[61]), .CK(clk), .RN(
        reset), .Q(out[61]) );
  SDFFR_X2 \out_reg[62]  ( .D(1'b0), .SI(n221), .SE(in[62]), .CK(clk), .RN(
        reset), .Q(out[62]) );
  SDFFR_X2 \out_reg[63]  ( .D(1'b0), .SI(n222), .SE(in[63]), .CK(clk), .RN(
        reset), .Q(out[63]) );
  SDFFR_X2 \out_reg[64]  ( .D(1'b0), .SI(n219), .SE(in[64]), .CK(clk), .RN(
        reset), .Q(out[64]) );
  SDFFR_X2 \out_reg[65]  ( .D(1'b0), .SI(n220), .SE(in[65]), .CK(clk), .RN(
        reset), .Q(out[65]) );
  SDFFR_X2 \out_reg[66]  ( .D(1'b0), .SI(n221), .SE(in[66]), .CK(clk), .RN(
        reset), .Q(out[66]) );
  SDFFR_X2 \out_reg[67]  ( .D(1'b0), .SI(n222), .SE(in[67]), .CK(clk), .RN(
        reset), .Q(out[67]) );
  SDFFR_X2 \out_reg[68]  ( .D(1'b0), .SI(n219), .SE(in[68]), .CK(clk), .RN(
        reset), .Q(out[68]) );
  SDFFR_X2 \out_reg[69]  ( .D(1'b0), .SI(n220), .SE(in[69]), .CK(clk), .RN(
        reset), .Q(out[69]) );
  SDFFR_X2 \out_reg[70]  ( .D(1'b0), .SI(n221), .SE(in[70]), .CK(clk), .RN(
        reset), .Q(out[70]) );
  SDFFR_X2 \out_reg[71]  ( .D(1'b0), .SI(n222), .SE(in[71]), .CK(clk), .RN(
        reset), .Q(out[71]) );
  SDFFR_X2 \out_reg[72]  ( .D(1'b0), .SI(n219), .SE(in[72]), .CK(clk), .RN(
        reset), .Q(out[72]) );
  SDFFR_X2 \out_reg[73]  ( .D(1'b0), .SI(n220), .SE(in[73]), .CK(clk), .RN(
        reset), .Q(out[73]) );
  SDFFR_X2 \out_reg[74]  ( .D(1'b0), .SI(n221), .SE(in[74]), .CK(clk), .RN(
        reset), .Q(out[74]) );
  SDFFR_X2 \out_reg[75]  ( .D(1'b0), .SI(n222), .SE(in[75]), .CK(clk), .RN(
        reset), .Q(out[75]) );
  SDFFR_X2 \out_reg[76]  ( .D(1'b0), .SI(n219), .SE(in[76]), .CK(clk), .RN(
        reset), .Q(out[76]) );
  SDFFR_X2 \out_reg[77]  ( .D(1'b0), .SI(n220), .SE(in[77]), .CK(clk), .RN(
        reset), .Q(out[77]) );
  SDFFR_X2 \out_reg[78]  ( .D(1'b0), .SI(n221), .SE(in[78]), .CK(clk), .RN(
        reset), .Q(out[78]) );
  SDFFR_X2 \out_reg[79]  ( .D(1'b0), .SI(n222), .SE(in[79]), .CK(clk), .RN(
        reset), .Q(out[79]) );
  SDFFR_X2 \out_reg[80]  ( .D(1'b0), .SI(n219), .SE(in[80]), .CK(clk), .RN(
        reset), .Q(out[80]) );
  SDFFR_X2 \out_reg[81]  ( .D(1'b0), .SI(n220), .SE(in[81]), .CK(clk), .RN(
        reset), .Q(out[81]) );
  SDFFR_X2 \out_reg[82]  ( .D(1'b0), .SI(n221), .SE(in[82]), .CK(clk), .RN(
        reset), .Q(out[82]) );
  SDFFR_X2 \out_reg[83]  ( .D(1'b0), .SI(n222), .SE(in[83]), .CK(clk), .RN(
        reset), .Q(out[83]) );
  SDFFR_X2 \out_reg[84]  ( .D(1'b0), .SI(n219), .SE(in[84]), .CK(clk), .RN(
        reset), .Q(out[84]) );
  SDFFR_X2 \out_reg[85]  ( .D(1'b0), .SI(n220), .SE(in[85]), .CK(clk), .RN(
        reset), .Q(out[85]) );
  SDFFR_X2 \out_reg[86]  ( .D(1'b0), .SI(n221), .SE(in[86]), .CK(clk), .RN(
        reset), .Q(out[86]) );
  SDFFR_X2 \out_reg[87]  ( .D(1'b0), .SI(n222), .SE(in[87]), .CK(clk), .RN(
        reset), .Q(out[87]) );
  SDFFR_X2 \out_reg[88]  ( .D(1'b0), .SI(n219), .SE(in[88]), .CK(clk), .RN(
        reset), .Q(out[88]) );
  SDFFR_X2 \out_reg[89]  ( .D(1'b0), .SI(n220), .SE(in[89]), .CK(clk), .RN(
        reset), .Q(out[89]) );
  SDFFR_X2 \out_reg[90]  ( .D(1'b0), .SI(n221), .SE(in[90]), .CK(clk), .RN(
        reset), .Q(out[90]) );
  SDFFR_X2 \out_reg[91]  ( .D(1'b0), .SI(n222), .SE(in[91]), .CK(clk), .RN(
        reset), .Q(out[91]) );
  SDFFR_X2 \out_reg[92]  ( .D(1'b0), .SI(n219), .SE(in[92]), .CK(clk), .RN(
        reset), .Q(out[92]) );
  SDFFR_X2 \out_reg[93]  ( .D(1'b0), .SI(n220), .SE(in[93]), .CK(clk), .RN(
        reset), .Q(out[93]) );
  SDFFR_X2 \out_reg[94]  ( .D(1'b0), .SI(n221), .SE(in[94]), .CK(clk), .RN(
        reset), .Q(out[94]) );
  SDFFR_X2 \out_reg[95]  ( .D(1'b0), .SI(n222), .SE(in[95]), .CK(clk), .RN(
        reset), .Q(out[95]) );
  SDFFR_X2 \out_reg[96]  ( .D(1'b0), .SI(n219), .SE(in[96]), .CK(clk), .RN(
        reset), .Q(out[96]) );
  SDFFR_X2 \out_reg[97]  ( .D(1'b0), .SI(n220), .SE(in[97]), .CK(clk), .RN(
        reset), .Q(out[97]) );
  SDFFR_X2 \out_reg[98]  ( .D(1'b0), .SI(n221), .SE(in[98]), .CK(clk), .RN(
        reset), .Q(out[98]) );
  SDFFR_X2 \out_reg[99]  ( .D(1'b0), .SI(n222), .SE(in[99]), .CK(clk), .RN(
        reset), .Q(out[99]) );
  SDFFR_X2 \out_reg[100]  ( .D(1'b0), .SI(n219), .SE(in[100]), .CK(clk), .RN(
        reset), .Q(out[100]) );
  SDFFR_X2 \out_reg[101]  ( .D(1'b0), .SI(n220), .SE(in[101]), .CK(clk), .RN(
        reset), .Q(out[101]) );
  SDFFR_X2 \out_reg[102]  ( .D(1'b0), .SI(n221), .SE(in[102]), .CK(clk), .RN(
        reset), .Q(out[102]) );
  SDFFR_X2 \out_reg[103]  ( .D(1'b0), .SI(n222), .SE(in[103]), .CK(clk), .RN(
        reset), .Q(out[103]) );
  SDFFR_X2 \out_reg[104]  ( .D(1'b0), .SI(n219), .SE(in[104]), .CK(clk), .RN(
        reset), .Q(out[104]) );
  SDFFR_X2 \out_reg[105]  ( .D(1'b0), .SI(n220), .SE(in[105]), .CK(clk), .RN(
        reset), .Q(out[105]) );
  SDFFR_X2 \out_reg[106]  ( .D(1'b0), .SI(n221), .SE(in[106]), .CK(clk), .RN(
        reset), .Q(out[106]) );
  SDFFR_X2 \out_reg[107]  ( .D(1'b0), .SI(n222), .SE(in[107]), .CK(clk), .RN(
        reset), .Q(out[107]) );
  INV_X1 U111 ( .A(ctl), .ZN(n217) );
  INV_X1 U112 ( .A(n217), .ZN(n218) );
  INV_X4 U113 ( .A(n218), .ZN(n219) );
  INV_X4 U114 ( .A(n218), .ZN(n220) );
  INV_X4 U115 ( .A(n218), .ZN(n221) );
  INV_X4 U116 ( .A(n218), .ZN(n222) );
endmodule

