
module mem_wb_reg ( in, flush, out, clk, reset, we );
  input [0:178] in;
  output [0:178] out;
  input flush, clk, reset, we;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396;

  DFFR_X1 MEM_WB_REG_out_reg_178_ ( .D(n359), .CK(clk), .RN(n392), .Q(out[178]) );
  DFFR_X1 MEM_WB_REG_out_reg_177_ ( .D(n358), .CK(clk), .RN(n385), .Q(out[177]) );
  DFFR_X1 MEM_WB_REG_out_reg_176_ ( .D(n357), .CK(clk), .RN(n391), .Q(out[176]) );
  DFFR_X1 MEM_WB_REG_out_reg_175_ ( .D(n356), .CK(clk), .RN(n385), .Q(out[175]) );
  DFFR_X1 MEM_WB_REG_out_reg_174_ ( .D(n355), .CK(clk), .RN(n391), .Q(out[174]) );
  DFFR_X1 MEM_WB_REG_out_reg_173_ ( .D(n354), .CK(clk), .RN(n386), .Q(out[173]) );
  DFFR_X1 MEM_WB_REG_out_reg_172_ ( .D(n353), .CK(clk), .RN(n391), .Q(out[172]) );
  DFFR_X1 MEM_WB_REG_out_reg_171_ ( .D(n352), .CK(clk), .RN(n386), .Q(out[171]) );
  DFFR_X1 MEM_WB_REG_out_reg_170_ ( .D(n351), .CK(clk), .RN(n391), .Q(out[170]) );
  DFFR_X1 MEM_WB_REG_out_reg_169_ ( .D(n350), .CK(clk), .RN(n391), .Q(out[169]) );
  DFFR_X1 MEM_WB_REG_out_reg_168_ ( .D(n349), .CK(clk), .RN(n386), .Q(out[168]) );
  DFFR_X1 MEM_WB_REG_out_reg_167_ ( .D(n348), .CK(clk), .RN(n391), .Q(out[167]) );
  DFFR_X1 MEM_WB_REG_out_reg_166_ ( .D(n347), .CK(clk), .RN(n386), .Q(out[166]) );
  DFFR_X1 MEM_WB_REG_out_reg_165_ ( .D(n346), .CK(clk), .RN(n391), .Q(out[165]) );
  DFFR_X1 MEM_WB_REG_out_reg_164_ ( .D(n345), .CK(clk), .RN(n386), .Q(out[164]) );
  DFFR_X1 MEM_WB_REG_out_reg_163_ ( .D(n344), .CK(clk), .RN(n391), .Q(out[163]) );
  DFFR_X1 MEM_WB_REG_out_reg_162_ ( .D(n343), .CK(clk), .RN(n386), .Q(out[162]) );
  DFFR_X1 MEM_WB_REG_out_reg_161_ ( .D(n342), .CK(clk), .RN(n391), .Q(out[161]) );
  DFFR_X1 MEM_WB_REG_out_reg_160_ ( .D(n341), .CK(clk), .RN(n386), .Q(out[160]) );
  DFFR_X1 MEM_WB_REG_out_reg_159_ ( .D(n340), .CK(clk), .RN(n386), .Q(out[159]) );
  DFFR_X1 MEM_WB_REG_out_reg_158_ ( .D(n339), .CK(clk), .RN(n391), .Q(out[158]) );
  DFFR_X1 MEM_WB_REG_out_reg_157_ ( .D(n338), .CK(clk), .RN(n386), .Q(out[157]) );
  DFFR_X1 MEM_WB_REG_out_reg_156_ ( .D(n337), .CK(clk), .RN(n391), .Q(out[156]) );
  DFFR_X1 MEM_WB_REG_out_reg_155_ ( .D(n336), .CK(clk), .RN(n386), .Q(out[155]) );
  DFFR_X1 MEM_WB_REG_out_reg_154_ ( .D(n335), .CK(clk), .RN(n390), .Q(out[154]) );
  DFFR_X1 MEM_WB_REG_out_reg_153_ ( .D(n334), .CK(clk), .RN(n386), .Q(out[153]) );
  DFFR_X1 MEM_WB_REG_out_reg_152_ ( .D(n333), .CK(clk), .RN(n390), .Q(out[152]) );
  DFFR_X1 MEM_WB_REG_out_reg_151_ ( .D(n332), .CK(clk), .RN(n387), .Q(out[151]) );
  DFFR_X1 MEM_WB_REG_out_reg_150_ ( .D(n331), .CK(clk), .RN(n390), .Q(out[150]) );
  DFFR_X1 MEM_WB_REG_out_reg_149_ ( .D(n330), .CK(clk), .RN(n390), .Q(out[149]) );
  DFFR_X1 MEM_WB_REG_out_reg_148_ ( .D(n329), .CK(clk), .RN(n387), .Q(out[148]) );
  DFFR_X1 MEM_WB_REG_out_reg_147_ ( .D(n328), .CK(clk), .RN(n390), .Q(out[147]) );
  DFFR_X1 MEM_WB_REG_out_reg_146_ ( .D(n327), .CK(clk), .RN(n387), .Q(out[146]) );
  DFFR_X1 MEM_WB_REG_out_reg_145_ ( .D(n326), .CK(clk), .RN(n390), .Q(out[145]) );
  DFFR_X1 MEM_WB_REG_out_reg_144_ ( .D(n325), .CK(clk), .RN(n387), .Q(out[144]) );
  DFFR_X1 MEM_WB_REG_out_reg_143_ ( .D(n324), .CK(clk), .RN(n390), .Q(out[143]) );
  DFFR_X1 MEM_WB_REG_out_reg_142_ ( .D(n323), .CK(clk), .RN(n387), .Q(out[142]) );
  DFFR_X1 MEM_WB_REG_out_reg_141_ ( .D(n322), .CK(clk), .RN(n390), .Q(out[141]) );
  DFFR_X1 MEM_WB_REG_out_reg_140_ ( .D(n321), .CK(clk), .RN(n387), .Q(out[140]) );
  DFFR_X1 MEM_WB_REG_out_reg_139_ ( .D(n320), .CK(clk), .RN(n387), .Q(out[139]) );
  DFFR_X1 MEM_WB_REG_out_reg_138_ ( .D(n319), .CK(clk), .RN(n390), .Q(out[138]) );
  DFFR_X1 MEM_WB_REG_out_reg_137_ ( .D(n318), .CK(clk), .RN(n387), .Q(out[137]) );
  DFFR_X1 MEM_WB_REG_out_reg_136_ ( .D(n317), .CK(clk), .RN(n390), .Q(out[136]) );
  DFFR_X1 MEM_WB_REG_out_reg_135_ ( .D(n316), .CK(clk), .RN(n387), .Q(out[135]) );
  DFFR_X1 MEM_WB_REG_out_reg_134_ ( .D(n315), .CK(clk), .RN(n390), .Q(out[134]) );
  DFFR_X1 MEM_WB_REG_out_reg_133_ ( .D(n314), .CK(clk), .RN(n387), .Q(out[133]) );
  DFFR_X1 MEM_WB_REG_out_reg_132_ ( .D(n313), .CK(clk), .RN(reset), .Q(
        out[132]) );
  DFFR_X1 MEM_WB_REG_out_reg_131_ ( .D(n312), .CK(clk), .RN(n387), .Q(out[131]) );
  DFFR_X1 MEM_WB_REG_out_reg_130_ ( .D(n311), .CK(clk), .RN(n390), .Q(out[130]) );
  DFFR_X1 MEM_WB_REG_out_reg_129_ ( .D(n310), .CK(clk), .RN(n391), .Q(out[129]) );
  DFFR_X1 MEM_WB_REG_out_reg_128_ ( .D(n309), .CK(clk), .RN(n388), .Q(out[128]) );
  DFFR_X1 MEM_WB_REG_out_reg_127_ ( .D(n308), .CK(clk), .RN(reset), .Q(
        out[127]) );
  DFFR_X1 MEM_WB_REG_out_reg_126_ ( .D(n307), .CK(clk), .RN(n388), .Q(out[126]) );
  DFFR_X1 MEM_WB_REG_out_reg_125_ ( .D(n306), .CK(clk), .RN(reset), .Q(
        out[125]) );
  DFFR_X1 MEM_WB_REG_out_reg_124_ ( .D(n305), .CK(clk), .RN(n388), .Q(out[124]) );
  DFFR_X1 MEM_WB_REG_out_reg_123_ ( .D(n304), .CK(clk), .RN(n390), .Q(out[123]) );
  DFFR_X1 MEM_WB_REG_out_reg_122_ ( .D(n303), .CK(clk), .RN(n388), .Q(out[122]) );
  DFFR_X1 MEM_WB_REG_out_reg_121_ ( .D(n302), .CK(clk), .RN(n391), .Q(out[121]) );
  DFFR_X1 MEM_WB_REG_out_reg_120_ ( .D(n301), .CK(clk), .RN(n388), .Q(out[120]) );
  DFFR_X1 MEM_WB_REG_out_reg_118_ ( .D(n299), .CK(clk), .RN(n384), .Q(out[118]) );
  DFFR_X1 MEM_WB_REG_out_reg_117_ ( .D(n298), .CK(clk), .RN(n388), .Q(out[117]) );
  DFFR_X1 MEM_WB_REG_out_reg_116_ ( .D(n297), .CK(clk), .RN(n383), .Q(out[116]) );
  DFFR_X1 MEM_WB_REG_out_reg_115_ ( .D(n296), .CK(clk), .RN(n388), .Q(out[115]) );
  DFFR_X1 MEM_WB_REG_out_reg_114_ ( .D(n295), .CK(clk), .RN(n382), .Q(out[114]) );
  DFFR_X1 MEM_WB_REG_out_reg_113_ ( .D(n294), .CK(clk), .RN(n388), .Q(out[113]) );
  DFFR_X1 MEM_WB_REG_out_reg_112_ ( .D(n293), .CK(clk), .RN(n392), .Q(out[112]) );
  DFFR_X1 MEM_WB_REG_out_reg_111_ ( .D(n292), .CK(clk), .RN(n388), .Q(out[111]) );
  DFFR_X1 MEM_WB_REG_out_reg_110_ ( .D(n291), .CK(clk), .RN(n389), .Q(out[110]) );
  DFFR_X1 MEM_WB_REG_out_reg_109_ ( .D(n290), .CK(clk), .RN(n389), .Q(out[109]) );
  DFFR_X1 MEM_WB_REG_out_reg_108_ ( .D(n289), .CK(clk), .RN(n389), .Q(out[108]) );
  DFFR_X1 MEM_WB_REG_out_reg_107_ ( .D(n288), .CK(clk), .RN(n389), .Q(out[107]) );
  DFFR_X1 MEM_WB_REG_out_reg_106_ ( .D(n287), .CK(clk), .RN(n389), .Q(out[106]) );
  DFFR_X1 MEM_WB_REG_out_reg_105_ ( .D(n286), .CK(clk), .RN(n389), .Q(out[105]) );
  DFFR_X1 MEM_WB_REG_out_reg_104_ ( .D(n285), .CK(clk), .RN(n389), .Q(out[104]) );
  DFFR_X1 MEM_WB_REG_out_reg_103_ ( .D(n284), .CK(clk), .RN(n389), .Q(out[103]) );
  DFFR_X1 MEM_WB_REG_out_reg_102_ ( .D(n283), .CK(clk), .RN(n389), .Q(out[102]) );
  DFFR_X1 MEM_WB_REG_out_reg_101_ ( .D(n282), .CK(clk), .RN(n389), .Q(out[101]) );
  DFFR_X1 MEM_WB_REG_out_reg_100_ ( .D(n281), .CK(clk), .RN(n389), .Q(out[100]) );
  DFFR_X1 MEM_WB_REG_out_reg_99_ ( .D(n280), .CK(clk), .RN(n382), .Q(out[99])
         );
  DFFR_X1 MEM_WB_REG_out_reg_98_ ( .D(n279), .CK(clk), .RN(n382), .Q(out[98])
         );
  DFFR_X1 MEM_WB_REG_out_reg_97_ ( .D(n278), .CK(clk), .RN(n382), .Q(out[97])
         );
  DFFR_X1 MEM_WB_REG_out_reg_96_ ( .D(n277), .CK(clk), .RN(n383), .Q(out[96])
         );
  DFFR_X1 MEM_WB_REG_out_reg_95_ ( .D(n276), .CK(clk), .RN(n382), .Q(out[95])
         );
  DFFR_X1 MEM_WB_REG_out_reg_94_ ( .D(n275), .CK(clk), .RN(n384), .Q(out[94])
         );
  DFFR_X1 MEM_WB_REG_out_reg_93_ ( .D(n274), .CK(clk), .RN(n382), .Q(out[93])
         );
  DFFR_X1 MEM_WB_REG_out_reg_92_ ( .D(n273), .CK(clk), .RN(n385), .Q(out[92])
         );
  DFFR_X1 MEM_WB_REG_out_reg_91_ ( .D(n272), .CK(clk), .RN(n382), .Q(out[91])
         );
  DFFR_X1 MEM_WB_REG_out_reg_90_ ( .D(n271), .CK(clk), .RN(n386), .Q(out[90])
         );
  DFFR_X1 MEM_WB_REG_out_reg_89_ ( .D(n270), .CK(clk), .RN(n387), .Q(out[89])
         );
  DFFR_X1 MEM_WB_REG_out_reg_88_ ( .D(n269), .CK(clk), .RN(n382), .Q(out[88])
         );
  DFFR_X1 MEM_WB_REG_out_reg_87_ ( .D(n268), .CK(clk), .RN(n388), .Q(out[87])
         );
  DFFR_X1 MEM_WB_REG_out_reg_86_ ( .D(n267), .CK(clk), .RN(n382), .Q(out[86])
         );
  DFFR_X1 MEM_WB_REG_out_reg_85_ ( .D(n266), .CK(clk), .RN(n389), .Q(out[85])
         );
  DFFR_X1 MEM_WB_REG_out_reg_84_ ( .D(n265), .CK(clk), .RN(n382), .Q(out[84])
         );
  DFFR_X1 MEM_WB_REG_out_reg_83_ ( .D(n264), .CK(clk), .RN(reset), .Q(out[83])
         );
  DFFR_X1 MEM_WB_REG_out_reg_82_ ( .D(n263), .CK(clk), .RN(n382), .Q(out[82])
         );
  DFFR_X1 MEM_WB_REG_out_reg_81_ ( .D(n262), .CK(clk), .RN(n390), .Q(out[81])
         );
  DFFR_X1 MEM_WB_REG_out_reg_80_ ( .D(n261), .CK(clk), .RN(n382), .Q(out[80])
         );
  DFFR_X1 MEM_WB_REG_out_reg_79_ ( .D(n260), .CK(clk), .RN(n382), .Q(out[79])
         );
  DFFR_X1 MEM_WB_REG_out_reg_78_ ( .D(n259), .CK(clk), .RN(n393), .Q(out[78])
         );
  DFFR_X1 MEM_WB_REG_out_reg_77_ ( .D(n258), .CK(clk), .RN(n383), .Q(out[77])
         );
  DFFR_X1 MEM_WB_REG_out_reg_76_ ( .D(n257), .CK(clk), .RN(n393), .Q(out[76])
         );
  DFFR_X1 MEM_WB_REG_out_reg_75_ ( .D(n256), .CK(clk), .RN(n383), .Q(out[75])
         );
  DFFR_X1 MEM_WB_REG_out_reg_74_ ( .D(n255), .CK(clk), .RN(n393), .Q(out[74])
         );
  DFFR_X1 MEM_WB_REG_out_reg_73_ ( .D(n254), .CK(clk), .RN(n383), .Q(out[73])
         );
  DFFR_X1 MEM_WB_REG_out_reg_72_ ( .D(n253), .CK(clk), .RN(n393), .Q(out[72])
         );
  DFFR_X1 MEM_WB_REG_out_reg_71_ ( .D(n252), .CK(clk), .RN(n383), .Q(out[71])
         );
  DFFR_X1 MEM_WB_REG_out_reg_70_ ( .D(n251), .CK(clk), .RN(n393), .Q(out[70])
         );
  DFFR_X1 MEM_WB_REG_out_reg_69_ ( .D(n250), .CK(clk), .RN(n393), .Q(out[69])
         );
  DFFR_X1 MEM_WB_REG_out_reg_68_ ( .D(n249), .CK(clk), .RN(n383), .Q(out[68])
         );
  DFFR_X1 MEM_WB_REG_out_reg_67_ ( .D(n248), .CK(clk), .RN(n393), .Q(out[67])
         );
  DFFR_X1 MEM_WB_REG_out_reg_66_ ( .D(n247), .CK(clk), .RN(n383), .Q(out[66])
         );
  DFFR_X1 MEM_WB_REG_out_reg_65_ ( .D(n246), .CK(clk), .RN(n393), .Q(out[65])
         );
  DFFR_X1 MEM_WB_REG_out_reg_64_ ( .D(n245), .CK(clk), .RN(n383), .Q(out[64])
         );
  DFFR_X1 MEM_WB_REG_out_reg_63_ ( .D(n244), .CK(clk), .RN(n393), .Q(out[63])
         );
  DFFR_X1 MEM_WB_REG_out_reg_62_ ( .D(n243), .CK(clk), .RN(n383), .Q(out[62])
         );
  DFFR_X1 MEM_WB_REG_out_reg_61_ ( .D(n242), .CK(clk), .RN(n393), .Q(out[61])
         );
  DFFR_X1 MEM_WB_REG_out_reg_60_ ( .D(n241), .CK(clk), .RN(n383), .Q(out[60])
         );
  DFFR_X1 MEM_WB_REG_out_reg_59_ ( .D(n240), .CK(clk), .RN(n383), .Q(out[59])
         );
  DFFR_X1 MEM_WB_REG_out_reg_58_ ( .D(n239), .CK(clk), .RN(n392), .Q(out[58])
         );
  DFFR_X1 MEM_WB_REG_out_reg_57_ ( .D(n238), .CK(clk), .RN(n383), .Q(out[57])
         );
  DFFR_X1 MEM_WB_REG_out_reg_56_ ( .D(n237), .CK(clk), .RN(n392), .Q(out[56])
         );
  DFFR_X1 MEM_WB_REG_out_reg_55_ ( .D(n236), .CK(clk), .RN(n384), .Q(out[55])
         );
  DFFR_X1 MEM_WB_REG_out_reg_54_ ( .D(n235), .CK(clk), .RN(n392), .Q(out[54])
         );
  DFFR_X1 MEM_WB_REG_out_reg_53_ ( .D(n234), .CK(clk), .RN(n384), .Q(out[53])
         );
  DFFR_X1 MEM_WB_REG_out_reg_52_ ( .D(n233), .CK(clk), .RN(n392), .Q(out[52])
         );
  DFFR_X1 MEM_WB_REG_out_reg_51_ ( .D(n232), .CK(clk), .RN(n384), .Q(out[51])
         );
  DFFR_X1 MEM_WB_REG_out_reg_50_ ( .D(n231), .CK(clk), .RN(n392), .Q(out[50])
         );
  DFFR_X1 MEM_WB_REG_out_reg_49_ ( .D(n230), .CK(clk), .RN(n392), .Q(out[49])
         );
  DFFR_X1 MEM_WB_REG_out_reg_48_ ( .D(n229), .CK(clk), .RN(n384), .Q(out[48])
         );
  DFFR_X1 MEM_WB_REG_out_reg_47_ ( .D(n228), .CK(clk), .RN(n392), .Q(out[47])
         );
  DFFR_X1 MEM_WB_REG_out_reg_46_ ( .D(n227), .CK(clk), .RN(n384), .Q(out[46])
         );
  DFFR_X1 MEM_WB_REG_out_reg_45_ ( .D(n226), .CK(clk), .RN(n392), .Q(out[45])
         );
  DFFR_X1 MEM_WB_REG_out_reg_44_ ( .D(n225), .CK(clk), .RN(n384), .Q(out[44])
         );
  DFFR_X1 MEM_WB_REG_out_reg_43_ ( .D(n224), .CK(clk), .RN(n392), .Q(out[43])
         );
  DFFR_X1 MEM_WB_REG_out_reg_42_ ( .D(n223), .CK(clk), .RN(n384), .Q(out[42])
         );
  DFFR_X1 MEM_WB_REG_out_reg_41_ ( .D(n222), .CK(clk), .RN(n392), .Q(out[41])
         );
  DFFR_X1 MEM_WB_REG_out_reg_40_ ( .D(n221), .CK(clk), .RN(n384), .Q(out[40])
         );
  DFFR_X1 MEM_WB_REG_out_reg_39_ ( .D(n220), .CK(clk), .RN(n384), .Q(out[39])
         );
  DFFR_X1 MEM_WB_REG_out_reg_38_ ( .D(n219), .CK(clk), .RN(n392), .Q(out[38])
         );
  DFFR_X1 MEM_WB_REG_out_reg_37_ ( .D(n218), .CK(clk), .RN(n384), .Q(out[37])
         );
  DFFR_X1 MEM_WB_REG_out_reg_36_ ( .D(n217), .CK(clk), .RN(n393), .Q(out[36])
         );
  DFFR_X1 MEM_WB_REG_out_reg_35_ ( .D(n216), .CK(clk), .RN(n384), .Q(out[35])
         );
  DFFR_X1 MEM_WB_REG_out_reg_34_ ( .D(n215), .CK(clk), .RN(n384), .Q(out[34])
         );
  DFFR_X1 MEM_WB_REG_out_reg_33_ ( .D(n214), .CK(clk), .RN(n385), .Q(out[33])
         );
  DFFR_X1 MEM_WB_REG_out_reg_32_ ( .D(n213), .CK(clk), .RN(n383), .Q(out[32])
         );
  DFFR_X1 MEM_WB_REG_out_reg_31_ ( .D(n212), .CK(clk), .RN(n385), .Q(out[31])
         );
  DFFR_X1 MEM_WB_REG_out_reg_30_ ( .D(n211), .CK(clk), .RN(n382), .Q(out[30])
         );
  DFFR_X1 MEM_WB_REG_out_reg_29_ ( .D(n210), .CK(clk), .RN(n392), .Q(out[29])
         );
  DFFR_X1 MEM_WB_REG_out_reg_28_ ( .D(n209), .CK(clk), .RN(n385), .Q(out[28])
         );
  DFFR_X1 MEM_WB_REG_out_reg_27_ ( .D(n208), .CK(clk), .RN(n393), .Q(out[27])
         );
  DFFR_X1 MEM_WB_REG_out_reg_26_ ( .D(n207), .CK(clk), .RN(n385), .Q(out[26])
         );
  DFFR_X1 MEM_WB_REG_out_reg_25_ ( .D(n206), .CK(clk), .RN(n385), .Q(out[25])
         );
  DFFR_X1 MEM_WB_REG_out_reg_24_ ( .D(n205), .CK(clk), .RN(n385), .Q(out[24])
         );
  DFFR_X1 MEM_WB_REG_out_reg_23_ ( .D(n204), .CK(clk), .RN(n386), .Q(out[23])
         );
  DFFR_X1 MEM_WB_REG_out_reg_22_ ( .D(n203), .CK(clk), .RN(n385), .Q(out[22])
         );
  DFFR_X1 MEM_WB_REG_out_reg_21_ ( .D(n202), .CK(clk), .RN(n387), .Q(out[21])
         );
  DFFR_X1 MEM_WB_REG_out_reg_20_ ( .D(n201), .CK(clk), .RN(n385), .Q(out[20])
         );
  DFFR_X1 MEM_WB_REG_out_reg_19_ ( .D(n200), .CK(clk), .RN(n385), .Q(out[19])
         );
  DFFR_X1 MEM_WB_REG_out_reg_18_ ( .D(n199), .CK(clk), .RN(n388), .Q(out[18])
         );
  DFFR_X1 MEM_WB_REG_out_reg_17_ ( .D(n198), .CK(clk), .RN(n385), .Q(out[17])
         );
  DFFR_X1 MEM_WB_REG_out_reg_16_ ( .D(n197), .CK(clk), .RN(n386), .Q(out[16])
         );
  DFFR_X1 MEM_WB_REG_out_reg_15_ ( .D(n196), .CK(clk), .RN(n391), .Q(out[15])
         );
  DFFR_X1 MEM_WB_REG_out_reg_14_ ( .D(n195), .CK(clk), .RN(n387), .Q(out[14])
         );
  DFFR_X1 MEM_WB_REG_out_reg_13_ ( .D(n194), .CK(clk), .RN(n390), .Q(out[13])
         );
  DFFR_X1 MEM_WB_REG_out_reg_12_ ( .D(n193), .CK(clk), .RN(n388), .Q(out[12])
         );
  DFFR_X1 MEM_WB_REG_out_reg_11_ ( .D(n192), .CK(clk), .RN(n393), .Q(out[11])
         );
  DFFR_X1 MEM_WB_REG_out_reg_10_ ( .D(n191), .CK(clk), .RN(n388), .Q(out[10])
         );
  DFFR_X1 MEM_WB_REG_out_reg_8_ ( .D(n189), .CK(clk), .RN(n382), .Q(out[8]) );
  DFFR_X1 MEM_WB_REG_out_reg_7_ ( .D(n188), .CK(clk), .RN(n393), .Q(out[7]) );
  DFFR_X1 MEM_WB_REG_out_reg_6_ ( .D(n187), .CK(clk), .RN(n383), .Q(out[6]) );
  DFFR_X1 MEM_WB_REG_out_reg_5_ ( .D(n186), .CK(clk), .RN(n393), .Q(out[5]) );
  DFFR_X1 MEM_WB_REG_out_reg_4_ ( .D(n185), .CK(clk), .RN(n384), .Q(out[4]) );
  DFFR_X1 MEM_WB_REG_out_reg_3_ ( .D(n184), .CK(clk), .RN(n392), .Q(out[3]) );
  DFFR_X1 MEM_WB_REG_out_reg_2_ ( .D(n183), .CK(clk), .RN(n385), .Q(out[2]) );
  DFFR_X1 MEM_WB_REG_out_reg_1_ ( .D(n182), .CK(clk), .RN(n389), .Q(out[1]) );
  DFFR_X1 MEM_WB_REG_out_reg_0_ ( .D(n181), .CK(clk), .RN(n389), .Q(out[0]) );
  INV_X1 U2 ( .A(n1), .ZN(n190) );
  AOI22_X1 U3 ( .A1(in[9]), .A2(n381), .B1(n360), .B2(out[9]), .ZN(n1) );
  INV_X1 U4 ( .A(n3), .ZN(n280) );
  AOI22_X1 U5 ( .A1(in[99]), .A2(n381), .B1(out[99]), .B2(n360), .ZN(n3) );
  INV_X1 U6 ( .A(n4), .ZN(n279) );
  AOI22_X1 U7 ( .A1(in[98]), .A2(n381), .B1(out[98]), .B2(n360), .ZN(n4) );
  INV_X1 U8 ( .A(n5), .ZN(n278) );
  AOI22_X1 U9 ( .A1(in[97]), .A2(n381), .B1(out[97]), .B2(n360), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(n277) );
  AOI22_X1 U11 ( .A1(in[96]), .A2(n381), .B1(out[96]), .B2(n360), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(n276) );
  AOI22_X1 U13 ( .A1(in[95]), .A2(n381), .B1(out[95]), .B2(n360), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(n275) );
  AOI22_X1 U15 ( .A1(in[94]), .A2(n381), .B1(out[94]), .B2(n360), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(n274) );
  AOI22_X1 U17 ( .A1(in[93]), .A2(n381), .B1(out[93]), .B2(n360), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(n273) );
  AOI22_X1 U19 ( .A1(in[92]), .A2(n381), .B1(out[92]), .B2(n360), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(n272) );
  AOI22_X1 U21 ( .A1(in[91]), .A2(n381), .B1(out[91]), .B2(n360), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(n271) );
  AOI22_X1 U23 ( .A1(in[90]), .A2(n381), .B1(out[90]), .B2(n360), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(n189) );
  AOI22_X1 U25 ( .A1(in[8]), .A2(n381), .B1(out[8]), .B2(n360), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(n270) );
  AOI22_X1 U27 ( .A1(in[89]), .A2(n381), .B1(out[89]), .B2(n361), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(n269) );
  AOI22_X1 U29 ( .A1(in[88]), .A2(n381), .B1(out[88]), .B2(n360), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(n268) );
  AOI22_X1 U31 ( .A1(in[87]), .A2(n381), .B1(out[87]), .B2(n361), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(n267) );
  AOI22_X1 U33 ( .A1(in[86]), .A2(n381), .B1(out[86]), .B2(n360), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(n266) );
  AOI22_X1 U35 ( .A1(in[85]), .A2(n381), .B1(out[85]), .B2(n361), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(n265) );
  AOI22_X1 U37 ( .A1(in[84]), .A2(n380), .B1(out[84]), .B2(n360), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(n264) );
  AOI22_X1 U39 ( .A1(in[83]), .A2(n380), .B1(out[83]), .B2(n361), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(n263) );
  AOI22_X1 U41 ( .A1(in[82]), .A2(n380), .B1(out[82]), .B2(n360), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(n262) );
  AOI22_X1 U43 ( .A1(in[81]), .A2(n380), .B1(out[81]), .B2(n361), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(n261) );
  AOI22_X1 U45 ( .A1(in[80]), .A2(n380), .B1(out[80]), .B2(n360), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(n188) );
  AOI22_X1 U47 ( .A1(in[7]), .A2(n380), .B1(out[7]), .B2(n361), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(n260) );
  AOI22_X1 U49 ( .A1(in[79]), .A2(n380), .B1(out[79]), .B2(n360), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(n259) );
  AOI22_X1 U51 ( .A1(in[78]), .A2(n380), .B1(out[78]), .B2(n361), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(n258) );
  AOI22_X1 U53 ( .A1(in[77]), .A2(n380), .B1(out[77]), .B2(n361), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(n257) );
  AOI22_X1 U55 ( .A1(in[76]), .A2(n380), .B1(out[76]), .B2(n361), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(n256) );
  AOI22_X1 U57 ( .A1(in[75]), .A2(n380), .B1(out[75]), .B2(n361), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(n255) );
  AOI22_X1 U59 ( .A1(in[74]), .A2(n380), .B1(out[74]), .B2(n361), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(n254) );
  AOI22_X1 U61 ( .A1(in[73]), .A2(n380), .B1(out[73]), .B2(n361), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(n253) );
  AOI22_X1 U63 ( .A1(in[72]), .A2(n380), .B1(out[72]), .B2(n361), .ZN(n32) );
  INV_X1 U64 ( .A(n33), .ZN(n252) );
  AOI22_X1 U65 ( .A1(in[71]), .A2(n380), .B1(out[71]), .B2(n361), .ZN(n33) );
  INV_X1 U66 ( .A(n34), .ZN(n251) );
  AOI22_X1 U67 ( .A1(in[70]), .A2(n380), .B1(out[70]), .B2(n361), .ZN(n34) );
  INV_X1 U68 ( .A(n35), .ZN(n187) );
  AOI22_X1 U69 ( .A1(in[6]), .A2(n380), .B1(out[6]), .B2(n361), .ZN(n35) );
  INV_X1 U70 ( .A(n36), .ZN(n250) );
  AOI22_X1 U71 ( .A1(in[69]), .A2(n380), .B1(out[69]), .B2(n361), .ZN(n36) );
  INV_X1 U72 ( .A(n37), .ZN(n249) );
  AOI22_X1 U73 ( .A1(in[68]), .A2(n380), .B1(out[68]), .B2(n361), .ZN(n37) );
  INV_X1 U74 ( .A(n38), .ZN(n248) );
  AOI22_X1 U75 ( .A1(in[67]), .A2(n380), .B1(out[67]), .B2(n363), .ZN(n38) );
  INV_X1 U76 ( .A(n39), .ZN(n247) );
  AOI22_X1 U77 ( .A1(in[66]), .A2(n380), .B1(out[66]), .B2(n362), .ZN(n39) );
  INV_X1 U78 ( .A(n40), .ZN(n246) );
  AOI22_X1 U79 ( .A1(in[65]), .A2(n380), .B1(out[65]), .B2(n363), .ZN(n40) );
  INV_X1 U80 ( .A(n41), .ZN(n245) );
  AOI22_X1 U81 ( .A1(in[64]), .A2(n380), .B1(out[64]), .B2(n362), .ZN(n41) );
  INV_X1 U82 ( .A(n42), .ZN(n244) );
  AOI22_X1 U83 ( .A1(in[63]), .A2(n380), .B1(out[63]), .B2(n363), .ZN(n42) );
  INV_X1 U84 ( .A(n43), .ZN(n243) );
  AOI22_X1 U85 ( .A1(in[62]), .A2(n380), .B1(out[62]), .B2(n362), .ZN(n43) );
  INV_X1 U86 ( .A(n44), .ZN(n242) );
  AOI22_X1 U87 ( .A1(in[61]), .A2(n380), .B1(out[61]), .B2(n363), .ZN(n44) );
  INV_X1 U88 ( .A(n45), .ZN(n241) );
  AOI22_X1 U89 ( .A1(in[60]), .A2(n380), .B1(out[60]), .B2(n362), .ZN(n45) );
  INV_X1 U90 ( .A(n46), .ZN(n186) );
  AOI22_X1 U91 ( .A1(in[5]), .A2(n379), .B1(out[5]), .B2(n363), .ZN(n46) );
  INV_X1 U92 ( .A(n47), .ZN(n240) );
  AOI22_X1 U93 ( .A1(in[59]), .A2(n379), .B1(out[59]), .B2(n362), .ZN(n47) );
  INV_X1 U94 ( .A(n48), .ZN(n239) );
  AOI22_X1 U95 ( .A1(in[58]), .A2(n379), .B1(out[58]), .B2(n363), .ZN(n48) );
  INV_X1 U96 ( .A(n49), .ZN(n238) );
  AOI22_X1 U97 ( .A1(in[57]), .A2(n379), .B1(out[57]), .B2(n362), .ZN(n49) );
  INV_X1 U98 ( .A(n50), .ZN(n237) );
  AOI22_X1 U99 ( .A1(in[56]), .A2(n379), .B1(out[56]), .B2(n362), .ZN(n50) );
  INV_X1 U100 ( .A(n51), .ZN(n236) );
  AOI22_X1 U101 ( .A1(in[55]), .A2(n379), .B1(out[55]), .B2(n362), .ZN(n51) );
  INV_X1 U102 ( .A(n52), .ZN(n235) );
  AOI22_X1 U103 ( .A1(in[54]), .A2(n379), .B1(out[54]), .B2(n362), .ZN(n52) );
  INV_X1 U104 ( .A(n53), .ZN(n234) );
  AOI22_X1 U105 ( .A1(in[53]), .A2(n379), .B1(out[53]), .B2(n362), .ZN(n53) );
  INV_X1 U106 ( .A(n54), .ZN(n233) );
  AOI22_X1 U107 ( .A1(in[52]), .A2(n379), .B1(out[52]), .B2(n362), .ZN(n54) );
  INV_X1 U108 ( .A(n55), .ZN(n232) );
  AOI22_X1 U109 ( .A1(in[51]), .A2(n379), .B1(out[51]), .B2(n362), .ZN(n55) );
  INV_X1 U110 ( .A(n56), .ZN(n231) );
  AOI22_X1 U111 ( .A1(in[50]), .A2(n379), .B1(out[50]), .B2(n362), .ZN(n56) );
  INV_X1 U112 ( .A(n57), .ZN(n185) );
  AOI22_X1 U113 ( .A1(in[4]), .A2(n379), .B1(out[4]), .B2(n362), .ZN(n57) );
  INV_X1 U114 ( .A(n58), .ZN(n230) );
  AOI22_X1 U115 ( .A1(in[49]), .A2(n379), .B1(out[49]), .B2(n362), .ZN(n58) );
  INV_X1 U116 ( .A(n59), .ZN(n229) );
  AOI22_X1 U117 ( .A1(in[48]), .A2(n379), .B1(out[48]), .B2(n362), .ZN(n59) );
  INV_X1 U118 ( .A(n60), .ZN(n228) );
  AOI22_X1 U119 ( .A1(in[47]), .A2(n379), .B1(out[47]), .B2(n362), .ZN(n60) );
  INV_X1 U120 ( .A(n61), .ZN(n227) );
  AOI22_X1 U121 ( .A1(in[46]), .A2(n379), .B1(out[46]), .B2(n362), .ZN(n61) );
  INV_X1 U122 ( .A(n62), .ZN(n226) );
  AOI22_X1 U123 ( .A1(in[45]), .A2(n379), .B1(out[45]), .B2(n363), .ZN(n62) );
  INV_X1 U124 ( .A(n63), .ZN(n225) );
  AOI22_X1 U125 ( .A1(in[44]), .A2(n379), .B1(out[44]), .B2(n363), .ZN(n63) );
  INV_X1 U126 ( .A(n64), .ZN(n224) );
  AOI22_X1 U127 ( .A1(in[43]), .A2(n379), .B1(out[43]), .B2(n363), .ZN(n64) );
  INV_X1 U128 ( .A(n65), .ZN(n223) );
  AOI22_X1 U129 ( .A1(in[42]), .A2(n379), .B1(out[42]), .B2(n363), .ZN(n65) );
  INV_X1 U130 ( .A(n66), .ZN(n222) );
  AOI22_X1 U131 ( .A1(in[41]), .A2(n379), .B1(out[41]), .B2(n363), .ZN(n66) );
  INV_X1 U132 ( .A(n67), .ZN(n221) );
  AOI22_X1 U133 ( .A1(in[40]), .A2(n379), .B1(out[40]), .B2(n363), .ZN(n67) );
  INV_X1 U134 ( .A(n68), .ZN(n184) );
  AOI22_X1 U135 ( .A1(in[3]), .A2(n379), .B1(out[3]), .B2(n363), .ZN(n68) );
  INV_X1 U136 ( .A(n69), .ZN(n220) );
  AOI22_X1 U137 ( .A1(in[39]), .A2(n379), .B1(out[39]), .B2(n363), .ZN(n69) );
  INV_X1 U138 ( .A(n70), .ZN(n219) );
  AOI22_X1 U139 ( .A1(in[38]), .A2(n379), .B1(out[38]), .B2(n363), .ZN(n70) );
  INV_X1 U140 ( .A(n71), .ZN(n218) );
  AOI22_X1 U141 ( .A1(in[37]), .A2(n379), .B1(out[37]), .B2(n363), .ZN(n71) );
  INV_X1 U142 ( .A(n72), .ZN(n217) );
  AOI22_X1 U143 ( .A1(in[36]), .A2(n379), .B1(out[36]), .B2(n363), .ZN(n72) );
  INV_X1 U144 ( .A(n73), .ZN(n216) );
  AOI22_X1 U145 ( .A1(in[35]), .A2(n378), .B1(out[35]), .B2(n363), .ZN(n73) );
  INV_X1 U146 ( .A(n74), .ZN(n215) );
  AOI22_X1 U147 ( .A1(in[34]), .A2(n378), .B1(out[34]), .B2(n365), .ZN(n74) );
  INV_X1 U148 ( .A(n75), .ZN(n214) );
  AOI22_X1 U149 ( .A1(in[33]), .A2(n378), .B1(out[33]), .B2(n364), .ZN(n75) );
  INV_X1 U150 ( .A(n76), .ZN(n213) );
  AOI22_X1 U151 ( .A1(in[32]), .A2(n378), .B1(out[32]), .B2(n365), .ZN(n76) );
  INV_X1 U152 ( .A(n77), .ZN(n212) );
  AOI22_X1 U153 ( .A1(in[31]), .A2(n378), .B1(out[31]), .B2(n364), .ZN(n77) );
  INV_X1 U154 ( .A(n78), .ZN(n211) );
  AOI22_X1 U155 ( .A1(in[30]), .A2(n378), .B1(out[30]), .B2(n365), .ZN(n78) );
  INV_X1 U156 ( .A(n79), .ZN(n183) );
  AOI22_X1 U157 ( .A1(in[2]), .A2(n378), .B1(out[2]), .B2(n364), .ZN(n79) );
  INV_X1 U158 ( .A(n80), .ZN(n210) );
  AOI22_X1 U159 ( .A1(in[29]), .A2(n378), .B1(out[29]), .B2(n365), .ZN(n80) );
  INV_X1 U160 ( .A(n81), .ZN(n209) );
  AOI22_X1 U161 ( .A1(in[28]), .A2(n378), .B1(out[28]), .B2(n364), .ZN(n81) );
  INV_X1 U162 ( .A(n82), .ZN(n208) );
  AOI22_X1 U163 ( .A1(in[27]), .A2(n378), .B1(out[27]), .B2(n365), .ZN(n82) );
  INV_X1 U164 ( .A(n83), .ZN(n207) );
  AOI22_X1 U165 ( .A1(in[26]), .A2(n378), .B1(out[26]), .B2(n364), .ZN(n83) );
  INV_X1 U166 ( .A(n84), .ZN(n206) );
  AOI22_X1 U167 ( .A1(in[25]), .A2(n378), .B1(out[25]), .B2(n365), .ZN(n84) );
  INV_X1 U168 ( .A(n85), .ZN(n205) );
  AOI22_X1 U169 ( .A1(in[24]), .A2(n378), .B1(out[24]), .B2(n364), .ZN(n85) );
  INV_X1 U170 ( .A(n86), .ZN(n204) );
  AOI22_X1 U171 ( .A1(in[23]), .A2(n378), .B1(out[23]), .B2(n364), .ZN(n86) );
  INV_X1 U172 ( .A(n87), .ZN(n203) );
  AOI22_X1 U173 ( .A1(in[22]), .A2(n378), .B1(out[22]), .B2(n364), .ZN(n87) );
  INV_X1 U174 ( .A(n88), .ZN(n202) );
  AOI22_X1 U175 ( .A1(in[21]), .A2(n378), .B1(out[21]), .B2(n364), .ZN(n88) );
  INV_X1 U176 ( .A(n89), .ZN(n201) );
  AOI22_X1 U177 ( .A1(in[20]), .A2(n378), .B1(out[20]), .B2(n364), .ZN(n89) );
  INV_X1 U178 ( .A(n90), .ZN(n182) );
  AOI22_X1 U179 ( .A1(in[1]), .A2(n378), .B1(out[1]), .B2(n364), .ZN(n90) );
  INV_X1 U180 ( .A(n91), .ZN(n200) );
  AOI22_X1 U181 ( .A1(in[19]), .A2(n378), .B1(out[19]), .B2(n364), .ZN(n91) );
  INV_X1 U182 ( .A(n92), .ZN(n199) );
  AOI22_X1 U183 ( .A1(in[18]), .A2(n378), .B1(out[18]), .B2(n364), .ZN(n92) );
  INV_X1 U184 ( .A(n93), .ZN(n198) );
  AOI22_X1 U185 ( .A1(in[17]), .A2(n378), .B1(out[17]), .B2(n364), .ZN(n93) );
  INV_X1 U186 ( .A(n94), .ZN(n359) );
  AOI22_X1 U187 ( .A1(in[178]), .A2(n378), .B1(out[178]), .B2(n364), .ZN(n94)
         );
  INV_X1 U188 ( .A(n95), .ZN(n358) );
  AOI22_X1 U189 ( .A1(in[177]), .A2(n378), .B1(out[177]), .B2(n364), .ZN(n95)
         );
  INV_X1 U190 ( .A(n96), .ZN(n357) );
  AOI22_X1 U191 ( .A1(in[176]), .A2(n378), .B1(out[176]), .B2(n364), .ZN(n96)
         );
  INV_X1 U192 ( .A(n97), .ZN(n356) );
  AOI22_X1 U193 ( .A1(in[175]), .A2(n378), .B1(out[175]), .B2(n364), .ZN(n97)
         );
  INV_X1 U194 ( .A(n98), .ZN(n355) );
  AOI22_X1 U195 ( .A1(in[174]), .A2(n378), .B1(out[174]), .B2(n365), .ZN(n98)
         );
  INV_X1 U196 ( .A(n99), .ZN(n354) );
  AOI22_X1 U197 ( .A1(in[173]), .A2(n378), .B1(out[173]), .B2(n365), .ZN(n99)
         );
  INV_X1 U198 ( .A(n100), .ZN(n353) );
  AOI22_X1 U199 ( .A1(in[172]), .A2(n377), .B1(out[172]), .B2(n365), .ZN(n100)
         );
  INV_X1 U200 ( .A(n101), .ZN(n352) );
  AOI22_X1 U201 ( .A1(in[171]), .A2(n377), .B1(out[171]), .B2(n365), .ZN(n101)
         );
  INV_X1 U202 ( .A(n102), .ZN(n351) );
  AOI22_X1 U203 ( .A1(in[170]), .A2(n377), .B1(out[170]), .B2(n365), .ZN(n102)
         );
  INV_X1 U204 ( .A(n103), .ZN(n197) );
  AOI22_X1 U205 ( .A1(in[16]), .A2(n377), .B1(out[16]), .B2(n365), .ZN(n103)
         );
  INV_X1 U206 ( .A(n104), .ZN(n350) );
  AOI22_X1 U207 ( .A1(in[169]), .A2(n377), .B1(out[169]), .B2(n365), .ZN(n104)
         );
  INV_X1 U208 ( .A(n105), .ZN(n349) );
  AOI22_X1 U209 ( .A1(in[168]), .A2(n377), .B1(out[168]), .B2(n365), .ZN(n105)
         );
  INV_X1 U210 ( .A(n106), .ZN(n348) );
  AOI22_X1 U211 ( .A1(in[167]), .A2(n377), .B1(out[167]), .B2(n365), .ZN(n106)
         );
  INV_X1 U212 ( .A(n107), .ZN(n347) );
  AOI22_X1 U213 ( .A1(in[166]), .A2(n377), .B1(out[166]), .B2(n365), .ZN(n107)
         );
  INV_X1 U214 ( .A(n108), .ZN(n346) );
  AOI22_X1 U215 ( .A1(in[165]), .A2(n377), .B1(out[165]), .B2(n365), .ZN(n108)
         );
  INV_X1 U216 ( .A(n109), .ZN(n345) );
  AOI22_X1 U217 ( .A1(in[164]), .A2(n377), .B1(out[164]), .B2(n365), .ZN(n109)
         );
  INV_X1 U218 ( .A(n110), .ZN(n344) );
  AOI22_X1 U219 ( .A1(in[163]), .A2(n377), .B1(out[163]), .B2(n367), .ZN(n110)
         );
  INV_X1 U220 ( .A(n111), .ZN(n343) );
  AOI22_X1 U221 ( .A1(in[162]), .A2(n377), .B1(out[162]), .B2(n366), .ZN(n111)
         );
  INV_X1 U222 ( .A(n112), .ZN(n342) );
  AOI22_X1 U223 ( .A1(in[161]), .A2(n377), .B1(out[161]), .B2(n367), .ZN(n112)
         );
  INV_X1 U224 ( .A(n113), .ZN(n341) );
  AOI22_X1 U225 ( .A1(in[160]), .A2(n377), .B1(out[160]), .B2(n366), .ZN(n113)
         );
  INV_X1 U226 ( .A(n114), .ZN(n196) );
  AOI22_X1 U227 ( .A1(in[15]), .A2(n377), .B1(out[15]), .B2(n367), .ZN(n114)
         );
  INV_X1 U228 ( .A(n115), .ZN(n340) );
  AOI22_X1 U229 ( .A1(in[159]), .A2(n377), .B1(out[159]), .B2(n366), .ZN(n115)
         );
  INV_X1 U230 ( .A(n116), .ZN(n339) );
  AOI22_X1 U231 ( .A1(in[158]), .A2(n377), .B1(out[158]), .B2(n367), .ZN(n116)
         );
  INV_X1 U232 ( .A(n117), .ZN(n338) );
  AOI22_X1 U233 ( .A1(in[157]), .A2(n377), .B1(out[157]), .B2(n366), .ZN(n117)
         );
  INV_X1 U234 ( .A(n118), .ZN(n337) );
  AOI22_X1 U235 ( .A1(in[156]), .A2(n377), .B1(out[156]), .B2(n367), .ZN(n118)
         );
  INV_X1 U236 ( .A(n119), .ZN(n336) );
  AOI22_X1 U237 ( .A1(in[155]), .A2(n377), .B1(out[155]), .B2(n366), .ZN(n119)
         );
  INV_X1 U238 ( .A(n120), .ZN(n335) );
  AOI22_X1 U239 ( .A1(in[154]), .A2(n377), .B1(out[154]), .B2(n367), .ZN(n120)
         );
  INV_X1 U240 ( .A(n121), .ZN(n334) );
  AOI22_X1 U241 ( .A1(in[153]), .A2(n377), .B1(out[153]), .B2(n366), .ZN(n121)
         );
  INV_X1 U242 ( .A(n122), .ZN(n333) );
  AOI22_X1 U243 ( .A1(in[152]), .A2(n377), .B1(out[152]), .B2(n366), .ZN(n122)
         );
  INV_X1 U244 ( .A(n123), .ZN(n332) );
  AOI22_X1 U245 ( .A1(in[151]), .A2(n377), .B1(out[151]), .B2(n366), .ZN(n123)
         );
  INV_X1 U246 ( .A(n124), .ZN(n331) );
  AOI22_X1 U247 ( .A1(in[150]), .A2(n377), .B1(out[150]), .B2(n366), .ZN(n124)
         );
  INV_X1 U248 ( .A(n125), .ZN(n195) );
  AOI22_X1 U249 ( .A1(in[14]), .A2(n377), .B1(out[14]), .B2(n366), .ZN(n125)
         );
  INV_X1 U250 ( .A(n126), .ZN(n330) );
  AOI22_X1 U251 ( .A1(in[149]), .A2(n377), .B1(out[149]), .B2(n366), .ZN(n126)
         );
  INV_X1 U252 ( .A(n127), .ZN(n329) );
  AOI22_X1 U253 ( .A1(in[148]), .A2(n376), .B1(out[148]), .B2(n366), .ZN(n127)
         );
  INV_X1 U254 ( .A(n128), .ZN(n328) );
  AOI22_X1 U255 ( .A1(in[147]), .A2(n376), .B1(out[147]), .B2(n366), .ZN(n128)
         );
  INV_X1 U256 ( .A(n129), .ZN(n327) );
  AOI22_X1 U257 ( .A1(in[146]), .A2(n376), .B1(out[146]), .B2(n366), .ZN(n129)
         );
  INV_X1 U258 ( .A(n130), .ZN(n326) );
  AOI22_X1 U259 ( .A1(in[145]), .A2(n376), .B1(out[145]), .B2(n366), .ZN(n130)
         );
  INV_X1 U260 ( .A(n131), .ZN(n325) );
  AOI22_X1 U261 ( .A1(in[144]), .A2(n376), .B1(out[144]), .B2(n366), .ZN(n131)
         );
  INV_X1 U262 ( .A(n132), .ZN(n324) );
  AOI22_X1 U263 ( .A1(in[143]), .A2(n376), .B1(out[143]), .B2(n366), .ZN(n132)
         );
  INV_X1 U264 ( .A(n133), .ZN(n323) );
  AOI22_X1 U265 ( .A1(in[142]), .A2(n376), .B1(out[142]), .B2(n366), .ZN(n133)
         );
  INV_X1 U266 ( .A(n134), .ZN(n322) );
  AOI22_X1 U267 ( .A1(in[141]), .A2(n376), .B1(out[141]), .B2(n367), .ZN(n134)
         );
  INV_X1 U268 ( .A(n135), .ZN(n321) );
  AOI22_X1 U269 ( .A1(in[140]), .A2(n376), .B1(out[140]), .B2(n367), .ZN(n135)
         );
  INV_X1 U270 ( .A(n136), .ZN(n194) );
  AOI22_X1 U271 ( .A1(in[13]), .A2(n376), .B1(out[13]), .B2(n367), .ZN(n136)
         );
  INV_X1 U272 ( .A(n137), .ZN(n320) );
  AOI22_X1 U273 ( .A1(in[139]), .A2(n376), .B1(out[139]), .B2(n367), .ZN(n137)
         );
  INV_X1 U274 ( .A(n138), .ZN(n319) );
  AOI22_X1 U275 ( .A1(in[138]), .A2(n376), .B1(out[138]), .B2(n367), .ZN(n138)
         );
  INV_X1 U276 ( .A(n139), .ZN(n318) );
  AOI22_X1 U277 ( .A1(in[137]), .A2(n376), .B1(out[137]), .B2(n367), .ZN(n139)
         );
  INV_X1 U278 ( .A(n140), .ZN(n317) );
  AOI22_X1 U279 ( .A1(in[136]), .A2(n376), .B1(out[136]), .B2(n367), .ZN(n140)
         );
  INV_X1 U280 ( .A(n141), .ZN(n316) );
  AOI22_X1 U281 ( .A1(in[135]), .A2(n376), .B1(out[135]), .B2(n367), .ZN(n141)
         );
  INV_X1 U282 ( .A(n142), .ZN(n315) );
  AOI22_X1 U283 ( .A1(in[134]), .A2(n376), .B1(out[134]), .B2(n367), .ZN(n142)
         );
  INV_X1 U284 ( .A(n143), .ZN(n314) );
  AOI22_X1 U285 ( .A1(in[133]), .A2(n376), .B1(out[133]), .B2(n367), .ZN(n143)
         );
  INV_X1 U286 ( .A(n144), .ZN(n313) );
  AOI22_X1 U287 ( .A1(in[132]), .A2(n376), .B1(out[132]), .B2(n367), .ZN(n144)
         );
  INV_X1 U288 ( .A(n145), .ZN(n312) );
  AOI22_X1 U289 ( .A1(in[131]), .A2(n376), .B1(out[131]), .B2(n367), .ZN(n145)
         );
  INV_X1 U290 ( .A(n146), .ZN(n311) );
  AOI22_X1 U291 ( .A1(in[130]), .A2(n376), .B1(out[130]), .B2(n368), .ZN(n146)
         );
  INV_X1 U292 ( .A(n147), .ZN(n193) );
  AOI22_X1 U293 ( .A1(in[12]), .A2(n376), .B1(out[12]), .B2(n368), .ZN(n147)
         );
  INV_X1 U294 ( .A(n148), .ZN(n310) );
  AOI22_X1 U295 ( .A1(in[129]), .A2(n376), .B1(out[129]), .B2(n368), .ZN(n148)
         );
  INV_X1 U296 ( .A(n149), .ZN(n309) );
  AOI22_X1 U297 ( .A1(in[128]), .A2(n376), .B1(out[128]), .B2(n368), .ZN(n149)
         );
  INV_X1 U298 ( .A(n150), .ZN(n308) );
  AOI22_X1 U299 ( .A1(in[127]), .A2(n376), .B1(out[127]), .B2(n368), .ZN(n150)
         );
  INV_X1 U300 ( .A(n151), .ZN(n307) );
  AOI22_X1 U301 ( .A1(in[126]), .A2(n376), .B1(out[126]), .B2(n368), .ZN(n151)
         );
  INV_X1 U302 ( .A(n152), .ZN(n306) );
  AOI22_X1 U303 ( .A1(in[125]), .A2(n376), .B1(out[125]), .B2(n368), .ZN(n152)
         );
  INV_X1 U304 ( .A(n153), .ZN(n305) );
  AOI22_X1 U305 ( .A1(in[124]), .A2(n376), .B1(out[124]), .B2(n368), .ZN(n153)
         );
  INV_X1 U306 ( .A(n154), .ZN(n304) );
  AOI22_X1 U307 ( .A1(in[123]), .A2(n375), .B1(out[123]), .B2(n368), .ZN(n154)
         );
  INV_X1 U308 ( .A(n155), .ZN(n303) );
  AOI22_X1 U309 ( .A1(in[122]), .A2(n375), .B1(out[122]), .B2(n368), .ZN(n155)
         );
  INV_X1 U310 ( .A(n156), .ZN(n302) );
  AOI22_X1 U311 ( .A1(in[121]), .A2(n375), .B1(out[121]), .B2(n368), .ZN(n156)
         );
  INV_X1 U312 ( .A(n157), .ZN(n301) );
  AOI22_X1 U313 ( .A1(in[120]), .A2(n375), .B1(out[120]), .B2(n368), .ZN(n157)
         );
  INV_X1 U314 ( .A(n158), .ZN(n192) );
  AOI22_X1 U315 ( .A1(in[11]), .A2(n375), .B1(out[11]), .B2(n369), .ZN(n158)
         );
  INV_X1 U316 ( .A(n159), .ZN(n300) );
  AOI22_X1 U317 ( .A1(in[119]), .A2(n375), .B1(out[119]), .B2(n369), .ZN(n159)
         );
  INV_X1 U318 ( .A(n160), .ZN(n299) );
  AOI22_X1 U319 ( .A1(in[118]), .A2(n375), .B1(out[118]), .B2(n369), .ZN(n160)
         );
  INV_X1 U320 ( .A(n161), .ZN(n298) );
  AOI22_X1 U321 ( .A1(in[117]), .A2(n375), .B1(out[117]), .B2(n369), .ZN(n161)
         );
  INV_X1 U322 ( .A(n162), .ZN(n297) );
  AOI22_X1 U323 ( .A1(in[116]), .A2(n375), .B1(out[116]), .B2(n369), .ZN(n162)
         );
  INV_X1 U324 ( .A(n163), .ZN(n296) );
  AOI22_X1 U325 ( .A1(in[115]), .A2(n375), .B1(out[115]), .B2(n369), .ZN(n163)
         );
  INV_X1 U326 ( .A(n164), .ZN(n295) );
  AOI22_X1 U327 ( .A1(in[114]), .A2(n375), .B1(out[114]), .B2(n369), .ZN(n164)
         );
  INV_X1 U328 ( .A(n165), .ZN(n294) );
  AOI22_X1 U329 ( .A1(in[113]), .A2(n375), .B1(out[113]), .B2(n369), .ZN(n165)
         );
  INV_X1 U330 ( .A(n166), .ZN(n293) );
  AOI22_X1 U331 ( .A1(in[112]), .A2(n375), .B1(out[112]), .B2(n369), .ZN(n166)
         );
  INV_X1 U332 ( .A(n167), .ZN(n292) );
  AOI22_X1 U333 ( .A1(in[111]), .A2(n375), .B1(out[111]), .B2(n369), .ZN(n167)
         );
  INV_X1 U334 ( .A(n168), .ZN(n291) );
  AOI22_X1 U335 ( .A1(in[110]), .A2(n375), .B1(out[110]), .B2(n369), .ZN(n168)
         );
  INV_X1 U336 ( .A(n169), .ZN(n191) );
  AOI22_X1 U337 ( .A1(in[10]), .A2(n375), .B1(out[10]), .B2(n369), .ZN(n169)
         );
  INV_X1 U338 ( .A(n170), .ZN(n290) );
  AOI22_X1 U339 ( .A1(in[109]), .A2(n375), .B1(out[109]), .B2(n368), .ZN(n170)
         );
  INV_X1 U340 ( .A(n171), .ZN(n289) );
  AOI22_X1 U341 ( .A1(in[108]), .A2(n375), .B1(out[108]), .B2(n369), .ZN(n171)
         );
  INV_X1 U342 ( .A(n172), .ZN(n288) );
  AOI22_X1 U343 ( .A1(in[107]), .A2(n375), .B1(out[107]), .B2(n368), .ZN(n172)
         );
  INV_X1 U344 ( .A(n173), .ZN(n287) );
  AOI22_X1 U345 ( .A1(in[106]), .A2(n375), .B1(out[106]), .B2(n369), .ZN(n173)
         );
  INV_X1 U346 ( .A(n174), .ZN(n286) );
  AOI22_X1 U347 ( .A1(in[105]), .A2(n375), .B1(out[105]), .B2(n368), .ZN(n174)
         );
  INV_X1 U348 ( .A(n175), .ZN(n285) );
  AOI22_X1 U349 ( .A1(in[104]), .A2(n375), .B1(out[104]), .B2(n369), .ZN(n175)
         );
  INV_X1 U350 ( .A(n176), .ZN(n284) );
  AOI22_X1 U351 ( .A1(in[103]), .A2(n375), .B1(out[103]), .B2(n368), .ZN(n176)
         );
  INV_X1 U352 ( .A(n177), .ZN(n283) );
  AOI22_X1 U353 ( .A1(in[102]), .A2(n375), .B1(out[102]), .B2(n369), .ZN(n177)
         );
  INV_X1 U354 ( .A(n178), .ZN(n282) );
  AOI22_X1 U355 ( .A1(in[101]), .A2(n375), .B1(out[101]), .B2(n368), .ZN(n178)
         );
  INV_X1 U356 ( .A(n179), .ZN(n281) );
  AOI22_X1 U357 ( .A1(in[100]), .A2(n375), .B1(out[100]), .B2(n369), .ZN(n179)
         );
  INV_X1 U358 ( .A(n180), .ZN(n181) );
  AOI22_X1 U359 ( .A1(in[0]), .A2(n375), .B1(out[0]), .B2(n368), .ZN(n180) );
  INV_X4 U361 ( .A(we), .ZN(n379) );
  INV_X4 U362 ( .A(we), .ZN(n380) );
  INV_X4 U363 ( .A(we), .ZN(n381) );
  INV_X4 U364 ( .A(we), .ZN(n375) );
  INV_X4 U365 ( .A(we), .ZN(n376) );
  INV_X4 U366 ( .A(we), .ZN(n377) );
  INV_X4 U367 ( .A(reset), .ZN(n396) );
  INV_X4 U368 ( .A(we), .ZN(n378) );
  INV_X4 U369 ( .A(n394), .ZN(n393) );
  INV_X4 U370 ( .A(n395), .ZN(n389) );
  INV_X4 U371 ( .A(n395), .ZN(n388) );
  INV_X4 U372 ( .A(n396), .ZN(n387) );
  INV_X4 U373 ( .A(n396), .ZN(n386) );
  INV_X4 U374 ( .A(n396), .ZN(n385) );
  INV_X4 U375 ( .A(n394), .ZN(n392) );
  INV_X4 U376 ( .A(we), .ZN(n371) );
  INV_X4 U377 ( .A(n371), .ZN(n366) );
  INV_X4 U378 ( .A(n371), .ZN(n367) );
  INV_X4 U379 ( .A(we), .ZN(n372) );
  INV_X4 U380 ( .A(n372), .ZN(n364) );
  INV_X4 U381 ( .A(n372), .ZN(n365) );
  INV_X4 U382 ( .A(reset), .ZN(n395) );
  INV_X4 U383 ( .A(n395), .ZN(n390) );
  INV_X4 U384 ( .A(n395), .ZN(n391) );
  INV_X4 U385 ( .A(we), .ZN(n373) );
  INV_X4 U386 ( .A(n373), .ZN(n362) );
  INV_X4 U387 ( .A(n373), .ZN(n363) );
  INV_X4 U388 ( .A(we), .ZN(n374) );
  INV_X4 U389 ( .A(n374), .ZN(n361) );
  INV_X4 U390 ( .A(n374), .ZN(n360) );
  INV_X4 U391 ( .A(we), .ZN(n370) );
  INV_X4 U392 ( .A(n370), .ZN(n368) );
  INV_X4 U393 ( .A(n370), .ZN(n369) );
  INV_X4 U394 ( .A(reset), .ZN(n394) );
  INV_X4 U395 ( .A(n394), .ZN(n382) );
  INV_X4 U396 ( .A(n394), .ZN(n383) );
  INV_X4 U397 ( .A(n394), .ZN(n384) );
  DFFR_X1 MEM_WB_REG_out_reg_9_ ( .D(n190), .CK(clk), .RN(reset), .Q(out[9])
         );
  DFFR_X1 MEM_WB_REG_out_reg_119_ ( .D(n300), .CK(clk), .RN(reset), .Q(
        out[119]) );
endmodule

