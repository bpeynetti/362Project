module write_back(
    
    
    );
    
    
    
    
    mux2to1_32bit MEM_OR_ALU(
        .X(),
        .Y(),
        .sel(),
        .Z()
    );