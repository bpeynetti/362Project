
module PipeCtlRegN_WIDTH108 ( out, in, ctl, clk, reset );
  output [0:107] out;
  input [0:107] in;
  input ctl, clk, reset;
  wire   n217, n218, n219, n220, n221, n222;

  SDFFR_X2 out_reg_0_ ( .D(1'b0), .SI(n219), .SE(in[0]), .CK(clk), .RN(reset), 
        .Q(out[0]) );
  SDFFR_X2 out_reg_1_ ( .D(1'b0), .SI(n220), .SE(in[1]), .CK(clk), .RN(reset), 
        .Q(out[1]) );
  SDFFR_X2 out_reg_2_ ( .D(1'b0), .SI(n221), .SE(in[2]), .CK(clk), .RN(reset), 
        .Q(out[2]) );
  SDFFR_X2 out_reg_3_ ( .D(1'b0), .SI(n222), .SE(in[3]), .CK(clk), .RN(reset), 
        .Q(out[3]) );
  SDFFR_X2 out_reg_4_ ( .D(1'b0), .SI(n219), .SE(in[4]), .CK(clk), .RN(reset), 
        .Q(out[4]) );
  SDFFR_X2 out_reg_5_ ( .D(1'b0), .SI(n220), .SE(in[5]), .CK(clk), .RN(reset), 
        .Q(out[5]) );
  SDFFR_X2 out_reg_6_ ( .D(1'b0), .SI(n221), .SE(in[6]), .CK(clk), .RN(reset), 
        .Q(out[6]) );
  SDFFR_X2 out_reg_7_ ( .D(1'b0), .SI(n222), .SE(in[7]), .CK(clk), .RN(reset), 
        .Q(out[7]) );
  SDFFR_X2 out_reg_8_ ( .D(1'b0), .SI(n219), .SE(in[8]), .CK(clk), .RN(reset), 
        .Q(out[8]) );
  SDFFR_X2 out_reg_9_ ( .D(1'b0), .SI(n220), .SE(in[9]), .CK(clk), .RN(reset), 
        .Q(out[9]) );
  SDFFR_X2 out_reg_10_ ( .D(1'b0), .SI(n221), .SE(in[10]), .CK(clk), .RN(reset), .Q(out[10]) );
  SDFFR_X2 out_reg_11_ ( .D(1'b0), .SI(n222), .SE(in[11]), .CK(clk), .RN(reset), .Q(out[11]) );
  SDFFR_X2 out_reg_12_ ( .D(1'b0), .SI(n219), .SE(in[12]), .CK(clk), .RN(reset), .Q(out[12]) );
  SDFFR_X2 out_reg_13_ ( .D(1'b0), .SI(n220), .SE(in[13]), .CK(clk), .RN(reset), .Q(out[13]) );
  SDFFR_X2 out_reg_14_ ( .D(1'b0), .SI(n221), .SE(in[14]), .CK(clk), .RN(reset), .Q(out[14]) );
  SDFFR_X2 out_reg_15_ ( .D(1'b0), .SI(n222), .SE(in[15]), .CK(clk), .RN(reset), .Q(out[15]) );
  SDFFR_X2 out_reg_16_ ( .D(1'b0), .SI(n219), .SE(in[16]), .CK(clk), .RN(reset), .Q(out[16]) );
  SDFFR_X2 out_reg_17_ ( .D(1'b0), .SI(n220), .SE(in[17]), .CK(clk), .RN(reset), .Q(out[17]) );
  SDFFR_X2 out_reg_18_ ( .D(1'b0), .SI(n221), .SE(in[18]), .CK(clk), .RN(reset), .Q(out[18]) );
  SDFFR_X2 out_reg_19_ ( .D(1'b0), .SI(n222), .SE(in[19]), .CK(clk), .RN(reset), .Q(out[19]) );
  SDFFR_X2 out_reg_20_ ( .D(1'b0), .SI(n219), .SE(in[20]), .CK(clk), .RN(reset), .Q(out[20]) );
  SDFFR_X2 out_reg_21_ ( .D(1'b0), .SI(n220), .SE(in[21]), .CK(clk), .RN(reset), .Q(out[21]) );
  SDFFR_X2 out_reg_22_ ( .D(1'b0), .SI(n221), .SE(in[22]), .CK(clk), .RN(reset), .Q(out[22]) );
  SDFFR_X2 out_reg_23_ ( .D(1'b0), .SI(n222), .SE(in[23]), .CK(clk), .RN(reset), .Q(out[23]) );
  SDFFR_X2 out_reg_24_ ( .D(1'b0), .SI(n219), .SE(in[24]), .CK(clk), .RN(reset), .Q(out[24]) );
  SDFFR_X2 out_reg_25_ ( .D(1'b0), .SI(n220), .SE(in[25]), .CK(clk), .RN(reset), .Q(out[25]) );
  SDFFR_X2 out_reg_26_ ( .D(1'b0), .SI(n221), .SE(in[26]), .CK(clk), .RN(reset), .Q(out[26]) );
  SDFFR_X2 out_reg_27_ ( .D(1'b0), .SI(n222), .SE(in[27]), .CK(clk), .RN(reset), .Q(out[27]) );
  SDFFR_X2 out_reg_28_ ( .D(1'b0), .SI(n219), .SE(in[28]), .CK(clk), .RN(reset), .Q(out[28]) );
  SDFFR_X2 out_reg_29_ ( .D(1'b0), .SI(n220), .SE(in[29]), .CK(clk), .RN(reset), .Q(out[29]) );
  SDFFR_X2 out_reg_30_ ( .D(1'b0), .SI(n221), .SE(in[30]), .CK(clk), .RN(reset), .Q(out[30]) );
  SDFFR_X2 out_reg_31_ ( .D(1'b0), .SI(n222), .SE(in[31]), .CK(clk), .RN(reset), .Q(out[31]) );
  SDFFR_X2 out_reg_32_ ( .D(1'b0), .SI(n219), .SE(in[32]), .CK(clk), .RN(reset), .Q(out[32]) );
  SDFFR_X2 out_reg_33_ ( .D(1'b0), .SI(n220), .SE(in[33]), .CK(clk), .RN(reset), .Q(out[33]) );
  SDFFR_X2 out_reg_34_ ( .D(1'b0), .SI(n221), .SE(in[34]), .CK(clk), .RN(reset), .Q(out[34]) );
  SDFFR_X2 out_reg_35_ ( .D(1'b0), .SI(n222), .SE(in[35]), .CK(clk), .RN(reset), .Q(out[35]) );
  SDFFR_X2 out_reg_36_ ( .D(1'b0), .SI(n219), .SE(in[36]), .CK(clk), .RN(reset), .Q(out[36]) );
  SDFFR_X2 out_reg_37_ ( .D(1'b0), .SI(n220), .SE(in[37]), .CK(clk), .RN(reset), .Q(out[37]) );
  SDFFR_X2 out_reg_38_ ( .D(1'b0), .SI(n221), .SE(in[38]), .CK(clk), .RN(reset), .Q(out[38]) );
  SDFFR_X2 out_reg_39_ ( .D(1'b0), .SI(n222), .SE(in[39]), .CK(clk), .RN(reset), .Q(out[39]) );
  SDFFR_X2 out_reg_40_ ( .D(1'b0), .SI(n219), .SE(in[40]), .CK(clk), .RN(reset), .Q(out[40]) );
  SDFFR_X2 out_reg_41_ ( .D(1'b0), .SI(n220), .SE(in[41]), .CK(clk), .RN(reset), .Q(out[41]) );
  SDFFR_X2 out_reg_42_ ( .D(1'b0), .SI(n221), .SE(in[42]), .CK(clk), .RN(reset), .Q(out[42]) );
  SDFFR_X2 out_reg_43_ ( .D(1'b0), .SI(n222), .SE(in[43]), .CK(clk), .RN(reset), .Q(out[43]) );
  SDFFR_X2 out_reg_44_ ( .D(1'b0), .SI(n219), .SE(in[44]), .CK(clk), .RN(reset), .Q(out[44]) );
  SDFFR_X2 out_reg_45_ ( .D(1'b0), .SI(n220), .SE(in[45]), .CK(clk), .RN(reset), .Q(out[45]) );
  SDFFR_X2 out_reg_46_ ( .D(1'b0), .SI(n221), .SE(in[46]), .CK(clk), .RN(reset), .Q(out[46]) );
  SDFFR_X2 out_reg_47_ ( .D(1'b0), .SI(n222), .SE(in[47]), .CK(clk), .RN(reset), .Q(out[47]) );
  SDFFR_X2 out_reg_48_ ( .D(1'b0), .SI(n219), .SE(in[48]), .CK(clk), .RN(reset), .Q(out[48]) );
  SDFFR_X2 out_reg_49_ ( .D(1'b0), .SI(n220), .SE(in[49]), .CK(clk), .RN(reset), .Q(out[49]) );
  SDFFR_X2 out_reg_50_ ( .D(1'b0), .SI(n221), .SE(in[50]), .CK(clk), .RN(reset), .Q(out[50]) );
  SDFFR_X2 out_reg_51_ ( .D(1'b0), .SI(n222), .SE(in[51]), .CK(clk), .RN(reset), .Q(out[51]) );
  SDFFR_X2 out_reg_52_ ( .D(1'b0), .SI(n219), .SE(in[52]), .CK(clk), .RN(reset), .Q(out[52]) );
  SDFFR_X2 out_reg_53_ ( .D(1'b0), .SI(n220), .SE(in[53]), .CK(clk), .RN(reset), .Q(out[53]) );
  SDFFR_X2 out_reg_54_ ( .D(1'b0), .SI(n221), .SE(in[54]), .CK(clk), .RN(reset), .Q(out[54]) );
  SDFFR_X2 out_reg_55_ ( .D(1'b0), .SI(n222), .SE(in[55]), .CK(clk), .RN(reset), .Q(out[55]) );
  SDFFR_X2 out_reg_56_ ( .D(1'b0), .SI(n219), .SE(in[56]), .CK(clk), .RN(reset), .Q(out[56]) );
  SDFFR_X2 out_reg_57_ ( .D(1'b0), .SI(n220), .SE(in[57]), .CK(clk), .RN(reset), .Q(out[57]) );
  SDFFR_X2 out_reg_58_ ( .D(1'b0), .SI(n221), .SE(in[58]), .CK(clk), .RN(reset), .Q(out[58]) );
  SDFFR_X2 out_reg_59_ ( .D(1'b0), .SI(n222), .SE(in[59]), .CK(clk), .RN(reset), .Q(out[59]) );
  SDFFR_X2 out_reg_60_ ( .D(1'b0), .SI(n219), .SE(in[60]), .CK(clk), .RN(reset), .Q(out[60]) );
  SDFFR_X2 out_reg_61_ ( .D(1'b0), .SI(n220), .SE(in[61]), .CK(clk), .RN(reset), .Q(out[61]) );
  SDFFR_X2 out_reg_62_ ( .D(1'b0), .SI(n221), .SE(in[62]), .CK(clk), .RN(reset), .Q(out[62]) );
  SDFFR_X2 out_reg_63_ ( .D(1'b0), .SI(n222), .SE(in[63]), .CK(clk), .RN(reset), .Q(out[63]) );
  SDFFR_X2 out_reg_64_ ( .D(1'b0), .SI(n219), .SE(in[64]), .CK(clk), .RN(reset), .Q(out[64]) );
  SDFFR_X2 out_reg_65_ ( .D(1'b0), .SI(n220), .SE(in[65]), .CK(clk), .RN(reset), .Q(out[65]) );
  SDFFR_X2 out_reg_66_ ( .D(1'b0), .SI(n221), .SE(in[66]), .CK(clk), .RN(reset), .Q(out[66]) );
  SDFFR_X2 out_reg_67_ ( .D(1'b0), .SI(n222), .SE(in[67]), .CK(clk), .RN(reset), .Q(out[67]) );
  SDFFR_X2 out_reg_68_ ( .D(1'b0), .SI(n219), .SE(in[68]), .CK(clk), .RN(reset), .Q(out[68]) );
  SDFFR_X2 out_reg_69_ ( .D(1'b0), .SI(n220), .SE(in[69]), .CK(clk), .RN(reset), .Q(out[69]) );
  SDFFR_X2 out_reg_70_ ( .D(1'b0), .SI(n221), .SE(in[70]), .CK(clk), .RN(reset), .Q(out[70]) );
  SDFFR_X2 out_reg_71_ ( .D(1'b0), .SI(n222), .SE(in[71]), .CK(clk), .RN(reset), .Q(out[71]) );
  SDFFR_X2 out_reg_72_ ( .D(1'b0), .SI(n219), .SE(in[72]), .CK(clk), .RN(reset), .Q(out[72]) );
  SDFFR_X2 out_reg_73_ ( .D(1'b0), .SI(n220), .SE(in[73]), .CK(clk), .RN(reset), .Q(out[73]) );
  SDFFR_X2 out_reg_74_ ( .D(1'b0), .SI(n221), .SE(in[74]), .CK(clk), .RN(reset), .Q(out[74]) );
  SDFFR_X2 out_reg_75_ ( .D(1'b0), .SI(n222), .SE(in[75]), .CK(clk), .RN(reset), .Q(out[75]) );
  SDFFR_X2 out_reg_76_ ( .D(1'b0), .SI(n219), .SE(in[76]), .CK(clk), .RN(reset), .Q(out[76]) );
  SDFFR_X2 out_reg_77_ ( .D(1'b0), .SI(n220), .SE(in[77]), .CK(clk), .RN(reset), .Q(out[77]) );
  SDFFR_X2 out_reg_78_ ( .D(1'b0), .SI(n221), .SE(in[78]), .CK(clk), .RN(reset), .Q(out[78]) );
  SDFFR_X2 out_reg_79_ ( .D(1'b0), .SI(n222), .SE(in[79]), .CK(clk), .RN(reset), .Q(out[79]) );
  SDFFR_X2 out_reg_80_ ( .D(1'b0), .SI(n219), .SE(in[80]), .CK(clk), .RN(reset), .Q(out[80]) );
  SDFFR_X2 out_reg_81_ ( .D(1'b0), .SI(n220), .SE(in[81]), .CK(clk), .RN(reset), .Q(out[81]) );
  SDFFR_X2 out_reg_82_ ( .D(1'b0), .SI(n221), .SE(in[82]), .CK(clk), .RN(reset), .Q(out[82]) );
  SDFFR_X2 out_reg_83_ ( .D(1'b0), .SI(n222), .SE(in[83]), .CK(clk), .RN(reset), .Q(out[83]) );
  SDFFR_X2 out_reg_84_ ( .D(1'b0), .SI(n219), .SE(in[84]), .CK(clk), .RN(reset), .Q(out[84]) );
  SDFFR_X2 out_reg_85_ ( .D(1'b0), .SI(n220), .SE(in[85]), .CK(clk), .RN(reset), .Q(out[85]) );
  SDFFR_X2 out_reg_86_ ( .D(1'b0), .SI(n221), .SE(in[86]), .CK(clk), .RN(reset), .Q(out[86]) );
  SDFFR_X2 out_reg_87_ ( .D(1'b0), .SI(n222), .SE(in[87]), .CK(clk), .RN(reset), .Q(out[87]) );
  SDFFR_X2 out_reg_88_ ( .D(1'b0), .SI(n219), .SE(in[88]), .CK(clk), .RN(reset), .Q(out[88]) );
  SDFFR_X2 out_reg_89_ ( .D(1'b0), .SI(n220), .SE(in[89]), .CK(clk), .RN(reset), .Q(out[89]) );
  SDFFR_X2 out_reg_90_ ( .D(1'b0), .SI(n221), .SE(in[90]), .CK(clk), .RN(reset), .Q(out[90]) );
  SDFFR_X2 out_reg_91_ ( .D(1'b0), .SI(n222), .SE(in[91]), .CK(clk), .RN(reset), .Q(out[91]) );
  SDFFR_X2 out_reg_92_ ( .D(1'b0), .SI(n219), .SE(in[92]), .CK(clk), .RN(reset), .Q(out[92]) );
  SDFFR_X2 out_reg_93_ ( .D(1'b0), .SI(n220), .SE(in[93]), .CK(clk), .RN(reset), .Q(out[93]) );
  SDFFR_X2 out_reg_94_ ( .D(1'b0), .SI(n221), .SE(in[94]), .CK(clk), .RN(reset), .Q(out[94]) );
  SDFFR_X2 out_reg_95_ ( .D(1'b0), .SI(n222), .SE(in[95]), .CK(clk), .RN(reset), .Q(out[95]) );
  SDFFR_X2 out_reg_96_ ( .D(1'b0), .SI(n219), .SE(in[96]), .CK(clk), .RN(reset), .Q(out[96]) );
  SDFFR_X2 out_reg_97_ ( .D(1'b0), .SI(n220), .SE(in[97]), .CK(clk), .RN(reset), .Q(out[97]) );
  SDFFR_X2 out_reg_98_ ( .D(1'b0), .SI(n221), .SE(in[98]), .CK(clk), .RN(reset), .Q(out[98]) );
  SDFFR_X2 out_reg_99_ ( .D(1'b0), .SI(n222), .SE(in[99]), .CK(clk), .RN(reset), .Q(out[99]) );
  SDFFR_X2 out_reg_100_ ( .D(1'b0), .SI(n219), .SE(in[100]), .CK(clk), .RN(
        reset), .Q(out[100]) );
  SDFFR_X2 out_reg_101_ ( .D(1'b0), .SI(n220), .SE(in[101]), .CK(clk), .RN(
        reset), .Q(out[101]) );
  SDFFR_X2 out_reg_102_ ( .D(1'b0), .SI(n221), .SE(in[102]), .CK(clk), .RN(
        reset), .Q(out[102]) );
  SDFFR_X2 out_reg_103_ ( .D(1'b0), .SI(n222), .SE(in[103]), .CK(clk), .RN(
        reset), .Q(out[103]) );
  SDFFR_X2 out_reg_104_ ( .D(1'b0), .SI(n219), .SE(in[104]), .CK(clk), .RN(
        reset), .Q(out[104]) );
  SDFFR_X2 out_reg_105_ ( .D(1'b0), .SI(n220), .SE(in[105]), .CK(clk), .RN(
        reset), .Q(out[105]) );
  SDFFR_X2 out_reg_106_ ( .D(1'b0), .SI(n221), .SE(in[106]), .CK(clk), .RN(
        reset), .Q(out[106]) );
  SDFFR_X2 out_reg_107_ ( .D(1'b0), .SI(n222), .SE(in[107]), .CK(clk), .RN(
        reset), .Q(out[107]) );
  INV_X1 U111 ( .A(ctl), .ZN(n217) );
  INV_X1 U112 ( .A(n217), .ZN(n218) );
  INV_X4 U113 ( .A(n218), .ZN(n219) );
  INV_X4 U114 ( .A(n218), .ZN(n220) );
  INV_X4 U115 ( .A(n218), .ZN(n221) );
  INV_X4 U116 ( .A(n218), .ZN(n222) );
endmodule

