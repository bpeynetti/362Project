
module multiplier_DW01_add_0 ( A, B, CI, SUM, CO );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [15:2] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(SUM[16]), .S(SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X2 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X4 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module multiplier_DW01_add_1 ( A, B, CI, SUM, CO );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [15:2] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(SUM[16]), .S(SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X2 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X4 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module multiplier_DW01_add_5 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16, n17,
         n33;
  wire   [32:18] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(n33), .CO(carry[18]), .S(SUM[17]) );
  XOR2_X2 U1 ( .A(B[33]), .B(n17), .Z(SUM[33]) );
  AND2_X4 U2 ( .A1(B[45]), .A2(n11), .ZN(n2) );
  AND2_X4 U3 ( .A1(B[43]), .A2(n12), .ZN(n3) );
  AND2_X4 U4 ( .A1(B[41]), .A2(n13), .ZN(n4) );
  AND2_X4 U5 ( .A1(B[39]), .A2(n14), .ZN(n5) );
  AND2_X4 U6 ( .A1(B[37]), .A2(n15), .ZN(n6) );
  AND2_X4 U7 ( .A1(B[35]), .A2(n16), .ZN(n7) );
  AND2_X4 U8 ( .A1(B[33]), .A2(n17), .ZN(n8) );
  XOR2_X2 U9 ( .A(B[32]), .B(carry[32]), .Z(SUM[32]) );
  AND2_X4 U10 ( .A1(B[46]), .A2(n2), .ZN(n10) );
  AND2_X4 U11 ( .A1(B[44]), .A2(n3), .ZN(n11) );
  AND2_X4 U12 ( .A1(B[42]), .A2(n4), .ZN(n12) );
  AND2_X4 U13 ( .A1(B[40]), .A2(n5), .ZN(n13) );
  AND2_X4 U14 ( .A1(B[38]), .A2(n6), .ZN(n14) );
  AND2_X4 U15 ( .A1(B[36]), .A2(n7), .ZN(n15) );
  AND2_X4 U16 ( .A1(B[34]), .A2(n8), .ZN(n16) );
  AND2_X4 U17 ( .A1(B[32]), .A2(carry[32]), .ZN(n17) );
  XOR2_X2 U18 ( .A(B[34]), .B(n8), .Z(SUM[34]) );
  XOR2_X2 U19 ( .A(B[35]), .B(n16), .Z(SUM[35]) );
  XOR2_X2 U20 ( .A(B[36]), .B(n7), .Z(SUM[36]) );
  XOR2_X2 U21 ( .A(B[37]), .B(n15), .Z(SUM[37]) );
  XOR2_X2 U22 ( .A(B[38]), .B(n6), .Z(SUM[38]) );
  XOR2_X2 U23 ( .A(B[39]), .B(n14), .Z(SUM[39]) );
  XOR2_X2 U24 ( .A(B[40]), .B(n5), .Z(SUM[40]) );
  XOR2_X2 U25 ( .A(B[41]), .B(n13), .Z(SUM[41]) );
  XOR2_X2 U26 ( .A(B[42]), .B(n4), .Z(SUM[42]) );
  XOR2_X2 U27 ( .A(B[43]), .B(n12), .Z(SUM[43]) );
  XOR2_X2 U28 ( .A(B[44]), .B(n3), .Z(SUM[44]) );
  XOR2_X2 U29 ( .A(B[45]), .B(n11), .Z(SUM[45]) );
  XOR2_X2 U30 ( .A(B[46]), .B(n2), .Z(SUM[46]) );
  XOR2_X2 U31 ( .A(B[47]), .B(n10), .Z(SUM[47]) );
  AND2_X4 U32 ( .A1(B[47]), .A2(n10), .ZN(SUM[48]) );
  AND2_X4 U33 ( .A1(B[16]), .A2(A[16]), .ZN(n33) );
  XOR2_X2 U34 ( .A(B[16]), .B(A[16]), .Z(SUM[16]) );
  BUF_X4 U35 ( .A(A[15]), .Z(SUM[15]) );
  BUF_X4 U36 ( .A(A[14]), .Z(SUM[14]) );
  BUF_X4 U37 ( .A(A[13]), .Z(SUM[13]) );
  BUF_X4 U38 ( .A(A[12]), .Z(SUM[12]) );
  BUF_X4 U39 ( .A(A[11]), .Z(SUM[11]) );
  BUF_X4 U40 ( .A(A[10]), .Z(SUM[10]) );
  BUF_X4 U41 ( .A(A[9]), .Z(SUM[9]) );
  BUF_X4 U42 ( .A(A[8]), .Z(SUM[8]) );
  BUF_X4 U43 ( .A(A[7]), .Z(SUM[7]) );
  BUF_X4 U44 ( .A(A[6]), .Z(SUM[6]) );
  BUF_X4 U45 ( .A(A[5]), .Z(SUM[5]) );
  BUF_X4 U46 ( .A(A[4]), .Z(SUM[4]) );
  BUF_X4 U47 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X4 U48 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X4 U49 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X4 U50 ( .A(A[0]), .Z(SUM[0]) );
endmodule


module multiplier_DW01_add_4 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;
  wire   [49:34] carry;

  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(n14), .CO(carry[34]), .S(SUM[33]) );
  AND2_X4 U1 ( .A1(A[60]), .A2(n8), .ZN(n1) );
  AND2_X4 U2 ( .A1(A[58]), .A2(n9), .ZN(n2) );
  AND2_X4 U3 ( .A1(A[56]), .A2(n10), .ZN(n3) );
  AND2_X4 U4 ( .A1(A[54]), .A2(n11), .ZN(n4) );
  AND2_X4 U5 ( .A1(A[52]), .A2(n12), .ZN(n5) );
  AND2_X4 U6 ( .A1(A[50]), .A2(n13), .ZN(n6) );
  AND2_X4 U7 ( .A1(A[61]), .A2(n1), .ZN(n7) );
  AND2_X4 U8 ( .A1(A[59]), .A2(n2), .ZN(n8) );
  AND2_X4 U9 ( .A1(A[57]), .A2(n3), .ZN(n9) );
  AND2_X4 U10 ( .A1(A[55]), .A2(n4), .ZN(n10) );
  AND2_X4 U11 ( .A1(A[53]), .A2(n5), .ZN(n11) );
  AND2_X4 U12 ( .A1(A[51]), .A2(n6), .ZN(n12) );
  AND2_X4 U13 ( .A1(A[49]), .A2(carry[49]), .ZN(n13) );
  AND2_X4 U14 ( .A1(B[32]), .A2(A[32]), .ZN(n14) );
  AND2_X4 U15 ( .A1(A[62]), .A2(n7), .ZN(n15) );
  XOR2_X2 U16 ( .A(A[49]), .B(carry[49]), .Z(SUM[49]) );
  XOR2_X2 U17 ( .A(B[32]), .B(A[32]), .Z(SUM[32]) );
  XOR2_X2 U18 ( .A(A[50]), .B(n13), .Z(SUM[50]) );
  XOR2_X2 U19 ( .A(A[51]), .B(n6), .Z(SUM[51]) );
  XOR2_X2 U20 ( .A(A[52]), .B(n12), .Z(SUM[52]) );
  XOR2_X2 U21 ( .A(A[53]), .B(n5), .Z(SUM[53]) );
  XOR2_X2 U22 ( .A(A[54]), .B(n11), .Z(SUM[54]) );
  XOR2_X2 U23 ( .A(A[55]), .B(n4), .Z(SUM[55]) );
  XOR2_X2 U24 ( .A(A[56]), .B(n10), .Z(SUM[56]) );
  XOR2_X2 U25 ( .A(A[57]), .B(n3), .Z(SUM[57]) );
  XOR2_X2 U26 ( .A(A[58]), .B(n9), .Z(SUM[58]) );
  XOR2_X2 U27 ( .A(A[59]), .B(n2), .Z(SUM[59]) );
  XOR2_X2 U28 ( .A(A[60]), .B(n8), .Z(SUM[60]) );
  XOR2_X2 U29 ( .A(A[61]), .B(n1), .Z(SUM[61]) );
  XOR2_X2 U30 ( .A(A[62]), .B(n7), .Z(SUM[62]) );
  XOR2_X2 U31 ( .A(A[63]), .B(n15), .Z(SUM[63]) );
  BUF_X4 U32 ( .A(B[31]), .Z(SUM[31]) );
  BUF_X4 U33 ( .A(B[30]), .Z(SUM[30]) );
  BUF_X4 U34 ( .A(B[29]), .Z(SUM[29]) );
  BUF_X4 U35 ( .A(B[28]), .Z(SUM[28]) );
  BUF_X4 U36 ( .A(B[27]), .Z(SUM[27]) );
  BUF_X4 U37 ( .A(B[26]), .Z(SUM[26]) );
  BUF_X4 U38 ( .A(B[25]), .Z(SUM[25]) );
  BUF_X32 U39 ( .A(B[0]), .Z(SUM[0]) );
  BUF_X32 U40 ( .A(B[1]), .Z(SUM[1]) );
  BUF_X32 U41 ( .A(B[2]), .Z(SUM[2]) );
  BUF_X32 U42 ( .A(B[3]), .Z(SUM[3]) );
  BUF_X32 U43 ( .A(B[4]), .Z(SUM[4]) );
  BUF_X32 U44 ( .A(B[5]), .Z(SUM[5]) );
  BUF_X32 U45 ( .A(B[6]), .Z(SUM[6]) );
  BUF_X32 U46 ( .A(B[7]), .Z(SUM[7]) );
  BUF_X32 U47 ( .A(B[8]), .Z(SUM[8]) );
  BUF_X32 U48 ( .A(B[9]), .Z(SUM[9]) );
  BUF_X32 U49 ( .A(B[10]), .Z(SUM[10]) );
  BUF_X32 U50 ( .A(B[11]), .Z(SUM[11]) );
  BUF_X32 U51 ( .A(B[12]), .Z(SUM[12]) );
  BUF_X32 U52 ( .A(B[13]), .Z(SUM[13]) );
  BUF_X32 U53 ( .A(B[14]), .Z(SUM[14]) );
  BUF_X32 U54 ( .A(B[15]), .Z(SUM[15]) );
  BUF_X32 U55 ( .A(B[16]), .Z(SUM[16]) );
  BUF_X32 U56 ( .A(B[17]), .Z(SUM[17]) );
  BUF_X32 U57 ( .A(B[18]), .Z(SUM[18]) );
  BUF_X32 U58 ( .A(B[19]), .Z(SUM[19]) );
  BUF_X32 U59 ( .A(B[20]), .Z(SUM[20]) );
  BUF_X32 U60 ( .A(B[21]), .Z(SUM[21]) );
  BUF_X32 U61 ( .A(B[22]), .Z(SUM[22]) );
  BUF_X32 U62 ( .A(B[23]), .Z(SUM[23]) );
  BUF_X32 U63 ( .A(B[24]), .Z(SUM[24]) );
endmodule


module multiplier_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [31:1] carry;

  FA_X1 U2_31 ( .A(A[31]), .B(n2), .CI(carry[31]), .S(DIFF[31]) );
  FA_X1 U2_30 ( .A(A[30]), .B(n3), .CI(carry[30]), .CO(carry[31]), .S(DIFF[30]) );
  FA_X1 U2_29 ( .A(A[29]), .B(n4), .CI(carry[29]), .CO(carry[30]), .S(DIFF[29]) );
  FA_X1 U2_28 ( .A(A[28]), .B(n5), .CI(carry[28]), .CO(carry[29]), .S(DIFF[28]) );
  FA_X1 U2_27 ( .A(A[27]), .B(n6), .CI(carry[27]), .CO(carry[28]), .S(DIFF[27]) );
  FA_X1 U2_26 ( .A(A[26]), .B(n7), .CI(carry[26]), .CO(carry[27]), .S(DIFF[26]) );
  FA_X1 U2_25 ( .A(A[25]), .B(n8), .CI(carry[25]), .CO(carry[26]), .S(DIFF[25]) );
  FA_X1 U2_24 ( .A(A[24]), .B(n9), .CI(carry[24]), .CO(carry[25]), .S(DIFF[24]) );
  FA_X1 U2_23 ( .A(A[23]), .B(n10), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FA_X1 U2_22 ( .A(A[22]), .B(n11), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FA_X1 U2_21 ( .A(A[21]), .B(n12), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FA_X1 U2_20 ( .A(A[20]), .B(n13), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FA_X1 U2_19 ( .A(A[19]), .B(n14), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FA_X1 U2_18 ( .A(A[18]), .B(n15), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FA_X1 U2_17 ( .A(A[17]), .B(n16), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FA_X1 U2_16 ( .A(A[16]), .B(n17), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FA_X1 U2_15 ( .A(A[15]), .B(n18), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FA_X1 U2_14 ( .A(A[14]), .B(n19), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(n20), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(n21), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(n22), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FA_X1 U2_10 ( .A(A[10]), .B(n23), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n24), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FA_X1 U2_8 ( .A(A[8]), .B(n25), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FA_X1 U2_7 ( .A(A[7]), .B(n26), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n27), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n28), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n29), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n30), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n31), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n32), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  NAND2_X2 U1 ( .A1(B[0]), .A2(n1), .ZN(carry[1]) );
  XNOR2_X2 U2 ( .A(n33), .B(A[0]), .ZN(DIFF[0]) );
  INV_X4 U3 ( .A(A[0]), .ZN(n1) );
  INV_X4 U4 ( .A(B[31]), .ZN(n2) );
  INV_X4 U5 ( .A(B[30]), .ZN(n3) );
  INV_X4 U6 ( .A(B[29]), .ZN(n4) );
  INV_X4 U7 ( .A(B[28]), .ZN(n5) );
  INV_X4 U8 ( .A(B[27]), .ZN(n6) );
  INV_X4 U9 ( .A(B[26]), .ZN(n7) );
  INV_X4 U10 ( .A(B[25]), .ZN(n8) );
  INV_X4 U11 ( .A(B[24]), .ZN(n9) );
  INV_X4 U12 ( .A(B[23]), .ZN(n10) );
  INV_X4 U13 ( .A(B[22]), .ZN(n11) );
  INV_X4 U14 ( .A(B[21]), .ZN(n12) );
  INV_X4 U15 ( .A(B[20]), .ZN(n13) );
  INV_X4 U16 ( .A(B[19]), .ZN(n14) );
  INV_X4 U17 ( .A(B[18]), .ZN(n15) );
  INV_X4 U18 ( .A(B[17]), .ZN(n16) );
  INV_X4 U19 ( .A(B[16]), .ZN(n17) );
  INV_X4 U20 ( .A(B[15]), .ZN(n18) );
  INV_X4 U21 ( .A(B[14]), .ZN(n19) );
  INV_X4 U22 ( .A(B[13]), .ZN(n20) );
  INV_X4 U23 ( .A(B[12]), .ZN(n21) );
  INV_X4 U24 ( .A(B[11]), .ZN(n22) );
  INV_X4 U25 ( .A(B[10]), .ZN(n23) );
  INV_X4 U26 ( .A(B[9]), .ZN(n24) );
  INV_X4 U27 ( .A(B[8]), .ZN(n25) );
  INV_X4 U28 ( .A(B[7]), .ZN(n26) );
  INV_X4 U29 ( .A(B[6]), .ZN(n27) );
  INV_X4 U30 ( .A(B[5]), .ZN(n28) );
  INV_X4 U31 ( .A(B[4]), .ZN(n29) );
  INV_X4 U32 ( .A(B[3]), .ZN(n30) );
  INV_X4 U33 ( .A(B[2]), .ZN(n31) );
  INV_X4 U34 ( .A(B[1]), .ZN(n32) );
  INV_X4 U35 ( .A(B[0]), .ZN(n33) );
endmodule


module multiplier_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [31:1] carry;

  FA_X1 U2_31 ( .A(A[31]), .B(n2), .CI(carry[31]), .S(DIFF[31]) );
  FA_X1 U2_30 ( .A(A[30]), .B(n3), .CI(carry[30]), .CO(carry[31]), .S(DIFF[30]) );
  FA_X1 U2_29 ( .A(A[29]), .B(n4), .CI(carry[29]), .CO(carry[30]), .S(DIFF[29]) );
  FA_X1 U2_28 ( .A(A[28]), .B(n5), .CI(carry[28]), .CO(carry[29]), .S(DIFF[28]) );
  FA_X1 U2_27 ( .A(A[27]), .B(n6), .CI(carry[27]), .CO(carry[28]), .S(DIFF[27]) );
  FA_X1 U2_26 ( .A(A[26]), .B(n7), .CI(carry[26]), .CO(carry[27]), .S(DIFF[26]) );
  FA_X1 U2_25 ( .A(A[25]), .B(n8), .CI(carry[25]), .CO(carry[26]), .S(DIFF[25]) );
  FA_X1 U2_24 ( .A(A[24]), .B(n9), .CI(carry[24]), .CO(carry[25]), .S(DIFF[24]) );
  FA_X1 U2_23 ( .A(A[23]), .B(n10), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FA_X1 U2_22 ( .A(A[22]), .B(n11), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FA_X1 U2_21 ( .A(A[21]), .B(n12), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FA_X1 U2_20 ( .A(A[20]), .B(n13), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FA_X1 U2_19 ( .A(A[19]), .B(n14), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FA_X1 U2_18 ( .A(A[18]), .B(n15), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FA_X1 U2_17 ( .A(A[17]), .B(n16), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FA_X1 U2_16 ( .A(A[16]), .B(n17), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FA_X1 U2_15 ( .A(A[15]), .B(n18), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FA_X1 U2_14 ( .A(A[14]), .B(n19), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(n20), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(n21), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(n22), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FA_X1 U2_10 ( .A(A[10]), .B(n23), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n24), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FA_X1 U2_8 ( .A(A[8]), .B(n25), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FA_X1 U2_7 ( .A(A[7]), .B(n26), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n27), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n28), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n29), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n30), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n31), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n32), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  NAND2_X2 U1 ( .A1(B[0]), .A2(n1), .ZN(carry[1]) );
  XNOR2_X2 U2 ( .A(n33), .B(A[0]), .ZN(DIFF[0]) );
  INV_X4 U3 ( .A(A[0]), .ZN(n1) );
  INV_X4 U4 ( .A(B[31]), .ZN(n2) );
  INV_X4 U5 ( .A(B[30]), .ZN(n3) );
  INV_X4 U6 ( .A(B[29]), .ZN(n4) );
  INV_X4 U7 ( .A(B[28]), .ZN(n5) );
  INV_X4 U8 ( .A(B[27]), .ZN(n6) );
  INV_X4 U9 ( .A(B[26]), .ZN(n7) );
  INV_X4 U10 ( .A(B[25]), .ZN(n8) );
  INV_X4 U11 ( .A(B[24]), .ZN(n9) );
  INV_X4 U12 ( .A(B[23]), .ZN(n10) );
  INV_X4 U13 ( .A(B[22]), .ZN(n11) );
  INV_X4 U14 ( .A(B[21]), .ZN(n12) );
  INV_X4 U15 ( .A(B[20]), .ZN(n13) );
  INV_X4 U16 ( .A(B[19]), .ZN(n14) );
  INV_X4 U17 ( .A(B[18]), .ZN(n15) );
  INV_X4 U18 ( .A(B[17]), .ZN(n16) );
  INV_X4 U19 ( .A(B[16]), .ZN(n17) );
  INV_X4 U20 ( .A(B[15]), .ZN(n18) );
  INV_X4 U21 ( .A(B[14]), .ZN(n19) );
  INV_X4 U22 ( .A(B[13]), .ZN(n20) );
  INV_X4 U23 ( .A(B[12]), .ZN(n21) );
  INV_X4 U24 ( .A(B[11]), .ZN(n22) );
  INV_X4 U25 ( .A(B[10]), .ZN(n23) );
  INV_X4 U26 ( .A(B[9]), .ZN(n24) );
  INV_X4 U27 ( .A(B[8]), .ZN(n25) );
  INV_X4 U28 ( .A(B[7]), .ZN(n26) );
  INV_X4 U29 ( .A(B[6]), .ZN(n27) );
  INV_X4 U30 ( .A(B[5]), .ZN(n28) );
  INV_X4 U31 ( .A(B[4]), .ZN(n29) );
  INV_X4 U32 ( .A(B[3]), .ZN(n30) );
  INV_X4 U33 ( .A(B[2]), .ZN(n31) );
  INV_X4 U34 ( .A(B[1]), .ZN(n32) );
  INV_X4 U35 ( .A(B[0]), .ZN(n33) );
endmodule


module multiplier_DW02_mult_2 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   \ab[16][15] , \ab[16][14] , \ab[16][13] , \ab[16][12] , \ab[16][11] ,
         \ab[16][10] , \ab[16][9] , \ab[16][8] , \ab[16][7] , \ab[16][6] ,
         \ab[16][5] , \ab[16][4] , \ab[16][3] , \ab[16][2] , \ab[16][1] ,
         \ab[16][0] , \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] ,
         \ab[15][11] , \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] ,
         \ab[15][6] , \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] ,
         \ab[15][1] , \ab[15][0] , \ab[14][15] , \ab[14][14] , \ab[14][13] ,
         \ab[14][12] , \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] ,
         \ab[14][7] , \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] ,
         \ab[14][2] , \ab[14][1] , \ab[14][0] , \ab[13][15] , \ab[13][14] ,
         \ab[13][13] , \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] ,
         \ab[13][8] , \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] ,
         \ab[13][3] , \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][15] ,
         \ab[12][14] , \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] ,
         \ab[12][9] , \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] ,
         \ab[12][4] , \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] ,
         \ab[11][15] , \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] ,
         \ab[11][10] , \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] ,
         \ab[11][5] , \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] ,
         \ab[11][0] , \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] ,
         \ab[10][11] , \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] ,
         \ab[10][6] , \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] ,
         \ab[10][1] , \ab[10][0] , \ab[9][15] , \ab[9][14] , \ab[9][13] ,
         \ab[9][12] , \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] ,
         \ab[9][7] , \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] ,
         \ab[9][2] , \ab[9][1] , \ab[9][0] , \ab[8][15] , \ab[8][14] ,
         \ab[8][13] , \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] ,
         \ab[8][8] , \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] ,
         \ab[8][3] , \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][15] ,
         \ab[7][14] , \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] ,
         \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] ,
         \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] ,
         \ab[6][15] , \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] ,
         \ab[6][10] , \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] ,
         \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] ,
         \ab[6][0] , \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] ,
         \ab[5][11] , \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] ,
         \ab[5][6] , \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] ,
         \ab[5][1] , \ab[5][0] , \ab[4][15] , \ab[4][14] , \ab[4][13] ,
         \ab[4][12] , \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] ,
         \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] ,
         \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][15] , \ab[3][14] ,
         \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] ,
         \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] ,
         \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][15] ,
         \ab[2][14] , \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] ,
         \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] ,
         \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] ,
         \ab[1][16] , \ab[1][15] , \ab[1][14] , \ab[1][13] , \ab[1][12] ,
         \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][8] , \ab[1][7] ,
         \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] ,
         \ab[1][1] , \ab[1][0] , \ab[0][16] , \ab[0][15] , \ab[0][14] ,
         \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] ,
         \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] ,
         \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[15][15] ,
         \CARRYB[15][14] , \CARRYB[15][13] , \CARRYB[15][12] ,
         \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] ,
         \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] ,
         \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] ,
         \CARRYB[14][15] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \CARRYB[13][15] , \CARRYB[13][14] , \CARRYB[13][13] ,
         \CARRYB[13][12] , \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] ,
         \CARRYB[13][8] , \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] ,
         \CARRYB[13][0] , \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][15] , \CARRYB[10][14] , \CARRYB[10][13] ,
         \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] ,
         \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] ,
         \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] ,
         \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] ,
         \CARRYB[9][0] , \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] ,
         \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] ,
         \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] ,
         \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] ,
         \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] ,
         \CARRYB[5][0] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][13] ,
         \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] ,
         \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[15][16] , \SUMB[15][15] , \SUMB[15][14] ,
         \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] , \SUMB[15][10] ,
         \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] , \SUMB[15][6] ,
         \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] , \SUMB[15][2] ,
         \SUMB[15][1] , \SUMB[14][16] , \SUMB[14][15] , \SUMB[14][14] ,
         \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] ,
         \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] ,
         \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] ,
         \SUMB[14][1] , \SUMB[13][16] , \SUMB[13][15] , \SUMB[13][14] ,
         \SUMB[13][13] , \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] ,
         \SUMB[13][9] , \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][6] ,
         \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] ,
         \SUMB[13][1] , \SUMB[12][16] , \SUMB[12][15] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][16] , \SUMB[11][15] , \SUMB[11][14] ,
         \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] , \SUMB[11][10] ,
         \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] , \SUMB[11][6] ,
         \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] , \SUMB[11][2] ,
         \SUMB[11][1] , \SUMB[10][16] , \SUMB[10][15] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][16] , \SUMB[9][15] , \SUMB[9][14] ,
         \SUMB[9][13] , \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] ,
         \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] ,
         \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][16] ,
         \SUMB[8][15] , \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] ,
         \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] ,
         \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] ,
         \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][16] , \SUMB[7][15] ,
         \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] , \SUMB[6][13] ,
         \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] , \SUMB[6][9] ,
         \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] ,
         \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][16] ,
         \SUMB[5][15] , \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] ,
         \SUMB[5][11] , \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] ,
         \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] ,
         \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][16] , \SUMB[4][15] ,
         \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] ,
         \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] , \SUMB[3][13] ,
         \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] , \SUMB[3][9] ,
         \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] ,
         \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][16] ,
         \SUMB[2][15] , \SUMB[2][14] , \SUMB[2][13] , \SUMB[2][12] ,
         \SUMB[2][11] , \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] ,
         \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , \CARRYB[30][0] , \CARRYB[29][1] ,
         \CARRYB[29][0] , \CARRYB[28][2] , \CARRYB[28][1] , \CARRYB[28][0] ,
         \CARRYB[27][3] , \CARRYB[27][2] , \CARRYB[27][1] , \CARRYB[27][0] ,
         \CARRYB[26][4] , \CARRYB[26][3] , \CARRYB[26][2] , \CARRYB[26][1] ,
         \CARRYB[26][0] , \CARRYB[25][5] , \CARRYB[25][4] , \CARRYB[25][3] ,
         \CARRYB[25][2] , \CARRYB[25][1] , \CARRYB[25][0] , \CARRYB[24][6] ,
         \CARRYB[24][5] , \CARRYB[24][4] , \CARRYB[24][3] , \CARRYB[24][2] ,
         \CARRYB[24][1] , \CARRYB[24][0] , \CARRYB[23][7] , \CARRYB[23][6] ,
         \CARRYB[23][5] , \CARRYB[23][4] , \CARRYB[23][3] , \CARRYB[23][2] ,
         \CARRYB[23][1] , \CARRYB[23][0] , \CARRYB[22][8] , \CARRYB[22][7] ,
         \CARRYB[22][6] , \CARRYB[22][5] , \CARRYB[22][4] , \CARRYB[22][3] ,
         \CARRYB[22][2] , \CARRYB[22][1] , \CARRYB[22][0] , \CARRYB[21][9] ,
         \CARRYB[21][8] , \CARRYB[21][7] , \CARRYB[21][6] , \CARRYB[21][5] ,
         \CARRYB[21][4] , \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] ,
         \CARRYB[21][0] , \CARRYB[20][10] , \CARRYB[20][9] , \CARRYB[20][8] ,
         \CARRYB[20][7] , \CARRYB[20][6] , \CARRYB[20][5] , \CARRYB[20][4] ,
         \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] , \CARRYB[20][0] ,
         \CARRYB[19][11] , \CARRYB[19][10] , \CARRYB[19][9] , \CARRYB[19][8] ,
         \CARRYB[19][7] , \CARRYB[19][6] , \CARRYB[19][5] , \CARRYB[19][4] ,
         \CARRYB[19][3] , \CARRYB[19][2] , \CARRYB[19][1] , \CARRYB[19][0] ,
         \CARRYB[18][12] , \CARRYB[18][11] , \CARRYB[18][10] , \CARRYB[18][9] ,
         \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][6] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] ,
         \CARRYB[18][0] , \CARRYB[17][13] , \CARRYB[17][12] , \CARRYB[17][11] ,
         \CARRYB[17][10] , \CARRYB[17][9] , \CARRYB[17][8] , \CARRYB[17][7] ,
         \CARRYB[17][6] , \CARRYB[17][5] , \CARRYB[17][4] , \CARRYB[17][3] ,
         \CARRYB[17][2] , \CARRYB[17][1] , \CARRYB[17][0] , \CARRYB[16][14] ,
         \CARRYB[16][13] , \CARRYB[16][12] , \CARRYB[16][11] ,
         \CARRYB[16][10] , \CARRYB[16][9] , \CARRYB[16][8] , \CARRYB[16][7] ,
         \CARRYB[16][6] , \CARRYB[16][5] , \CARRYB[16][4] , \CARRYB[16][3] ,
         \CARRYB[16][2] , \CARRYB[16][1] , \CARRYB[16][0] , \SUMB[30][1] ,
         \SUMB[29][2] , \SUMB[29][1] , \SUMB[28][3] , \SUMB[28][2] ,
         \SUMB[28][1] , \SUMB[27][4] , \SUMB[27][3] , \SUMB[27][2] ,
         \SUMB[27][1] , \SUMB[26][5] , \SUMB[26][4] , \SUMB[26][3] ,
         \SUMB[26][2] , \SUMB[26][1] , \SUMB[25][6] , \SUMB[25][5] ,
         \SUMB[25][4] , \SUMB[25][3] , \SUMB[25][2] , \SUMB[25][1] ,
         \SUMB[24][7] , \SUMB[24][6] , \SUMB[24][5] , \SUMB[24][4] ,
         \SUMB[24][3] , \SUMB[24][2] , \SUMB[24][1] , \SUMB[23][8] ,
         \SUMB[23][7] , \SUMB[23][6] , \SUMB[23][5] , \SUMB[23][4] ,
         \SUMB[23][3] , \SUMB[23][2] , \SUMB[23][1] , \SUMB[22][9] ,
         \SUMB[22][8] , \SUMB[22][7] , \SUMB[22][6] , \SUMB[22][5] ,
         \SUMB[22][4] , \SUMB[22][3] , \SUMB[22][2] , \SUMB[22][1] ,
         \SUMB[21][10] , \SUMB[21][9] , \SUMB[21][8] , \SUMB[21][7] ,
         \SUMB[21][6] , \SUMB[21][5] , \SUMB[21][4] , \SUMB[21][3] ,
         \SUMB[21][2] , \SUMB[21][1] , \SUMB[20][11] , \SUMB[20][10] ,
         \SUMB[20][9] , \SUMB[20][8] , \SUMB[20][7] , \SUMB[20][6] ,
         \SUMB[20][5] , \SUMB[20][4] , \SUMB[20][3] , \SUMB[20][2] ,
         \SUMB[20][1] , \SUMB[19][12] , \SUMB[19][11] , \SUMB[19][10] ,
         \SUMB[19][9] , \SUMB[19][8] , \SUMB[19][7] , \SUMB[19][6] ,
         \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] , \SUMB[19][2] ,
         \SUMB[19][1] , \SUMB[18][13] , \SUMB[18][12] , \SUMB[18][11] ,
         \SUMB[18][10] , \SUMB[18][9] , \SUMB[18][8] , \SUMB[18][7] ,
         \SUMB[18][6] , \SUMB[18][5] , \SUMB[18][4] , \SUMB[18][3] ,
         \SUMB[18][2] , \SUMB[18][1] , \SUMB[17][14] , \SUMB[17][13] ,
         \SUMB[17][12] , \SUMB[17][11] , \SUMB[17][10] , \SUMB[17][9] ,
         \SUMB[17][8] , \SUMB[17][7] , \SUMB[17][6] , \SUMB[17][5] ,
         \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] , \SUMB[17][1] ,
         \SUMB[16][15] , \SUMB[16][14] , \SUMB[16][13] , \SUMB[16][12] ,
         \SUMB[16][11] , \SUMB[16][10] , \SUMB[16][9] , \SUMB[16][8] ,
         \SUMB[16][7] , \SUMB[16][6] , \SUMB[16][5] , \SUMB[16][4] ,
         \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] , n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300;

  FA_X1 S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(PRODUCT[16]) );
  FA_X1 S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA_X1 S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), 
        .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA_X1 S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), 
        .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA_X1 S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA_X1 S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), 
        .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA_X1 S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), 
        .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA_X1 S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA_X1 S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA_X1 S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA_X1 S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), 
        .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA_X1 S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(\SUMB[15][12] ), 
        .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FA_X1 S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), 
        .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FA_X1 S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(\SUMB[15][14] ), 
        .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FA_X1 S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(\SUMB[15][15] ), 
        .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FA_X1 S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), 
        .S(\SUMB[16][15] ) );
  FA_X1 S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), 
        .CO(\CARRYB[15][0] ), .S(PRODUCT[15]) );
  FA_X1 S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), 
        .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA_X1 S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), 
        .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA_X1 S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), 
        .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA_X1 S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA_X1 S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA_X1 S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), 
        .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA_X1 S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), 
        .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA_X1 S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), 
        .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA_X1 S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA_X1 S2_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA_X1 S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA_X1 S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA_X1 S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA_X1 S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA_X1 S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), 
        .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FA_X1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(PRODUCT[14]) );
  FA_X1 S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA_X1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA_X1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA_X1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA_X1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA_X1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA_X1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA_X1 S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA_X1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA_X1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA_X1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA_X1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA_X1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA_X1 S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA_X1 S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\SUMB[13][16] ), 
        .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA_X1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(PRODUCT[13]) );
  FA_X1 S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA_X1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA_X1 S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA_X1 S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA_X1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA_X1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA_X1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA_X1 S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA_X1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA_X1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA_X1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA_X1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA_X1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA_X1 S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA_X1 S2_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\SUMB[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA_X1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(PRODUCT[12]) );
  FA_X1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA_X1 S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA_X1 S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA_X1 S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA_X1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA_X1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA_X1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA_X1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA_X1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA_X1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA_X1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA_X1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA_X1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA_X1 S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA_X1 S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\SUMB[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA_X1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(PRODUCT[11]) );
  FA_X1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA_X1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA_X1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA_X1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA_X1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA_X1 S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA_X1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA_X1 S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA_X1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA_X1 S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA_X1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA_X1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA_X1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA_X1 S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA_X1 S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA_X1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(PRODUCT[10]) );
  FA_X1 S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA_X1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA_X1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA_X1 S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA_X1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA_X1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA_X1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA_X1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA_X1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA_X1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA_X1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA_X1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA_X1 S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA_X1 S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA_X1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(PRODUCT[9]) );
  FA_X1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA_X1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA_X1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA_X1 S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA_X1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA_X1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA_X1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA_X1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA_X1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA_X1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA_X1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA_X1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA_X1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA_X1 S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA_X1 S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), 
        .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA_X1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(PRODUCT[8]) );
  FA_X1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA_X1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA_X1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA_X1 S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA_X1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA_X1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA_X1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA_X1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA_X1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA_X1 S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA_X1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA_X1 S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA_X1 S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA_X1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(PRODUCT[7]) );
  FA_X1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA_X1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA_X1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA_X1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA_X1 S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA_X1 S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA_X1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA_X1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA_X1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA_X1 S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA_X1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA_X1 S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA_X1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA_X1 S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA_X1 S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA_X1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(PRODUCT[6]) );
  FA_X1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA_X1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA_X1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA_X1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA_X1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA_X1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA_X1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA_X1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA_X1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA_X1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA_X1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA_X1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA_X1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA_X1 S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA_X1 S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA_X1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(PRODUCT[5]) );
  FA_X1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA_X1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA_X1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA_X1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA_X1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA_X1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA_X1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA_X1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA_X1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA_X1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA_X1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA_X1 S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA_X1 S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA_X1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(PRODUCT[4]) );
  FA_X1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA_X1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA_X1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA_X1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA_X1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA_X1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA_X1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA_X1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA_X1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA_X1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA_X1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA_X1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA_X1 S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA_X1 S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA_X1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(PRODUCT[3]) );
  FA_X1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA_X1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA_X1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA_X1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA_X1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA_X1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA_X1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA_X1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA_X1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA_X1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA_X1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA_X1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA_X1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA_X1 S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA_X1 S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), 
        .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(n235), .CI(n258), .CO(\CARRYB[2][0] ), .S(
        PRODUCT[2]) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(n243), .CI(n257), .CO(\CARRYB[2][1] ), .S(
        \SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(n242), .CI(n256), .CO(\CARRYB[2][2] ), .S(
        \SUMB[2][2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2][3] ), .B(n241), .CI(n255), .CO(\CARRYB[2][3] ), .S(
        \SUMB[2][3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2][4] ), .B(n240), .CI(n254), .CO(\CARRYB[2][4] ), .S(
        \SUMB[2][4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2][5] ), .B(n239), .CI(n253), .CO(\CARRYB[2][5] ), .S(
        \SUMB[2][5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2][6] ), .B(n238), .CI(n252), .CO(\CARRYB[2][6] ), .S(
        \SUMB[2][6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(n237), .CI(n251), .CO(\CARRYB[2][7] ), .S(
        \SUMB[2][7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(n236), .CI(n250), .CO(\CARRYB[2][8] ), .S(
        \SUMB[2][8] ) );
  FA_X1 S2_2_9 ( .A(\ab[2][9] ), .B(n234), .CI(n248), .CO(\CARRYB[2][9] ), .S(
        \SUMB[2][9] ) );
  FA_X1 S2_2_10 ( .A(\ab[2][10] ), .B(n233), .CI(n247), .CO(\CARRYB[2][10] ), 
        .S(\SUMB[2][10] ) );
  FA_X1 S2_2_11 ( .A(\ab[2][11] ), .B(n232), .CI(n246), .CO(\CARRYB[2][11] ), 
        .S(\SUMB[2][11] ) );
  FA_X1 S2_2_12 ( .A(\ab[2][12] ), .B(n231), .CI(n245), .CO(\CARRYB[2][12] ), 
        .S(\SUMB[2][12] ) );
  FA_X1 S2_2_13 ( .A(\ab[2][13] ), .B(n230), .CI(n244), .CO(\CARRYB[2][13] ), 
        .S(\SUMB[2][13] ) );
  FA_X1 S2_2_14 ( .A(\ab[2][14] ), .B(n229), .CI(n249), .CO(\CARRYB[2][14] ), 
        .S(\SUMB[2][14] ) );
  FA_X1 S2_2_15 ( .A(\ab[2][15] ), .B(n228), .CI(\ab[1][16] ), .CO(
        \CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  NAND2_X2 U2 ( .A1(\SUMB[20][10] ), .A2(\CARRYB[20][9] ), .ZN(n3) );
  INV_X4 U3 ( .A(n3), .ZN(\CARRYB[21][9] ) );
  XNOR2_X2 U4 ( .A(\CARRYB[20][9] ), .B(\SUMB[20][10] ), .ZN(n4) );
  INV_X4 U5 ( .A(n4), .ZN(\SUMB[21][9] ) );
  NAND2_X2 U6 ( .A1(\SUMB[20][1] ), .A2(\CARRYB[20][0] ), .ZN(n5) );
  INV_X4 U7 ( .A(n5), .ZN(\CARRYB[21][0] ) );
  XNOR2_X2 U8 ( .A(\CARRYB[20][0] ), .B(\SUMB[20][1] ), .ZN(n6) );
  INV_X4 U9 ( .A(n6), .ZN(PRODUCT[21]) );
  XNOR2_X2 U10 ( .A(\CARRYB[20][10] ), .B(\SUMB[20][11] ), .ZN(n7) );
  INV_X4 U11 ( .A(n7), .ZN(\SUMB[21][10] ) );
  NAND2_X2 U12 ( .A1(\SUMB[20][2] ), .A2(\CARRYB[20][1] ), .ZN(n8) );
  INV_X4 U13 ( .A(n8), .ZN(\CARRYB[21][1] ) );
  XNOR2_X2 U14 ( .A(\CARRYB[20][1] ), .B(\SUMB[20][2] ), .ZN(n9) );
  INV_X4 U15 ( .A(n9), .ZN(\SUMB[21][1] ) );
  NAND2_X2 U16 ( .A1(\SUMB[20][3] ), .A2(\CARRYB[20][2] ), .ZN(n10) );
  INV_X4 U17 ( .A(n10), .ZN(\CARRYB[21][2] ) );
  XNOR2_X2 U18 ( .A(\CARRYB[20][2] ), .B(\SUMB[20][3] ), .ZN(n11) );
  INV_X4 U19 ( .A(n11), .ZN(\SUMB[21][2] ) );
  NAND2_X2 U20 ( .A1(\SUMB[20][4] ), .A2(\CARRYB[20][3] ), .ZN(n12) );
  INV_X4 U21 ( .A(n12), .ZN(\CARRYB[21][3] ) );
  XNOR2_X2 U22 ( .A(\CARRYB[20][3] ), .B(\SUMB[20][4] ), .ZN(n13) );
  INV_X4 U23 ( .A(n13), .ZN(\SUMB[21][3] ) );
  NAND2_X2 U24 ( .A1(\SUMB[20][5] ), .A2(\CARRYB[20][4] ), .ZN(n14) );
  INV_X4 U25 ( .A(n14), .ZN(\CARRYB[21][4] ) );
  XNOR2_X2 U26 ( .A(\CARRYB[20][4] ), .B(\SUMB[20][5] ), .ZN(n15) );
  INV_X4 U27 ( .A(n15), .ZN(\SUMB[21][4] ) );
  NAND2_X2 U28 ( .A1(\SUMB[20][6] ), .A2(\CARRYB[20][5] ), .ZN(n16) );
  INV_X4 U29 ( .A(n16), .ZN(\CARRYB[21][5] ) );
  XNOR2_X2 U30 ( .A(\CARRYB[20][5] ), .B(\SUMB[20][6] ), .ZN(n17) );
  INV_X4 U31 ( .A(n17), .ZN(\SUMB[21][5] ) );
  NAND2_X2 U32 ( .A1(\SUMB[20][7] ), .A2(\CARRYB[20][6] ), .ZN(n18) );
  INV_X4 U33 ( .A(n18), .ZN(\CARRYB[21][6] ) );
  XNOR2_X2 U34 ( .A(\CARRYB[20][6] ), .B(\SUMB[20][7] ), .ZN(n19) );
  INV_X4 U35 ( .A(n19), .ZN(\SUMB[21][6] ) );
  NAND2_X2 U36 ( .A1(\SUMB[20][8] ), .A2(\CARRYB[20][7] ), .ZN(n20) );
  INV_X4 U37 ( .A(n20), .ZN(\CARRYB[21][7] ) );
  XNOR2_X2 U38 ( .A(\CARRYB[20][7] ), .B(\SUMB[20][8] ), .ZN(n21) );
  INV_X4 U39 ( .A(n21), .ZN(\SUMB[21][7] ) );
  NAND2_X2 U40 ( .A1(\SUMB[20][9] ), .A2(\CARRYB[20][8] ), .ZN(n22) );
  INV_X4 U41 ( .A(n22), .ZN(\CARRYB[21][8] ) );
  XNOR2_X2 U42 ( .A(\CARRYB[20][8] ), .B(\SUMB[20][9] ), .ZN(n23) );
  INV_X4 U43 ( .A(n23), .ZN(\SUMB[21][8] ) );
  NAND2_X2 U44 ( .A1(\SUMB[19][10] ), .A2(\CARRYB[19][9] ), .ZN(n24) );
  INV_X4 U45 ( .A(n24), .ZN(\CARRYB[20][9] ) );
  XNOR2_X2 U46 ( .A(\CARRYB[19][9] ), .B(\SUMB[19][10] ), .ZN(n25) );
  INV_X4 U47 ( .A(n25), .ZN(\SUMB[20][9] ) );
  NAND2_X2 U48 ( .A1(\SUMB[19][1] ), .A2(\CARRYB[19][0] ), .ZN(n26) );
  INV_X4 U49 ( .A(n26), .ZN(\CARRYB[20][0] ) );
  XNOR2_X2 U50 ( .A(\CARRYB[19][0] ), .B(\SUMB[19][1] ), .ZN(n27) );
  INV_X4 U51 ( .A(n27), .ZN(PRODUCT[20]) );
  NAND2_X2 U52 ( .A1(\SUMB[19][11] ), .A2(\CARRYB[19][10] ), .ZN(n28) );
  INV_X4 U53 ( .A(n28), .ZN(\CARRYB[20][10] ) );
  XNOR2_X2 U54 ( .A(\CARRYB[19][10] ), .B(\SUMB[19][11] ), .ZN(n29) );
  INV_X4 U55 ( .A(n29), .ZN(\SUMB[20][10] ) );
  XNOR2_X2 U56 ( .A(\CARRYB[19][11] ), .B(\SUMB[19][12] ), .ZN(n30) );
  INV_X4 U57 ( .A(n30), .ZN(\SUMB[20][11] ) );
  NAND2_X2 U58 ( .A1(\SUMB[19][2] ), .A2(\CARRYB[19][1] ), .ZN(n31) );
  INV_X4 U59 ( .A(n31), .ZN(\CARRYB[20][1] ) );
  XNOR2_X2 U60 ( .A(\CARRYB[19][1] ), .B(\SUMB[19][2] ), .ZN(n32) );
  INV_X4 U61 ( .A(n32), .ZN(\SUMB[20][1] ) );
  NAND2_X2 U62 ( .A1(\SUMB[19][3] ), .A2(\CARRYB[19][2] ), .ZN(n33) );
  INV_X4 U63 ( .A(n33), .ZN(\CARRYB[20][2] ) );
  XNOR2_X2 U64 ( .A(\CARRYB[19][2] ), .B(\SUMB[19][3] ), .ZN(n34) );
  INV_X4 U65 ( .A(n34), .ZN(\SUMB[20][2] ) );
  NAND2_X2 U66 ( .A1(\SUMB[19][4] ), .A2(\CARRYB[19][3] ), .ZN(n35) );
  INV_X4 U67 ( .A(n35), .ZN(\CARRYB[20][3] ) );
  XNOR2_X2 U68 ( .A(\CARRYB[19][3] ), .B(\SUMB[19][4] ), .ZN(n36) );
  INV_X4 U69 ( .A(n36), .ZN(\SUMB[20][3] ) );
  NAND2_X2 U70 ( .A1(\SUMB[19][5] ), .A2(\CARRYB[19][4] ), .ZN(n37) );
  INV_X4 U71 ( .A(n37), .ZN(\CARRYB[20][4] ) );
  XNOR2_X2 U72 ( .A(\CARRYB[19][4] ), .B(\SUMB[19][5] ), .ZN(n38) );
  INV_X4 U73 ( .A(n38), .ZN(\SUMB[20][4] ) );
  NAND2_X2 U74 ( .A1(\SUMB[19][6] ), .A2(\CARRYB[19][5] ), .ZN(n39) );
  INV_X4 U75 ( .A(n39), .ZN(\CARRYB[20][5] ) );
  XNOR2_X2 U76 ( .A(\CARRYB[19][5] ), .B(\SUMB[19][6] ), .ZN(n40) );
  INV_X4 U77 ( .A(n40), .ZN(\SUMB[20][5] ) );
  NAND2_X2 U78 ( .A1(\SUMB[19][7] ), .A2(\CARRYB[19][6] ), .ZN(n41) );
  INV_X4 U79 ( .A(n41), .ZN(\CARRYB[20][6] ) );
  XNOR2_X2 U80 ( .A(\CARRYB[19][6] ), .B(\SUMB[19][7] ), .ZN(n42) );
  INV_X4 U81 ( .A(n42), .ZN(\SUMB[20][6] ) );
  NAND2_X2 U82 ( .A1(\SUMB[19][8] ), .A2(\CARRYB[19][7] ), .ZN(n43) );
  INV_X4 U83 ( .A(n43), .ZN(\CARRYB[20][7] ) );
  XNOR2_X2 U84 ( .A(\CARRYB[19][7] ), .B(\SUMB[19][8] ), .ZN(n44) );
  INV_X4 U85 ( .A(n44), .ZN(\SUMB[20][7] ) );
  NAND2_X2 U86 ( .A1(\SUMB[19][9] ), .A2(\CARRYB[19][8] ), .ZN(n45) );
  INV_X4 U87 ( .A(n45), .ZN(\CARRYB[20][8] ) );
  XNOR2_X2 U88 ( .A(\CARRYB[19][8] ), .B(\SUMB[19][9] ), .ZN(n46) );
  INV_X4 U89 ( .A(n46), .ZN(\SUMB[20][8] ) );
  NAND2_X2 U90 ( .A1(\SUMB[18][10] ), .A2(\CARRYB[18][9] ), .ZN(n47) );
  INV_X4 U91 ( .A(n47), .ZN(\CARRYB[19][9] ) );
  XNOR2_X2 U92 ( .A(\CARRYB[18][9] ), .B(\SUMB[18][10] ), .ZN(n48) );
  INV_X4 U93 ( .A(n48), .ZN(\SUMB[19][9] ) );
  NAND2_X2 U94 ( .A1(\SUMB[18][1] ), .A2(\CARRYB[18][0] ), .ZN(n49) );
  INV_X4 U95 ( .A(n49), .ZN(\CARRYB[19][0] ) );
  XNOR2_X2 U96 ( .A(\CARRYB[18][0] ), .B(\SUMB[18][1] ), .ZN(n50) );
  INV_X4 U97 ( .A(n50), .ZN(PRODUCT[19]) );
  NAND2_X2 U98 ( .A1(\SUMB[18][11] ), .A2(\CARRYB[18][10] ), .ZN(n51) );
  INV_X4 U99 ( .A(n51), .ZN(\CARRYB[19][10] ) );
  XNOR2_X2 U100 ( .A(\CARRYB[18][10] ), .B(\SUMB[18][11] ), .ZN(n52) );
  INV_X4 U101 ( .A(n52), .ZN(\SUMB[19][10] ) );
  NAND2_X2 U102 ( .A1(\SUMB[18][12] ), .A2(\CARRYB[18][11] ), .ZN(n53) );
  INV_X4 U103 ( .A(n53), .ZN(\CARRYB[19][11] ) );
  XNOR2_X2 U104 ( .A(\CARRYB[18][11] ), .B(\SUMB[18][12] ), .ZN(n54) );
  INV_X4 U105 ( .A(n54), .ZN(\SUMB[19][11] ) );
  XNOR2_X2 U106 ( .A(\CARRYB[18][12] ), .B(\SUMB[18][13] ), .ZN(n55) );
  INV_X4 U107 ( .A(n55), .ZN(\SUMB[19][12] ) );
  NAND2_X2 U108 ( .A1(\SUMB[18][2] ), .A2(\CARRYB[18][1] ), .ZN(n56) );
  INV_X4 U109 ( .A(n56), .ZN(\CARRYB[19][1] ) );
  XNOR2_X2 U110 ( .A(\CARRYB[18][1] ), .B(\SUMB[18][2] ), .ZN(n57) );
  INV_X4 U111 ( .A(n57), .ZN(\SUMB[19][1] ) );
  NAND2_X2 U112 ( .A1(\SUMB[18][3] ), .A2(\CARRYB[18][2] ), .ZN(n58) );
  INV_X4 U113 ( .A(n58), .ZN(\CARRYB[19][2] ) );
  XNOR2_X2 U114 ( .A(\CARRYB[18][2] ), .B(\SUMB[18][3] ), .ZN(n59) );
  INV_X4 U115 ( .A(n59), .ZN(\SUMB[19][2] ) );
  NAND2_X2 U116 ( .A1(\SUMB[18][4] ), .A2(\CARRYB[18][3] ), .ZN(n60) );
  INV_X4 U117 ( .A(n60), .ZN(\CARRYB[19][3] ) );
  XNOR2_X2 U118 ( .A(\CARRYB[18][3] ), .B(\SUMB[18][4] ), .ZN(n61) );
  INV_X4 U119 ( .A(n61), .ZN(\SUMB[19][3] ) );
  NAND2_X2 U120 ( .A1(\SUMB[18][5] ), .A2(\CARRYB[18][4] ), .ZN(n62) );
  INV_X4 U121 ( .A(n62), .ZN(\CARRYB[19][4] ) );
  XNOR2_X2 U122 ( .A(\CARRYB[18][4] ), .B(\SUMB[18][5] ), .ZN(n63) );
  INV_X4 U123 ( .A(n63), .ZN(\SUMB[19][4] ) );
  NAND2_X2 U124 ( .A1(\SUMB[18][6] ), .A2(\CARRYB[18][5] ), .ZN(n64) );
  INV_X4 U125 ( .A(n64), .ZN(\CARRYB[19][5] ) );
  XNOR2_X2 U126 ( .A(\CARRYB[18][5] ), .B(\SUMB[18][6] ), .ZN(n65) );
  INV_X4 U127 ( .A(n65), .ZN(\SUMB[19][5] ) );
  NAND2_X2 U128 ( .A1(\SUMB[18][7] ), .A2(\CARRYB[18][6] ), .ZN(n66) );
  INV_X4 U129 ( .A(n66), .ZN(\CARRYB[19][6] ) );
  XNOR2_X2 U130 ( .A(\CARRYB[18][6] ), .B(\SUMB[18][7] ), .ZN(n67) );
  INV_X4 U131 ( .A(n67), .ZN(\SUMB[19][6] ) );
  NAND2_X2 U132 ( .A1(\SUMB[18][8] ), .A2(\CARRYB[18][7] ), .ZN(n68) );
  INV_X4 U133 ( .A(n68), .ZN(\CARRYB[19][7] ) );
  XNOR2_X2 U134 ( .A(\CARRYB[18][7] ), .B(\SUMB[18][8] ), .ZN(n69) );
  INV_X4 U135 ( .A(n69), .ZN(\SUMB[19][7] ) );
  NAND2_X2 U136 ( .A1(\SUMB[18][9] ), .A2(\CARRYB[18][8] ), .ZN(n70) );
  INV_X4 U137 ( .A(n70), .ZN(\CARRYB[19][8] ) );
  XNOR2_X2 U138 ( .A(\CARRYB[18][8] ), .B(\SUMB[18][9] ), .ZN(n71) );
  INV_X4 U139 ( .A(n71), .ZN(\SUMB[19][8] ) );
  NAND2_X2 U140 ( .A1(\SUMB[17][10] ), .A2(\CARRYB[17][9] ), .ZN(n72) );
  INV_X4 U141 ( .A(n72), .ZN(\CARRYB[18][9] ) );
  XNOR2_X2 U142 ( .A(\CARRYB[17][9] ), .B(\SUMB[17][10] ), .ZN(n73) );
  INV_X4 U143 ( .A(n73), .ZN(\SUMB[18][9] ) );
  NAND2_X2 U144 ( .A1(\SUMB[17][1] ), .A2(\CARRYB[17][0] ), .ZN(n74) );
  INV_X4 U145 ( .A(n74), .ZN(\CARRYB[18][0] ) );
  XNOR2_X2 U146 ( .A(\CARRYB[17][0] ), .B(\SUMB[17][1] ), .ZN(n75) );
  INV_X4 U147 ( .A(n75), .ZN(PRODUCT[18]) );
  NAND2_X2 U148 ( .A1(\SUMB[17][11] ), .A2(\CARRYB[17][10] ), .ZN(n76) );
  INV_X4 U149 ( .A(n76), .ZN(\CARRYB[18][10] ) );
  XNOR2_X2 U150 ( .A(\CARRYB[17][10] ), .B(\SUMB[17][11] ), .ZN(n77) );
  INV_X4 U151 ( .A(n77), .ZN(\SUMB[18][10] ) );
  NAND2_X2 U152 ( .A1(\SUMB[17][12] ), .A2(\CARRYB[17][11] ), .ZN(n78) );
  INV_X4 U153 ( .A(n78), .ZN(\CARRYB[18][11] ) );
  XNOR2_X2 U154 ( .A(\CARRYB[17][11] ), .B(\SUMB[17][12] ), .ZN(n79) );
  INV_X4 U155 ( .A(n79), .ZN(\SUMB[18][11] ) );
  NAND2_X2 U156 ( .A1(\SUMB[17][13] ), .A2(\CARRYB[17][12] ), .ZN(n80) );
  INV_X4 U157 ( .A(n80), .ZN(\CARRYB[18][12] ) );
  XNOR2_X2 U158 ( .A(\CARRYB[17][12] ), .B(\SUMB[17][13] ), .ZN(n81) );
  INV_X4 U159 ( .A(n81), .ZN(\SUMB[18][12] ) );
  XNOR2_X2 U160 ( .A(\CARRYB[17][13] ), .B(\SUMB[17][14] ), .ZN(n82) );
  INV_X4 U161 ( .A(n82), .ZN(\SUMB[18][13] ) );
  NAND2_X2 U162 ( .A1(\SUMB[17][2] ), .A2(\CARRYB[17][1] ), .ZN(n83) );
  INV_X4 U163 ( .A(n83), .ZN(\CARRYB[18][1] ) );
  XNOR2_X2 U164 ( .A(\CARRYB[17][1] ), .B(\SUMB[17][2] ), .ZN(n84) );
  INV_X4 U165 ( .A(n84), .ZN(\SUMB[18][1] ) );
  NAND2_X2 U166 ( .A1(\SUMB[17][3] ), .A2(\CARRYB[17][2] ), .ZN(n85) );
  INV_X4 U167 ( .A(n85), .ZN(\CARRYB[18][2] ) );
  XNOR2_X2 U168 ( .A(\CARRYB[17][2] ), .B(\SUMB[17][3] ), .ZN(n86) );
  INV_X4 U169 ( .A(n86), .ZN(\SUMB[18][2] ) );
  NAND2_X2 U170 ( .A1(\SUMB[17][4] ), .A2(\CARRYB[17][3] ), .ZN(n87) );
  INV_X4 U171 ( .A(n87), .ZN(\CARRYB[18][3] ) );
  XNOR2_X2 U172 ( .A(\CARRYB[17][3] ), .B(\SUMB[17][4] ), .ZN(n88) );
  INV_X4 U173 ( .A(n88), .ZN(\SUMB[18][3] ) );
  NAND2_X2 U174 ( .A1(\SUMB[17][5] ), .A2(\CARRYB[17][4] ), .ZN(n89) );
  INV_X4 U175 ( .A(n89), .ZN(\CARRYB[18][4] ) );
  XNOR2_X2 U176 ( .A(\CARRYB[17][4] ), .B(\SUMB[17][5] ), .ZN(n90) );
  INV_X4 U177 ( .A(n90), .ZN(\SUMB[18][4] ) );
  NAND2_X2 U178 ( .A1(\SUMB[17][6] ), .A2(\CARRYB[17][5] ), .ZN(n91) );
  INV_X4 U179 ( .A(n91), .ZN(\CARRYB[18][5] ) );
  XNOR2_X2 U180 ( .A(\CARRYB[17][5] ), .B(\SUMB[17][6] ), .ZN(n92) );
  INV_X4 U181 ( .A(n92), .ZN(\SUMB[18][5] ) );
  NAND2_X2 U182 ( .A1(\SUMB[17][7] ), .A2(\CARRYB[17][6] ), .ZN(n93) );
  INV_X4 U183 ( .A(n93), .ZN(\CARRYB[18][6] ) );
  XNOR2_X2 U184 ( .A(\CARRYB[17][6] ), .B(\SUMB[17][7] ), .ZN(n94) );
  INV_X4 U185 ( .A(n94), .ZN(\SUMB[18][6] ) );
  NAND2_X2 U186 ( .A1(\SUMB[17][8] ), .A2(\CARRYB[17][7] ), .ZN(n95) );
  INV_X4 U187 ( .A(n95), .ZN(\CARRYB[18][7] ) );
  XNOR2_X2 U188 ( .A(\CARRYB[17][7] ), .B(\SUMB[17][8] ), .ZN(n96) );
  INV_X4 U189 ( .A(n96), .ZN(\SUMB[18][7] ) );
  NAND2_X2 U190 ( .A1(\SUMB[17][9] ), .A2(\CARRYB[17][8] ), .ZN(n97) );
  INV_X4 U191 ( .A(n97), .ZN(\CARRYB[18][8] ) );
  XNOR2_X2 U192 ( .A(\CARRYB[17][8] ), .B(\SUMB[17][9] ), .ZN(n98) );
  INV_X4 U193 ( .A(n98), .ZN(\SUMB[18][8] ) );
  NAND2_X2 U194 ( .A1(\SUMB[16][10] ), .A2(\CARRYB[16][9] ), .ZN(n99) );
  INV_X4 U195 ( .A(n99), .ZN(\CARRYB[17][9] ) );
  XNOR2_X2 U196 ( .A(\CARRYB[16][9] ), .B(\SUMB[16][10] ), .ZN(n100) );
  INV_X4 U197 ( .A(n100), .ZN(\SUMB[17][9] ) );
  NAND2_X2 U198 ( .A1(\SUMB[16][1] ), .A2(\CARRYB[16][0] ), .ZN(n101) );
  INV_X4 U199 ( .A(n101), .ZN(\CARRYB[17][0] ) );
  XNOR2_X2 U200 ( .A(\CARRYB[16][0] ), .B(\SUMB[16][1] ), .ZN(n102) );
  INV_X4 U201 ( .A(n102), .ZN(PRODUCT[17]) );
  NAND2_X2 U202 ( .A1(\SUMB[16][11] ), .A2(\CARRYB[16][10] ), .ZN(n103) );
  INV_X4 U203 ( .A(n103), .ZN(\CARRYB[17][10] ) );
  XNOR2_X2 U204 ( .A(\CARRYB[16][10] ), .B(\SUMB[16][11] ), .ZN(n104) );
  INV_X4 U205 ( .A(n104), .ZN(\SUMB[17][10] ) );
  NAND2_X2 U206 ( .A1(\SUMB[16][12] ), .A2(\CARRYB[16][11] ), .ZN(n105) );
  INV_X4 U207 ( .A(n105), .ZN(\CARRYB[17][11] ) );
  XNOR2_X2 U208 ( .A(\CARRYB[16][11] ), .B(\SUMB[16][12] ), .ZN(n106) );
  INV_X4 U209 ( .A(n106), .ZN(\SUMB[17][11] ) );
  NAND2_X2 U210 ( .A1(\SUMB[16][13] ), .A2(\CARRYB[16][12] ), .ZN(n107) );
  INV_X4 U211 ( .A(n107), .ZN(\CARRYB[17][12] ) );
  XNOR2_X2 U212 ( .A(\CARRYB[16][12] ), .B(\SUMB[16][13] ), .ZN(n108) );
  INV_X4 U213 ( .A(n108), .ZN(\SUMB[17][12] ) );
  NAND2_X2 U214 ( .A1(\SUMB[16][14] ), .A2(\CARRYB[16][13] ), .ZN(n109) );
  INV_X4 U215 ( .A(n109), .ZN(\CARRYB[17][13] ) );
  XNOR2_X2 U216 ( .A(\CARRYB[16][13] ), .B(\SUMB[16][14] ), .ZN(n110) );
  INV_X4 U217 ( .A(n110), .ZN(\SUMB[17][13] ) );
  XNOR2_X2 U218 ( .A(\CARRYB[16][14] ), .B(\SUMB[16][15] ), .ZN(n111) );
  INV_X4 U219 ( .A(n111), .ZN(\SUMB[17][14] ) );
  NAND2_X2 U220 ( .A1(\SUMB[16][2] ), .A2(\CARRYB[16][1] ), .ZN(n112) );
  INV_X4 U221 ( .A(n112), .ZN(\CARRYB[17][1] ) );
  XNOR2_X2 U222 ( .A(\CARRYB[16][1] ), .B(\SUMB[16][2] ), .ZN(n113) );
  INV_X4 U223 ( .A(n113), .ZN(\SUMB[17][1] ) );
  NAND2_X2 U224 ( .A1(\SUMB[16][3] ), .A2(\CARRYB[16][2] ), .ZN(n114) );
  INV_X4 U225 ( .A(n114), .ZN(\CARRYB[17][2] ) );
  XNOR2_X2 U226 ( .A(\CARRYB[16][2] ), .B(\SUMB[16][3] ), .ZN(n115) );
  INV_X4 U227 ( .A(n115), .ZN(\SUMB[17][2] ) );
  NAND2_X2 U228 ( .A1(\SUMB[16][4] ), .A2(\CARRYB[16][3] ), .ZN(n116) );
  INV_X4 U229 ( .A(n116), .ZN(\CARRYB[17][3] ) );
  XNOR2_X2 U230 ( .A(\CARRYB[16][3] ), .B(\SUMB[16][4] ), .ZN(n117) );
  INV_X4 U231 ( .A(n117), .ZN(\SUMB[17][3] ) );
  NAND2_X2 U232 ( .A1(\SUMB[16][5] ), .A2(\CARRYB[16][4] ), .ZN(n118) );
  INV_X4 U233 ( .A(n118), .ZN(\CARRYB[17][4] ) );
  XNOR2_X2 U234 ( .A(\CARRYB[16][4] ), .B(\SUMB[16][5] ), .ZN(n119) );
  INV_X4 U235 ( .A(n119), .ZN(\SUMB[17][4] ) );
  NAND2_X2 U236 ( .A1(\SUMB[16][6] ), .A2(\CARRYB[16][5] ), .ZN(n120) );
  INV_X4 U237 ( .A(n120), .ZN(\CARRYB[17][5] ) );
  XNOR2_X2 U238 ( .A(\CARRYB[16][5] ), .B(\SUMB[16][6] ), .ZN(n121) );
  INV_X4 U239 ( .A(n121), .ZN(\SUMB[17][5] ) );
  NAND2_X2 U240 ( .A1(\SUMB[16][7] ), .A2(\CARRYB[16][6] ), .ZN(n122) );
  INV_X4 U241 ( .A(n122), .ZN(\CARRYB[17][6] ) );
  XNOR2_X2 U242 ( .A(\CARRYB[16][6] ), .B(\SUMB[16][7] ), .ZN(n123) );
  INV_X4 U243 ( .A(n123), .ZN(\SUMB[17][6] ) );
  NAND2_X2 U244 ( .A1(\SUMB[16][8] ), .A2(\CARRYB[16][7] ), .ZN(n124) );
  INV_X4 U245 ( .A(n124), .ZN(\CARRYB[17][7] ) );
  XNOR2_X2 U246 ( .A(\CARRYB[16][7] ), .B(\SUMB[16][8] ), .ZN(n125) );
  INV_X4 U247 ( .A(n125), .ZN(\SUMB[17][7] ) );
  NAND2_X2 U248 ( .A1(\SUMB[16][9] ), .A2(\CARRYB[16][8] ), .ZN(n126) );
  INV_X4 U249 ( .A(n126), .ZN(\CARRYB[17][8] ) );
  XNOR2_X2 U250 ( .A(\CARRYB[16][8] ), .B(\SUMB[16][9] ), .ZN(n127) );
  INV_X4 U251 ( .A(n127), .ZN(\SUMB[17][8] ) );
  XNOR2_X2 U252 ( .A(\CARRYB[29][1] ), .B(\SUMB[29][2] ), .ZN(n128) );
  INV_X4 U253 ( .A(n128), .ZN(\SUMB[30][1] ) );
  NAND2_X2 U254 ( .A1(\SUMB[29][1] ), .A2(\CARRYB[29][0] ), .ZN(n129) );
  INV_X4 U255 ( .A(n129), .ZN(\CARRYB[30][0] ) );
  XNOR2_X2 U256 ( .A(\CARRYB[29][0] ), .B(\SUMB[29][1] ), .ZN(n130) );
  INV_X4 U257 ( .A(n130), .ZN(PRODUCT[30]) );
  XNOR2_X2 U258 ( .A(\CARRYB[28][2] ), .B(\SUMB[28][3] ), .ZN(n131) );
  INV_X4 U259 ( .A(n131), .ZN(\SUMB[29][2] ) );
  NAND2_X2 U260 ( .A1(\SUMB[28][1] ), .A2(\CARRYB[28][0] ), .ZN(n132) );
  INV_X4 U261 ( .A(n132), .ZN(\CARRYB[29][0] ) );
  XNOR2_X2 U262 ( .A(\CARRYB[28][0] ), .B(\SUMB[28][1] ), .ZN(n133) );
  INV_X4 U263 ( .A(n133), .ZN(PRODUCT[29]) );
  NAND2_X2 U264 ( .A1(\SUMB[28][2] ), .A2(\CARRYB[28][1] ), .ZN(n134) );
  INV_X4 U265 ( .A(n134), .ZN(\CARRYB[29][1] ) );
  XNOR2_X2 U266 ( .A(\CARRYB[28][1] ), .B(\SUMB[28][2] ), .ZN(n135) );
  INV_X4 U267 ( .A(n135), .ZN(\SUMB[29][1] ) );
  XNOR2_X2 U268 ( .A(\CARRYB[27][3] ), .B(\SUMB[27][4] ), .ZN(n136) );
  INV_X4 U269 ( .A(n136), .ZN(\SUMB[28][3] ) );
  NAND2_X2 U270 ( .A1(\SUMB[27][1] ), .A2(\CARRYB[27][0] ), .ZN(n137) );
  INV_X4 U271 ( .A(n137), .ZN(\CARRYB[28][0] ) );
  XNOR2_X2 U272 ( .A(\CARRYB[27][0] ), .B(\SUMB[27][1] ), .ZN(n138) );
  INV_X4 U273 ( .A(n138), .ZN(PRODUCT[28]) );
  NAND2_X2 U274 ( .A1(\SUMB[27][2] ), .A2(\CARRYB[27][1] ), .ZN(n139) );
  INV_X4 U275 ( .A(n139), .ZN(\CARRYB[28][1] ) );
  XNOR2_X2 U276 ( .A(\CARRYB[27][1] ), .B(\SUMB[27][2] ), .ZN(n140) );
  INV_X4 U277 ( .A(n140), .ZN(\SUMB[28][1] ) );
  NAND2_X2 U278 ( .A1(\SUMB[27][3] ), .A2(\CARRYB[27][2] ), .ZN(n141) );
  INV_X4 U279 ( .A(n141), .ZN(\CARRYB[28][2] ) );
  XNOR2_X2 U280 ( .A(\CARRYB[27][2] ), .B(\SUMB[27][3] ), .ZN(n142) );
  INV_X4 U281 ( .A(n142), .ZN(\SUMB[28][2] ) );
  XNOR2_X2 U282 ( .A(\CARRYB[26][4] ), .B(\SUMB[26][5] ), .ZN(n143) );
  INV_X4 U283 ( .A(n143), .ZN(\SUMB[27][4] ) );
  NAND2_X2 U284 ( .A1(\SUMB[26][1] ), .A2(\CARRYB[26][0] ), .ZN(n144) );
  INV_X4 U285 ( .A(n144), .ZN(\CARRYB[27][0] ) );
  XNOR2_X2 U286 ( .A(\CARRYB[26][0] ), .B(\SUMB[26][1] ), .ZN(n145) );
  INV_X4 U287 ( .A(n145), .ZN(PRODUCT[27]) );
  NAND2_X2 U288 ( .A1(\SUMB[26][2] ), .A2(\CARRYB[26][1] ), .ZN(n146) );
  INV_X4 U289 ( .A(n146), .ZN(\CARRYB[27][1] ) );
  XNOR2_X2 U290 ( .A(\CARRYB[26][1] ), .B(\SUMB[26][2] ), .ZN(n147) );
  INV_X4 U291 ( .A(n147), .ZN(\SUMB[27][1] ) );
  NAND2_X2 U292 ( .A1(\SUMB[26][3] ), .A2(\CARRYB[26][2] ), .ZN(n148) );
  INV_X4 U293 ( .A(n148), .ZN(\CARRYB[27][2] ) );
  XNOR2_X2 U294 ( .A(\CARRYB[26][2] ), .B(\SUMB[26][3] ), .ZN(n149) );
  INV_X4 U295 ( .A(n149), .ZN(\SUMB[27][2] ) );
  NAND2_X2 U296 ( .A1(\SUMB[26][4] ), .A2(\CARRYB[26][3] ), .ZN(n150) );
  INV_X4 U297 ( .A(n150), .ZN(\CARRYB[27][3] ) );
  XNOR2_X2 U298 ( .A(\CARRYB[26][3] ), .B(\SUMB[26][4] ), .ZN(n151) );
  INV_X4 U299 ( .A(n151), .ZN(\SUMB[27][3] ) );
  XNOR2_X2 U300 ( .A(\CARRYB[25][5] ), .B(\SUMB[25][6] ), .ZN(n152) );
  INV_X4 U301 ( .A(n152), .ZN(\SUMB[26][5] ) );
  NAND2_X2 U302 ( .A1(\SUMB[25][1] ), .A2(\CARRYB[25][0] ), .ZN(n153) );
  INV_X4 U303 ( .A(n153), .ZN(\CARRYB[26][0] ) );
  XNOR2_X2 U304 ( .A(\CARRYB[25][0] ), .B(\SUMB[25][1] ), .ZN(n154) );
  INV_X4 U305 ( .A(n154), .ZN(PRODUCT[26]) );
  NAND2_X2 U306 ( .A1(\SUMB[25][2] ), .A2(\CARRYB[25][1] ), .ZN(n155) );
  INV_X4 U307 ( .A(n155), .ZN(\CARRYB[26][1] ) );
  XNOR2_X2 U308 ( .A(\CARRYB[25][1] ), .B(\SUMB[25][2] ), .ZN(n156) );
  INV_X4 U309 ( .A(n156), .ZN(\SUMB[26][1] ) );
  NAND2_X2 U310 ( .A1(\SUMB[25][3] ), .A2(\CARRYB[25][2] ), .ZN(n157) );
  INV_X4 U311 ( .A(n157), .ZN(\CARRYB[26][2] ) );
  XNOR2_X2 U312 ( .A(\CARRYB[25][2] ), .B(\SUMB[25][3] ), .ZN(n158) );
  INV_X4 U313 ( .A(n158), .ZN(\SUMB[26][2] ) );
  NAND2_X2 U314 ( .A1(\SUMB[25][4] ), .A2(\CARRYB[25][3] ), .ZN(n159) );
  INV_X4 U315 ( .A(n159), .ZN(\CARRYB[26][3] ) );
  XNOR2_X2 U316 ( .A(\CARRYB[25][3] ), .B(\SUMB[25][4] ), .ZN(n160) );
  INV_X4 U317 ( .A(n160), .ZN(\SUMB[26][3] ) );
  NAND2_X2 U318 ( .A1(\SUMB[25][5] ), .A2(\CARRYB[25][4] ), .ZN(n161) );
  INV_X4 U319 ( .A(n161), .ZN(\CARRYB[26][4] ) );
  XNOR2_X2 U320 ( .A(\CARRYB[25][4] ), .B(\SUMB[25][5] ), .ZN(n162) );
  INV_X4 U321 ( .A(n162), .ZN(\SUMB[26][4] ) );
  XNOR2_X2 U322 ( .A(\CARRYB[24][6] ), .B(\SUMB[24][7] ), .ZN(n163) );
  INV_X4 U323 ( .A(n163), .ZN(\SUMB[25][6] ) );
  NAND2_X2 U324 ( .A1(\SUMB[24][1] ), .A2(\CARRYB[24][0] ), .ZN(n164) );
  INV_X4 U325 ( .A(n164), .ZN(\CARRYB[25][0] ) );
  XNOR2_X2 U326 ( .A(\CARRYB[24][0] ), .B(\SUMB[24][1] ), .ZN(n165) );
  INV_X4 U327 ( .A(n165), .ZN(PRODUCT[25]) );
  NAND2_X2 U328 ( .A1(\SUMB[24][2] ), .A2(\CARRYB[24][1] ), .ZN(n166) );
  INV_X4 U329 ( .A(n166), .ZN(\CARRYB[25][1] ) );
  XNOR2_X2 U330 ( .A(\CARRYB[24][1] ), .B(\SUMB[24][2] ), .ZN(n167) );
  INV_X4 U331 ( .A(n167), .ZN(\SUMB[25][1] ) );
  NAND2_X2 U332 ( .A1(\SUMB[24][3] ), .A2(\CARRYB[24][2] ), .ZN(n168) );
  INV_X4 U333 ( .A(n168), .ZN(\CARRYB[25][2] ) );
  XNOR2_X2 U334 ( .A(\CARRYB[24][2] ), .B(\SUMB[24][3] ), .ZN(n169) );
  INV_X4 U335 ( .A(n169), .ZN(\SUMB[25][2] ) );
  NAND2_X2 U336 ( .A1(\SUMB[24][4] ), .A2(\CARRYB[24][3] ), .ZN(n170) );
  INV_X4 U337 ( .A(n170), .ZN(\CARRYB[25][3] ) );
  XNOR2_X2 U338 ( .A(\CARRYB[24][3] ), .B(\SUMB[24][4] ), .ZN(n171) );
  INV_X4 U339 ( .A(n171), .ZN(\SUMB[25][3] ) );
  NAND2_X2 U340 ( .A1(\SUMB[24][5] ), .A2(\CARRYB[24][4] ), .ZN(n172) );
  INV_X4 U341 ( .A(n172), .ZN(\CARRYB[25][4] ) );
  XNOR2_X2 U342 ( .A(\CARRYB[24][4] ), .B(\SUMB[24][5] ), .ZN(n173) );
  INV_X4 U343 ( .A(n173), .ZN(\SUMB[25][4] ) );
  NAND2_X2 U344 ( .A1(\SUMB[24][6] ), .A2(\CARRYB[24][5] ), .ZN(n174) );
  INV_X4 U345 ( .A(n174), .ZN(\CARRYB[25][5] ) );
  XNOR2_X2 U346 ( .A(\CARRYB[24][5] ), .B(\SUMB[24][6] ), .ZN(n175) );
  INV_X4 U347 ( .A(n175), .ZN(\SUMB[25][5] ) );
  XNOR2_X2 U348 ( .A(\CARRYB[23][7] ), .B(\SUMB[23][8] ), .ZN(n176) );
  INV_X4 U349 ( .A(n176), .ZN(\SUMB[24][7] ) );
  NAND2_X2 U350 ( .A1(\SUMB[23][1] ), .A2(\CARRYB[23][0] ), .ZN(n177) );
  INV_X4 U351 ( .A(n177), .ZN(\CARRYB[24][0] ) );
  XNOR2_X2 U352 ( .A(\CARRYB[23][0] ), .B(\SUMB[23][1] ), .ZN(n178) );
  INV_X4 U353 ( .A(n178), .ZN(PRODUCT[24]) );
  NAND2_X2 U354 ( .A1(\SUMB[23][2] ), .A2(\CARRYB[23][1] ), .ZN(n179) );
  INV_X4 U355 ( .A(n179), .ZN(\CARRYB[24][1] ) );
  XNOR2_X2 U356 ( .A(\CARRYB[23][1] ), .B(\SUMB[23][2] ), .ZN(n180) );
  INV_X4 U357 ( .A(n180), .ZN(\SUMB[24][1] ) );
  NAND2_X2 U358 ( .A1(\SUMB[23][3] ), .A2(\CARRYB[23][2] ), .ZN(n181) );
  INV_X4 U359 ( .A(n181), .ZN(\CARRYB[24][2] ) );
  XNOR2_X2 U360 ( .A(\CARRYB[23][2] ), .B(\SUMB[23][3] ), .ZN(n182) );
  INV_X4 U361 ( .A(n182), .ZN(\SUMB[24][2] ) );
  NAND2_X2 U362 ( .A1(\SUMB[23][4] ), .A2(\CARRYB[23][3] ), .ZN(n183) );
  INV_X4 U363 ( .A(n183), .ZN(\CARRYB[24][3] ) );
  XNOR2_X2 U364 ( .A(\CARRYB[23][3] ), .B(\SUMB[23][4] ), .ZN(n184) );
  INV_X4 U365 ( .A(n184), .ZN(\SUMB[24][3] ) );
  NAND2_X2 U366 ( .A1(\SUMB[23][5] ), .A2(\CARRYB[23][4] ), .ZN(n185) );
  INV_X4 U367 ( .A(n185), .ZN(\CARRYB[24][4] ) );
  XNOR2_X2 U368 ( .A(\CARRYB[23][4] ), .B(\SUMB[23][5] ), .ZN(n186) );
  INV_X4 U369 ( .A(n186), .ZN(\SUMB[24][4] ) );
  NAND2_X2 U370 ( .A1(\SUMB[23][6] ), .A2(\CARRYB[23][5] ), .ZN(n187) );
  INV_X4 U371 ( .A(n187), .ZN(\CARRYB[24][5] ) );
  XNOR2_X2 U372 ( .A(\CARRYB[23][5] ), .B(\SUMB[23][6] ), .ZN(n188) );
  INV_X4 U373 ( .A(n188), .ZN(\SUMB[24][5] ) );
  NAND2_X2 U374 ( .A1(\SUMB[23][7] ), .A2(\CARRYB[23][6] ), .ZN(n189) );
  INV_X4 U375 ( .A(n189), .ZN(\CARRYB[24][6] ) );
  XNOR2_X2 U376 ( .A(\CARRYB[23][6] ), .B(\SUMB[23][7] ), .ZN(n190) );
  INV_X4 U377 ( .A(n190), .ZN(\SUMB[24][6] ) );
  XNOR2_X2 U378 ( .A(\CARRYB[22][8] ), .B(\SUMB[22][9] ), .ZN(n191) );
  INV_X4 U379 ( .A(n191), .ZN(\SUMB[23][8] ) );
  NAND2_X2 U380 ( .A1(\SUMB[22][1] ), .A2(\CARRYB[22][0] ), .ZN(n192) );
  INV_X4 U381 ( .A(n192), .ZN(\CARRYB[23][0] ) );
  XNOR2_X2 U382 ( .A(\CARRYB[22][0] ), .B(\SUMB[22][1] ), .ZN(n193) );
  INV_X4 U383 ( .A(n193), .ZN(PRODUCT[23]) );
  NAND2_X2 U384 ( .A1(\SUMB[22][2] ), .A2(\CARRYB[22][1] ), .ZN(n194) );
  INV_X4 U385 ( .A(n194), .ZN(\CARRYB[23][1] ) );
  XNOR2_X2 U386 ( .A(\CARRYB[22][1] ), .B(\SUMB[22][2] ), .ZN(n195) );
  INV_X4 U387 ( .A(n195), .ZN(\SUMB[23][1] ) );
  NAND2_X2 U388 ( .A1(\SUMB[22][3] ), .A2(\CARRYB[22][2] ), .ZN(n196) );
  INV_X4 U389 ( .A(n196), .ZN(\CARRYB[23][2] ) );
  XNOR2_X2 U390 ( .A(\CARRYB[22][2] ), .B(\SUMB[22][3] ), .ZN(n197) );
  INV_X4 U391 ( .A(n197), .ZN(\SUMB[23][2] ) );
  NAND2_X2 U392 ( .A1(\SUMB[22][4] ), .A2(\CARRYB[22][3] ), .ZN(n198) );
  INV_X4 U393 ( .A(n198), .ZN(\CARRYB[23][3] ) );
  XNOR2_X2 U394 ( .A(\CARRYB[22][3] ), .B(\SUMB[22][4] ), .ZN(n199) );
  INV_X4 U395 ( .A(n199), .ZN(\SUMB[23][3] ) );
  NAND2_X2 U396 ( .A1(\SUMB[22][5] ), .A2(\CARRYB[22][4] ), .ZN(n200) );
  INV_X4 U397 ( .A(n200), .ZN(\CARRYB[23][4] ) );
  XNOR2_X2 U398 ( .A(\CARRYB[22][4] ), .B(\SUMB[22][5] ), .ZN(n201) );
  INV_X4 U399 ( .A(n201), .ZN(\SUMB[23][4] ) );
  NAND2_X2 U400 ( .A1(\SUMB[22][6] ), .A2(\CARRYB[22][5] ), .ZN(n202) );
  INV_X4 U401 ( .A(n202), .ZN(\CARRYB[23][5] ) );
  XNOR2_X2 U402 ( .A(\CARRYB[22][5] ), .B(\SUMB[22][6] ), .ZN(n203) );
  INV_X4 U403 ( .A(n203), .ZN(\SUMB[23][5] ) );
  NAND2_X2 U404 ( .A1(\SUMB[22][7] ), .A2(\CARRYB[22][6] ), .ZN(n204) );
  INV_X4 U405 ( .A(n204), .ZN(\CARRYB[23][6] ) );
  XNOR2_X2 U406 ( .A(\CARRYB[22][6] ), .B(\SUMB[22][7] ), .ZN(n205) );
  INV_X4 U407 ( .A(n205), .ZN(\SUMB[23][6] ) );
  NAND2_X2 U408 ( .A1(\SUMB[22][8] ), .A2(\CARRYB[22][7] ), .ZN(n206) );
  INV_X4 U409 ( .A(n206), .ZN(\CARRYB[23][7] ) );
  XNOR2_X2 U410 ( .A(\CARRYB[22][7] ), .B(\SUMB[22][8] ), .ZN(n207) );
  INV_X4 U411 ( .A(n207), .ZN(\SUMB[23][7] ) );
  XNOR2_X2 U412 ( .A(\CARRYB[21][9] ), .B(\SUMB[21][10] ), .ZN(n208) );
  INV_X4 U413 ( .A(n208), .ZN(\SUMB[22][9] ) );
  NAND2_X2 U414 ( .A1(\SUMB[21][1] ), .A2(\CARRYB[21][0] ), .ZN(n209) );
  INV_X4 U415 ( .A(n209), .ZN(\CARRYB[22][0] ) );
  XNOR2_X2 U416 ( .A(\CARRYB[21][0] ), .B(\SUMB[21][1] ), .ZN(n210) );
  INV_X4 U417 ( .A(n210), .ZN(PRODUCT[22]) );
  NAND2_X2 U418 ( .A1(\SUMB[21][2] ), .A2(\CARRYB[21][1] ), .ZN(n211) );
  INV_X4 U419 ( .A(n211), .ZN(\CARRYB[22][1] ) );
  XNOR2_X2 U420 ( .A(\CARRYB[21][1] ), .B(\SUMB[21][2] ), .ZN(n212) );
  INV_X4 U421 ( .A(n212), .ZN(\SUMB[22][1] ) );
  NAND2_X2 U422 ( .A1(\SUMB[21][3] ), .A2(\CARRYB[21][2] ), .ZN(n213) );
  INV_X4 U423 ( .A(n213), .ZN(\CARRYB[22][2] ) );
  XNOR2_X2 U424 ( .A(\CARRYB[21][2] ), .B(\SUMB[21][3] ), .ZN(n214) );
  INV_X4 U425 ( .A(n214), .ZN(\SUMB[22][2] ) );
  NAND2_X2 U426 ( .A1(\SUMB[21][4] ), .A2(\CARRYB[21][3] ), .ZN(n215) );
  INV_X4 U427 ( .A(n215), .ZN(\CARRYB[22][3] ) );
  XNOR2_X2 U428 ( .A(\CARRYB[21][3] ), .B(\SUMB[21][4] ), .ZN(n216) );
  INV_X4 U429 ( .A(n216), .ZN(\SUMB[22][3] ) );
  NAND2_X2 U430 ( .A1(\SUMB[21][5] ), .A2(\CARRYB[21][4] ), .ZN(n217) );
  INV_X4 U431 ( .A(n217), .ZN(\CARRYB[22][4] ) );
  XNOR2_X2 U432 ( .A(\CARRYB[21][4] ), .B(\SUMB[21][5] ), .ZN(n218) );
  INV_X4 U433 ( .A(n218), .ZN(\SUMB[22][4] ) );
  NAND2_X2 U434 ( .A1(\SUMB[21][6] ), .A2(\CARRYB[21][5] ), .ZN(n219) );
  INV_X4 U435 ( .A(n219), .ZN(\CARRYB[22][5] ) );
  XNOR2_X2 U436 ( .A(\CARRYB[21][5] ), .B(\SUMB[21][6] ), .ZN(n220) );
  INV_X4 U437 ( .A(n220), .ZN(\SUMB[22][5] ) );
  NAND2_X2 U438 ( .A1(\SUMB[21][7] ), .A2(\CARRYB[21][6] ), .ZN(n221) );
  INV_X4 U439 ( .A(n221), .ZN(\CARRYB[22][6] ) );
  XNOR2_X2 U440 ( .A(\CARRYB[21][6] ), .B(\SUMB[21][7] ), .ZN(n222) );
  INV_X4 U441 ( .A(n222), .ZN(\SUMB[22][6] ) );
  NAND2_X2 U442 ( .A1(\SUMB[21][8] ), .A2(\CARRYB[21][7] ), .ZN(n223) );
  INV_X4 U443 ( .A(n223), .ZN(\CARRYB[22][7] ) );
  XNOR2_X2 U444 ( .A(\CARRYB[21][7] ), .B(\SUMB[21][8] ), .ZN(n224) );
  INV_X4 U445 ( .A(n224), .ZN(\SUMB[22][7] ) );
  NAND2_X2 U446 ( .A1(\SUMB[21][9] ), .A2(\CARRYB[21][8] ), .ZN(n225) );
  INV_X4 U447 ( .A(n225), .ZN(\CARRYB[22][8] ) );
  XNOR2_X2 U448 ( .A(\CARRYB[21][8] ), .B(\SUMB[21][9] ), .ZN(n226) );
  INV_X4 U449 ( .A(n226), .ZN(\SUMB[22][8] ) );
  XNOR2_X2 U450 ( .A(\CARRYB[30][0] ), .B(\SUMB[30][1] ), .ZN(n227) );
  INV_X4 U451 ( .A(n227), .ZN(PRODUCT[31]) );
  INV_X4 U452 ( .A(B[8]), .ZN(n277) );
  INV_X4 U453 ( .A(B[9]), .ZN(n276) );
  INV_X4 U454 ( .A(B[7]), .ZN(n278) );
  INV_X4 U455 ( .A(B[10]), .ZN(n275) );
  INV_X4 U456 ( .A(B[11]), .ZN(n274) );
  INV_X4 U457 ( .A(B[6]), .ZN(n279) );
  INV_X4 U458 ( .A(B[12]), .ZN(n273) );
  INV_X4 U459 ( .A(B[5]), .ZN(n280) );
  INV_X4 U460 ( .A(B[16]), .ZN(n269) );
  INV_X4 U461 ( .A(B[13]), .ZN(n272) );
  INV_X4 U462 ( .A(B[4]), .ZN(n281) );
  INV_X4 U463 ( .A(B[14]), .ZN(n271) );
  INV_X4 U464 ( .A(B[15]), .ZN(n270) );
  INV_X4 U465 ( .A(A[4]), .ZN(n297) );
  INV_X4 U466 ( .A(A[5]), .ZN(n296) );
  INV_X4 U467 ( .A(A[6]), .ZN(n295) );
  INV_X4 U468 ( .A(A[7]), .ZN(n294) );
  INV_X4 U469 ( .A(A[8]), .ZN(n293) );
  INV_X4 U470 ( .A(A[9]), .ZN(n292) );
  INV_X4 U471 ( .A(A[10]), .ZN(n291) );
  INV_X4 U472 ( .A(A[11]), .ZN(n290) );
  INV_X4 U473 ( .A(A[12]), .ZN(n289) );
  INV_X4 U474 ( .A(A[13]), .ZN(n288) );
  INV_X4 U475 ( .A(A[14]), .ZN(n287) );
  INV_X4 U476 ( .A(A[15]), .ZN(n286) );
  INV_X4 U477 ( .A(A[16]), .ZN(n285) );
  INV_X4 U478 ( .A(B[1]), .ZN(n262) );
  AND2_X4 U479 ( .A1(\ab[0][16] ), .A2(\ab[1][15] ), .ZN(n228) );
  AND2_X4 U480 ( .A1(\ab[0][15] ), .A2(\ab[1][14] ), .ZN(n229) );
  AND2_X4 U481 ( .A1(\ab[0][14] ), .A2(\ab[1][13] ), .ZN(n230) );
  AND2_X4 U482 ( .A1(\ab[0][13] ), .A2(\ab[1][12] ), .ZN(n231) );
  AND2_X4 U483 ( .A1(\ab[0][12] ), .A2(\ab[1][11] ), .ZN(n232) );
  AND2_X4 U484 ( .A1(\ab[0][11] ), .A2(\ab[1][10] ), .ZN(n233) );
  AND2_X4 U485 ( .A1(\ab[0][10] ), .A2(\ab[1][9] ), .ZN(n234) );
  AND2_X4 U486 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .ZN(n235) );
  AND2_X4 U487 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .ZN(n236) );
  AND2_X4 U488 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .ZN(n237) );
  AND2_X4 U489 ( .A1(\ab[0][7] ), .A2(\ab[1][6] ), .ZN(n238) );
  AND2_X4 U490 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .ZN(n239) );
  AND2_X4 U491 ( .A1(\ab[0][5] ), .A2(\ab[1][4] ), .ZN(n240) );
  AND2_X4 U492 ( .A1(\ab[0][4] ), .A2(\ab[1][3] ), .ZN(n241) );
  AND2_X4 U493 ( .A1(\ab[0][3] ), .A2(\ab[1][2] ), .ZN(n242) );
  AND2_X4 U494 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .ZN(n243) );
  XOR2_X2 U495 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(n244) );
  XOR2_X2 U496 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(n245) );
  XOR2_X2 U497 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(n246) );
  XOR2_X2 U498 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(n247) );
  XOR2_X2 U499 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(n248) );
  XOR2_X2 U500 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(n249) );
  XOR2_X2 U501 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(n250) );
  XOR2_X2 U502 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(n251) );
  XOR2_X2 U503 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(n252) );
  XOR2_X2 U504 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(n253) );
  XOR2_X2 U505 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(n254) );
  XOR2_X2 U506 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(n255) );
  XOR2_X2 U507 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(n256) );
  XOR2_X2 U508 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(n257) );
  XOR2_X2 U509 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(n258) );
  XOR2_X2 U510 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  INV_X4 U511 ( .A(B[3]), .ZN(n260) );
  INV_X4 U512 ( .A(A[3]), .ZN(n265) );
  INV_X4 U513 ( .A(A[3]), .ZN(n264) );
  INV_X4 U514 ( .A(B[2]), .ZN(n261) );
  INV_X4 U515 ( .A(B[0]), .ZN(n263) );
  INV_X4 U516 ( .A(A[2]), .ZN(n266) );
  INV_X4 U517 ( .A(A[1]), .ZN(n267) );
  INV_X4 U518 ( .A(A[0]), .ZN(n268) );
  INV_X4 U519 ( .A(B[3]), .ZN(n282) );
  INV_X4 U520 ( .A(B[2]), .ZN(n283) );
  INV_X4 U521 ( .A(B[0]), .ZN(n284) );
  INV_X4 U522 ( .A(A[2]), .ZN(n298) );
  INV_X4 U523 ( .A(A[1]), .ZN(n299) );
  INV_X4 U524 ( .A(A[0]), .ZN(n300) );
  NOR2_X1 U525 ( .A1(n292), .A2(n276), .ZN(\ab[9][9] ) );
  NOR2_X1 U526 ( .A1(n292), .A2(n277), .ZN(\ab[9][8] ) );
  NOR2_X1 U527 ( .A1(n292), .A2(n278), .ZN(\ab[9][7] ) );
  NOR2_X1 U528 ( .A1(n292), .A2(n279), .ZN(\ab[9][6] ) );
  NOR2_X1 U529 ( .A1(n292), .A2(n280), .ZN(\ab[9][5] ) );
  NOR2_X1 U530 ( .A1(n292), .A2(n281), .ZN(\ab[9][4] ) );
  NOR2_X1 U531 ( .A1(n292), .A2(n260), .ZN(\ab[9][3] ) );
  NOR2_X1 U532 ( .A1(n292), .A2(n261), .ZN(\ab[9][2] ) );
  NOR2_X1 U533 ( .A1(n292), .A2(n262), .ZN(\ab[9][1] ) );
  NOR2_X1 U534 ( .A1(n292), .A2(n269), .ZN(\SUMB[9][16] ) );
  NOR2_X1 U535 ( .A1(n292), .A2(n270), .ZN(\ab[9][15] ) );
  NOR2_X1 U536 ( .A1(n292), .A2(n271), .ZN(\ab[9][14] ) );
  NOR2_X1 U537 ( .A1(n292), .A2(n272), .ZN(\ab[9][13] ) );
  NOR2_X1 U538 ( .A1(n292), .A2(n273), .ZN(\ab[9][12] ) );
  NOR2_X1 U539 ( .A1(n292), .A2(n274), .ZN(\ab[9][11] ) );
  NOR2_X1 U540 ( .A1(n292), .A2(n275), .ZN(\ab[9][10] ) );
  NOR2_X1 U541 ( .A1(n292), .A2(n263), .ZN(\ab[9][0] ) );
  NOR2_X1 U542 ( .A1(n276), .A2(n293), .ZN(\ab[8][9] ) );
  NOR2_X1 U543 ( .A1(n277), .A2(n293), .ZN(\ab[8][8] ) );
  NOR2_X1 U544 ( .A1(n278), .A2(n293), .ZN(\ab[8][7] ) );
  NOR2_X1 U545 ( .A1(n279), .A2(n293), .ZN(\ab[8][6] ) );
  NOR2_X1 U546 ( .A1(n280), .A2(n293), .ZN(\ab[8][5] ) );
  NOR2_X1 U547 ( .A1(n281), .A2(n293), .ZN(\ab[8][4] ) );
  NOR2_X1 U548 ( .A1(n260), .A2(n293), .ZN(\ab[8][3] ) );
  NOR2_X1 U549 ( .A1(n261), .A2(n293), .ZN(\ab[8][2] ) );
  NOR2_X1 U550 ( .A1(n262), .A2(n293), .ZN(\ab[8][1] ) );
  NOR2_X1 U551 ( .A1(n269), .A2(n293), .ZN(\SUMB[8][16] ) );
  NOR2_X1 U552 ( .A1(n270), .A2(n293), .ZN(\ab[8][15] ) );
  NOR2_X1 U553 ( .A1(n271), .A2(n293), .ZN(\ab[8][14] ) );
  NOR2_X1 U554 ( .A1(n272), .A2(n293), .ZN(\ab[8][13] ) );
  NOR2_X1 U555 ( .A1(n273), .A2(n293), .ZN(\ab[8][12] ) );
  NOR2_X1 U556 ( .A1(n274), .A2(n293), .ZN(\ab[8][11] ) );
  NOR2_X1 U557 ( .A1(n275), .A2(n293), .ZN(\ab[8][10] ) );
  NOR2_X1 U558 ( .A1(n263), .A2(n293), .ZN(\ab[8][0] ) );
  NOR2_X1 U559 ( .A1(n276), .A2(n294), .ZN(\ab[7][9] ) );
  NOR2_X1 U560 ( .A1(n277), .A2(n294), .ZN(\ab[7][8] ) );
  NOR2_X1 U561 ( .A1(n278), .A2(n294), .ZN(\ab[7][7] ) );
  NOR2_X1 U562 ( .A1(n279), .A2(n294), .ZN(\ab[7][6] ) );
  NOR2_X1 U563 ( .A1(n280), .A2(n294), .ZN(\ab[7][5] ) );
  NOR2_X1 U564 ( .A1(n281), .A2(n294), .ZN(\ab[7][4] ) );
  NOR2_X1 U565 ( .A1(n260), .A2(n294), .ZN(\ab[7][3] ) );
  NOR2_X1 U566 ( .A1(n261), .A2(n294), .ZN(\ab[7][2] ) );
  NOR2_X1 U567 ( .A1(n262), .A2(n294), .ZN(\ab[7][1] ) );
  NOR2_X1 U568 ( .A1(n269), .A2(n294), .ZN(\SUMB[7][16] ) );
  NOR2_X1 U569 ( .A1(n270), .A2(n294), .ZN(\ab[7][15] ) );
  NOR2_X1 U570 ( .A1(n271), .A2(n294), .ZN(\ab[7][14] ) );
  NOR2_X1 U571 ( .A1(n272), .A2(n294), .ZN(\ab[7][13] ) );
  NOR2_X1 U572 ( .A1(n273), .A2(n294), .ZN(\ab[7][12] ) );
  NOR2_X1 U573 ( .A1(n274), .A2(n294), .ZN(\ab[7][11] ) );
  NOR2_X1 U574 ( .A1(n275), .A2(n294), .ZN(\ab[7][10] ) );
  NOR2_X1 U575 ( .A1(n263), .A2(n294), .ZN(\ab[7][0] ) );
  NOR2_X1 U576 ( .A1(n276), .A2(n295), .ZN(\ab[6][9] ) );
  NOR2_X1 U577 ( .A1(n277), .A2(n295), .ZN(\ab[6][8] ) );
  NOR2_X1 U578 ( .A1(n278), .A2(n295), .ZN(\ab[6][7] ) );
  NOR2_X1 U579 ( .A1(n279), .A2(n295), .ZN(\ab[6][6] ) );
  NOR2_X1 U580 ( .A1(n280), .A2(n295), .ZN(\ab[6][5] ) );
  NOR2_X1 U581 ( .A1(n281), .A2(n295), .ZN(\ab[6][4] ) );
  NOR2_X1 U582 ( .A1(n260), .A2(n295), .ZN(\ab[6][3] ) );
  NOR2_X1 U583 ( .A1(n261), .A2(n295), .ZN(\ab[6][2] ) );
  NOR2_X1 U584 ( .A1(n262), .A2(n295), .ZN(\ab[6][1] ) );
  NOR2_X1 U585 ( .A1(n269), .A2(n295), .ZN(\SUMB[6][16] ) );
  NOR2_X1 U586 ( .A1(n270), .A2(n295), .ZN(\ab[6][15] ) );
  NOR2_X1 U587 ( .A1(n271), .A2(n295), .ZN(\ab[6][14] ) );
  NOR2_X1 U588 ( .A1(n272), .A2(n295), .ZN(\ab[6][13] ) );
  NOR2_X1 U589 ( .A1(n273), .A2(n295), .ZN(\ab[6][12] ) );
  NOR2_X1 U590 ( .A1(n274), .A2(n295), .ZN(\ab[6][11] ) );
  NOR2_X1 U591 ( .A1(n275), .A2(n295), .ZN(\ab[6][10] ) );
  NOR2_X1 U592 ( .A1(n263), .A2(n295), .ZN(\ab[6][0] ) );
  NOR2_X1 U593 ( .A1(n276), .A2(n296), .ZN(\ab[5][9] ) );
  NOR2_X1 U594 ( .A1(n277), .A2(n296), .ZN(\ab[5][8] ) );
  NOR2_X1 U595 ( .A1(n278), .A2(n296), .ZN(\ab[5][7] ) );
  NOR2_X1 U596 ( .A1(n279), .A2(n296), .ZN(\ab[5][6] ) );
  NOR2_X1 U597 ( .A1(n280), .A2(n296), .ZN(\ab[5][5] ) );
  NOR2_X1 U598 ( .A1(n281), .A2(n296), .ZN(\ab[5][4] ) );
  NOR2_X1 U599 ( .A1(n260), .A2(n296), .ZN(\ab[5][3] ) );
  NOR2_X1 U600 ( .A1(n261), .A2(n296), .ZN(\ab[5][2] ) );
  NOR2_X1 U601 ( .A1(n262), .A2(n296), .ZN(\ab[5][1] ) );
  NOR2_X1 U602 ( .A1(n269), .A2(n296), .ZN(\SUMB[5][16] ) );
  NOR2_X1 U603 ( .A1(n270), .A2(n296), .ZN(\ab[5][15] ) );
  NOR2_X1 U604 ( .A1(n271), .A2(n296), .ZN(\ab[5][14] ) );
  NOR2_X1 U605 ( .A1(n272), .A2(n296), .ZN(\ab[5][13] ) );
  NOR2_X1 U606 ( .A1(n273), .A2(n296), .ZN(\ab[5][12] ) );
  NOR2_X1 U607 ( .A1(n274), .A2(n296), .ZN(\ab[5][11] ) );
  NOR2_X1 U608 ( .A1(n275), .A2(n296), .ZN(\ab[5][10] ) );
  NOR2_X1 U609 ( .A1(n263), .A2(n296), .ZN(\ab[5][0] ) );
  NOR2_X1 U610 ( .A1(n276), .A2(n297), .ZN(\ab[4][9] ) );
  NOR2_X1 U611 ( .A1(n277), .A2(n297), .ZN(\ab[4][8] ) );
  NOR2_X1 U612 ( .A1(n278), .A2(n297), .ZN(\ab[4][7] ) );
  NOR2_X1 U613 ( .A1(n279), .A2(n297), .ZN(\ab[4][6] ) );
  NOR2_X1 U614 ( .A1(n280), .A2(n297), .ZN(\ab[4][5] ) );
  NOR2_X1 U615 ( .A1(n281), .A2(n297), .ZN(\ab[4][4] ) );
  NOR2_X1 U616 ( .A1(n260), .A2(n297), .ZN(\ab[4][3] ) );
  NOR2_X1 U617 ( .A1(n261), .A2(n297), .ZN(\ab[4][2] ) );
  NOR2_X1 U618 ( .A1(n262), .A2(n297), .ZN(\ab[4][1] ) );
  NOR2_X1 U619 ( .A1(n269), .A2(n297), .ZN(\SUMB[4][16] ) );
  NOR2_X1 U620 ( .A1(n270), .A2(n297), .ZN(\ab[4][15] ) );
  NOR2_X1 U621 ( .A1(n271), .A2(n297), .ZN(\ab[4][14] ) );
  NOR2_X1 U622 ( .A1(n272), .A2(n297), .ZN(\ab[4][13] ) );
  NOR2_X1 U623 ( .A1(n273), .A2(n297), .ZN(\ab[4][12] ) );
  NOR2_X1 U624 ( .A1(n274), .A2(n297), .ZN(\ab[4][11] ) );
  NOR2_X1 U625 ( .A1(n275), .A2(n297), .ZN(\ab[4][10] ) );
  NOR2_X1 U626 ( .A1(n263), .A2(n297), .ZN(\ab[4][0] ) );
  NOR2_X1 U627 ( .A1(n276), .A2(n265), .ZN(\ab[3][9] ) );
  NOR2_X1 U628 ( .A1(n277), .A2(n265), .ZN(\ab[3][8] ) );
  NOR2_X1 U629 ( .A1(n278), .A2(n265), .ZN(\ab[3][7] ) );
  NOR2_X1 U630 ( .A1(n279), .A2(n265), .ZN(\ab[3][6] ) );
  NOR2_X1 U631 ( .A1(n280), .A2(n265), .ZN(\ab[3][5] ) );
  NOR2_X1 U632 ( .A1(n281), .A2(n265), .ZN(\ab[3][4] ) );
  NOR2_X1 U633 ( .A1(n260), .A2(n265), .ZN(\ab[3][3] ) );
  NOR2_X1 U634 ( .A1(n261), .A2(n265), .ZN(\ab[3][2] ) );
  NOR2_X1 U635 ( .A1(n262), .A2(n264), .ZN(\ab[3][1] ) );
  NOR2_X1 U636 ( .A1(n269), .A2(n264), .ZN(\SUMB[3][16] ) );
  NOR2_X1 U637 ( .A1(n270), .A2(n264), .ZN(\ab[3][15] ) );
  NOR2_X1 U638 ( .A1(n271), .A2(n264), .ZN(\ab[3][14] ) );
  NOR2_X1 U639 ( .A1(n272), .A2(n264), .ZN(\ab[3][13] ) );
  NOR2_X1 U640 ( .A1(n273), .A2(n264), .ZN(\ab[3][12] ) );
  NOR2_X1 U641 ( .A1(n274), .A2(n264), .ZN(\ab[3][11] ) );
  NOR2_X1 U642 ( .A1(n275), .A2(n264), .ZN(\ab[3][10] ) );
  NOR2_X1 U643 ( .A1(n263), .A2(n264), .ZN(\ab[3][0] ) );
  NOR2_X1 U644 ( .A1(n276), .A2(n298), .ZN(\ab[2][9] ) );
  NOR2_X1 U645 ( .A1(n277), .A2(n298), .ZN(\ab[2][8] ) );
  NOR2_X1 U646 ( .A1(n278), .A2(n298), .ZN(\ab[2][7] ) );
  NOR2_X1 U647 ( .A1(n279), .A2(n298), .ZN(\ab[2][6] ) );
  NOR2_X1 U648 ( .A1(n280), .A2(n298), .ZN(\ab[2][5] ) );
  NOR2_X1 U649 ( .A1(n281), .A2(n298), .ZN(\ab[2][4] ) );
  NOR2_X1 U650 ( .A1(n260), .A2(n298), .ZN(\ab[2][3] ) );
  NOR2_X1 U651 ( .A1(n261), .A2(n266), .ZN(\ab[2][2] ) );
  NOR2_X1 U652 ( .A1(n262), .A2(n266), .ZN(\ab[2][1] ) );
  NOR2_X1 U653 ( .A1(n269), .A2(n266), .ZN(\SUMB[2][16] ) );
  NOR2_X1 U654 ( .A1(n270), .A2(n266), .ZN(\ab[2][15] ) );
  NOR2_X1 U655 ( .A1(n271), .A2(n266), .ZN(\ab[2][14] ) );
  NOR2_X1 U656 ( .A1(n272), .A2(n266), .ZN(\ab[2][13] ) );
  NOR2_X1 U657 ( .A1(n273), .A2(n266), .ZN(\ab[2][12] ) );
  NOR2_X1 U658 ( .A1(n274), .A2(n266), .ZN(\ab[2][11] ) );
  NOR2_X1 U659 ( .A1(n275), .A2(n266), .ZN(\ab[2][10] ) );
  NOR2_X1 U660 ( .A1(n263), .A2(n266), .ZN(\ab[2][0] ) );
  NOR2_X1 U661 ( .A1(n276), .A2(n299), .ZN(\ab[1][9] ) );
  NOR2_X1 U662 ( .A1(n277), .A2(n299), .ZN(\ab[1][8] ) );
  NOR2_X1 U663 ( .A1(n278), .A2(n299), .ZN(\ab[1][7] ) );
  NOR2_X1 U664 ( .A1(n279), .A2(n299), .ZN(\ab[1][6] ) );
  NOR2_X1 U665 ( .A1(n280), .A2(n299), .ZN(\ab[1][5] ) );
  NOR2_X1 U666 ( .A1(n281), .A2(n299), .ZN(\ab[1][4] ) );
  NOR2_X1 U667 ( .A1(n260), .A2(n299), .ZN(\ab[1][3] ) );
  NOR2_X1 U668 ( .A1(n261), .A2(n267), .ZN(\ab[1][2] ) );
  NOR2_X1 U669 ( .A1(n262), .A2(n267), .ZN(\ab[1][1] ) );
  NOR2_X1 U670 ( .A1(n269), .A2(n267), .ZN(\ab[1][16] ) );
  NOR2_X1 U671 ( .A1(n270), .A2(n267), .ZN(\ab[1][15] ) );
  NOR2_X1 U672 ( .A1(n271), .A2(n267), .ZN(\ab[1][14] ) );
  NOR2_X1 U673 ( .A1(n272), .A2(n267), .ZN(\ab[1][13] ) );
  NOR2_X1 U674 ( .A1(n273), .A2(n267), .ZN(\ab[1][12] ) );
  NOR2_X1 U675 ( .A1(n274), .A2(n267), .ZN(\ab[1][11] ) );
  NOR2_X1 U676 ( .A1(n275), .A2(n267), .ZN(\ab[1][10] ) );
  NOR2_X1 U677 ( .A1(n263), .A2(n267), .ZN(\ab[1][0] ) );
  NOR2_X1 U678 ( .A1(n276), .A2(n285), .ZN(\ab[16][9] ) );
  NOR2_X1 U679 ( .A1(n277), .A2(n285), .ZN(\ab[16][8] ) );
  NOR2_X1 U680 ( .A1(n278), .A2(n285), .ZN(\ab[16][7] ) );
  NOR2_X1 U681 ( .A1(n279), .A2(n285), .ZN(\ab[16][6] ) );
  NOR2_X1 U682 ( .A1(n280), .A2(n285), .ZN(\ab[16][5] ) );
  NOR2_X1 U683 ( .A1(n281), .A2(n285), .ZN(\ab[16][4] ) );
  NOR2_X1 U684 ( .A1(n282), .A2(n285), .ZN(\ab[16][3] ) );
  NOR2_X1 U685 ( .A1(n283), .A2(n285), .ZN(\ab[16][2] ) );
  NOR2_X1 U686 ( .A1(n262), .A2(n285), .ZN(\ab[16][1] ) );
  NOR2_X1 U687 ( .A1(n270), .A2(n285), .ZN(\ab[16][15] ) );
  NOR2_X1 U688 ( .A1(n271), .A2(n285), .ZN(\ab[16][14] ) );
  NOR2_X1 U689 ( .A1(n272), .A2(n285), .ZN(\ab[16][13] ) );
  NOR2_X1 U690 ( .A1(n273), .A2(n285), .ZN(\ab[16][12] ) );
  NOR2_X1 U691 ( .A1(n274), .A2(n285), .ZN(\ab[16][11] ) );
  NOR2_X1 U692 ( .A1(n275), .A2(n285), .ZN(\ab[16][10] ) );
  NOR2_X1 U693 ( .A1(n284), .A2(n285), .ZN(\ab[16][0] ) );
  NOR2_X1 U694 ( .A1(n276), .A2(n286), .ZN(\ab[15][9] ) );
  NOR2_X1 U695 ( .A1(n277), .A2(n286), .ZN(\ab[15][8] ) );
  NOR2_X1 U696 ( .A1(n278), .A2(n286), .ZN(\ab[15][7] ) );
  NOR2_X1 U697 ( .A1(n279), .A2(n286), .ZN(\ab[15][6] ) );
  NOR2_X1 U698 ( .A1(n280), .A2(n286), .ZN(\ab[15][5] ) );
  NOR2_X1 U699 ( .A1(n281), .A2(n286), .ZN(\ab[15][4] ) );
  NOR2_X1 U700 ( .A1(n282), .A2(n286), .ZN(\ab[15][3] ) );
  NOR2_X1 U701 ( .A1(n283), .A2(n286), .ZN(\ab[15][2] ) );
  NOR2_X1 U702 ( .A1(n262), .A2(n286), .ZN(\ab[15][1] ) );
  NOR2_X1 U703 ( .A1(n269), .A2(n286), .ZN(\SUMB[15][16] ) );
  NOR2_X1 U704 ( .A1(n270), .A2(n286), .ZN(\ab[15][15] ) );
  NOR2_X1 U705 ( .A1(n271), .A2(n286), .ZN(\ab[15][14] ) );
  NOR2_X1 U706 ( .A1(n272), .A2(n286), .ZN(\ab[15][13] ) );
  NOR2_X1 U707 ( .A1(n273), .A2(n286), .ZN(\ab[15][12] ) );
  NOR2_X1 U708 ( .A1(n274), .A2(n286), .ZN(\ab[15][11] ) );
  NOR2_X1 U709 ( .A1(n275), .A2(n286), .ZN(\ab[15][10] ) );
  NOR2_X1 U710 ( .A1(n284), .A2(n286), .ZN(\ab[15][0] ) );
  NOR2_X1 U711 ( .A1(n276), .A2(n287), .ZN(\ab[14][9] ) );
  NOR2_X1 U712 ( .A1(n277), .A2(n287), .ZN(\ab[14][8] ) );
  NOR2_X1 U713 ( .A1(n278), .A2(n287), .ZN(\ab[14][7] ) );
  NOR2_X1 U714 ( .A1(n279), .A2(n287), .ZN(\ab[14][6] ) );
  NOR2_X1 U715 ( .A1(n280), .A2(n287), .ZN(\ab[14][5] ) );
  NOR2_X1 U716 ( .A1(n281), .A2(n287), .ZN(\ab[14][4] ) );
  NOR2_X1 U717 ( .A1(n282), .A2(n287), .ZN(\ab[14][3] ) );
  NOR2_X1 U718 ( .A1(n283), .A2(n287), .ZN(\ab[14][2] ) );
  NOR2_X1 U719 ( .A1(n262), .A2(n287), .ZN(\ab[14][1] ) );
  NOR2_X1 U720 ( .A1(n269), .A2(n287), .ZN(\SUMB[14][16] ) );
  NOR2_X1 U721 ( .A1(n270), .A2(n287), .ZN(\ab[14][15] ) );
  NOR2_X1 U722 ( .A1(n271), .A2(n287), .ZN(\ab[14][14] ) );
  NOR2_X1 U723 ( .A1(n272), .A2(n287), .ZN(\ab[14][13] ) );
  NOR2_X1 U724 ( .A1(n273), .A2(n287), .ZN(\ab[14][12] ) );
  NOR2_X1 U725 ( .A1(n274), .A2(n287), .ZN(\ab[14][11] ) );
  NOR2_X1 U726 ( .A1(n275), .A2(n287), .ZN(\ab[14][10] ) );
  NOR2_X1 U727 ( .A1(n284), .A2(n287), .ZN(\ab[14][0] ) );
  NOR2_X1 U728 ( .A1(n276), .A2(n288), .ZN(\ab[13][9] ) );
  NOR2_X1 U729 ( .A1(n277), .A2(n288), .ZN(\ab[13][8] ) );
  NOR2_X1 U730 ( .A1(n278), .A2(n288), .ZN(\ab[13][7] ) );
  NOR2_X1 U731 ( .A1(n279), .A2(n288), .ZN(\ab[13][6] ) );
  NOR2_X1 U732 ( .A1(n280), .A2(n288), .ZN(\ab[13][5] ) );
  NOR2_X1 U733 ( .A1(n281), .A2(n288), .ZN(\ab[13][4] ) );
  NOR2_X1 U734 ( .A1(n282), .A2(n288), .ZN(\ab[13][3] ) );
  NOR2_X1 U735 ( .A1(n283), .A2(n288), .ZN(\ab[13][2] ) );
  NOR2_X1 U736 ( .A1(n262), .A2(n288), .ZN(\ab[13][1] ) );
  NOR2_X1 U737 ( .A1(n269), .A2(n288), .ZN(\SUMB[13][16] ) );
  NOR2_X1 U738 ( .A1(n270), .A2(n288), .ZN(\ab[13][15] ) );
  NOR2_X1 U739 ( .A1(n271), .A2(n288), .ZN(\ab[13][14] ) );
  NOR2_X1 U740 ( .A1(n272), .A2(n288), .ZN(\ab[13][13] ) );
  NOR2_X1 U741 ( .A1(n273), .A2(n288), .ZN(\ab[13][12] ) );
  NOR2_X1 U742 ( .A1(n274), .A2(n288), .ZN(\ab[13][11] ) );
  NOR2_X1 U743 ( .A1(n275), .A2(n288), .ZN(\ab[13][10] ) );
  NOR2_X1 U744 ( .A1(n284), .A2(n288), .ZN(\ab[13][0] ) );
  NOR2_X1 U745 ( .A1(n276), .A2(n289), .ZN(\ab[12][9] ) );
  NOR2_X1 U746 ( .A1(n277), .A2(n289), .ZN(\ab[12][8] ) );
  NOR2_X1 U747 ( .A1(n278), .A2(n289), .ZN(\ab[12][7] ) );
  NOR2_X1 U748 ( .A1(n279), .A2(n289), .ZN(\ab[12][6] ) );
  NOR2_X1 U749 ( .A1(n280), .A2(n289), .ZN(\ab[12][5] ) );
  NOR2_X1 U750 ( .A1(n281), .A2(n289), .ZN(\ab[12][4] ) );
  NOR2_X1 U751 ( .A1(n282), .A2(n289), .ZN(\ab[12][3] ) );
  NOR2_X1 U752 ( .A1(n283), .A2(n289), .ZN(\ab[12][2] ) );
  NOR2_X1 U753 ( .A1(n262), .A2(n289), .ZN(\ab[12][1] ) );
  NOR2_X1 U754 ( .A1(n269), .A2(n289), .ZN(\SUMB[12][16] ) );
  NOR2_X1 U755 ( .A1(n270), .A2(n289), .ZN(\ab[12][15] ) );
  NOR2_X1 U756 ( .A1(n271), .A2(n289), .ZN(\ab[12][14] ) );
  NOR2_X1 U757 ( .A1(n272), .A2(n289), .ZN(\ab[12][13] ) );
  NOR2_X1 U758 ( .A1(n273), .A2(n289), .ZN(\ab[12][12] ) );
  NOR2_X1 U759 ( .A1(n274), .A2(n289), .ZN(\ab[12][11] ) );
  NOR2_X1 U760 ( .A1(n275), .A2(n289), .ZN(\ab[12][10] ) );
  NOR2_X1 U761 ( .A1(n284), .A2(n289), .ZN(\ab[12][0] ) );
  NOR2_X1 U762 ( .A1(n276), .A2(n290), .ZN(\ab[11][9] ) );
  NOR2_X1 U763 ( .A1(n277), .A2(n290), .ZN(\ab[11][8] ) );
  NOR2_X1 U764 ( .A1(n278), .A2(n290), .ZN(\ab[11][7] ) );
  NOR2_X1 U765 ( .A1(n279), .A2(n290), .ZN(\ab[11][6] ) );
  NOR2_X1 U766 ( .A1(n280), .A2(n290), .ZN(\ab[11][5] ) );
  NOR2_X1 U767 ( .A1(n281), .A2(n290), .ZN(\ab[11][4] ) );
  NOR2_X1 U768 ( .A1(n282), .A2(n290), .ZN(\ab[11][3] ) );
  NOR2_X1 U769 ( .A1(n283), .A2(n290), .ZN(\ab[11][2] ) );
  NOR2_X1 U770 ( .A1(n262), .A2(n290), .ZN(\ab[11][1] ) );
  NOR2_X1 U771 ( .A1(n269), .A2(n290), .ZN(\SUMB[11][16] ) );
  NOR2_X1 U772 ( .A1(n270), .A2(n290), .ZN(\ab[11][15] ) );
  NOR2_X1 U773 ( .A1(n271), .A2(n290), .ZN(\ab[11][14] ) );
  NOR2_X1 U774 ( .A1(n272), .A2(n290), .ZN(\ab[11][13] ) );
  NOR2_X1 U775 ( .A1(n273), .A2(n290), .ZN(\ab[11][12] ) );
  NOR2_X1 U776 ( .A1(n274), .A2(n290), .ZN(\ab[11][11] ) );
  NOR2_X1 U777 ( .A1(n275), .A2(n290), .ZN(\ab[11][10] ) );
  NOR2_X1 U778 ( .A1(n284), .A2(n290), .ZN(\ab[11][0] ) );
  NOR2_X1 U779 ( .A1(n276), .A2(n291), .ZN(\ab[10][9] ) );
  NOR2_X1 U780 ( .A1(n277), .A2(n291), .ZN(\ab[10][8] ) );
  NOR2_X1 U781 ( .A1(n278), .A2(n291), .ZN(\ab[10][7] ) );
  NOR2_X1 U782 ( .A1(n279), .A2(n291), .ZN(\ab[10][6] ) );
  NOR2_X1 U783 ( .A1(n280), .A2(n291), .ZN(\ab[10][5] ) );
  NOR2_X1 U784 ( .A1(n281), .A2(n291), .ZN(\ab[10][4] ) );
  NOR2_X1 U785 ( .A1(n282), .A2(n291), .ZN(\ab[10][3] ) );
  NOR2_X1 U786 ( .A1(n283), .A2(n291), .ZN(\ab[10][2] ) );
  NOR2_X1 U787 ( .A1(n262), .A2(n291), .ZN(\ab[10][1] ) );
  NOR2_X1 U788 ( .A1(n269), .A2(n291), .ZN(\SUMB[10][16] ) );
  NOR2_X1 U789 ( .A1(n270), .A2(n291), .ZN(\ab[10][15] ) );
  NOR2_X1 U790 ( .A1(n271), .A2(n291), .ZN(\ab[10][14] ) );
  NOR2_X1 U791 ( .A1(n272), .A2(n291), .ZN(\ab[10][13] ) );
  NOR2_X1 U792 ( .A1(n273), .A2(n291), .ZN(\ab[10][12] ) );
  NOR2_X1 U793 ( .A1(n274), .A2(n291), .ZN(\ab[10][11] ) );
  NOR2_X1 U794 ( .A1(n275), .A2(n291), .ZN(\ab[10][10] ) );
  NOR2_X1 U795 ( .A1(n284), .A2(n291), .ZN(\ab[10][0] ) );
  NOR2_X1 U796 ( .A1(n276), .A2(n300), .ZN(\ab[0][9] ) );
  NOR2_X1 U797 ( .A1(n277), .A2(n300), .ZN(\ab[0][8] ) );
  NOR2_X1 U798 ( .A1(n278), .A2(n300), .ZN(\ab[0][7] ) );
  NOR2_X1 U799 ( .A1(n279), .A2(n300), .ZN(\ab[0][6] ) );
  NOR2_X1 U800 ( .A1(n280), .A2(n300), .ZN(\ab[0][5] ) );
  NOR2_X1 U801 ( .A1(n281), .A2(n300), .ZN(\ab[0][4] ) );
  NOR2_X1 U802 ( .A1(n260), .A2(n300), .ZN(\ab[0][3] ) );
  NOR2_X1 U803 ( .A1(n261), .A2(n268), .ZN(\ab[0][2] ) );
  NOR2_X1 U804 ( .A1(n262), .A2(n268), .ZN(\ab[0][1] ) );
  NOR2_X1 U805 ( .A1(n269), .A2(n268), .ZN(\ab[0][16] ) );
  NOR2_X1 U806 ( .A1(n270), .A2(n268), .ZN(\ab[0][15] ) );
  NOR2_X1 U807 ( .A1(n271), .A2(n268), .ZN(\ab[0][14] ) );
  NOR2_X1 U808 ( .A1(n272), .A2(n268), .ZN(\ab[0][13] ) );
  NOR2_X1 U809 ( .A1(n273), .A2(n268), .ZN(\ab[0][12] ) );
  NOR2_X1 U810 ( .A1(n274), .A2(n268), .ZN(\ab[0][11] ) );
  NOR2_X1 U811 ( .A1(n275), .A2(n268), .ZN(\ab[0][10] ) );
  NOR2_X1 U812 ( .A1(n263), .A2(n268), .ZN(PRODUCT[0]) );
endmodule


module multiplier_DW01_add_2 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70;

  OR2_X4 U2 ( .A1(B[15]), .A2(A[15]), .ZN(n1) );
  AND2_X4 U3 ( .A1(n1), .A2(n70), .ZN(SUM[15]) );
  INV_X4 U4 ( .A(B[29]), .ZN(n3) );
  INV_X4 U5 ( .A(n21), .ZN(n4) );
  INV_X4 U6 ( .A(n23), .ZN(n5) );
  INV_X4 U7 ( .A(n29), .ZN(n6) );
  INV_X4 U8 ( .A(n31), .ZN(n7) );
  INV_X4 U9 ( .A(n37), .ZN(n8) );
  INV_X4 U10 ( .A(n39), .ZN(n9) );
  INV_X4 U11 ( .A(n45), .ZN(n10) );
  INV_X4 U12 ( .A(n47), .ZN(n11) );
  INV_X4 U13 ( .A(n53), .ZN(n12) );
  INV_X4 U14 ( .A(n55), .ZN(n13) );
  INV_X4 U15 ( .A(n61), .ZN(n14) );
  INV_X4 U16 ( .A(n63), .ZN(n15) );
  INV_X4 U17 ( .A(n68), .ZN(n16) );
  INV_X4 U18 ( .A(n70), .ZN(n17) );
  XOR2_X1 U19 ( .A(n3), .B(n18), .Z(SUM[29]) );
  AOI21_X1 U20 ( .B1(n19), .B2(n4), .A(n20), .ZN(n18) );
  XOR2_X1 U21 ( .A(n19), .B(n22), .Z(SUM[28]) );
  NOR2_X1 U22 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U23 ( .A1(B[28]), .A2(A[28]), .ZN(n21) );
  AND2_X1 U24 ( .A1(B[28]), .A2(A[28]), .ZN(n20) );
  OAI21_X1 U25 ( .B1(n23), .B2(n24), .A(n25), .ZN(n19) );
  XOR2_X1 U26 ( .A(n26), .B(n24), .Z(SUM[27]) );
  AOI21_X1 U27 ( .B1(n6), .B2(n27), .A(n28), .ZN(n24) );
  NAND2_X1 U28 ( .A1(n5), .A2(n25), .ZN(n26) );
  NAND2_X1 U29 ( .A1(B[27]), .A2(A[27]), .ZN(n25) );
  NOR2_X1 U30 ( .A1(B[27]), .A2(A[27]), .ZN(n23) );
  XOR2_X1 U31 ( .A(n27), .B(n30), .Z(SUM[26]) );
  NOR2_X1 U32 ( .A1(n28), .A2(n29), .ZN(n30) );
  NOR2_X1 U33 ( .A1(B[26]), .A2(A[26]), .ZN(n29) );
  AND2_X1 U34 ( .A1(B[26]), .A2(A[26]), .ZN(n28) );
  OAI21_X1 U35 ( .B1(n31), .B2(n32), .A(n33), .ZN(n27) );
  XOR2_X1 U36 ( .A(n34), .B(n32), .Z(SUM[25]) );
  AOI21_X1 U37 ( .B1(n8), .B2(n35), .A(n36), .ZN(n32) );
  NAND2_X1 U38 ( .A1(n7), .A2(n33), .ZN(n34) );
  NAND2_X1 U39 ( .A1(B[25]), .A2(A[25]), .ZN(n33) );
  NOR2_X1 U40 ( .A1(B[25]), .A2(A[25]), .ZN(n31) );
  XOR2_X1 U41 ( .A(n35), .B(n38), .Z(SUM[24]) );
  NOR2_X1 U42 ( .A1(n36), .A2(n37), .ZN(n38) );
  NOR2_X1 U43 ( .A1(B[24]), .A2(A[24]), .ZN(n37) );
  AND2_X1 U44 ( .A1(B[24]), .A2(A[24]), .ZN(n36) );
  OAI21_X1 U45 ( .B1(n39), .B2(n40), .A(n41), .ZN(n35) );
  XOR2_X1 U46 ( .A(n42), .B(n40), .Z(SUM[23]) );
  AOI21_X1 U47 ( .B1(n10), .B2(n43), .A(n44), .ZN(n40) );
  NAND2_X1 U48 ( .A1(n9), .A2(n41), .ZN(n42) );
  NAND2_X1 U49 ( .A1(B[23]), .A2(A[23]), .ZN(n41) );
  NOR2_X1 U50 ( .A1(B[23]), .A2(A[23]), .ZN(n39) );
  XOR2_X1 U51 ( .A(n43), .B(n46), .Z(SUM[22]) );
  NOR2_X1 U52 ( .A1(n44), .A2(n45), .ZN(n46) );
  NOR2_X1 U53 ( .A1(B[22]), .A2(A[22]), .ZN(n45) );
  AND2_X1 U54 ( .A1(B[22]), .A2(A[22]), .ZN(n44) );
  OAI21_X1 U55 ( .B1(n47), .B2(n48), .A(n49), .ZN(n43) );
  XOR2_X1 U56 ( .A(n50), .B(n48), .Z(SUM[21]) );
  AOI21_X1 U57 ( .B1(n12), .B2(n51), .A(n52), .ZN(n48) );
  NAND2_X1 U58 ( .A1(n11), .A2(n49), .ZN(n50) );
  NAND2_X1 U59 ( .A1(B[21]), .A2(A[21]), .ZN(n49) );
  NOR2_X1 U60 ( .A1(B[21]), .A2(A[21]), .ZN(n47) );
  XOR2_X1 U61 ( .A(n51), .B(n54), .Z(SUM[20]) );
  NOR2_X1 U62 ( .A1(n52), .A2(n53), .ZN(n54) );
  NOR2_X1 U63 ( .A1(B[20]), .A2(A[20]), .ZN(n53) );
  AND2_X1 U64 ( .A1(B[20]), .A2(A[20]), .ZN(n52) );
  OAI21_X1 U65 ( .B1(n55), .B2(n56), .A(n57), .ZN(n51) );
  XOR2_X1 U66 ( .A(n58), .B(n56), .Z(SUM[19]) );
  AOI21_X1 U67 ( .B1(n14), .B2(n59), .A(n60), .ZN(n56) );
  NAND2_X1 U68 ( .A1(n13), .A2(n57), .ZN(n58) );
  NAND2_X1 U69 ( .A1(B[19]), .A2(A[19]), .ZN(n57) );
  NOR2_X1 U70 ( .A1(B[19]), .A2(A[19]), .ZN(n55) );
  XOR2_X1 U71 ( .A(n59), .B(n62), .Z(SUM[18]) );
  NOR2_X1 U72 ( .A1(n60), .A2(n61), .ZN(n62) );
  NOR2_X1 U73 ( .A1(B[18]), .A2(A[18]), .ZN(n61) );
  AND2_X1 U74 ( .A1(B[18]), .A2(A[18]), .ZN(n60) );
  OAI21_X1 U75 ( .B1(n63), .B2(n64), .A(n65), .ZN(n59) );
  XOR2_X1 U76 ( .A(n66), .B(n64), .Z(SUM[17]) );
  AOI21_X1 U77 ( .B1(n16), .B2(n17), .A(n67), .ZN(n64) );
  NAND2_X1 U78 ( .A1(n15), .A2(n65), .ZN(n66) );
  NAND2_X1 U79 ( .A1(B[17]), .A2(A[17]), .ZN(n65) );
  NOR2_X1 U80 ( .A1(B[17]), .A2(A[17]), .ZN(n63) );
  XOR2_X1 U81 ( .A(n17), .B(n69), .Z(SUM[16]) );
  NOR2_X1 U82 ( .A1(n67), .A2(n68), .ZN(n69) );
  NOR2_X1 U83 ( .A1(B[16]), .A2(A[16]), .ZN(n68) );
  AND2_X1 U84 ( .A1(B[16]), .A2(A[16]), .ZN(n67) );
  NAND2_X1 U85 ( .A1(B[15]), .A2(A[15]), .ZN(n70) );
  BUF_X32 U86 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X32 U87 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X32 U88 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X32 U89 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X32 U90 ( .A(A[4]), .Z(SUM[4]) );
  BUF_X32 U91 ( .A(A[5]), .Z(SUM[5]) );
  BUF_X32 U92 ( .A(A[6]), .Z(SUM[6]) );
  BUF_X32 U93 ( .A(A[7]), .Z(SUM[7]) );
  BUF_X32 U94 ( .A(A[8]), .Z(SUM[8]) );
  BUF_X32 U95 ( .A(A[9]), .Z(SUM[9]) );
  BUF_X32 U96 ( .A(A[10]), .Z(SUM[10]) );
  BUF_X32 U97 ( .A(A[11]), .Z(SUM[11]) );
  BUF_X32 U98 ( .A(A[12]), .Z(SUM[12]) );
  BUF_X32 U99 ( .A(A[13]), .Z(SUM[13]) );
  BUF_X32 U100 ( .A(A[14]), .Z(SUM[14]) );
endmodule


module multiplier_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [15:0] A;
  input [15:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] ,
         \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] ,
         \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] ,
         \ab[15][0] , \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] ,
         \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] ,
         \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][15] , \ab[13][14] , \ab[13][13] ,
         \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] ,
         \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] ,
         \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][15] , \ab[12][14] ,
         \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] ,
         \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] ,
         \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][15] ,
         \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] ,
         \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] ,
         \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] ,
         \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] ,
         \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][15] , \ab[8][14] , \ab[8][13] ,
         \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][15] , \ab[7][14] ,
         \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] , \ab[7][9] ,
         \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] ,
         \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][15] ,
         \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] ,
         \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] ,
         \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][15] , \ab[3][14] , \ab[3][13] ,
         \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][15] , \ab[2][14] ,
         \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] , \ab[2][9] ,
         \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] ,
         \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][15] ,
         \ab[1][14] , \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] ,
         \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] ,
         \ab[0][15] , \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] ,
         \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] ,
         \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] ,
         \CARRYB[15][14] , \CARRYB[15][13] , \CARRYB[15][12] ,
         \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] ,
         \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] ,
         \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] ,
         \CARRYB[14][14] , \CARRYB[14][13] , \CARRYB[14][12] ,
         \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] ,
         \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] ,
         \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][14] , \CARRYB[12][13] , \CARRYB[12][12] ,
         \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] ,
         \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] ,
         \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] ,
         \CARRYB[11][14] , \CARRYB[11][13] , \CARRYB[11][12] ,
         \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] ,
         \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] ,
         \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] ,
         \CARRYB[10][14] , \CARRYB[10][13] , \CARRYB[10][12] ,
         \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] ,
         \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] ,
         \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] ,
         \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] ,
         \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] ,
         \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][14] ,
         \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] ,
         \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] ,
         \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] ,
         \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] ,
         \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] ,
         \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] ,
         \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] ,
         \CARRYB[5][14] , \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] ,
         \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] ,
         \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] ,
         \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][14] ,
         \CARRYB[4][13] , \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] ,
         \CARRYB[4][9] , \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] ,
         \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] ,
         \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][14] , \CARRYB[3][13] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] ,
         \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] ,
         \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] ,
         \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[15][0] , \SUMB[14][14] ,
         \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] ,
         \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] ,
         \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] ,
         \SUMB[14][1] , \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] ,
         \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] ,
         \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] ,
         \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] ,
         \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] ,
         \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] ,
         \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][14] , \SUMB[8][13] ,
         \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] ,
         \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] ,
         \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \A1[12] ,
         \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] ,
         \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] , n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94;

  FA_X1 S4_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), .CO(
        \CARRYB[15][0] ), .S(\SUMB[15][0] ) );
  FA_X1 S4_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), .CO(
        \CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA_X1 S4_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), .CO(
        \CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA_X1 S4_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), .CO(
        \CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA_X1 S4_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), .CO(
        \CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA_X1 S4_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), .CO(
        \CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA_X1 S4_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), .CO(
        \CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA_X1 S4_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), .CO(
        \CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA_X1 S4_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), .CO(
        \CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA_X1 S4_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), .CO(
        \CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA_X1 S4_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA_X1 S4_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA_X1 S4_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA_X1 S4_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA_X1 S5_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\ab[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA_X1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FA_X1 S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA_X1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA_X1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA_X1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA_X1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA_X1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA_X1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA_X1 S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA_X1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA_X1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA_X1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA_X1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA_X1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA_X1 S3_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\ab[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA_X1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA_X1 S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA_X1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA_X1 S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA_X1 S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA_X1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA_X1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA_X1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA_X1 S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA_X1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA_X1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA_X1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA_X1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA_X1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA_X1 S3_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\ab[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA_X1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA_X1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA_X1 S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA_X1 S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA_X1 S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA_X1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA_X1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA_X1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA_X1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA_X1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA_X1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA_X1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA_X1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA_X1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA_X1 S3_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\ab[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA_X1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA_X1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA_X1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA_X1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA_X1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA_X1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA_X1 S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA_X1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA_X1 S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA_X1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA_X1 S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA_X1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA_X1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA_X1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA_X1 S3_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\ab[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA_X1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA_X1 S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA_X1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA_X1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA_X1 S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA_X1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA_X1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA_X1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA_X1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA_X1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA_X1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA_X1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA_X1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA_X1 S3_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\ab[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA_X1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA_X1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA_X1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA_X1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA_X1 S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA_X1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA_X1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA_X1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA_X1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA_X1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA_X1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA_X1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA_X1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA_X1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA_X1 S3_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\ab[8][15] ), .CO(
        \CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA_X1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA_X1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA_X1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA_X1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA_X1 S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA_X1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA_X1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA_X1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA_X1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA_X1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA_X1 S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA_X1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA_X1 S3_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\ab[7][15] ), .CO(
        \CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA_X1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA_X1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA_X1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA_X1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA_X1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA_X1 S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA_X1 S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA_X1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA_X1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA_X1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA_X1 S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA_X1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA_X1 S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA_X1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA_X1 S3_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\ab[6][15] ), .CO(
        \CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA_X1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA_X1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA_X1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA_X1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA_X1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA_X1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA_X1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA_X1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA_X1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA_X1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA_X1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA_X1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA_X1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA_X1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA_X1 S3_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\ab[5][15] ), .CO(
        \CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA_X1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA_X1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA_X1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA_X1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA_X1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA_X1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA_X1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA_X1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA_X1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA_X1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA_X1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA_X1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA_X1 S3_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\ab[4][15] ), .CO(
        \CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA_X1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA_X1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA_X1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA_X1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA_X1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA_X1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA_X1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA_X1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA_X1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA_X1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA_X1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA_X1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA_X1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA_X1 S3_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\ab[3][15] ), .CO(
        \CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA_X1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA_X1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA_X1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA_X1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA_X1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA_X1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA_X1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA_X1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA_X1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA_X1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA_X1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA_X1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA_X1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA_X1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA_X1 S3_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\ab[2][15] ), .CO(
        \CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(n16), .CI(n45), .CO(\CARRYB[2][0] ), .S(
        \A1[0] ) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(n15), .CI(n44), .CO(\CARRYB[2][1] ), .S(
        \SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(n14), .CI(n43), .CO(\CARRYB[2][2] ), .S(
        \SUMB[2][2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2][3] ), .B(n13), .CI(n42), .CO(\CARRYB[2][3] ), .S(
        \SUMB[2][3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2][4] ), .B(n12), .CI(n41), .CO(\CARRYB[2][4] ), .S(
        \SUMB[2][4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2][5] ), .B(n11), .CI(n40), .CO(\CARRYB[2][5] ), .S(
        \SUMB[2][5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2][6] ), .B(n10), .CI(n39), .CO(\CARRYB[2][6] ), .S(
        \SUMB[2][6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(n9), .CI(n38), .CO(\CARRYB[2][7] ), .S(
        \SUMB[2][7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(n8), .CI(n37), .CO(\CARRYB[2][8] ), .S(
        \SUMB[2][8] ) );
  FA_X1 S2_2_9 ( .A(\ab[2][9] ), .B(n7), .CI(n36), .CO(\CARRYB[2][9] ), .S(
        \SUMB[2][9] ) );
  FA_X1 S2_2_10 ( .A(\ab[2][10] ), .B(n6), .CI(n35), .CO(\CARRYB[2][10] ), .S(
        \SUMB[2][10] ) );
  FA_X1 S2_2_11 ( .A(\ab[2][11] ), .B(n5), .CI(n34), .CO(\CARRYB[2][11] ), .S(
        \SUMB[2][11] ) );
  FA_X1 S2_2_12 ( .A(\ab[2][12] ), .B(n4), .CI(n33), .CO(\CARRYB[2][12] ), .S(
        \SUMB[2][12] ) );
  FA_X1 S2_2_13 ( .A(\ab[2][13] ), .B(n3), .CI(n32), .CO(\CARRYB[2][13] ), .S(
        \SUMB[2][13] ) );
  FA_X1 S3_2_14 ( .A(\ab[2][14] ), .B(n31), .CI(\ab[1][15] ), .CO(
        \CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  INV_X4 U2 ( .A(B[4]), .ZN(n90) );
  INV_X4 U3 ( .A(B[5]), .ZN(n89) );
  INV_X4 U4 ( .A(B[6]), .ZN(n88) );
  INV_X4 U5 ( .A(B[7]), .ZN(n87) );
  INV_X4 U6 ( .A(B[8]), .ZN(n86) );
  INV_X4 U7 ( .A(B[9]), .ZN(n85) );
  INV_X4 U8 ( .A(B[10]), .ZN(n84) );
  INV_X4 U9 ( .A(B[11]), .ZN(n83) );
  INV_X4 U10 ( .A(B[12]), .ZN(n82) );
  INV_X4 U11 ( .A(B[13]), .ZN(n81) );
  INV_X4 U12 ( .A(B[3]), .ZN(n91) );
  INV_X4 U13 ( .A(B[2]), .ZN(n92) );
  INV_X4 U14 ( .A(A[1]), .ZN(n77) );
  INV_X4 U15 ( .A(B[1]), .ZN(n93) );
  INV_X4 U16 ( .A(B[14]), .ZN(n80) );
  INV_X4 U17 ( .A(B[15]), .ZN(n79) );
  INV_X4 U18 ( .A(A[0]), .ZN(n78) );
  INV_X4 U19 ( .A(A[2]), .ZN(n76) );
  INV_X4 U20 ( .A(A[3]), .ZN(n75) );
  INV_X4 U21 ( .A(A[4]), .ZN(n74) );
  INV_X4 U22 ( .A(A[5]), .ZN(n73) );
  INV_X4 U23 ( .A(A[6]), .ZN(n72) );
  INV_X4 U24 ( .A(A[7]), .ZN(n71) );
  INV_X4 U25 ( .A(A[8]), .ZN(n70) );
  INV_X4 U26 ( .A(A[9]), .ZN(n69) );
  INV_X4 U27 ( .A(A[10]), .ZN(n68) );
  INV_X4 U28 ( .A(A[11]), .ZN(n67) );
  INV_X4 U29 ( .A(A[12]), .ZN(n66) );
  INV_X4 U30 ( .A(A[13]), .ZN(n65) );
  INV_X4 U31 ( .A(A[14]), .ZN(n64) );
  INV_X4 U32 ( .A(A[15]), .ZN(n63) );
  INV_X4 U33 ( .A(B[0]), .ZN(n94) );
  AND2_X4 U34 ( .A1(\ab[0][14] ), .A2(\ab[1][13] ), .ZN(n3) );
  AND2_X4 U35 ( .A1(\ab[0][13] ), .A2(\ab[1][12] ), .ZN(n4) );
  AND2_X4 U36 ( .A1(\ab[0][12] ), .A2(\ab[1][11] ), .ZN(n5) );
  AND2_X4 U37 ( .A1(\ab[0][11] ), .A2(\ab[1][10] ), .ZN(n6) );
  AND2_X4 U38 ( .A1(\ab[0][10] ), .A2(\ab[1][9] ), .ZN(n7) );
  AND2_X4 U39 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .ZN(n8) );
  AND2_X4 U40 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .ZN(n9) );
  AND2_X4 U41 ( .A1(\ab[0][7] ), .A2(\ab[1][6] ), .ZN(n10) );
  AND2_X4 U42 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .ZN(n11) );
  AND2_X4 U43 ( .A1(\ab[0][5] ), .A2(\ab[1][4] ), .ZN(n12) );
  AND2_X4 U44 ( .A1(\ab[0][4] ), .A2(\ab[1][3] ), .ZN(n13) );
  AND2_X4 U45 ( .A1(\ab[0][3] ), .A2(\ab[1][2] ), .ZN(n14) );
  AND2_X4 U46 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .ZN(n15) );
  AND2_X4 U47 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .ZN(n16) );
  XOR2_X2 U48 ( .A(\CARRYB[15][14] ), .B(\ab[15][15] ), .Z(n17) );
  XOR2_X2 U49 ( .A(\CARRYB[15][12] ), .B(\SUMB[15][13] ), .Z(n18) );
  XOR2_X2 U50 ( .A(\CARRYB[15][10] ), .B(\SUMB[15][11] ), .Z(n19) );
  XOR2_X2 U51 ( .A(\CARRYB[15][8] ), .B(\SUMB[15][9] ), .Z(n20) );
  XOR2_X2 U52 ( .A(\CARRYB[15][6] ), .B(\SUMB[15][7] ), .Z(n21) );
  XOR2_X2 U53 ( .A(\CARRYB[15][4] ), .B(\SUMB[15][5] ), .Z(n22) );
  XOR2_X2 U54 ( .A(\CARRYB[15][2] ), .B(\SUMB[15][3] ), .Z(n23) );
  XOR2_X2 U55 ( .A(\CARRYB[15][1] ), .B(\SUMB[15][2] ), .Z(n24) );
  XOR2_X2 U56 ( .A(\CARRYB[15][13] ), .B(\SUMB[15][14] ), .Z(n25) );
  XOR2_X2 U57 ( .A(\CARRYB[15][11] ), .B(\SUMB[15][12] ), .Z(n26) );
  XOR2_X2 U58 ( .A(\CARRYB[15][9] ), .B(\SUMB[15][10] ), .Z(n27) );
  XOR2_X2 U59 ( .A(\CARRYB[15][7] ), .B(\SUMB[15][8] ), .Z(n28) );
  XOR2_X2 U60 ( .A(\CARRYB[15][5] ), .B(\SUMB[15][6] ), .Z(n29) );
  XOR2_X2 U61 ( .A(\CARRYB[15][3] ), .B(\SUMB[15][4] ), .Z(n30) );
  AND2_X4 U62 ( .A1(\ab[0][15] ), .A2(\ab[1][14] ), .ZN(n31) );
  XOR2_X2 U63 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(n32) );
  XOR2_X2 U64 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(n33) );
  XOR2_X2 U65 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(n34) );
  XOR2_X2 U66 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(n35) );
  XOR2_X2 U67 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(n36) );
  XOR2_X2 U68 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(n37) );
  XOR2_X2 U69 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(n38) );
  XOR2_X2 U70 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(n39) );
  XOR2_X2 U71 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(n40) );
  XOR2_X2 U72 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(n41) );
  XOR2_X2 U73 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(n42) );
  XOR2_X2 U74 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(n43) );
  XOR2_X2 U75 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(n44) );
  XOR2_X2 U76 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(n45) );
  XOR2_X2 U77 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  AND2_X4 U78 ( .A1(\CARRYB[15][13] ), .A2(\SUMB[15][14] ), .ZN(n47) );
  AND2_X4 U79 ( .A1(\CARRYB[15][11] ), .A2(\SUMB[15][12] ), .ZN(n48) );
  AND2_X4 U80 ( .A1(\CARRYB[15][9] ), .A2(\SUMB[15][10] ), .ZN(n49) );
  AND2_X4 U81 ( .A1(\CARRYB[15][7] ), .A2(\SUMB[15][8] ), .ZN(n50) );
  AND2_X4 U82 ( .A1(\CARRYB[15][5] ), .A2(\SUMB[15][6] ), .ZN(n51) );
  AND2_X4 U83 ( .A1(\CARRYB[15][3] ), .A2(\SUMB[15][4] ), .ZN(n52) );
  AND2_X4 U84 ( .A1(\CARRYB[15][1] ), .A2(\SUMB[15][2] ), .ZN(n53) );
  AND2_X4 U85 ( .A1(\CARRYB[15][12] ), .A2(\SUMB[15][13] ), .ZN(n54) );
  AND2_X4 U86 ( .A1(\CARRYB[15][10] ), .A2(\SUMB[15][11] ), .ZN(n55) );
  AND2_X4 U87 ( .A1(\CARRYB[15][8] ), .A2(\SUMB[15][9] ), .ZN(n56) );
  AND2_X4 U88 ( .A1(\CARRYB[15][6] ), .A2(\SUMB[15][7] ), .ZN(n57) );
  AND2_X4 U89 ( .A1(\CARRYB[15][4] ), .A2(\SUMB[15][5] ), .ZN(n58) );
  AND2_X4 U90 ( .A1(\CARRYB[15][2] ), .A2(\SUMB[15][3] ), .ZN(n59) );
  AND2_X4 U91 ( .A1(\CARRYB[15][0] ), .A2(\SUMB[15][1] ), .ZN(n60) );
  XOR2_X2 U92 ( .A(\CARRYB[15][0] ), .B(\SUMB[15][1] ), .Z(n61) );
  AND2_X4 U93 ( .A1(\CARRYB[15][14] ), .A2(\ab[15][15] ), .ZN(n62) );
  NOR2_X1 U95 ( .A1(n69), .A2(n85), .ZN(\ab[9][9] ) );
  NOR2_X1 U96 ( .A1(n69), .A2(n86), .ZN(\ab[9][8] ) );
  NOR2_X1 U97 ( .A1(n69), .A2(n87), .ZN(\ab[9][7] ) );
  NOR2_X1 U98 ( .A1(n69), .A2(n88), .ZN(\ab[9][6] ) );
  NOR2_X1 U99 ( .A1(n69), .A2(n89), .ZN(\ab[9][5] ) );
  NOR2_X1 U100 ( .A1(n69), .A2(n90), .ZN(\ab[9][4] ) );
  NOR2_X1 U101 ( .A1(n69), .A2(n91), .ZN(\ab[9][3] ) );
  NOR2_X1 U102 ( .A1(n69), .A2(n92), .ZN(\ab[9][2] ) );
  NOR2_X1 U103 ( .A1(n69), .A2(n93), .ZN(\ab[9][1] ) );
  NOR2_X1 U104 ( .A1(n69), .A2(n79), .ZN(\ab[9][15] ) );
  NOR2_X1 U105 ( .A1(n69), .A2(n80), .ZN(\ab[9][14] ) );
  NOR2_X1 U106 ( .A1(n69), .A2(n81), .ZN(\ab[9][13] ) );
  NOR2_X1 U107 ( .A1(n69), .A2(n82), .ZN(\ab[9][12] ) );
  NOR2_X1 U108 ( .A1(n69), .A2(n83), .ZN(\ab[9][11] ) );
  NOR2_X1 U109 ( .A1(n69), .A2(n84), .ZN(\ab[9][10] ) );
  NOR2_X1 U110 ( .A1(n69), .A2(n94), .ZN(\ab[9][0] ) );
  NOR2_X1 U111 ( .A1(n85), .A2(n70), .ZN(\ab[8][9] ) );
  NOR2_X1 U112 ( .A1(n86), .A2(n70), .ZN(\ab[8][8] ) );
  NOR2_X1 U113 ( .A1(n87), .A2(n70), .ZN(\ab[8][7] ) );
  NOR2_X1 U114 ( .A1(n88), .A2(n70), .ZN(\ab[8][6] ) );
  NOR2_X1 U115 ( .A1(n89), .A2(n70), .ZN(\ab[8][5] ) );
  NOR2_X1 U116 ( .A1(n90), .A2(n70), .ZN(\ab[8][4] ) );
  NOR2_X1 U117 ( .A1(n91), .A2(n70), .ZN(\ab[8][3] ) );
  NOR2_X1 U118 ( .A1(n92), .A2(n70), .ZN(\ab[8][2] ) );
  NOR2_X1 U119 ( .A1(n93), .A2(n70), .ZN(\ab[8][1] ) );
  NOR2_X1 U120 ( .A1(n79), .A2(n70), .ZN(\ab[8][15] ) );
  NOR2_X1 U121 ( .A1(n80), .A2(n70), .ZN(\ab[8][14] ) );
  NOR2_X1 U122 ( .A1(n81), .A2(n70), .ZN(\ab[8][13] ) );
  NOR2_X1 U123 ( .A1(n82), .A2(n70), .ZN(\ab[8][12] ) );
  NOR2_X1 U124 ( .A1(n83), .A2(n70), .ZN(\ab[8][11] ) );
  NOR2_X1 U125 ( .A1(n84), .A2(n70), .ZN(\ab[8][10] ) );
  NOR2_X1 U126 ( .A1(n94), .A2(n70), .ZN(\ab[8][0] ) );
  NOR2_X1 U127 ( .A1(n85), .A2(n71), .ZN(\ab[7][9] ) );
  NOR2_X1 U128 ( .A1(n86), .A2(n71), .ZN(\ab[7][8] ) );
  NOR2_X1 U129 ( .A1(n87), .A2(n71), .ZN(\ab[7][7] ) );
  NOR2_X1 U130 ( .A1(n88), .A2(n71), .ZN(\ab[7][6] ) );
  NOR2_X1 U131 ( .A1(n89), .A2(n71), .ZN(\ab[7][5] ) );
  NOR2_X1 U132 ( .A1(n90), .A2(n71), .ZN(\ab[7][4] ) );
  NOR2_X1 U133 ( .A1(n91), .A2(n71), .ZN(\ab[7][3] ) );
  NOR2_X1 U134 ( .A1(n92), .A2(n71), .ZN(\ab[7][2] ) );
  NOR2_X1 U135 ( .A1(n93), .A2(n71), .ZN(\ab[7][1] ) );
  NOR2_X1 U136 ( .A1(n79), .A2(n71), .ZN(\ab[7][15] ) );
  NOR2_X1 U137 ( .A1(n80), .A2(n71), .ZN(\ab[7][14] ) );
  NOR2_X1 U138 ( .A1(n81), .A2(n71), .ZN(\ab[7][13] ) );
  NOR2_X1 U139 ( .A1(n82), .A2(n71), .ZN(\ab[7][12] ) );
  NOR2_X1 U140 ( .A1(n83), .A2(n71), .ZN(\ab[7][11] ) );
  NOR2_X1 U141 ( .A1(n84), .A2(n71), .ZN(\ab[7][10] ) );
  NOR2_X1 U142 ( .A1(n94), .A2(n71), .ZN(\ab[7][0] ) );
  NOR2_X1 U143 ( .A1(n85), .A2(n72), .ZN(\ab[6][9] ) );
  NOR2_X1 U144 ( .A1(n86), .A2(n72), .ZN(\ab[6][8] ) );
  NOR2_X1 U145 ( .A1(n87), .A2(n72), .ZN(\ab[6][7] ) );
  NOR2_X1 U146 ( .A1(n88), .A2(n72), .ZN(\ab[6][6] ) );
  NOR2_X1 U147 ( .A1(n89), .A2(n72), .ZN(\ab[6][5] ) );
  NOR2_X1 U148 ( .A1(n90), .A2(n72), .ZN(\ab[6][4] ) );
  NOR2_X1 U149 ( .A1(n91), .A2(n72), .ZN(\ab[6][3] ) );
  NOR2_X1 U150 ( .A1(n92), .A2(n72), .ZN(\ab[6][2] ) );
  NOR2_X1 U151 ( .A1(n93), .A2(n72), .ZN(\ab[6][1] ) );
  NOR2_X1 U152 ( .A1(n79), .A2(n72), .ZN(\ab[6][15] ) );
  NOR2_X1 U153 ( .A1(n80), .A2(n72), .ZN(\ab[6][14] ) );
  NOR2_X1 U154 ( .A1(n81), .A2(n72), .ZN(\ab[6][13] ) );
  NOR2_X1 U155 ( .A1(n82), .A2(n72), .ZN(\ab[6][12] ) );
  NOR2_X1 U156 ( .A1(n83), .A2(n72), .ZN(\ab[6][11] ) );
  NOR2_X1 U157 ( .A1(n84), .A2(n72), .ZN(\ab[6][10] ) );
  NOR2_X1 U158 ( .A1(n94), .A2(n72), .ZN(\ab[6][0] ) );
  NOR2_X1 U159 ( .A1(n85), .A2(n73), .ZN(\ab[5][9] ) );
  NOR2_X1 U160 ( .A1(n86), .A2(n73), .ZN(\ab[5][8] ) );
  NOR2_X1 U161 ( .A1(n87), .A2(n73), .ZN(\ab[5][7] ) );
  NOR2_X1 U162 ( .A1(n88), .A2(n73), .ZN(\ab[5][6] ) );
  NOR2_X1 U163 ( .A1(n89), .A2(n73), .ZN(\ab[5][5] ) );
  NOR2_X1 U164 ( .A1(n90), .A2(n73), .ZN(\ab[5][4] ) );
  NOR2_X1 U165 ( .A1(n91), .A2(n73), .ZN(\ab[5][3] ) );
  NOR2_X1 U166 ( .A1(n92), .A2(n73), .ZN(\ab[5][2] ) );
  NOR2_X1 U167 ( .A1(n93), .A2(n73), .ZN(\ab[5][1] ) );
  NOR2_X1 U168 ( .A1(n79), .A2(n73), .ZN(\ab[5][15] ) );
  NOR2_X1 U169 ( .A1(n80), .A2(n73), .ZN(\ab[5][14] ) );
  NOR2_X1 U170 ( .A1(n81), .A2(n73), .ZN(\ab[5][13] ) );
  NOR2_X1 U171 ( .A1(n82), .A2(n73), .ZN(\ab[5][12] ) );
  NOR2_X1 U172 ( .A1(n83), .A2(n73), .ZN(\ab[5][11] ) );
  NOR2_X1 U173 ( .A1(n84), .A2(n73), .ZN(\ab[5][10] ) );
  NOR2_X1 U174 ( .A1(n94), .A2(n73), .ZN(\ab[5][0] ) );
  NOR2_X1 U175 ( .A1(n85), .A2(n74), .ZN(\ab[4][9] ) );
  NOR2_X1 U176 ( .A1(n86), .A2(n74), .ZN(\ab[4][8] ) );
  NOR2_X1 U177 ( .A1(n87), .A2(n74), .ZN(\ab[4][7] ) );
  NOR2_X1 U178 ( .A1(n88), .A2(n74), .ZN(\ab[4][6] ) );
  NOR2_X1 U179 ( .A1(n89), .A2(n74), .ZN(\ab[4][5] ) );
  NOR2_X1 U180 ( .A1(n90), .A2(n74), .ZN(\ab[4][4] ) );
  NOR2_X1 U181 ( .A1(n91), .A2(n74), .ZN(\ab[4][3] ) );
  NOR2_X1 U182 ( .A1(n92), .A2(n74), .ZN(\ab[4][2] ) );
  NOR2_X1 U183 ( .A1(n93), .A2(n74), .ZN(\ab[4][1] ) );
  NOR2_X1 U184 ( .A1(n79), .A2(n74), .ZN(\ab[4][15] ) );
  NOR2_X1 U185 ( .A1(n80), .A2(n74), .ZN(\ab[4][14] ) );
  NOR2_X1 U186 ( .A1(n81), .A2(n74), .ZN(\ab[4][13] ) );
  NOR2_X1 U187 ( .A1(n82), .A2(n74), .ZN(\ab[4][12] ) );
  NOR2_X1 U188 ( .A1(n83), .A2(n74), .ZN(\ab[4][11] ) );
  NOR2_X1 U189 ( .A1(n84), .A2(n74), .ZN(\ab[4][10] ) );
  NOR2_X1 U190 ( .A1(n94), .A2(n74), .ZN(\ab[4][0] ) );
  NOR2_X1 U191 ( .A1(n85), .A2(n75), .ZN(\ab[3][9] ) );
  NOR2_X1 U192 ( .A1(n86), .A2(n75), .ZN(\ab[3][8] ) );
  NOR2_X1 U193 ( .A1(n87), .A2(n75), .ZN(\ab[3][7] ) );
  NOR2_X1 U194 ( .A1(n88), .A2(n75), .ZN(\ab[3][6] ) );
  NOR2_X1 U195 ( .A1(n89), .A2(n75), .ZN(\ab[3][5] ) );
  NOR2_X1 U196 ( .A1(n90), .A2(n75), .ZN(\ab[3][4] ) );
  NOR2_X1 U197 ( .A1(n91), .A2(n75), .ZN(\ab[3][3] ) );
  NOR2_X1 U198 ( .A1(n92), .A2(n75), .ZN(\ab[3][2] ) );
  NOR2_X1 U199 ( .A1(n93), .A2(n75), .ZN(\ab[3][1] ) );
  NOR2_X1 U200 ( .A1(n79), .A2(n75), .ZN(\ab[3][15] ) );
  NOR2_X1 U201 ( .A1(n80), .A2(n75), .ZN(\ab[3][14] ) );
  NOR2_X1 U202 ( .A1(n81), .A2(n75), .ZN(\ab[3][13] ) );
  NOR2_X1 U203 ( .A1(n82), .A2(n75), .ZN(\ab[3][12] ) );
  NOR2_X1 U204 ( .A1(n83), .A2(n75), .ZN(\ab[3][11] ) );
  NOR2_X1 U205 ( .A1(n84), .A2(n75), .ZN(\ab[3][10] ) );
  NOR2_X1 U206 ( .A1(n94), .A2(n75), .ZN(\ab[3][0] ) );
  NOR2_X1 U207 ( .A1(n85), .A2(n76), .ZN(\ab[2][9] ) );
  NOR2_X1 U208 ( .A1(n86), .A2(n76), .ZN(\ab[2][8] ) );
  NOR2_X1 U209 ( .A1(n87), .A2(n76), .ZN(\ab[2][7] ) );
  NOR2_X1 U210 ( .A1(n88), .A2(n76), .ZN(\ab[2][6] ) );
  NOR2_X1 U211 ( .A1(n89), .A2(n76), .ZN(\ab[2][5] ) );
  NOR2_X1 U212 ( .A1(n90), .A2(n76), .ZN(\ab[2][4] ) );
  NOR2_X1 U213 ( .A1(n91), .A2(n76), .ZN(\ab[2][3] ) );
  NOR2_X1 U214 ( .A1(n92), .A2(n76), .ZN(\ab[2][2] ) );
  NOR2_X1 U215 ( .A1(n93), .A2(n76), .ZN(\ab[2][1] ) );
  NOR2_X1 U216 ( .A1(n79), .A2(n76), .ZN(\ab[2][15] ) );
  NOR2_X1 U217 ( .A1(n80), .A2(n76), .ZN(\ab[2][14] ) );
  NOR2_X1 U218 ( .A1(n81), .A2(n76), .ZN(\ab[2][13] ) );
  NOR2_X1 U219 ( .A1(n82), .A2(n76), .ZN(\ab[2][12] ) );
  NOR2_X1 U220 ( .A1(n83), .A2(n76), .ZN(\ab[2][11] ) );
  NOR2_X1 U221 ( .A1(n84), .A2(n76), .ZN(\ab[2][10] ) );
  NOR2_X1 U222 ( .A1(n94), .A2(n76), .ZN(\ab[2][0] ) );
  NOR2_X1 U223 ( .A1(n85), .A2(n77), .ZN(\ab[1][9] ) );
  NOR2_X1 U224 ( .A1(n86), .A2(n77), .ZN(\ab[1][8] ) );
  NOR2_X1 U225 ( .A1(n87), .A2(n77), .ZN(\ab[1][7] ) );
  NOR2_X1 U226 ( .A1(n88), .A2(n77), .ZN(\ab[1][6] ) );
  NOR2_X1 U227 ( .A1(n89), .A2(n77), .ZN(\ab[1][5] ) );
  NOR2_X1 U228 ( .A1(n90), .A2(n77), .ZN(\ab[1][4] ) );
  NOR2_X1 U229 ( .A1(n91), .A2(n77), .ZN(\ab[1][3] ) );
  NOR2_X1 U230 ( .A1(n92), .A2(n77), .ZN(\ab[1][2] ) );
  NOR2_X1 U231 ( .A1(n93), .A2(n77), .ZN(\ab[1][1] ) );
  NOR2_X1 U232 ( .A1(n79), .A2(n77), .ZN(\ab[1][15] ) );
  NOR2_X1 U233 ( .A1(n80), .A2(n77), .ZN(\ab[1][14] ) );
  NOR2_X1 U234 ( .A1(n81), .A2(n77), .ZN(\ab[1][13] ) );
  NOR2_X1 U235 ( .A1(n82), .A2(n77), .ZN(\ab[1][12] ) );
  NOR2_X1 U236 ( .A1(n83), .A2(n77), .ZN(\ab[1][11] ) );
  NOR2_X1 U237 ( .A1(n84), .A2(n77), .ZN(\ab[1][10] ) );
  NOR2_X1 U238 ( .A1(n94), .A2(n77), .ZN(\ab[1][0] ) );
  NOR2_X1 U239 ( .A1(n85), .A2(n63), .ZN(\ab[15][9] ) );
  NOR2_X1 U240 ( .A1(n86), .A2(n63), .ZN(\ab[15][8] ) );
  NOR2_X1 U241 ( .A1(n87), .A2(n63), .ZN(\ab[15][7] ) );
  NOR2_X1 U242 ( .A1(n88), .A2(n63), .ZN(\ab[15][6] ) );
  NOR2_X1 U243 ( .A1(n89), .A2(n63), .ZN(\ab[15][5] ) );
  NOR2_X1 U244 ( .A1(n90), .A2(n63), .ZN(\ab[15][4] ) );
  NOR2_X1 U245 ( .A1(n91), .A2(n63), .ZN(\ab[15][3] ) );
  NOR2_X1 U246 ( .A1(n92), .A2(n63), .ZN(\ab[15][2] ) );
  NOR2_X1 U247 ( .A1(n93), .A2(n63), .ZN(\ab[15][1] ) );
  NOR2_X1 U248 ( .A1(n79), .A2(n63), .ZN(\ab[15][15] ) );
  NOR2_X1 U249 ( .A1(n80), .A2(n63), .ZN(\ab[15][14] ) );
  NOR2_X1 U250 ( .A1(n81), .A2(n63), .ZN(\ab[15][13] ) );
  NOR2_X1 U251 ( .A1(n82), .A2(n63), .ZN(\ab[15][12] ) );
  NOR2_X1 U252 ( .A1(n83), .A2(n63), .ZN(\ab[15][11] ) );
  NOR2_X1 U253 ( .A1(n84), .A2(n63), .ZN(\ab[15][10] ) );
  NOR2_X1 U254 ( .A1(n94), .A2(n63), .ZN(\ab[15][0] ) );
  NOR2_X1 U255 ( .A1(n85), .A2(n64), .ZN(\ab[14][9] ) );
  NOR2_X1 U256 ( .A1(n86), .A2(n64), .ZN(\ab[14][8] ) );
  NOR2_X1 U257 ( .A1(n87), .A2(n64), .ZN(\ab[14][7] ) );
  NOR2_X1 U258 ( .A1(n88), .A2(n64), .ZN(\ab[14][6] ) );
  NOR2_X1 U259 ( .A1(n89), .A2(n64), .ZN(\ab[14][5] ) );
  NOR2_X1 U260 ( .A1(n90), .A2(n64), .ZN(\ab[14][4] ) );
  NOR2_X1 U261 ( .A1(n91), .A2(n64), .ZN(\ab[14][3] ) );
  NOR2_X1 U262 ( .A1(n92), .A2(n64), .ZN(\ab[14][2] ) );
  NOR2_X1 U263 ( .A1(n93), .A2(n64), .ZN(\ab[14][1] ) );
  NOR2_X1 U264 ( .A1(n79), .A2(n64), .ZN(\ab[14][15] ) );
  NOR2_X1 U265 ( .A1(n80), .A2(n64), .ZN(\ab[14][14] ) );
  NOR2_X1 U266 ( .A1(n81), .A2(n64), .ZN(\ab[14][13] ) );
  NOR2_X1 U267 ( .A1(n82), .A2(n64), .ZN(\ab[14][12] ) );
  NOR2_X1 U268 ( .A1(n83), .A2(n64), .ZN(\ab[14][11] ) );
  NOR2_X1 U269 ( .A1(n84), .A2(n64), .ZN(\ab[14][10] ) );
  NOR2_X1 U270 ( .A1(n94), .A2(n64), .ZN(\ab[14][0] ) );
  NOR2_X1 U271 ( .A1(n85), .A2(n65), .ZN(\ab[13][9] ) );
  NOR2_X1 U272 ( .A1(n86), .A2(n65), .ZN(\ab[13][8] ) );
  NOR2_X1 U273 ( .A1(n87), .A2(n65), .ZN(\ab[13][7] ) );
  NOR2_X1 U274 ( .A1(n88), .A2(n65), .ZN(\ab[13][6] ) );
  NOR2_X1 U275 ( .A1(n89), .A2(n65), .ZN(\ab[13][5] ) );
  NOR2_X1 U276 ( .A1(n90), .A2(n65), .ZN(\ab[13][4] ) );
  NOR2_X1 U277 ( .A1(n91), .A2(n65), .ZN(\ab[13][3] ) );
  NOR2_X1 U278 ( .A1(n92), .A2(n65), .ZN(\ab[13][2] ) );
  NOR2_X1 U279 ( .A1(n93), .A2(n65), .ZN(\ab[13][1] ) );
  NOR2_X1 U280 ( .A1(n79), .A2(n65), .ZN(\ab[13][15] ) );
  NOR2_X1 U281 ( .A1(n80), .A2(n65), .ZN(\ab[13][14] ) );
  NOR2_X1 U282 ( .A1(n81), .A2(n65), .ZN(\ab[13][13] ) );
  NOR2_X1 U283 ( .A1(n82), .A2(n65), .ZN(\ab[13][12] ) );
  NOR2_X1 U284 ( .A1(n83), .A2(n65), .ZN(\ab[13][11] ) );
  NOR2_X1 U285 ( .A1(n84), .A2(n65), .ZN(\ab[13][10] ) );
  NOR2_X1 U286 ( .A1(n94), .A2(n65), .ZN(\ab[13][0] ) );
  NOR2_X1 U287 ( .A1(n85), .A2(n66), .ZN(\ab[12][9] ) );
  NOR2_X1 U288 ( .A1(n86), .A2(n66), .ZN(\ab[12][8] ) );
  NOR2_X1 U289 ( .A1(n87), .A2(n66), .ZN(\ab[12][7] ) );
  NOR2_X1 U290 ( .A1(n88), .A2(n66), .ZN(\ab[12][6] ) );
  NOR2_X1 U291 ( .A1(n89), .A2(n66), .ZN(\ab[12][5] ) );
  NOR2_X1 U292 ( .A1(n90), .A2(n66), .ZN(\ab[12][4] ) );
  NOR2_X1 U293 ( .A1(n91), .A2(n66), .ZN(\ab[12][3] ) );
  NOR2_X1 U294 ( .A1(n92), .A2(n66), .ZN(\ab[12][2] ) );
  NOR2_X1 U295 ( .A1(n93), .A2(n66), .ZN(\ab[12][1] ) );
  NOR2_X1 U296 ( .A1(n79), .A2(n66), .ZN(\ab[12][15] ) );
  NOR2_X1 U297 ( .A1(n80), .A2(n66), .ZN(\ab[12][14] ) );
  NOR2_X1 U298 ( .A1(n81), .A2(n66), .ZN(\ab[12][13] ) );
  NOR2_X1 U299 ( .A1(n82), .A2(n66), .ZN(\ab[12][12] ) );
  NOR2_X1 U300 ( .A1(n83), .A2(n66), .ZN(\ab[12][11] ) );
  NOR2_X1 U301 ( .A1(n84), .A2(n66), .ZN(\ab[12][10] ) );
  NOR2_X1 U302 ( .A1(n94), .A2(n66), .ZN(\ab[12][0] ) );
  NOR2_X1 U303 ( .A1(n85), .A2(n67), .ZN(\ab[11][9] ) );
  NOR2_X1 U304 ( .A1(n86), .A2(n67), .ZN(\ab[11][8] ) );
  NOR2_X1 U305 ( .A1(n87), .A2(n67), .ZN(\ab[11][7] ) );
  NOR2_X1 U306 ( .A1(n88), .A2(n67), .ZN(\ab[11][6] ) );
  NOR2_X1 U307 ( .A1(n89), .A2(n67), .ZN(\ab[11][5] ) );
  NOR2_X1 U308 ( .A1(n90), .A2(n67), .ZN(\ab[11][4] ) );
  NOR2_X1 U309 ( .A1(n91), .A2(n67), .ZN(\ab[11][3] ) );
  NOR2_X1 U310 ( .A1(n92), .A2(n67), .ZN(\ab[11][2] ) );
  NOR2_X1 U311 ( .A1(n93), .A2(n67), .ZN(\ab[11][1] ) );
  NOR2_X1 U312 ( .A1(n79), .A2(n67), .ZN(\ab[11][15] ) );
  NOR2_X1 U313 ( .A1(n80), .A2(n67), .ZN(\ab[11][14] ) );
  NOR2_X1 U314 ( .A1(n81), .A2(n67), .ZN(\ab[11][13] ) );
  NOR2_X1 U315 ( .A1(n82), .A2(n67), .ZN(\ab[11][12] ) );
  NOR2_X1 U316 ( .A1(n83), .A2(n67), .ZN(\ab[11][11] ) );
  NOR2_X1 U317 ( .A1(n84), .A2(n67), .ZN(\ab[11][10] ) );
  NOR2_X1 U318 ( .A1(n94), .A2(n67), .ZN(\ab[11][0] ) );
  NOR2_X1 U319 ( .A1(n85), .A2(n68), .ZN(\ab[10][9] ) );
  NOR2_X1 U320 ( .A1(n86), .A2(n68), .ZN(\ab[10][8] ) );
  NOR2_X1 U321 ( .A1(n87), .A2(n68), .ZN(\ab[10][7] ) );
  NOR2_X1 U322 ( .A1(n88), .A2(n68), .ZN(\ab[10][6] ) );
  NOR2_X1 U323 ( .A1(n89), .A2(n68), .ZN(\ab[10][5] ) );
  NOR2_X1 U324 ( .A1(n90), .A2(n68), .ZN(\ab[10][4] ) );
  NOR2_X1 U325 ( .A1(n91), .A2(n68), .ZN(\ab[10][3] ) );
  NOR2_X1 U326 ( .A1(n92), .A2(n68), .ZN(\ab[10][2] ) );
  NOR2_X1 U327 ( .A1(n93), .A2(n68), .ZN(\ab[10][1] ) );
  NOR2_X1 U328 ( .A1(n79), .A2(n68), .ZN(\ab[10][15] ) );
  NOR2_X1 U329 ( .A1(n80), .A2(n68), .ZN(\ab[10][14] ) );
  NOR2_X1 U330 ( .A1(n81), .A2(n68), .ZN(\ab[10][13] ) );
  NOR2_X1 U331 ( .A1(n82), .A2(n68), .ZN(\ab[10][12] ) );
  NOR2_X1 U332 ( .A1(n83), .A2(n68), .ZN(\ab[10][11] ) );
  NOR2_X1 U333 ( .A1(n84), .A2(n68), .ZN(\ab[10][10] ) );
  NOR2_X1 U334 ( .A1(n94), .A2(n68), .ZN(\ab[10][0] ) );
  NOR2_X1 U335 ( .A1(n85), .A2(n78), .ZN(\ab[0][9] ) );
  NOR2_X1 U336 ( .A1(n86), .A2(n78), .ZN(\ab[0][8] ) );
  NOR2_X1 U337 ( .A1(n87), .A2(n78), .ZN(\ab[0][7] ) );
  NOR2_X1 U338 ( .A1(n88), .A2(n78), .ZN(\ab[0][6] ) );
  NOR2_X1 U339 ( .A1(n89), .A2(n78), .ZN(\ab[0][5] ) );
  NOR2_X1 U340 ( .A1(n90), .A2(n78), .ZN(\ab[0][4] ) );
  NOR2_X1 U341 ( .A1(n91), .A2(n78), .ZN(\ab[0][3] ) );
  NOR2_X1 U342 ( .A1(n92), .A2(n78), .ZN(\ab[0][2] ) );
  NOR2_X1 U343 ( .A1(n93), .A2(n78), .ZN(\ab[0][1] ) );
  NOR2_X1 U344 ( .A1(n79), .A2(n78), .ZN(\ab[0][15] ) );
  NOR2_X1 U345 ( .A1(n80), .A2(n78), .ZN(\ab[0][14] ) );
  NOR2_X1 U346 ( .A1(n81), .A2(n78), .ZN(\ab[0][13] ) );
  NOR2_X1 U347 ( .A1(n82), .A2(n78), .ZN(\ab[0][12] ) );
  NOR2_X1 U348 ( .A1(n83), .A2(n78), .ZN(\ab[0][11] ) );
  NOR2_X1 U349 ( .A1(n84), .A2(n78), .ZN(\ab[0][10] ) );
  NOR2_X1 U350 ( .A1(n94), .A2(n78), .ZN(PRODUCT[0]) );
  multiplier_DW01_add_2 FS_1 ( .A({1'b0, n17, n25, n18, n26, n19, n27, n20, 
        n28, n21, n29, n22, n30, n23, n24, n61, \SUMB[15][0] , \A1[12] , 
        \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , 
        \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({n62, n47, n54, n48, 
        n55, n49, n56, n50, n57, n51, n58, n52, n59, n53, n60, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .CI(1'b0), .SUM(PRODUCT[31:2]) );
endmodule


module multiplier_DW01_add_3 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70;

  OR2_X4 U2 ( .A1(B[15]), .A2(A[15]), .ZN(n1) );
  AND2_X4 U3 ( .A1(n1), .A2(n70), .ZN(SUM[15]) );
  INV_X4 U4 ( .A(B[29]), .ZN(n3) );
  INV_X4 U5 ( .A(n21), .ZN(n4) );
  INV_X4 U6 ( .A(n23), .ZN(n5) );
  INV_X4 U7 ( .A(n29), .ZN(n6) );
  INV_X4 U8 ( .A(n31), .ZN(n7) );
  INV_X4 U9 ( .A(n37), .ZN(n8) );
  INV_X4 U10 ( .A(n39), .ZN(n9) );
  INV_X4 U11 ( .A(n45), .ZN(n10) );
  INV_X4 U12 ( .A(n47), .ZN(n11) );
  INV_X4 U13 ( .A(n53), .ZN(n12) );
  INV_X4 U14 ( .A(n55), .ZN(n13) );
  INV_X4 U15 ( .A(n61), .ZN(n14) );
  INV_X4 U16 ( .A(n63), .ZN(n15) );
  INV_X4 U17 ( .A(n68), .ZN(n16) );
  INV_X4 U18 ( .A(n70), .ZN(n17) );
  XOR2_X1 U19 ( .A(n3), .B(n18), .Z(SUM[29]) );
  AOI21_X1 U20 ( .B1(n19), .B2(n4), .A(n20), .ZN(n18) );
  XOR2_X1 U21 ( .A(n19), .B(n22), .Z(SUM[28]) );
  NOR2_X1 U22 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U23 ( .A1(B[28]), .A2(A[28]), .ZN(n21) );
  AND2_X1 U24 ( .A1(B[28]), .A2(A[28]), .ZN(n20) );
  OAI21_X1 U25 ( .B1(n23), .B2(n24), .A(n25), .ZN(n19) );
  XOR2_X1 U26 ( .A(n26), .B(n24), .Z(SUM[27]) );
  AOI21_X1 U27 ( .B1(n6), .B2(n27), .A(n28), .ZN(n24) );
  NAND2_X1 U28 ( .A1(n5), .A2(n25), .ZN(n26) );
  NAND2_X1 U29 ( .A1(B[27]), .A2(A[27]), .ZN(n25) );
  NOR2_X1 U30 ( .A1(B[27]), .A2(A[27]), .ZN(n23) );
  XOR2_X1 U31 ( .A(n27), .B(n30), .Z(SUM[26]) );
  NOR2_X1 U32 ( .A1(n28), .A2(n29), .ZN(n30) );
  NOR2_X1 U33 ( .A1(B[26]), .A2(A[26]), .ZN(n29) );
  AND2_X1 U34 ( .A1(B[26]), .A2(A[26]), .ZN(n28) );
  OAI21_X1 U35 ( .B1(n31), .B2(n32), .A(n33), .ZN(n27) );
  XOR2_X1 U36 ( .A(n34), .B(n32), .Z(SUM[25]) );
  AOI21_X1 U37 ( .B1(n8), .B2(n35), .A(n36), .ZN(n32) );
  NAND2_X1 U38 ( .A1(n7), .A2(n33), .ZN(n34) );
  NAND2_X1 U39 ( .A1(B[25]), .A2(A[25]), .ZN(n33) );
  NOR2_X1 U40 ( .A1(B[25]), .A2(A[25]), .ZN(n31) );
  XOR2_X1 U41 ( .A(n35), .B(n38), .Z(SUM[24]) );
  NOR2_X1 U42 ( .A1(n36), .A2(n37), .ZN(n38) );
  NOR2_X1 U43 ( .A1(B[24]), .A2(A[24]), .ZN(n37) );
  AND2_X1 U44 ( .A1(B[24]), .A2(A[24]), .ZN(n36) );
  OAI21_X1 U45 ( .B1(n39), .B2(n40), .A(n41), .ZN(n35) );
  XOR2_X1 U46 ( .A(n42), .B(n40), .Z(SUM[23]) );
  AOI21_X1 U47 ( .B1(n10), .B2(n43), .A(n44), .ZN(n40) );
  NAND2_X1 U48 ( .A1(n9), .A2(n41), .ZN(n42) );
  NAND2_X1 U49 ( .A1(B[23]), .A2(A[23]), .ZN(n41) );
  NOR2_X1 U50 ( .A1(B[23]), .A2(A[23]), .ZN(n39) );
  XOR2_X1 U51 ( .A(n43), .B(n46), .Z(SUM[22]) );
  NOR2_X1 U52 ( .A1(n44), .A2(n45), .ZN(n46) );
  NOR2_X1 U53 ( .A1(B[22]), .A2(A[22]), .ZN(n45) );
  AND2_X1 U54 ( .A1(B[22]), .A2(A[22]), .ZN(n44) );
  OAI21_X1 U55 ( .B1(n47), .B2(n48), .A(n49), .ZN(n43) );
  XOR2_X1 U56 ( .A(n50), .B(n48), .Z(SUM[21]) );
  AOI21_X1 U57 ( .B1(n12), .B2(n51), .A(n52), .ZN(n48) );
  NAND2_X1 U58 ( .A1(n11), .A2(n49), .ZN(n50) );
  NAND2_X1 U59 ( .A1(B[21]), .A2(A[21]), .ZN(n49) );
  NOR2_X1 U60 ( .A1(B[21]), .A2(A[21]), .ZN(n47) );
  XOR2_X1 U61 ( .A(n51), .B(n54), .Z(SUM[20]) );
  NOR2_X1 U62 ( .A1(n52), .A2(n53), .ZN(n54) );
  NOR2_X1 U63 ( .A1(B[20]), .A2(A[20]), .ZN(n53) );
  AND2_X1 U64 ( .A1(B[20]), .A2(A[20]), .ZN(n52) );
  OAI21_X1 U65 ( .B1(n55), .B2(n56), .A(n57), .ZN(n51) );
  XOR2_X1 U66 ( .A(n58), .B(n56), .Z(SUM[19]) );
  AOI21_X1 U67 ( .B1(n14), .B2(n59), .A(n60), .ZN(n56) );
  NAND2_X1 U68 ( .A1(n13), .A2(n57), .ZN(n58) );
  NAND2_X1 U69 ( .A1(B[19]), .A2(A[19]), .ZN(n57) );
  NOR2_X1 U70 ( .A1(B[19]), .A2(A[19]), .ZN(n55) );
  XOR2_X1 U71 ( .A(n59), .B(n62), .Z(SUM[18]) );
  NOR2_X1 U72 ( .A1(n60), .A2(n61), .ZN(n62) );
  NOR2_X1 U73 ( .A1(B[18]), .A2(A[18]), .ZN(n61) );
  AND2_X1 U74 ( .A1(B[18]), .A2(A[18]), .ZN(n60) );
  OAI21_X1 U75 ( .B1(n63), .B2(n64), .A(n65), .ZN(n59) );
  XOR2_X1 U76 ( .A(n66), .B(n64), .Z(SUM[17]) );
  AOI21_X1 U77 ( .B1(n16), .B2(n17), .A(n67), .ZN(n64) );
  NAND2_X1 U78 ( .A1(n15), .A2(n65), .ZN(n66) );
  NAND2_X1 U79 ( .A1(B[17]), .A2(A[17]), .ZN(n65) );
  NOR2_X1 U80 ( .A1(B[17]), .A2(A[17]), .ZN(n63) );
  XOR2_X1 U81 ( .A(n17), .B(n69), .Z(SUM[16]) );
  NOR2_X1 U82 ( .A1(n67), .A2(n68), .ZN(n69) );
  NOR2_X1 U83 ( .A1(B[16]), .A2(A[16]), .ZN(n68) );
  AND2_X1 U84 ( .A1(B[16]), .A2(A[16]), .ZN(n67) );
  NAND2_X1 U85 ( .A1(B[15]), .A2(A[15]), .ZN(n70) );
  BUF_X32 U86 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X32 U87 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X32 U88 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X32 U89 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X32 U90 ( .A(A[4]), .Z(SUM[4]) );
  BUF_X32 U91 ( .A(A[5]), .Z(SUM[5]) );
  BUF_X32 U92 ( .A(A[6]), .Z(SUM[6]) );
  BUF_X32 U93 ( .A(A[7]), .Z(SUM[7]) );
  BUF_X32 U94 ( .A(A[8]), .Z(SUM[8]) );
  BUF_X32 U95 ( .A(A[9]), .Z(SUM[9]) );
  BUF_X32 U96 ( .A(A[10]), .Z(SUM[10]) );
  BUF_X32 U97 ( .A(A[11]), .Z(SUM[11]) );
  BUF_X32 U98 ( .A(A[12]), .Z(SUM[12]) );
  BUF_X32 U99 ( .A(A[13]), .Z(SUM[13]) );
  BUF_X32 U100 ( .A(A[14]), .Z(SUM[14]) );
endmodule


module multiplier_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [15:0] A;
  input [15:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] ,
         \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] ,
         \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] ,
         \ab[15][0] , \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] ,
         \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] ,
         \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][15] , \ab[13][14] , \ab[13][13] ,
         \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] ,
         \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] ,
         \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][15] , \ab[12][14] ,
         \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] ,
         \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] ,
         \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][15] ,
         \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] ,
         \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] ,
         \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] ,
         \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] ,
         \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][15] , \ab[8][14] , \ab[8][13] ,
         \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][15] , \ab[7][14] ,
         \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] , \ab[7][9] ,
         \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] ,
         \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][15] ,
         \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] ,
         \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] ,
         \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][15] , \ab[3][14] , \ab[3][13] ,
         \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][15] , \ab[2][14] ,
         \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] , \ab[2][9] ,
         \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] ,
         \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][15] ,
         \ab[1][14] , \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] ,
         \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] ,
         \ab[0][15] , \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] ,
         \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] ,
         \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] ,
         \CARRYB[15][14] , \CARRYB[15][13] , \CARRYB[15][12] ,
         \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] ,
         \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] ,
         \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] ,
         \CARRYB[14][14] , \CARRYB[14][13] , \CARRYB[14][12] ,
         \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] ,
         \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] ,
         \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][14] , \CARRYB[12][13] , \CARRYB[12][12] ,
         \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] ,
         \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] ,
         \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] ,
         \CARRYB[11][14] , \CARRYB[11][13] , \CARRYB[11][12] ,
         \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] ,
         \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] ,
         \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] ,
         \CARRYB[10][14] , \CARRYB[10][13] , \CARRYB[10][12] ,
         \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] ,
         \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] ,
         \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] ,
         \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] ,
         \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] ,
         \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][14] ,
         \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] ,
         \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] ,
         \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] ,
         \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] ,
         \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] ,
         \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] ,
         \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] ,
         \CARRYB[5][14] , \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] ,
         \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] ,
         \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] ,
         \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][14] ,
         \CARRYB[4][13] , \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] ,
         \CARRYB[4][9] , \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] ,
         \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] ,
         \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][14] , \CARRYB[3][13] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] ,
         \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] ,
         \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] ,
         \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[15][0] , \SUMB[14][14] ,
         \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] ,
         \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] ,
         \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] ,
         \SUMB[14][1] , \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] ,
         \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] ,
         \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] ,
         \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] ,
         \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] ,
         \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] ,
         \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][14] , \SUMB[8][13] ,
         \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] ,
         \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] ,
         \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \A1[12] ,
         \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] ,
         \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] , n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94;

  FA_X1 S4_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), .CO(
        \CARRYB[15][0] ), .S(\SUMB[15][0] ) );
  FA_X1 S4_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), .CO(
        \CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA_X1 S4_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), .CO(
        \CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA_X1 S4_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), .CO(
        \CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA_X1 S4_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), .CO(
        \CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA_X1 S4_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), .CO(
        \CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA_X1 S4_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), .CO(
        \CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA_X1 S4_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), .CO(
        \CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA_X1 S4_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), .CO(
        \CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA_X1 S4_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), .CO(
        \CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA_X1 S4_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA_X1 S4_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA_X1 S4_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA_X1 S4_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA_X1 S5_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\ab[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA_X1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FA_X1 S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA_X1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA_X1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA_X1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA_X1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA_X1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA_X1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA_X1 S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA_X1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA_X1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA_X1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA_X1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA_X1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA_X1 S3_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\ab[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA_X1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA_X1 S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA_X1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA_X1 S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA_X1 S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA_X1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA_X1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA_X1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA_X1 S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA_X1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA_X1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA_X1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA_X1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA_X1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA_X1 S3_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\ab[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA_X1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA_X1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA_X1 S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA_X1 S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA_X1 S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA_X1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA_X1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA_X1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA_X1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA_X1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA_X1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA_X1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA_X1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA_X1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA_X1 S3_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\ab[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA_X1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA_X1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA_X1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA_X1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA_X1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA_X1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA_X1 S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA_X1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA_X1 S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA_X1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA_X1 S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA_X1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA_X1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA_X1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA_X1 S3_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\ab[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA_X1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA_X1 S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA_X1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA_X1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA_X1 S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA_X1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA_X1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA_X1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA_X1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA_X1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA_X1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA_X1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA_X1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA_X1 S3_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\ab[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA_X1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA_X1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA_X1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA_X1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA_X1 S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA_X1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA_X1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA_X1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA_X1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA_X1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA_X1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA_X1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA_X1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA_X1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA_X1 S3_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\ab[8][15] ), .CO(
        \CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA_X1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA_X1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA_X1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA_X1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA_X1 S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA_X1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA_X1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA_X1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA_X1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA_X1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA_X1 S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA_X1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA_X1 S3_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\ab[7][15] ), .CO(
        \CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA_X1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA_X1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA_X1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA_X1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA_X1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA_X1 S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA_X1 S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA_X1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA_X1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA_X1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA_X1 S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA_X1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA_X1 S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA_X1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA_X1 S3_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\ab[6][15] ), .CO(
        \CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA_X1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA_X1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA_X1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA_X1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA_X1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA_X1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA_X1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA_X1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA_X1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA_X1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA_X1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA_X1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA_X1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA_X1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA_X1 S3_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\ab[5][15] ), .CO(
        \CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA_X1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA_X1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA_X1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA_X1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA_X1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA_X1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA_X1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA_X1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA_X1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA_X1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA_X1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA_X1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA_X1 S3_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\ab[4][15] ), .CO(
        \CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA_X1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA_X1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA_X1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA_X1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA_X1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA_X1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA_X1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA_X1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA_X1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA_X1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA_X1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA_X1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA_X1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA_X1 S3_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\ab[3][15] ), .CO(
        \CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA_X1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA_X1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA_X1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA_X1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA_X1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA_X1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA_X1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA_X1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA_X1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA_X1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA_X1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA_X1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA_X1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA_X1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA_X1 S3_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\ab[2][15] ), .CO(
        \CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(n16), .CI(n45), .CO(\CARRYB[2][0] ), .S(
        \A1[0] ) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(n15), .CI(n44), .CO(\CARRYB[2][1] ), .S(
        \SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(n14), .CI(n43), .CO(\CARRYB[2][2] ), .S(
        \SUMB[2][2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2][3] ), .B(n13), .CI(n42), .CO(\CARRYB[2][3] ), .S(
        \SUMB[2][3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2][4] ), .B(n12), .CI(n41), .CO(\CARRYB[2][4] ), .S(
        \SUMB[2][4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2][5] ), .B(n11), .CI(n40), .CO(\CARRYB[2][5] ), .S(
        \SUMB[2][5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2][6] ), .B(n10), .CI(n39), .CO(\CARRYB[2][6] ), .S(
        \SUMB[2][6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(n9), .CI(n38), .CO(\CARRYB[2][7] ), .S(
        \SUMB[2][7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(n8), .CI(n37), .CO(\CARRYB[2][8] ), .S(
        \SUMB[2][8] ) );
  FA_X1 S2_2_9 ( .A(\ab[2][9] ), .B(n7), .CI(n36), .CO(\CARRYB[2][9] ), .S(
        \SUMB[2][9] ) );
  FA_X1 S2_2_10 ( .A(\ab[2][10] ), .B(n6), .CI(n35), .CO(\CARRYB[2][10] ), .S(
        \SUMB[2][10] ) );
  FA_X1 S2_2_11 ( .A(\ab[2][11] ), .B(n5), .CI(n34), .CO(\CARRYB[2][11] ), .S(
        \SUMB[2][11] ) );
  FA_X1 S2_2_12 ( .A(\ab[2][12] ), .B(n4), .CI(n33), .CO(\CARRYB[2][12] ), .S(
        \SUMB[2][12] ) );
  FA_X1 S2_2_13 ( .A(\ab[2][13] ), .B(n3), .CI(n32), .CO(\CARRYB[2][13] ), .S(
        \SUMB[2][13] ) );
  FA_X1 S3_2_14 ( .A(\ab[2][14] ), .B(n31), .CI(\ab[1][15] ), .CO(
        \CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  INV_X4 U2 ( .A(B[3]), .ZN(n91) );
  INV_X4 U3 ( .A(B[4]), .ZN(n90) );
  INV_X4 U4 ( .A(B[5]), .ZN(n89) );
  INV_X4 U5 ( .A(B[6]), .ZN(n88) );
  INV_X4 U6 ( .A(B[7]), .ZN(n87) );
  INV_X4 U7 ( .A(B[8]), .ZN(n86) );
  INV_X4 U8 ( .A(B[9]), .ZN(n85) );
  INV_X4 U9 ( .A(B[10]), .ZN(n84) );
  INV_X4 U10 ( .A(B[11]), .ZN(n83) );
  INV_X4 U11 ( .A(B[12]), .ZN(n82) );
  INV_X4 U12 ( .A(B[13]), .ZN(n81) );
  INV_X4 U13 ( .A(B[2]), .ZN(n92) );
  INV_X4 U14 ( .A(B[14]), .ZN(n80) );
  INV_X4 U15 ( .A(B[15]), .ZN(n79) );
  INV_X4 U16 ( .A(A[1]), .ZN(n77) );
  INV_X4 U17 ( .A(A[2]), .ZN(n76) );
  INV_X4 U18 ( .A(A[3]), .ZN(n75) );
  INV_X4 U19 ( .A(A[4]), .ZN(n74) );
  INV_X4 U20 ( .A(A[5]), .ZN(n73) );
  INV_X4 U21 ( .A(A[6]), .ZN(n72) );
  INV_X4 U22 ( .A(A[7]), .ZN(n71) );
  INV_X4 U23 ( .A(A[8]), .ZN(n70) );
  INV_X4 U24 ( .A(A[9]), .ZN(n69) );
  INV_X4 U25 ( .A(A[10]), .ZN(n68) );
  INV_X4 U26 ( .A(A[11]), .ZN(n67) );
  INV_X4 U27 ( .A(A[12]), .ZN(n66) );
  INV_X4 U28 ( .A(A[13]), .ZN(n65) );
  INV_X4 U29 ( .A(A[14]), .ZN(n64) );
  INV_X4 U30 ( .A(B[1]), .ZN(n93) );
  INV_X4 U31 ( .A(A[15]), .ZN(n63) );
  INV_X4 U32 ( .A(A[0]), .ZN(n78) );
  INV_X4 U33 ( .A(B[0]), .ZN(n94) );
  AND2_X4 U34 ( .A1(\ab[0][14] ), .A2(\ab[1][13] ), .ZN(n3) );
  AND2_X4 U35 ( .A1(\ab[0][13] ), .A2(\ab[1][12] ), .ZN(n4) );
  AND2_X4 U36 ( .A1(\ab[0][12] ), .A2(\ab[1][11] ), .ZN(n5) );
  AND2_X4 U37 ( .A1(\ab[0][11] ), .A2(\ab[1][10] ), .ZN(n6) );
  AND2_X4 U38 ( .A1(\ab[0][10] ), .A2(\ab[1][9] ), .ZN(n7) );
  AND2_X4 U39 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .ZN(n8) );
  AND2_X4 U40 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .ZN(n9) );
  AND2_X4 U41 ( .A1(\ab[0][7] ), .A2(\ab[1][6] ), .ZN(n10) );
  AND2_X4 U42 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .ZN(n11) );
  AND2_X4 U43 ( .A1(\ab[0][5] ), .A2(\ab[1][4] ), .ZN(n12) );
  AND2_X4 U44 ( .A1(\ab[0][4] ), .A2(\ab[1][3] ), .ZN(n13) );
  AND2_X4 U45 ( .A1(\ab[0][3] ), .A2(\ab[1][2] ), .ZN(n14) );
  AND2_X4 U46 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .ZN(n15) );
  AND2_X4 U47 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .ZN(n16) );
  XOR2_X2 U48 ( .A(\CARRYB[15][14] ), .B(\ab[15][15] ), .Z(n17) );
  XOR2_X2 U49 ( .A(\CARRYB[15][12] ), .B(\SUMB[15][13] ), .Z(n18) );
  XOR2_X2 U50 ( .A(\CARRYB[15][10] ), .B(\SUMB[15][11] ), .Z(n19) );
  XOR2_X2 U51 ( .A(\CARRYB[15][8] ), .B(\SUMB[15][9] ), .Z(n20) );
  XOR2_X2 U52 ( .A(\CARRYB[15][6] ), .B(\SUMB[15][7] ), .Z(n21) );
  XOR2_X2 U53 ( .A(\CARRYB[15][4] ), .B(\SUMB[15][5] ), .Z(n22) );
  XOR2_X2 U54 ( .A(\CARRYB[15][2] ), .B(\SUMB[15][3] ), .Z(n23) );
  XOR2_X2 U55 ( .A(\CARRYB[15][1] ), .B(\SUMB[15][2] ), .Z(n24) );
  XOR2_X2 U56 ( .A(\CARRYB[15][13] ), .B(\SUMB[15][14] ), .Z(n25) );
  XOR2_X2 U57 ( .A(\CARRYB[15][11] ), .B(\SUMB[15][12] ), .Z(n26) );
  XOR2_X2 U58 ( .A(\CARRYB[15][9] ), .B(\SUMB[15][10] ), .Z(n27) );
  XOR2_X2 U59 ( .A(\CARRYB[15][7] ), .B(\SUMB[15][8] ), .Z(n28) );
  XOR2_X2 U60 ( .A(\CARRYB[15][5] ), .B(\SUMB[15][6] ), .Z(n29) );
  XOR2_X2 U61 ( .A(\CARRYB[15][3] ), .B(\SUMB[15][4] ), .Z(n30) );
  AND2_X4 U62 ( .A1(\ab[0][15] ), .A2(\ab[1][14] ), .ZN(n31) );
  XOR2_X2 U63 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(n32) );
  XOR2_X2 U64 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(n33) );
  XOR2_X2 U65 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(n34) );
  XOR2_X2 U66 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(n35) );
  XOR2_X2 U67 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(n36) );
  XOR2_X2 U68 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(n37) );
  XOR2_X2 U69 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(n38) );
  XOR2_X2 U70 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(n39) );
  XOR2_X2 U71 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(n40) );
  XOR2_X2 U72 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(n41) );
  XOR2_X2 U73 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(n42) );
  XOR2_X2 U74 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(n43) );
  XOR2_X2 U75 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(n44) );
  XOR2_X2 U76 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(n45) );
  AND2_X4 U77 ( .A1(\CARRYB[15][13] ), .A2(\SUMB[15][14] ), .ZN(n46) );
  AND2_X4 U78 ( .A1(\CARRYB[15][11] ), .A2(\SUMB[15][12] ), .ZN(n47) );
  AND2_X4 U79 ( .A1(\CARRYB[15][9] ), .A2(\SUMB[15][10] ), .ZN(n48) );
  AND2_X4 U80 ( .A1(\CARRYB[15][7] ), .A2(\SUMB[15][8] ), .ZN(n49) );
  AND2_X4 U81 ( .A1(\CARRYB[15][5] ), .A2(\SUMB[15][6] ), .ZN(n50) );
  AND2_X4 U82 ( .A1(\CARRYB[15][3] ), .A2(\SUMB[15][4] ), .ZN(n51) );
  AND2_X4 U83 ( .A1(\CARRYB[15][1] ), .A2(\SUMB[15][2] ), .ZN(n52) );
  AND2_X4 U84 ( .A1(\CARRYB[15][12] ), .A2(\SUMB[15][13] ), .ZN(n53) );
  AND2_X4 U85 ( .A1(\CARRYB[15][10] ), .A2(\SUMB[15][11] ), .ZN(n54) );
  AND2_X4 U86 ( .A1(\CARRYB[15][8] ), .A2(\SUMB[15][9] ), .ZN(n55) );
  AND2_X4 U87 ( .A1(\CARRYB[15][6] ), .A2(\SUMB[15][7] ), .ZN(n56) );
  AND2_X4 U88 ( .A1(\CARRYB[15][4] ), .A2(\SUMB[15][5] ), .ZN(n57) );
  AND2_X4 U89 ( .A1(\CARRYB[15][2] ), .A2(\SUMB[15][3] ), .ZN(n58) );
  AND2_X4 U90 ( .A1(\CARRYB[15][0] ), .A2(\SUMB[15][1] ), .ZN(n59) );
  XOR2_X2 U91 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  XOR2_X2 U92 ( .A(\CARRYB[15][0] ), .B(\SUMB[15][1] ), .Z(n61) );
  AND2_X4 U93 ( .A1(\CARRYB[15][14] ), .A2(\ab[15][15] ), .ZN(n62) );
  NOR2_X1 U95 ( .A1(n69), .A2(n85), .ZN(\ab[9][9] ) );
  NOR2_X1 U96 ( .A1(n69), .A2(n86), .ZN(\ab[9][8] ) );
  NOR2_X1 U97 ( .A1(n69), .A2(n87), .ZN(\ab[9][7] ) );
  NOR2_X1 U98 ( .A1(n69), .A2(n88), .ZN(\ab[9][6] ) );
  NOR2_X1 U99 ( .A1(n69), .A2(n89), .ZN(\ab[9][5] ) );
  NOR2_X1 U100 ( .A1(n69), .A2(n90), .ZN(\ab[9][4] ) );
  NOR2_X1 U101 ( .A1(n69), .A2(n91), .ZN(\ab[9][3] ) );
  NOR2_X1 U102 ( .A1(n69), .A2(n92), .ZN(\ab[9][2] ) );
  NOR2_X1 U103 ( .A1(n69), .A2(n93), .ZN(\ab[9][1] ) );
  NOR2_X1 U104 ( .A1(n69), .A2(n79), .ZN(\ab[9][15] ) );
  NOR2_X1 U105 ( .A1(n69), .A2(n80), .ZN(\ab[9][14] ) );
  NOR2_X1 U106 ( .A1(n69), .A2(n81), .ZN(\ab[9][13] ) );
  NOR2_X1 U107 ( .A1(n69), .A2(n82), .ZN(\ab[9][12] ) );
  NOR2_X1 U108 ( .A1(n69), .A2(n83), .ZN(\ab[9][11] ) );
  NOR2_X1 U109 ( .A1(n69), .A2(n84), .ZN(\ab[9][10] ) );
  NOR2_X1 U110 ( .A1(n69), .A2(n94), .ZN(\ab[9][0] ) );
  NOR2_X1 U111 ( .A1(n85), .A2(n70), .ZN(\ab[8][9] ) );
  NOR2_X1 U112 ( .A1(n86), .A2(n70), .ZN(\ab[8][8] ) );
  NOR2_X1 U113 ( .A1(n87), .A2(n70), .ZN(\ab[8][7] ) );
  NOR2_X1 U114 ( .A1(n88), .A2(n70), .ZN(\ab[8][6] ) );
  NOR2_X1 U115 ( .A1(n89), .A2(n70), .ZN(\ab[8][5] ) );
  NOR2_X1 U116 ( .A1(n90), .A2(n70), .ZN(\ab[8][4] ) );
  NOR2_X1 U117 ( .A1(n91), .A2(n70), .ZN(\ab[8][3] ) );
  NOR2_X1 U118 ( .A1(n92), .A2(n70), .ZN(\ab[8][2] ) );
  NOR2_X1 U119 ( .A1(n93), .A2(n70), .ZN(\ab[8][1] ) );
  NOR2_X1 U120 ( .A1(n79), .A2(n70), .ZN(\ab[8][15] ) );
  NOR2_X1 U121 ( .A1(n80), .A2(n70), .ZN(\ab[8][14] ) );
  NOR2_X1 U122 ( .A1(n81), .A2(n70), .ZN(\ab[8][13] ) );
  NOR2_X1 U123 ( .A1(n82), .A2(n70), .ZN(\ab[8][12] ) );
  NOR2_X1 U124 ( .A1(n83), .A2(n70), .ZN(\ab[8][11] ) );
  NOR2_X1 U125 ( .A1(n84), .A2(n70), .ZN(\ab[8][10] ) );
  NOR2_X1 U126 ( .A1(n94), .A2(n70), .ZN(\ab[8][0] ) );
  NOR2_X1 U127 ( .A1(n85), .A2(n71), .ZN(\ab[7][9] ) );
  NOR2_X1 U128 ( .A1(n86), .A2(n71), .ZN(\ab[7][8] ) );
  NOR2_X1 U129 ( .A1(n87), .A2(n71), .ZN(\ab[7][7] ) );
  NOR2_X1 U130 ( .A1(n88), .A2(n71), .ZN(\ab[7][6] ) );
  NOR2_X1 U131 ( .A1(n89), .A2(n71), .ZN(\ab[7][5] ) );
  NOR2_X1 U132 ( .A1(n90), .A2(n71), .ZN(\ab[7][4] ) );
  NOR2_X1 U133 ( .A1(n91), .A2(n71), .ZN(\ab[7][3] ) );
  NOR2_X1 U134 ( .A1(n92), .A2(n71), .ZN(\ab[7][2] ) );
  NOR2_X1 U135 ( .A1(n93), .A2(n71), .ZN(\ab[7][1] ) );
  NOR2_X1 U136 ( .A1(n79), .A2(n71), .ZN(\ab[7][15] ) );
  NOR2_X1 U137 ( .A1(n80), .A2(n71), .ZN(\ab[7][14] ) );
  NOR2_X1 U138 ( .A1(n81), .A2(n71), .ZN(\ab[7][13] ) );
  NOR2_X1 U139 ( .A1(n82), .A2(n71), .ZN(\ab[7][12] ) );
  NOR2_X1 U140 ( .A1(n83), .A2(n71), .ZN(\ab[7][11] ) );
  NOR2_X1 U141 ( .A1(n84), .A2(n71), .ZN(\ab[7][10] ) );
  NOR2_X1 U142 ( .A1(n94), .A2(n71), .ZN(\ab[7][0] ) );
  NOR2_X1 U143 ( .A1(n85), .A2(n72), .ZN(\ab[6][9] ) );
  NOR2_X1 U144 ( .A1(n86), .A2(n72), .ZN(\ab[6][8] ) );
  NOR2_X1 U145 ( .A1(n87), .A2(n72), .ZN(\ab[6][7] ) );
  NOR2_X1 U146 ( .A1(n88), .A2(n72), .ZN(\ab[6][6] ) );
  NOR2_X1 U147 ( .A1(n89), .A2(n72), .ZN(\ab[6][5] ) );
  NOR2_X1 U148 ( .A1(n90), .A2(n72), .ZN(\ab[6][4] ) );
  NOR2_X1 U149 ( .A1(n91), .A2(n72), .ZN(\ab[6][3] ) );
  NOR2_X1 U150 ( .A1(n92), .A2(n72), .ZN(\ab[6][2] ) );
  NOR2_X1 U151 ( .A1(n93), .A2(n72), .ZN(\ab[6][1] ) );
  NOR2_X1 U152 ( .A1(n79), .A2(n72), .ZN(\ab[6][15] ) );
  NOR2_X1 U153 ( .A1(n80), .A2(n72), .ZN(\ab[6][14] ) );
  NOR2_X1 U154 ( .A1(n81), .A2(n72), .ZN(\ab[6][13] ) );
  NOR2_X1 U155 ( .A1(n82), .A2(n72), .ZN(\ab[6][12] ) );
  NOR2_X1 U156 ( .A1(n83), .A2(n72), .ZN(\ab[6][11] ) );
  NOR2_X1 U157 ( .A1(n84), .A2(n72), .ZN(\ab[6][10] ) );
  NOR2_X1 U158 ( .A1(n94), .A2(n72), .ZN(\ab[6][0] ) );
  NOR2_X1 U159 ( .A1(n85), .A2(n73), .ZN(\ab[5][9] ) );
  NOR2_X1 U160 ( .A1(n86), .A2(n73), .ZN(\ab[5][8] ) );
  NOR2_X1 U161 ( .A1(n87), .A2(n73), .ZN(\ab[5][7] ) );
  NOR2_X1 U162 ( .A1(n88), .A2(n73), .ZN(\ab[5][6] ) );
  NOR2_X1 U163 ( .A1(n89), .A2(n73), .ZN(\ab[5][5] ) );
  NOR2_X1 U164 ( .A1(n90), .A2(n73), .ZN(\ab[5][4] ) );
  NOR2_X1 U165 ( .A1(n91), .A2(n73), .ZN(\ab[5][3] ) );
  NOR2_X1 U166 ( .A1(n92), .A2(n73), .ZN(\ab[5][2] ) );
  NOR2_X1 U167 ( .A1(n93), .A2(n73), .ZN(\ab[5][1] ) );
  NOR2_X1 U168 ( .A1(n79), .A2(n73), .ZN(\ab[5][15] ) );
  NOR2_X1 U169 ( .A1(n80), .A2(n73), .ZN(\ab[5][14] ) );
  NOR2_X1 U170 ( .A1(n81), .A2(n73), .ZN(\ab[5][13] ) );
  NOR2_X1 U171 ( .A1(n82), .A2(n73), .ZN(\ab[5][12] ) );
  NOR2_X1 U172 ( .A1(n83), .A2(n73), .ZN(\ab[5][11] ) );
  NOR2_X1 U173 ( .A1(n84), .A2(n73), .ZN(\ab[5][10] ) );
  NOR2_X1 U174 ( .A1(n94), .A2(n73), .ZN(\ab[5][0] ) );
  NOR2_X1 U175 ( .A1(n85), .A2(n74), .ZN(\ab[4][9] ) );
  NOR2_X1 U176 ( .A1(n86), .A2(n74), .ZN(\ab[4][8] ) );
  NOR2_X1 U177 ( .A1(n87), .A2(n74), .ZN(\ab[4][7] ) );
  NOR2_X1 U178 ( .A1(n88), .A2(n74), .ZN(\ab[4][6] ) );
  NOR2_X1 U179 ( .A1(n89), .A2(n74), .ZN(\ab[4][5] ) );
  NOR2_X1 U180 ( .A1(n90), .A2(n74), .ZN(\ab[4][4] ) );
  NOR2_X1 U181 ( .A1(n91), .A2(n74), .ZN(\ab[4][3] ) );
  NOR2_X1 U182 ( .A1(n92), .A2(n74), .ZN(\ab[4][2] ) );
  NOR2_X1 U183 ( .A1(n93), .A2(n74), .ZN(\ab[4][1] ) );
  NOR2_X1 U184 ( .A1(n79), .A2(n74), .ZN(\ab[4][15] ) );
  NOR2_X1 U185 ( .A1(n80), .A2(n74), .ZN(\ab[4][14] ) );
  NOR2_X1 U186 ( .A1(n81), .A2(n74), .ZN(\ab[4][13] ) );
  NOR2_X1 U187 ( .A1(n82), .A2(n74), .ZN(\ab[4][12] ) );
  NOR2_X1 U188 ( .A1(n83), .A2(n74), .ZN(\ab[4][11] ) );
  NOR2_X1 U189 ( .A1(n84), .A2(n74), .ZN(\ab[4][10] ) );
  NOR2_X1 U190 ( .A1(n94), .A2(n74), .ZN(\ab[4][0] ) );
  NOR2_X1 U191 ( .A1(n85), .A2(n75), .ZN(\ab[3][9] ) );
  NOR2_X1 U192 ( .A1(n86), .A2(n75), .ZN(\ab[3][8] ) );
  NOR2_X1 U193 ( .A1(n87), .A2(n75), .ZN(\ab[3][7] ) );
  NOR2_X1 U194 ( .A1(n88), .A2(n75), .ZN(\ab[3][6] ) );
  NOR2_X1 U195 ( .A1(n89), .A2(n75), .ZN(\ab[3][5] ) );
  NOR2_X1 U196 ( .A1(n90), .A2(n75), .ZN(\ab[3][4] ) );
  NOR2_X1 U197 ( .A1(n91), .A2(n75), .ZN(\ab[3][3] ) );
  NOR2_X1 U198 ( .A1(n92), .A2(n75), .ZN(\ab[3][2] ) );
  NOR2_X1 U199 ( .A1(n93), .A2(n75), .ZN(\ab[3][1] ) );
  NOR2_X1 U200 ( .A1(n79), .A2(n75), .ZN(\ab[3][15] ) );
  NOR2_X1 U201 ( .A1(n80), .A2(n75), .ZN(\ab[3][14] ) );
  NOR2_X1 U202 ( .A1(n81), .A2(n75), .ZN(\ab[3][13] ) );
  NOR2_X1 U203 ( .A1(n82), .A2(n75), .ZN(\ab[3][12] ) );
  NOR2_X1 U204 ( .A1(n83), .A2(n75), .ZN(\ab[3][11] ) );
  NOR2_X1 U205 ( .A1(n84), .A2(n75), .ZN(\ab[3][10] ) );
  NOR2_X1 U206 ( .A1(n94), .A2(n75), .ZN(\ab[3][0] ) );
  NOR2_X1 U207 ( .A1(n85), .A2(n76), .ZN(\ab[2][9] ) );
  NOR2_X1 U208 ( .A1(n86), .A2(n76), .ZN(\ab[2][8] ) );
  NOR2_X1 U209 ( .A1(n87), .A2(n76), .ZN(\ab[2][7] ) );
  NOR2_X1 U210 ( .A1(n88), .A2(n76), .ZN(\ab[2][6] ) );
  NOR2_X1 U211 ( .A1(n89), .A2(n76), .ZN(\ab[2][5] ) );
  NOR2_X1 U212 ( .A1(n90), .A2(n76), .ZN(\ab[2][4] ) );
  NOR2_X1 U213 ( .A1(n91), .A2(n76), .ZN(\ab[2][3] ) );
  NOR2_X1 U214 ( .A1(n92), .A2(n76), .ZN(\ab[2][2] ) );
  NOR2_X1 U215 ( .A1(n93), .A2(n76), .ZN(\ab[2][1] ) );
  NOR2_X1 U216 ( .A1(n79), .A2(n76), .ZN(\ab[2][15] ) );
  NOR2_X1 U217 ( .A1(n80), .A2(n76), .ZN(\ab[2][14] ) );
  NOR2_X1 U218 ( .A1(n81), .A2(n76), .ZN(\ab[2][13] ) );
  NOR2_X1 U219 ( .A1(n82), .A2(n76), .ZN(\ab[2][12] ) );
  NOR2_X1 U220 ( .A1(n83), .A2(n76), .ZN(\ab[2][11] ) );
  NOR2_X1 U221 ( .A1(n84), .A2(n76), .ZN(\ab[2][10] ) );
  NOR2_X1 U222 ( .A1(n94), .A2(n76), .ZN(\ab[2][0] ) );
  NOR2_X1 U223 ( .A1(n85), .A2(n77), .ZN(\ab[1][9] ) );
  NOR2_X1 U224 ( .A1(n86), .A2(n77), .ZN(\ab[1][8] ) );
  NOR2_X1 U225 ( .A1(n87), .A2(n77), .ZN(\ab[1][7] ) );
  NOR2_X1 U226 ( .A1(n88), .A2(n77), .ZN(\ab[1][6] ) );
  NOR2_X1 U227 ( .A1(n89), .A2(n77), .ZN(\ab[1][5] ) );
  NOR2_X1 U228 ( .A1(n90), .A2(n77), .ZN(\ab[1][4] ) );
  NOR2_X1 U229 ( .A1(n91), .A2(n77), .ZN(\ab[1][3] ) );
  NOR2_X1 U230 ( .A1(n92), .A2(n77), .ZN(\ab[1][2] ) );
  NOR2_X1 U231 ( .A1(n93), .A2(n77), .ZN(\ab[1][1] ) );
  NOR2_X1 U232 ( .A1(n79), .A2(n77), .ZN(\ab[1][15] ) );
  NOR2_X1 U233 ( .A1(n80), .A2(n77), .ZN(\ab[1][14] ) );
  NOR2_X1 U234 ( .A1(n81), .A2(n77), .ZN(\ab[1][13] ) );
  NOR2_X1 U235 ( .A1(n82), .A2(n77), .ZN(\ab[1][12] ) );
  NOR2_X1 U236 ( .A1(n83), .A2(n77), .ZN(\ab[1][11] ) );
  NOR2_X1 U237 ( .A1(n84), .A2(n77), .ZN(\ab[1][10] ) );
  NOR2_X1 U238 ( .A1(n94), .A2(n77), .ZN(\ab[1][0] ) );
  NOR2_X1 U239 ( .A1(n85), .A2(n63), .ZN(\ab[15][9] ) );
  NOR2_X1 U240 ( .A1(n86), .A2(n63), .ZN(\ab[15][8] ) );
  NOR2_X1 U241 ( .A1(n87), .A2(n63), .ZN(\ab[15][7] ) );
  NOR2_X1 U242 ( .A1(n88), .A2(n63), .ZN(\ab[15][6] ) );
  NOR2_X1 U243 ( .A1(n89), .A2(n63), .ZN(\ab[15][5] ) );
  NOR2_X1 U244 ( .A1(n90), .A2(n63), .ZN(\ab[15][4] ) );
  NOR2_X1 U245 ( .A1(n91), .A2(n63), .ZN(\ab[15][3] ) );
  NOR2_X1 U246 ( .A1(n92), .A2(n63), .ZN(\ab[15][2] ) );
  NOR2_X1 U247 ( .A1(n93), .A2(n63), .ZN(\ab[15][1] ) );
  NOR2_X1 U248 ( .A1(n79), .A2(n63), .ZN(\ab[15][15] ) );
  NOR2_X1 U249 ( .A1(n80), .A2(n63), .ZN(\ab[15][14] ) );
  NOR2_X1 U250 ( .A1(n81), .A2(n63), .ZN(\ab[15][13] ) );
  NOR2_X1 U251 ( .A1(n82), .A2(n63), .ZN(\ab[15][12] ) );
  NOR2_X1 U252 ( .A1(n83), .A2(n63), .ZN(\ab[15][11] ) );
  NOR2_X1 U253 ( .A1(n84), .A2(n63), .ZN(\ab[15][10] ) );
  NOR2_X1 U254 ( .A1(n94), .A2(n63), .ZN(\ab[15][0] ) );
  NOR2_X1 U255 ( .A1(n85), .A2(n64), .ZN(\ab[14][9] ) );
  NOR2_X1 U256 ( .A1(n86), .A2(n64), .ZN(\ab[14][8] ) );
  NOR2_X1 U257 ( .A1(n87), .A2(n64), .ZN(\ab[14][7] ) );
  NOR2_X1 U258 ( .A1(n88), .A2(n64), .ZN(\ab[14][6] ) );
  NOR2_X1 U259 ( .A1(n89), .A2(n64), .ZN(\ab[14][5] ) );
  NOR2_X1 U260 ( .A1(n90), .A2(n64), .ZN(\ab[14][4] ) );
  NOR2_X1 U261 ( .A1(n91), .A2(n64), .ZN(\ab[14][3] ) );
  NOR2_X1 U262 ( .A1(n92), .A2(n64), .ZN(\ab[14][2] ) );
  NOR2_X1 U263 ( .A1(n93), .A2(n64), .ZN(\ab[14][1] ) );
  NOR2_X1 U264 ( .A1(n79), .A2(n64), .ZN(\ab[14][15] ) );
  NOR2_X1 U265 ( .A1(n80), .A2(n64), .ZN(\ab[14][14] ) );
  NOR2_X1 U266 ( .A1(n81), .A2(n64), .ZN(\ab[14][13] ) );
  NOR2_X1 U267 ( .A1(n82), .A2(n64), .ZN(\ab[14][12] ) );
  NOR2_X1 U268 ( .A1(n83), .A2(n64), .ZN(\ab[14][11] ) );
  NOR2_X1 U269 ( .A1(n84), .A2(n64), .ZN(\ab[14][10] ) );
  NOR2_X1 U270 ( .A1(n94), .A2(n64), .ZN(\ab[14][0] ) );
  NOR2_X1 U271 ( .A1(n85), .A2(n65), .ZN(\ab[13][9] ) );
  NOR2_X1 U272 ( .A1(n86), .A2(n65), .ZN(\ab[13][8] ) );
  NOR2_X1 U273 ( .A1(n87), .A2(n65), .ZN(\ab[13][7] ) );
  NOR2_X1 U274 ( .A1(n88), .A2(n65), .ZN(\ab[13][6] ) );
  NOR2_X1 U275 ( .A1(n89), .A2(n65), .ZN(\ab[13][5] ) );
  NOR2_X1 U276 ( .A1(n90), .A2(n65), .ZN(\ab[13][4] ) );
  NOR2_X1 U277 ( .A1(n91), .A2(n65), .ZN(\ab[13][3] ) );
  NOR2_X1 U278 ( .A1(n92), .A2(n65), .ZN(\ab[13][2] ) );
  NOR2_X1 U279 ( .A1(n93), .A2(n65), .ZN(\ab[13][1] ) );
  NOR2_X1 U280 ( .A1(n79), .A2(n65), .ZN(\ab[13][15] ) );
  NOR2_X1 U281 ( .A1(n80), .A2(n65), .ZN(\ab[13][14] ) );
  NOR2_X1 U282 ( .A1(n81), .A2(n65), .ZN(\ab[13][13] ) );
  NOR2_X1 U283 ( .A1(n82), .A2(n65), .ZN(\ab[13][12] ) );
  NOR2_X1 U284 ( .A1(n83), .A2(n65), .ZN(\ab[13][11] ) );
  NOR2_X1 U285 ( .A1(n84), .A2(n65), .ZN(\ab[13][10] ) );
  NOR2_X1 U286 ( .A1(n94), .A2(n65), .ZN(\ab[13][0] ) );
  NOR2_X1 U287 ( .A1(n85), .A2(n66), .ZN(\ab[12][9] ) );
  NOR2_X1 U288 ( .A1(n86), .A2(n66), .ZN(\ab[12][8] ) );
  NOR2_X1 U289 ( .A1(n87), .A2(n66), .ZN(\ab[12][7] ) );
  NOR2_X1 U290 ( .A1(n88), .A2(n66), .ZN(\ab[12][6] ) );
  NOR2_X1 U291 ( .A1(n89), .A2(n66), .ZN(\ab[12][5] ) );
  NOR2_X1 U292 ( .A1(n90), .A2(n66), .ZN(\ab[12][4] ) );
  NOR2_X1 U293 ( .A1(n91), .A2(n66), .ZN(\ab[12][3] ) );
  NOR2_X1 U294 ( .A1(n92), .A2(n66), .ZN(\ab[12][2] ) );
  NOR2_X1 U295 ( .A1(n93), .A2(n66), .ZN(\ab[12][1] ) );
  NOR2_X1 U296 ( .A1(n79), .A2(n66), .ZN(\ab[12][15] ) );
  NOR2_X1 U297 ( .A1(n80), .A2(n66), .ZN(\ab[12][14] ) );
  NOR2_X1 U298 ( .A1(n81), .A2(n66), .ZN(\ab[12][13] ) );
  NOR2_X1 U299 ( .A1(n82), .A2(n66), .ZN(\ab[12][12] ) );
  NOR2_X1 U300 ( .A1(n83), .A2(n66), .ZN(\ab[12][11] ) );
  NOR2_X1 U301 ( .A1(n84), .A2(n66), .ZN(\ab[12][10] ) );
  NOR2_X1 U302 ( .A1(n94), .A2(n66), .ZN(\ab[12][0] ) );
  NOR2_X1 U303 ( .A1(n85), .A2(n67), .ZN(\ab[11][9] ) );
  NOR2_X1 U304 ( .A1(n86), .A2(n67), .ZN(\ab[11][8] ) );
  NOR2_X1 U305 ( .A1(n87), .A2(n67), .ZN(\ab[11][7] ) );
  NOR2_X1 U306 ( .A1(n88), .A2(n67), .ZN(\ab[11][6] ) );
  NOR2_X1 U307 ( .A1(n89), .A2(n67), .ZN(\ab[11][5] ) );
  NOR2_X1 U308 ( .A1(n90), .A2(n67), .ZN(\ab[11][4] ) );
  NOR2_X1 U309 ( .A1(n91), .A2(n67), .ZN(\ab[11][3] ) );
  NOR2_X1 U310 ( .A1(n92), .A2(n67), .ZN(\ab[11][2] ) );
  NOR2_X1 U311 ( .A1(n93), .A2(n67), .ZN(\ab[11][1] ) );
  NOR2_X1 U312 ( .A1(n79), .A2(n67), .ZN(\ab[11][15] ) );
  NOR2_X1 U313 ( .A1(n80), .A2(n67), .ZN(\ab[11][14] ) );
  NOR2_X1 U314 ( .A1(n81), .A2(n67), .ZN(\ab[11][13] ) );
  NOR2_X1 U315 ( .A1(n82), .A2(n67), .ZN(\ab[11][12] ) );
  NOR2_X1 U316 ( .A1(n83), .A2(n67), .ZN(\ab[11][11] ) );
  NOR2_X1 U317 ( .A1(n84), .A2(n67), .ZN(\ab[11][10] ) );
  NOR2_X1 U318 ( .A1(n94), .A2(n67), .ZN(\ab[11][0] ) );
  NOR2_X1 U319 ( .A1(n85), .A2(n68), .ZN(\ab[10][9] ) );
  NOR2_X1 U320 ( .A1(n86), .A2(n68), .ZN(\ab[10][8] ) );
  NOR2_X1 U321 ( .A1(n87), .A2(n68), .ZN(\ab[10][7] ) );
  NOR2_X1 U322 ( .A1(n88), .A2(n68), .ZN(\ab[10][6] ) );
  NOR2_X1 U323 ( .A1(n89), .A2(n68), .ZN(\ab[10][5] ) );
  NOR2_X1 U324 ( .A1(n90), .A2(n68), .ZN(\ab[10][4] ) );
  NOR2_X1 U325 ( .A1(n91), .A2(n68), .ZN(\ab[10][3] ) );
  NOR2_X1 U326 ( .A1(n92), .A2(n68), .ZN(\ab[10][2] ) );
  NOR2_X1 U327 ( .A1(n93), .A2(n68), .ZN(\ab[10][1] ) );
  NOR2_X1 U328 ( .A1(n79), .A2(n68), .ZN(\ab[10][15] ) );
  NOR2_X1 U329 ( .A1(n80), .A2(n68), .ZN(\ab[10][14] ) );
  NOR2_X1 U330 ( .A1(n81), .A2(n68), .ZN(\ab[10][13] ) );
  NOR2_X1 U331 ( .A1(n82), .A2(n68), .ZN(\ab[10][12] ) );
  NOR2_X1 U332 ( .A1(n83), .A2(n68), .ZN(\ab[10][11] ) );
  NOR2_X1 U333 ( .A1(n84), .A2(n68), .ZN(\ab[10][10] ) );
  NOR2_X1 U334 ( .A1(n94), .A2(n68), .ZN(\ab[10][0] ) );
  NOR2_X1 U335 ( .A1(n85), .A2(n78), .ZN(\ab[0][9] ) );
  NOR2_X1 U336 ( .A1(n86), .A2(n78), .ZN(\ab[0][8] ) );
  NOR2_X1 U337 ( .A1(n87), .A2(n78), .ZN(\ab[0][7] ) );
  NOR2_X1 U338 ( .A1(n88), .A2(n78), .ZN(\ab[0][6] ) );
  NOR2_X1 U339 ( .A1(n89), .A2(n78), .ZN(\ab[0][5] ) );
  NOR2_X1 U340 ( .A1(n90), .A2(n78), .ZN(\ab[0][4] ) );
  NOR2_X1 U341 ( .A1(n91), .A2(n78), .ZN(\ab[0][3] ) );
  NOR2_X1 U342 ( .A1(n92), .A2(n78), .ZN(\ab[0][2] ) );
  NOR2_X1 U343 ( .A1(n93), .A2(n78), .ZN(\ab[0][1] ) );
  NOR2_X1 U344 ( .A1(n79), .A2(n78), .ZN(\ab[0][15] ) );
  NOR2_X1 U345 ( .A1(n80), .A2(n78), .ZN(\ab[0][14] ) );
  NOR2_X1 U346 ( .A1(n81), .A2(n78), .ZN(\ab[0][13] ) );
  NOR2_X1 U347 ( .A1(n82), .A2(n78), .ZN(\ab[0][12] ) );
  NOR2_X1 U348 ( .A1(n83), .A2(n78), .ZN(\ab[0][11] ) );
  NOR2_X1 U349 ( .A1(n84), .A2(n78), .ZN(\ab[0][10] ) );
  NOR2_X1 U350 ( .A1(n94), .A2(n78), .ZN(PRODUCT[0]) );
  multiplier_DW01_add_3 FS_1 ( .A({1'b0, n17, n25, n18, n26, n19, n27, n20, 
        n28, n21, n29, n22, n30, n23, n24, n61, \SUMB[15][0] , \A1[12] , 
        \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , 
        \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({n62, n46, n53, n47, 
        n54, n48, n55, n49, n56, n50, n57, n51, n58, n52, n59, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .CI(1'b0), .SUM(PRODUCT[31:2]) );
endmodule


module multiplier ( clk, reset, mul, a, b, done, working, result );
  input [0:31] a;
  input [0:31] b;
  output [0:63] result;
  input clk, reset, mul;
  output done, working;
  wire   N14, N15, N16, N43, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93,
         N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160,
         N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171,
         N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182,
         N183, N184, N185, N218, N219, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N314, N315, N316, N317, N318, N319, N320, N321, N322,
         N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333,
         N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344,
         N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366,
         N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377,
         N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410,
         N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421,
         N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432,
         N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443,
         N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454,
         N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465,
         N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476,
         N477, N478, n32, n33, n34, n35, n36, n37, n38, N298, N297, N296, N295,
         N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284,
         N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273,
         N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262,
         N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251,
         N250, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208,
         N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197,
         N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n66, n67;
  wire   [0:2] CurrentState;
  wire   [0:31] L;
  wire   [0:31] Z;
  wire   [0:31] H;
  wire   [0:31] P1;
  wire   [0:31] P;
  wire   [0:31] P2;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46;

  OAI211_X2 U3 ( .C1(n59), .C2(n63), .A(n33), .B(n34), .ZN(N478) );
  AND2_X2 U9 ( .A1(N185), .A2(n40), .ZN(N476) );
  AND2_X2 U10 ( .A1(N184), .A2(n40), .ZN(N475) );
  AND2_X2 U11 ( .A1(N183), .A2(n40), .ZN(N474) );
  AND2_X2 U12 ( .A1(N182), .A2(n40), .ZN(N473) );
  AND2_X2 U13 ( .A1(N181), .A2(n40), .ZN(N472) );
  AND2_X2 U14 ( .A1(N180), .A2(n64), .ZN(N471) );
  AND2_X2 U15 ( .A1(N179), .A2(n64), .ZN(N470) );
  AND2_X2 U16 ( .A1(N178), .A2(n64), .ZN(N469) );
  AND2_X2 U17 ( .A1(N177), .A2(n64), .ZN(N468) );
  AND2_X2 U18 ( .A1(N176), .A2(n64), .ZN(N467) );
  AND2_X2 U19 ( .A1(N175), .A2(n40), .ZN(N466) );
  AND2_X2 U20 ( .A1(N174), .A2(n40), .ZN(N465) );
  AND2_X2 U21 ( .A1(N173), .A2(n40), .ZN(N464) );
  AND2_X2 U22 ( .A1(N172), .A2(n40), .ZN(N463) );
  AND2_X2 U23 ( .A1(N171), .A2(n40), .ZN(N462) );
  AND2_X2 U24 ( .A1(N170), .A2(n40), .ZN(N461) );
  AND2_X2 U25 ( .A1(N169), .A2(n40), .ZN(N460) );
  AND2_X2 U26 ( .A1(N168), .A2(n40), .ZN(N459) );
  AND2_X2 U27 ( .A1(N167), .A2(n40), .ZN(N458) );
  AND2_X2 U28 ( .A1(N166), .A2(n40), .ZN(N457) );
  AND2_X2 U29 ( .A1(N165), .A2(n40), .ZN(N456) );
  AND2_X2 U30 ( .A1(N164), .A2(n40), .ZN(N455) );
  AND2_X2 U31 ( .A1(N163), .A2(n40), .ZN(N454) );
  AND2_X2 U32 ( .A1(N162), .A2(n40), .ZN(N453) );
  AND2_X2 U33 ( .A1(N161), .A2(n40), .ZN(N452) );
  AND2_X2 U34 ( .A1(N160), .A2(n40), .ZN(N451) );
  AND2_X2 U35 ( .A1(N159), .A2(n40), .ZN(N450) );
  AND2_X2 U36 ( .A1(N158), .A2(n40), .ZN(N449) );
  AND2_X2 U37 ( .A1(N157), .A2(n40), .ZN(N448) );
  AND2_X2 U38 ( .A1(N156), .A2(n40), .ZN(N447) );
  AND2_X2 U39 ( .A1(N155), .A2(n40), .ZN(N446) );
  AND2_X2 U40 ( .A1(N154), .A2(n40), .ZN(N445) );
  NAND2_X2 U41 ( .A1(n59), .A2(n35), .ZN(N444) );
  AND2_X2 U42 ( .A1(N249), .A2(n41), .ZN(N443) );
  AND2_X2 U43 ( .A1(N248), .A2(n41), .ZN(N442) );
  AND2_X2 U44 ( .A1(N247), .A2(n41), .ZN(N441) );
  AND2_X2 U45 ( .A1(N246), .A2(n41), .ZN(N440) );
  AND2_X2 U46 ( .A1(N245), .A2(n41), .ZN(N439) );
  AND2_X2 U47 ( .A1(N244), .A2(n41), .ZN(N438) );
  AND2_X2 U48 ( .A1(N243), .A2(n41), .ZN(N437) );
  AND2_X2 U49 ( .A1(N242), .A2(n41), .ZN(N436) );
  AND2_X2 U50 ( .A1(N241), .A2(n41), .ZN(N435) );
  AND2_X2 U51 ( .A1(N240), .A2(n41), .ZN(N434) );
  AND2_X2 U52 ( .A1(N239), .A2(n41), .ZN(N433) );
  AND2_X2 U53 ( .A1(N238), .A2(n42), .ZN(N432) );
  AND2_X2 U54 ( .A1(N237), .A2(n42), .ZN(N431) );
  AND2_X2 U55 ( .A1(N236), .A2(n42), .ZN(N430) );
  AND2_X2 U56 ( .A1(N235), .A2(n42), .ZN(N429) );
  AND2_X2 U57 ( .A1(N234), .A2(n42), .ZN(N428) );
  AND2_X2 U58 ( .A1(N233), .A2(n42), .ZN(N427) );
  AND2_X2 U59 ( .A1(N232), .A2(n42), .ZN(N426) );
  AND2_X2 U60 ( .A1(N231), .A2(n42), .ZN(N425) );
  AND2_X2 U61 ( .A1(N230), .A2(n42), .ZN(N424) );
  AND2_X2 U62 ( .A1(N229), .A2(n42), .ZN(N423) );
  AND2_X2 U63 ( .A1(N228), .A2(n42), .ZN(N422) );
  AND2_X2 U64 ( .A1(N227), .A2(n42), .ZN(N421) );
  AND2_X2 U65 ( .A1(N226), .A2(n41), .ZN(N420) );
  AND2_X2 U66 ( .A1(N225), .A2(n66), .ZN(N419) );
  AND2_X2 U67 ( .A1(N224), .A2(n66), .ZN(N418) );
  AND2_X2 U68 ( .A1(N223), .A2(n42), .ZN(N417) );
  AND2_X2 U69 ( .A1(N222), .A2(n41), .ZN(N416) );
  AND2_X2 U70 ( .A1(N221), .A2(n66), .ZN(N415) );
  AND2_X2 U71 ( .A1(N220), .A2(n42), .ZN(N414) );
  AND2_X2 U72 ( .A1(N219), .A2(n41), .ZN(N413) );
  AND2_X2 U73 ( .A1(N218), .A2(n66), .ZN(N412) );
  NAND2_X2 U74 ( .A1(n59), .A2(n33), .ZN(N411) );
  AND2_X2 U75 ( .A1(N153), .A2(n38), .ZN(N410) );
  AND2_X2 U76 ( .A1(N152), .A2(n38), .ZN(N409) );
  AND2_X2 U77 ( .A1(N151), .A2(n38), .ZN(N408) );
  AND2_X2 U78 ( .A1(N150), .A2(n38), .ZN(N407) );
  AND2_X2 U79 ( .A1(N149), .A2(n38), .ZN(N406) );
  AND2_X2 U80 ( .A1(N148), .A2(n38), .ZN(N405) );
  AND2_X2 U81 ( .A1(N147), .A2(n38), .ZN(N404) );
  AND2_X2 U82 ( .A1(N146), .A2(n38), .ZN(N403) );
  AND2_X2 U83 ( .A1(N145), .A2(n38), .ZN(N402) );
  AND2_X2 U84 ( .A1(N144), .A2(n38), .ZN(N401) );
  AND2_X2 U85 ( .A1(N143), .A2(n45), .ZN(N400) );
  AND2_X2 U86 ( .A1(N142), .A2(n43), .ZN(N399) );
  AND2_X2 U87 ( .A1(N141), .A2(n43), .ZN(N398) );
  AND2_X2 U88 ( .A1(N140), .A2(n38), .ZN(N397) );
  AND2_X2 U89 ( .A1(N139), .A2(n38), .ZN(N396) );
  AND2_X2 U90 ( .A1(N138), .A2(n38), .ZN(N395) );
  AND2_X2 U91 ( .A1(N137), .A2(n38), .ZN(N394) );
  AND2_X2 U92 ( .A1(N136), .A2(n43), .ZN(N393) );
  AND2_X2 U93 ( .A1(N135), .A2(n38), .ZN(N392) );
  AND2_X2 U94 ( .A1(N134), .A2(n38), .ZN(N391) );
  AND2_X2 U95 ( .A1(N133), .A2(n38), .ZN(N390) );
  AND2_X2 U96 ( .A1(N132), .A2(n38), .ZN(N389) );
  AND2_X2 U97 ( .A1(N131), .A2(n38), .ZN(N388) );
  AND2_X2 U98 ( .A1(N130), .A2(n38), .ZN(N387) );
  AND2_X2 U99 ( .A1(N129), .A2(n38), .ZN(N386) );
  AND2_X2 U100 ( .A1(N128), .A2(n38), .ZN(N385) );
  AND2_X2 U101 ( .A1(N127), .A2(n38), .ZN(N384) );
  AND2_X2 U102 ( .A1(N126), .A2(n38), .ZN(N383) );
  AND2_X2 U103 ( .A1(N125), .A2(n38), .ZN(N382) );
  AND2_X2 U104 ( .A1(N124), .A2(n43), .ZN(N381) );
  AND2_X2 U105 ( .A1(N123), .A2(n38), .ZN(N380) );
  AND2_X2 U106 ( .A1(N122), .A2(n38), .ZN(N379) );
  OR2_X2 U107 ( .A1(N43), .A2(n45), .ZN(N378) );
  DFF_X2 \CurrentState_reg[0]  ( .D(N16), .CK(clk), .Q(CurrentState[0]), .QN(
        n39) );
  DLH_X2 \P2_reg[15]  ( .G(n45), .D(N121), .Q(P2[15]) );
  DLH_X2 \P2_reg[16]  ( .G(n45), .D(N120), .Q(P2[16]) );
  DLH_X2 \P2_reg[17]  ( .G(n45), .D(N119), .Q(P2[17]) );
  DLH_X2 \P2_reg[18]  ( .G(n45), .D(N118), .Q(P2[18]) );
  DLH_X2 \P2_reg[19]  ( .G(n45), .D(N117), .Q(P2[19]) );
  DLH_X2 \P2_reg[20]  ( .G(n45), .D(N116), .Q(P2[20]) );
  DLH_X2 \P2_reg[21]  ( .G(n45), .D(N115), .Q(P2[21]) );
  DLH_X2 \P2_reg[22]  ( .G(n45), .D(N114), .Q(P2[22]) );
  DLH_X2 \P2_reg[23]  ( .G(n45), .D(N113), .Q(P2[23]) );
  DLH_X2 \P2_reg[24]  ( .G(n45), .D(N112), .Q(P2[24]) );
  DLH_X2 \P2_reg[25]  ( .G(n45), .D(N111), .Q(P2[25]) );
  DLH_X2 \P2_reg[26]  ( .G(n45), .D(N110), .Q(P2[26]) );
  DLH_X2 \P2_reg[27]  ( .G(n45), .D(N109), .Q(P2[27]) );
  DLH_X2 \P2_reg[28]  ( .G(n45), .D(N108), .Q(P2[28]) );
  DLH_X2 \P2_reg[29]  ( .G(n45), .D(N107), .Q(P2[29]) );
  DLH_X2 \P2_reg[30]  ( .G(n45), .D(N106), .Q(P2[30]) );
  DLH_X2 \P2_reg[31]  ( .G(n45), .D(N105), .Q(P2[31]) );
  DLH_X2 done_reg ( .G(n67), .D(n37), .Q(done) );
  DLH_X2 \P_reg[0]  ( .G(n49), .D(N476), .Q(P[0]) );
  DLH_X2 \P_reg[1]  ( .G(n49), .D(N475), .Q(P[1]) );
  DLH_X2 \P_reg[2]  ( .G(n49), .D(N474), .Q(P[2]) );
  DLH_X2 \P_reg[3]  ( .G(n49), .D(N473), .Q(P[3]) );
  DLH_X2 \P_reg[4]  ( .G(n49), .D(N472), .Q(P[4]) );
  DLH_X2 \P_reg[5]  ( .G(n49), .D(N471), .Q(P[5]) );
  DLH_X2 \P_reg[6]  ( .G(n49), .D(N470), .Q(P[6]) );
  DLH_X2 \P_reg[7]  ( .G(n49), .D(N469), .Q(P[7]) );
  DLH_X2 \P_reg[8]  ( .G(n49), .D(N468), .Q(P[8]) );
  DLH_X2 \P_reg[9]  ( .G(n49), .D(N467), .Q(P[9]) );
  DLH_X2 \P_reg[10]  ( .G(n49), .D(N466), .Q(P[10]) );
  DLH_X2 \P_reg[11]  ( .G(n50), .D(N465), .Q(P[11]) );
  DLH_X2 \P_reg[12]  ( .G(n50), .D(N464), .Q(P[12]) );
  DLH_X2 \P_reg[13]  ( .G(n50), .D(N463), .Q(P[13]) );
  DLH_X2 \P_reg[14]  ( .G(n50), .D(N462), .Q(P[14]) );
  DLH_X2 \P_reg[15]  ( .G(n50), .D(N461), .Q(P[15]) );
  DLH_X2 \P_reg[16]  ( .G(n50), .D(N460), .Q(P[16]) );
  DLH_X2 \P_reg[17]  ( .G(n50), .D(N459), .Q(P[17]) );
  DLH_X2 \P_reg[18]  ( .G(n50), .D(N458), .Q(P[18]) );
  DLH_X2 \P_reg[19]  ( .G(n50), .D(N457), .Q(P[19]) );
  DLH_X2 \P_reg[20]  ( .G(n50), .D(N456), .Q(P[20]) );
  DLH_X2 \P_reg[21]  ( .G(n50), .D(N455), .Q(P[21]) );
  DLH_X2 \P_reg[22]  ( .G(N444), .D(N454), .Q(P[22]) );
  DLH_X2 \P_reg[23]  ( .G(n50), .D(N453), .Q(P[23]) );
  DLH_X2 \P_reg[24]  ( .G(n49), .D(N452), .Q(P[24]) );
  DLH_X2 \P_reg[25]  ( .G(N444), .D(N451), .Q(P[25]) );
  DLH_X2 \P_reg[26]  ( .G(n50), .D(N450), .Q(P[26]) );
  DLH_X2 \P_reg[27]  ( .G(n49), .D(N449), .Q(P[27]) );
  DLH_X2 \P_reg[28]  ( .G(N444), .D(N448), .Q(P[28]) );
  DLH_X2 \P_reg[29]  ( .G(N444), .D(N447), .Q(P[29]) );
  DLH_X2 \P_reg[30]  ( .G(N444), .D(N446), .Q(P[30]) );
  DLH_X2 \P_reg[31]  ( .G(N444), .D(N445), .Q(P[31]) );
  DLH_X2 \P1_reg[15]  ( .G(N43), .D(N104), .Q(P1[15]) );
  DLH_X2 \P1_reg[16]  ( .G(N43), .D(N103), .Q(P1[16]) );
  DLH_X2 \P1_reg[17]  ( .G(N43), .D(N102), .Q(P1[17]) );
  DLH_X2 \P1_reg[18]  ( .G(N43), .D(N101), .Q(P1[18]) );
  DLH_X2 \P1_reg[19]  ( .G(N43), .D(N100), .Q(P1[19]) );
  DLH_X2 \P1_reg[20]  ( .G(N43), .D(N99), .Q(P1[20]) );
  DLH_X2 \P1_reg[21]  ( .G(N43), .D(N98), .Q(P1[21]) );
  DLH_X2 \P1_reg[22]  ( .G(N43), .D(N97), .Q(P1[22]) );
  DLH_X2 \P1_reg[23]  ( .G(N43), .D(N96), .Q(P1[23]) );
  DLH_X2 \P1_reg[24]  ( .G(N43), .D(N95), .Q(P1[24]) );
  DLH_X2 \P1_reg[25]  ( .G(n58), .D(N94), .Q(P1[25]) );
  DLH_X2 \P1_reg[26]  ( .G(N43), .D(N93), .Q(P1[26]) );
  DLH_X2 \P1_reg[27]  ( .G(n58), .D(N92), .Q(P1[27]) );
  DLH_X2 \P1_reg[28]  ( .G(N43), .D(N91), .Q(P1[28]) );
  DLH_X2 \P1_reg[29]  ( .G(N43), .D(N90), .Q(P1[29]) );
  DLH_X2 \P1_reg[30]  ( .G(N43), .D(N89), .Q(P1[30]) );
  DLH_X2 \P1_reg[31]  ( .G(N43), .D(N88), .Q(P1[31]) );
  DLH_X2 working_reg ( .G(N477), .D(N478), .Q(working) );
  DLH_X2 \L_reg[0]  ( .G(n55), .D(N410), .Q(L[0]) );
  DLH_X2 \L_reg[1]  ( .G(n55), .D(N409), .Q(L[1]) );
  DLH_X2 \L_reg[2]  ( .G(n55), .D(N408), .Q(L[2]) );
  DLH_X2 \L_reg[3]  ( .G(n55), .D(N407), .Q(L[3]) );
  DLH_X2 \L_reg[4]  ( .G(n55), .D(N406), .Q(L[4]) );
  DLH_X2 \L_reg[5]  ( .G(n55), .D(N405), .Q(L[5]) );
  DLH_X2 \L_reg[6]  ( .G(n55), .D(N404), .Q(L[6]) );
  DLH_X2 \L_reg[7]  ( .G(n55), .D(N403), .Q(L[7]) );
  DLH_X2 \L_reg[8]  ( .G(n55), .D(N402), .Q(L[8]) );
  DLH_X2 \L_reg[9]  ( .G(n55), .D(N401), .Q(L[9]) );
  DLH_X2 \L_reg[10]  ( .G(n55), .D(N400), .Q(L[10]) );
  DLH_X2 \L_reg[11]  ( .G(n56), .D(N399), .Q(L[11]) );
  DLH_X2 \L_reg[12]  ( .G(n56), .D(N398), .Q(L[12]) );
  DLH_X2 \L_reg[13]  ( .G(n56), .D(N397), .Q(L[13]) );
  DLH_X2 \L_reg[14]  ( .G(n56), .D(N396), .Q(L[14]) );
  DLH_X2 \L_reg[15]  ( .G(n56), .D(N395), .Q(L[15]) );
  DLH_X2 \L_reg[16]  ( .G(n56), .D(N394), .Q(L[16]) );
  DLH_X2 \L_reg[17]  ( .G(n56), .D(N393), .Q(L[17]) );
  DLH_X2 \L_reg[18]  ( .G(n56), .D(N392), .Q(L[18]) );
  DLH_X2 \L_reg[19]  ( .G(n56), .D(N391), .Q(L[19]) );
  DLH_X2 \L_reg[20]  ( .G(n56), .D(N390), .Q(L[20]) );
  DLH_X2 \L_reg[21]  ( .G(n56), .D(N389), .Q(L[21]) );
  DLH_X2 \L_reg[22]  ( .G(N378), .D(N388), .Q(L[22]) );
  DLH_X2 \L_reg[23]  ( .G(n56), .D(N387), .Q(L[23]) );
  DLH_X2 \L_reg[24]  ( .G(n55), .D(N386), .Q(L[24]) );
  DLH_X2 \L_reg[25]  ( .G(N378), .D(N385), .Q(L[25]) );
  DLH_X2 \L_reg[26]  ( .G(n56), .D(N384), .Q(L[26]) );
  DLH_X2 \L_reg[27]  ( .G(n55), .D(N383), .Q(L[27]) );
  DLH_X2 \L_reg[28]  ( .G(N378), .D(N382), .Q(L[28]) );
  DLH_X2 \L_reg[29]  ( .G(N378), .D(N381), .Q(L[29]) );
  DLH_X2 \L_reg[30]  ( .G(N378), .D(N380), .Q(L[30]) );
  DLH_X2 \L_reg[31]  ( .G(N378), .D(N379), .Q(L[31]) );
  DLH_X2 \Z_reg[0]  ( .G(n52), .D(N443), .Q(Z[0]) );
  DLH_X2 \Z_reg[1]  ( .G(n52), .D(N442), .Q(Z[1]) );
  DLH_X2 \Z_reg[2]  ( .G(n52), .D(N441), .Q(Z[2]) );
  DLH_X2 \Z_reg[3]  ( .G(n52), .D(N440), .Q(Z[3]) );
  DLH_X2 \Z_reg[4]  ( .G(n52), .D(N439), .Q(Z[4]) );
  DLH_X2 \Z_reg[5]  ( .G(n52), .D(N438), .Q(Z[5]) );
  DLH_X2 \Z_reg[6]  ( .G(n52), .D(N437), .Q(Z[6]) );
  DLH_X2 \Z_reg[7]  ( .G(n52), .D(N436), .Q(Z[7]) );
  DLH_X2 \Z_reg[8]  ( .G(n52), .D(N435), .Q(Z[8]) );
  DLH_X2 \Z_reg[9]  ( .G(n52), .D(N434), .Q(Z[9]) );
  DLH_X2 \Z_reg[10]  ( .G(n52), .D(N433), .Q(Z[10]) );
  DLH_X2 \Z_reg[11]  ( .G(n53), .D(N432), .Q(Z[11]) );
  DLH_X2 \Z_reg[12]  ( .G(n53), .D(N431), .Q(Z[12]) );
  DLH_X2 \Z_reg[13]  ( .G(n53), .D(N430), .Q(Z[13]) );
  DLH_X2 \Z_reg[14]  ( .G(n53), .D(N429), .Q(Z[14]) );
  DLH_X2 \Z_reg[15]  ( .G(n53), .D(N428), .Q(Z[15]) );
  DLH_X2 \Z_reg[16]  ( .G(n53), .D(N427), .Q(Z[16]) );
  DLH_X2 \Z_reg[17]  ( .G(n53), .D(N426), .Q(Z[17]) );
  DLH_X2 \Z_reg[18]  ( .G(n53), .D(N425), .Q(Z[18]) );
  DLH_X2 \Z_reg[19]  ( .G(n53), .D(N424), .Q(Z[19]) );
  DLH_X2 \Z_reg[20]  ( .G(n53), .D(N423), .Q(Z[20]) );
  DLH_X2 \Z_reg[21]  ( .G(n53), .D(N422), .Q(Z[21]) );
  DLH_X2 \Z_reg[22]  ( .G(N411), .D(N421), .Q(Z[22]) );
  DLH_X2 \Z_reg[23]  ( .G(N411), .D(N420), .Q(Z[23]) );
  DLH_X2 \Z_reg[24]  ( .G(N411), .D(N419), .Q(Z[24]) );
  DLH_X2 \Z_reg[25]  ( .G(N411), .D(N418), .Q(Z[25]) );
  DLH_X2 \Z_reg[26]  ( .G(n53), .D(N417), .Q(Z[26]) );
  DLH_X2 \Z_reg[27]  ( .G(n52), .D(N416), .Q(Z[27]) );
  DLH_X2 \Z_reg[28]  ( .G(n52), .D(N415), .Q(Z[28]) );
  DLH_X2 \Z_reg[29]  ( .G(N411), .D(N414), .Q(Z[29]) );
  DLH_X2 \Z_reg[30]  ( .G(n53), .D(N413), .Q(Z[30]) );
  DLH_X2 \Z_reg[31]  ( .G(N411), .D(N412), .Q(Z[31]) );
  DLH_X2 \result_reg[0]  ( .G(n37), .D(N377), .Q(result[0]) );
  DLH_X2 \result_reg[1]  ( .G(n47), .D(N376), .Q(result[1]) );
  DLH_X2 \result_reg[2]  ( .G(n46), .D(N375), .Q(result[2]) );
  DLH_X2 \result_reg[3]  ( .G(n37), .D(N374), .Q(result[3]) );
  DLH_X2 \result_reg[4]  ( .G(n47), .D(N373), .Q(result[4]) );
  DLH_X2 \result_reg[5]  ( .G(n46), .D(N372), .Q(result[5]) );
  DLH_X2 \result_reg[6]  ( .G(n37), .D(N371), .Q(result[6]) );
  DLH_X2 \result_reg[7]  ( .G(n47), .D(N370), .Q(result[7]) );
  DLH_X2 \result_reg[8]  ( .G(n46), .D(N369), .Q(result[8]) );
  DLH_X2 \result_reg[9]  ( .G(n37), .D(N368), .Q(result[9]) );
  DLH_X2 \result_reg[10]  ( .G(n47), .D(N367), .Q(result[10]) );
  DLH_X2 \result_reg[11]  ( .G(n46), .D(N366), .Q(result[11]) );
  DLH_X2 \result_reg[12]  ( .G(n37), .D(N365), .Q(result[12]) );
  DLH_X2 \result_reg[13]  ( .G(n47), .D(N364), .Q(result[13]) );
  DLH_X2 \result_reg[14]  ( .G(n46), .D(N363), .Q(result[14]) );
  DLH_X2 \result_reg[15]  ( .G(n37), .D(N362), .Q(result[15]) );
  DLH_X2 \result_reg[16]  ( .G(n47), .D(N361), .Q(result[16]) );
  DLH_X2 \result_reg[17]  ( .G(n47), .D(N360), .Q(result[17]) );
  DLH_X2 \result_reg[18]  ( .G(n47), .D(N359), .Q(result[18]) );
  DLH_X2 \result_reg[19]  ( .G(n47), .D(N358), .Q(result[19]) );
  DLH_X2 \result_reg[20]  ( .G(n47), .D(N357), .Q(result[20]) );
  DLH_X2 \result_reg[21]  ( .G(n47), .D(N356), .Q(result[21]) );
  DLH_X2 \result_reg[22]  ( .G(n47), .D(N355), .Q(result[22]) );
  DLH_X2 \result_reg[23]  ( .G(n47), .D(N354), .Q(result[23]) );
  DLH_X2 \result_reg[24]  ( .G(n47), .D(N353), .Q(result[24]) );
  DLH_X2 \result_reg[25]  ( .G(n47), .D(N352), .Q(result[25]) );
  DLH_X2 \result_reg[26]  ( .G(n47), .D(N351), .Q(result[26]) );
  DLH_X2 \result_reg[27]  ( .G(n47), .D(N350), .Q(result[27]) );
  DLH_X2 \result_reg[28]  ( .G(n47), .D(N349), .Q(result[28]) );
  DLH_X2 \result_reg[29]  ( .G(n47), .D(N348), .Q(result[29]) );
  DLH_X2 \result_reg[30]  ( .G(n47), .D(N347), .Q(result[30]) );
  DLH_X2 \result_reg[31]  ( .G(n47), .D(N346), .Q(result[31]) );
  DLH_X2 \result_reg[32]  ( .G(n47), .D(N345), .Q(result[32]) );
  DLH_X2 \result_reg[33]  ( .G(n46), .D(N344), .Q(result[33]) );
  DLH_X2 \result_reg[34]  ( .G(n46), .D(N343), .Q(result[34]) );
  DLH_X2 \result_reg[35]  ( .G(n46), .D(N342), .Q(result[35]) );
  DLH_X2 \result_reg[36]  ( .G(n46), .D(N341), .Q(result[36]) );
  DLH_X2 \result_reg[37]  ( .G(n46), .D(N340), .Q(result[37]) );
  DLH_X2 \result_reg[38]  ( .G(n46), .D(N339), .Q(result[38]) );
  DLH_X2 \result_reg[39]  ( .G(n46), .D(N338), .Q(result[39]) );
  DLH_X2 \result_reg[40]  ( .G(n46), .D(N337), .Q(result[40]) );
  DLH_X2 \result_reg[41]  ( .G(n46), .D(N336), .Q(result[41]) );
  DLH_X2 \result_reg[42]  ( .G(n46), .D(N335), .Q(result[42]) );
  DLH_X2 \result_reg[43]  ( .G(n46), .D(N334), .Q(result[43]) );
  DLH_X2 \result_reg[44]  ( .G(n46), .D(N333), .Q(result[44]) );
  DLH_X2 \result_reg[45]  ( .G(n46), .D(N332), .Q(result[45]) );
  DLH_X2 \result_reg[46]  ( .G(n46), .D(N331), .Q(result[46]) );
  DLH_X2 \result_reg[47]  ( .G(n46), .D(N330), .Q(result[47]) );
  DLH_X2 \result_reg[48]  ( .G(n46), .D(N329), .Q(result[48]) );
  DLH_X2 \result_reg[49]  ( .G(n46), .D(N328), .Q(result[49]) );
  DLH_X2 \result_reg[50]  ( .G(n37), .D(N327), .Q(result[50]) );
  DLH_X2 \result_reg[51]  ( .G(n37), .D(N326), .Q(result[51]) );
  DLH_X2 \result_reg[52]  ( .G(n37), .D(N325), .Q(result[52]) );
  DLH_X2 \result_reg[53]  ( .G(n37), .D(N324), .Q(result[53]) );
  DLH_X2 \result_reg[54]  ( .G(n37), .D(N323), .Q(result[54]) );
  DLH_X2 \result_reg[55]  ( .G(n37), .D(N322), .Q(result[55]) );
  DLH_X2 \result_reg[56]  ( .G(n47), .D(N321), .Q(result[56]) );
  DLH_X2 \result_reg[57]  ( .G(n37), .D(N320), .Q(result[57]) );
  DLH_X2 \result_reg[58]  ( .G(n37), .D(N319), .Q(result[58]) );
  DLH_X2 \result_reg[59]  ( .G(n46), .D(N318), .Q(result[59]) );
  DLH_X2 \result_reg[60]  ( .G(n37), .D(N317), .Q(result[60]) );
  DLH_X2 \result_reg[61]  ( .G(n37), .D(N316), .Q(result[61]) );
  DLH_X2 \result_reg[62]  ( .G(n46), .D(N315), .Q(result[62]) );
  DLH_X2 \result_reg[63]  ( .G(n47), .D(N314), .Q(result[63]) );
  DLH_X2 \H_reg[0]  ( .G(N43), .D(N87), .Q(H[0]) );
  DLH_X2 \H_reg[1]  ( .G(N43), .D(N86), .Q(H[1]) );
  DLH_X2 \H_reg[2]  ( .G(n58), .D(N85), .Q(H[2]) );
  DLH_X2 \H_reg[3]  ( .G(N43), .D(N84), .Q(H[3]) );
  DLH_X2 \H_reg[4]  ( .G(n58), .D(N83), .Q(H[4]) );
  DLH_X2 \H_reg[5]  ( .G(N43), .D(N82), .Q(H[5]) );
  DLH_X2 \H_reg[6]  ( .G(n58), .D(N81), .Q(H[6]) );
  DLH_X2 \H_reg[7]  ( .G(N43), .D(N80), .Q(H[7]) );
  DLH_X2 \H_reg[8]  ( .G(n58), .D(N79), .Q(H[8]) );
  DLH_X2 \H_reg[9]  ( .G(N43), .D(N78), .Q(H[9]) );
  DLH_X2 \H_reg[10]  ( .G(n58), .D(N77), .Q(H[10]) );
  DLH_X2 \H_reg[11]  ( .G(N43), .D(N76), .Q(H[11]) );
  DLH_X2 \H_reg[12]  ( .G(n58), .D(N75), .Q(H[12]) );
  DLH_X2 \H_reg[13]  ( .G(N43), .D(N74), .Q(H[13]) );
  DLH_X2 \H_reg[14]  ( .G(n58), .D(N73), .Q(H[14]) );
  DLH_X2 \H_reg[15]  ( .G(n58), .D(N72), .Q(H[15]) );
  DLH_X2 \H_reg[16]  ( .G(n58), .D(N71), .Q(H[16]) );
  DLH_X2 \H_reg[17]  ( .G(N43), .D(N70), .Q(H[17]) );
  DLH_X2 \H_reg[18]  ( .G(n58), .D(N69), .Q(H[18]) );
  DLH_X2 \H_reg[19]  ( .G(n58), .D(N68), .Q(H[19]) );
  DLH_X2 \H_reg[20]  ( .G(n58), .D(N67), .Q(H[20]) );
  DLH_X2 \H_reg[21]  ( .G(n58), .D(N66), .Q(H[21]) );
  DLH_X2 \H_reg[22]  ( .G(n58), .D(N65), .Q(H[22]) );
  DLH_X2 \H_reg[23]  ( .G(n58), .D(N64), .Q(H[23]) );
  DLH_X2 \H_reg[24]  ( .G(n58), .D(N63), .Q(H[24]) );
  DLH_X2 \H_reg[25]  ( .G(n58), .D(N62), .Q(H[25]) );
  DLH_X2 \H_reg[26]  ( .G(n58), .D(N61), .Q(H[26]) );
  DLH_X2 \H_reg[27]  ( .G(n58), .D(N60), .Q(H[27]) );
  DLH_X2 \H_reg[28]  ( .G(n58), .D(N59), .Q(H[28]) );
  DLH_X2 \H_reg[29]  ( .G(n58), .D(N58), .Q(H[29]) );
  DLH_X2 \H_reg[30]  ( .G(n58), .D(N57), .Q(H[30]) );
  DLH_X2 \H_reg[31]  ( .G(n58), .D(N56), .Q(H[31]) );
  NOR2_X2 U125 ( .A1(n37), .A2(n58), .ZN(n32) );
  NOR2_X2 U126 ( .A1(n45), .A2(n40), .ZN(n34) );
  NAND3_X2 U127 ( .A1(n33), .A2(n32), .A3(n34), .ZN(N477) );
  NOR2_X2 U128 ( .A1(n34), .A2(n62), .ZN(N15) );
  NOR2_X2 U129 ( .A1(n33), .A2(n62), .ZN(N16) );
  AOI21_X2 U130 ( .B1(n35), .B2(n36), .A(n62), .ZN(N14) );
  NAND3_X2 U131 ( .A1(n39), .A2(n65), .A3(mul), .ZN(n36) );
  INV_X4 U132 ( .A(n38), .ZN(n44) );
  INV_X4 U133 ( .A(n44), .ZN(n45) );
  NOR3_X2 U134 ( .A1(CurrentState[0]), .A2(CurrentState[1]), .A3(n65), .ZN(n38) );
  INV_X4 U135 ( .A(N43), .ZN(n59) );
  INV_X4 U136 ( .A(n37), .ZN(n48) );
  INV_X4 U137 ( .A(n59), .ZN(n58) );
  INV_X4 U138 ( .A(n44), .ZN(n43) );
  NAND3_X2 U139 ( .A1(n39), .A2(n65), .A3(CurrentState[1]), .ZN(n35) );
  INV_X4 U140 ( .A(n48), .ZN(n46) );
  INV_X4 U141 ( .A(n48), .ZN(n47) );
  NAND3_X2 U142 ( .A1(CurrentState[2]), .A2(n39), .A3(CurrentState[1]), .ZN(
        n33) );
  INV_X4 U143 ( .A(N378), .ZN(n57) );
  INV_X4 U144 ( .A(n57), .ZN(n55) );
  INV_X4 U145 ( .A(n57), .ZN(n56) );
  NOR3_X2 U146 ( .A1(CurrentState[1]), .A2(CurrentState[2]), .A3(n39), .ZN(n37) );
  INV_X4 U147 ( .A(N411), .ZN(n54) );
  INV_X4 U148 ( .A(n54), .ZN(n52) );
  INV_X4 U149 ( .A(n54), .ZN(n53) );
  INV_X4 U150 ( .A(N444), .ZN(n51) );
  INV_X4 U151 ( .A(n51), .ZN(n49) );
  INV_X4 U152 ( .A(n51), .ZN(n50) );
  INV_X4 U153 ( .A(n33), .ZN(n41) );
  INV_X4 U154 ( .A(n33), .ZN(n42) );
  INV_X4 U155 ( .A(n35), .ZN(n40) );
  NOR3_X2 U156 ( .A1(CurrentState[1]), .A2(CurrentState[2]), .A3(
        CurrentState[0]), .ZN(N43) );
  INV_X4 U187 ( .A(reset), .ZN(n62) );
  INV_X4 U188 ( .A(mul), .ZN(n63) );
  INV_X4 U189 ( .A(n35), .ZN(n64) );
  INV_X4 U191 ( .A(n33), .ZN(n66) );
  INV_X4 U192 ( .A(n32), .ZN(n67) );
  multiplier_DW01_add_0 add_85 ( .A({1'b0, b[0:15]}), .B({1'b0, b[16:31]}), 
        .CI(1'b0), .SUM({N121, N120, N119, N118, N117, N116, N115, N114, N113, 
        N112, N111, N110, N109, N108, N107, N106, N105}) );
  multiplier_DW01_add_1 add_77 ( .A({1'b0, a[0:15]}), .B({1'b0, a[16:31]}), 
        .CI(1'b0), .SUM({N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, 
        N94, N93, N92, N91, N90, N89, N88}) );
  multiplier_DW01_add_5 add_1_root_add_0_root_add_98_2 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, L}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, Z, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, N298, N297, N296, 
        N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, 
        N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, 
        N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, 
        N259, N258, N257, N256, N255, N254, N253, N252, N251, N250}) );
  multiplier_DW01_add_4 add_0_root_add_0_root_add_98_2 ( .A({Z, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N298, N297, 
        N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, 
        N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, 
        N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, 
        N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250}), 
        .CI(1'b0), .SUM({N377, N376, N375, N374, N373, N372, N371, N370, N369, 
        N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, 
        N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, 
        N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, 
        N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, 
        N320, N319, N318, N317, N316, N315, N314}) );
  multiplier_DW01_sub_1 sub_1_root_sub_0_root_sub_94_2 ( .A(P), .B(L), .CI(
        1'b0), .DIFF({N217, N216, N215, N214, N213, N212, N211, N210, N209, 
        N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, 
        N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186}) );
  multiplier_DW01_sub_0 sub_0_root_sub_0_root_sub_94_2 ( .A({N217, N216, N215, 
        N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, 
        N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, 
        N190, N189, N188, N187, N186}), .B(H), .CI(1'b0), .DIFF({N249, N248, 
        N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, 
        N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, 
        N223, N222, N221, N220, N219, N218}) );
  multiplier_DW02_mult_2 mult_90 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, P1[15:31]}), .B(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, P2[15:31]}), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, N185, N184, N183, 
        N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, 
        N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, 
        N158, N157, N156, N155, N154}) );
  multiplier_DW02_mult_0 mult_76 ( .A(a[0:15]), .B(b[0:15]), .TC(1'b0), 
        .PRODUCT({N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, 
        N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, 
        N61, N60, N59, N58, N57, N56}) );
  multiplier_DW02_mult_1 mult_86 ( .A(a[16:31]), .B(b[16:31]), .TC(1'b0), 
        .PRODUCT({N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, 
        N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, 
        N131, N130, N129, N128, N127, N126, N125, N124, N123, N122}) );
  DFF_X1 \CurrentState_reg[1]  ( .D(N15), .CK(clk), .Q(CurrentState[1]) );
  DFF_X1 \CurrentState_reg[2]  ( .D(N14), .CK(clk), .Q(CurrentState[2]), .QN(
        n65) );
endmodule

