module register1(inData, clk, writeEnable, outData);
    
    input inData, clk, writeEnable;
    output outData;
    
    

endmodule