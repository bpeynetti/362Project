
module id_ex_reg ( in, flush, out, clk, reset, we );
  input [0:276] in;
  output [0:276] out;
  input flush, clk, reset, we;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623;

  DFFR_X1 ID_EX_REG_out_reg_276_ ( .D(n555), .CK(clk), .RN(reset), .Q(out[276]) );
  DFFR_X1 ID_EX_REG_out_reg_275_ ( .D(n554), .CK(clk), .RN(n620), .Q(out[275])
         );
  DFFR_X1 ID_EX_REG_out_reg_274_ ( .D(n553), .CK(clk), .RN(n623), .Q(out[274])
         );
  DFFR_X1 ID_EX_REG_out_reg_273_ ( .D(n552), .CK(clk), .RN(n620), .Q(out[273])
         );
  DFFR_X1 ID_EX_REG_out_reg_272_ ( .D(n551), .CK(clk), .RN(n622), .Q(out[272])
         );
  DFFR_X1 ID_EX_REG_out_reg_271_ ( .D(n550), .CK(clk), .RN(n620), .Q(out[271])
         );
  DFFR_X1 ID_EX_REG_out_reg_270_ ( .D(n549), .CK(clk), .RN(n621), .Q(out[270])
         );
  DFFR_X1 ID_EX_REG_out_reg_269_ ( .D(n548), .CK(clk), .RN(n620), .Q(out[269])
         );
  DFFR_X1 ID_EX_REG_out_reg_268_ ( .D(n547), .CK(clk), .RN(n620), .Q(out[268])
         );
  DFFR_X1 ID_EX_REG_out_reg_267_ ( .D(n546), .CK(clk), .RN(reset), .Q(out[267]) );
  DFFR_X1 ID_EX_REG_out_reg_266_ ( .D(n545), .CK(clk), .RN(n620), .Q(out[266])
         );
  DFFR_X1 ID_EX_REG_out_reg_265_ ( .D(n544), .CK(clk), .RN(n619), .Q(out[265])
         );
  DFFR_X1 ID_EX_REG_out_reg_264_ ( .D(n543), .CK(clk), .RN(n620), .Q(out[264])
         );
  DFFR_X1 ID_EX_REG_out_reg_263_ ( .D(n542), .CK(clk), .RN(n618), .Q(out[263])
         );
  DFFR_X1 ID_EX_REG_out_reg_262_ ( .D(n541), .CK(clk), .RN(n620), .Q(out[262])
         );
  DFFR_X1 ID_EX_REG_out_reg_261_ ( .D(n540), .CK(clk), .RN(n613), .Q(out[261])
         );
  DFFR_X1 ID_EX_REG_out_reg_260_ ( .D(n539), .CK(clk), .RN(n611), .Q(out[260])
         );
  DFFR_X1 ID_EX_REG_out_reg_259_ ( .D(n538), .CK(clk), .RN(n612), .Q(out[259])
         );
  DFFR_X1 ID_EX_REG_out_reg_258_ ( .D(n537), .CK(clk), .RN(n612), .Q(out[258])
         );
  DFFR_X1 ID_EX_REG_out_reg_257_ ( .D(n536), .CK(clk), .RN(n613), .Q(out[257])
         );
  DFFR_X1 ID_EX_REG_out_reg_256_ ( .D(n535), .CK(clk), .RN(n611), .Q(out[256])
         );
  DFFR_X1 ID_EX_REG_out_reg_255_ ( .D(n534), .CK(clk), .RN(n621), .Q(out[255])
         );
  DFFR_X1 ID_EX_REG_out_reg_254_ ( .D(n533), .CK(clk), .RN(n610), .Q(out[254])
         );
  DFFR_X1 ID_EX_REG_out_reg_253_ ( .D(n532), .CK(clk), .RN(n622), .Q(out[253])
         );
  DFFR_X1 ID_EX_REG_out_reg_252_ ( .D(n531), .CK(clk), .RN(n609), .Q(out[252])
         );
  DFFR_X1 ID_EX_REG_out_reg_251_ ( .D(n530), .CK(clk), .RN(n623), .Q(out[251])
         );
  DFFR_X1 ID_EX_REG_out_reg_250_ ( .D(n529), .CK(clk), .RN(n608), .Q(out[250])
         );
  DFFR_X1 ID_EX_REG_out_reg_249_ ( .D(n528), .CK(clk), .RN(n610), .Q(out[249])
         );
  DFFR_X1 ID_EX_REG_out_reg_248_ ( .D(n527), .CK(clk), .RN(n619), .Q(out[248])
         );
  DFFR_X1 ID_EX_REG_out_reg_247_ ( .D(n526), .CK(clk), .RN(n607), .Q(out[247])
         );
  DFFR_X1 ID_EX_REG_out_reg_246_ ( .D(n525), .CK(clk), .RN(n618), .Q(out[246])
         );
  DFFR_X1 ID_EX_REG_out_reg_245_ ( .D(n524), .CK(clk), .RN(n606), .Q(out[245])
         );
  DFFR_X1 ID_EX_REG_out_reg_244_ ( .D(n523), .CK(clk), .RN(n617), .Q(out[244])
         );
  DFFR_X1 ID_EX_REG_out_reg_243_ ( .D(n522), .CK(clk), .RN(n605), .Q(out[243])
         );
  DFFR_X1 ID_EX_REG_out_reg_242_ ( .D(n521), .CK(clk), .RN(n616), .Q(out[242])
         );
  DFFR_X1 ID_EX_REG_out_reg_241_ ( .D(n520), .CK(clk), .RN(reset), .Q(out[241]) );
  DFFR_X1 ID_EX_REG_out_reg_240_ ( .D(n519), .CK(clk), .RN(n615), .Q(out[240])
         );
  DFFR_X1 ID_EX_REG_out_reg_239_ ( .D(n518), .CK(clk), .RN(n619), .Q(out[239])
         );
  DFFR_X1 ID_EX_REG_out_reg_238_ ( .D(n517), .CK(clk), .RN(n609), .Q(out[238])
         );
  DFFR_X1 ID_EX_REG_out_reg_237_ ( .D(n516), .CK(clk), .RN(n619), .Q(out[237])
         );
  DFFR_X1 ID_EX_REG_out_reg_236_ ( .D(n515), .CK(clk), .RN(n608), .Q(out[236])
         );
  DFFR_X1 ID_EX_REG_out_reg_235_ ( .D(n514), .CK(clk), .RN(n619), .Q(out[235])
         );
  DFFR_X1 ID_EX_REG_out_reg_234_ ( .D(n513), .CK(clk), .RN(n607), .Q(out[234])
         );
  DFFR_X1 ID_EX_REG_out_reg_233_ ( .D(n512), .CK(clk), .RN(n619), .Q(out[233])
         );
  DFFR_X1 ID_EX_REG_out_reg_232_ ( .D(n511), .CK(clk), .RN(n606), .Q(out[232])
         );
  DFFR_X1 ID_EX_REG_out_reg_231_ ( .D(n510), .CK(clk), .RN(n619), .Q(out[231])
         );
  DFFR_X1 ID_EX_REG_out_reg_230_ ( .D(n509), .CK(clk), .RN(n605), .Q(out[230])
         );
  DFFR_X1 ID_EX_REG_out_reg_229_ ( .D(n508), .CK(clk), .RN(reset), .Q(out[229]) );
  DFFR_X1 ID_EX_REG_out_reg_228_ ( .D(n507), .CK(clk), .RN(n619), .Q(out[228])
         );
  DFFR_X1 ID_EX_REG_out_reg_227_ ( .D(n506), .CK(clk), .RN(n611), .Q(out[227])
         );
  DFFR_X1 ID_EX_REG_out_reg_226_ ( .D(n505), .CK(clk), .RN(n619), .Q(out[226])
         );
  DFFR_X1 ID_EX_REG_out_reg_225_ ( .D(n504), .CK(clk), .RN(n612), .Q(out[225])
         );
  DFFR_X1 ID_EX_REG_out_reg_224_ ( .D(n503), .CK(clk), .RN(n619), .Q(out[224])
         );
  DFFR_X1 ID_EX_REG_out_reg_223_ ( .D(n502), .CK(clk), .RN(n613), .Q(out[223])
         );
  DFFR_X1 ID_EX_REG_out_reg_222_ ( .D(n501), .CK(clk), .RN(n619), .Q(out[222])
         );
  DFFR_X1 ID_EX_REG_out_reg_221_ ( .D(n500), .CK(clk), .RN(n620), .Q(out[221])
         );
  DFFR_X1 ID_EX_REG_out_reg_220_ ( .D(n499), .CK(clk), .RN(n619), .Q(out[220])
         );
  DFFR_X1 ID_EX_REG_out_reg_219_ ( .D(n498), .CK(clk), .RN(n619), .Q(out[219])
         );
  DFFR_X1 ID_EX_REG_out_reg_218_ ( .D(n497), .CK(clk), .RN(n608), .Q(out[218])
         );
  DFFR_X1 ID_EX_REG_out_reg_217_ ( .D(n496), .CK(clk), .RN(n618), .Q(out[217])
         );
  DFFR_X1 ID_EX_REG_out_reg_216_ ( .D(n495), .CK(clk), .RN(n608), .Q(out[216])
         );
  DFFR_X1 ID_EX_REG_out_reg_215_ ( .D(n494), .CK(clk), .RN(n618), .Q(out[215])
         );
  DFFR_X1 ID_EX_REG_out_reg_214_ ( .D(n493), .CK(clk), .RN(n608), .Q(out[214])
         );
  DFFR_X1 ID_EX_REG_out_reg_213_ ( .D(n492), .CK(clk), .RN(n618), .Q(out[213])
         );
  DFFR_X1 ID_EX_REG_out_reg_212_ ( .D(n491), .CK(clk), .RN(n608), .Q(out[212])
         );
  DFFR_X1 ID_EX_REG_out_reg_211_ ( .D(n490), .CK(clk), .RN(n618), .Q(out[211])
         );
  DFFR_X1 ID_EX_REG_out_reg_210_ ( .D(n489), .CK(clk), .RN(n608), .Q(out[210])
         );
  DFFR_X1 ID_EX_REG_out_reg_209_ ( .D(n488), .CK(clk), .RN(n608), .Q(out[209])
         );
  DFFR_X1 ID_EX_REG_out_reg_208_ ( .D(n487), .CK(clk), .RN(n618), .Q(out[208])
         );
  DFFR_X1 ID_EX_REG_out_reg_207_ ( .D(n486), .CK(clk), .RN(n608), .Q(out[207])
         );
  DFFR_X1 ID_EX_REG_out_reg_206_ ( .D(n485), .CK(clk), .RN(n618), .Q(out[206])
         );
  DFFR_X1 ID_EX_REG_out_reg_205_ ( .D(n484), .CK(clk), .RN(n608), .Q(out[205])
         );
  DFFR_X1 ID_EX_REG_out_reg_204_ ( .D(n483), .CK(clk), .RN(n618), .Q(out[204])
         );
  DFFR_X1 ID_EX_REG_out_reg_203_ ( .D(n482), .CK(clk), .RN(n608), .Q(out[203])
         );
  DFFR_X1 ID_EX_REG_out_reg_202_ ( .D(n481), .CK(clk), .RN(n618), .Q(out[202])
         );
  DFFR_X1 ID_EX_REG_out_reg_201_ ( .D(n480), .CK(clk), .RN(n608), .Q(out[201])
         );
  DFFR_X1 ID_EX_REG_out_reg_200_ ( .D(n479), .CK(clk), .RN(n618), .Q(out[200])
         );
  DFFR_X1 ID_EX_REG_out_reg_199_ ( .D(n478), .CK(clk), .RN(n608), .Q(out[199])
         );
  DFFR_X1 ID_EX_REG_out_reg_198_ ( .D(n477), .CK(clk), .RN(n618), .Q(out[198])
         );
  DFFR_X1 ID_EX_REG_out_reg_197_ ( .D(n476), .CK(clk), .RN(n609), .Q(out[197])
         );
  DFFR_X1 ID_EX_REG_out_reg_196_ ( .D(n475), .CK(clk), .RN(n617), .Q(out[196])
         );
  DFFR_X1 ID_EX_REG_out_reg_195_ ( .D(n474), .CK(clk), .RN(n609), .Q(out[195])
         );
  DFFR_X1 ID_EX_REG_out_reg_194_ ( .D(n473), .CK(clk), .RN(n617), .Q(out[194])
         );
  DFFR_X1 ID_EX_REG_out_reg_193_ ( .D(n472), .CK(clk), .RN(n609), .Q(out[193])
         );
  DFFR_X1 ID_EX_REG_out_reg_192_ ( .D(n471), .CK(clk), .RN(n617), .Q(out[192])
         );
  DFFR_X1 ID_EX_REG_out_reg_191_ ( .D(n470), .CK(clk), .RN(n609), .Q(out[191])
         );
  DFFR_X1 ID_EX_REG_out_reg_190_ ( .D(n469), .CK(clk), .RN(n617), .Q(out[190])
         );
  DFFR_X1 ID_EX_REG_out_reg_189_ ( .D(n468), .CK(clk), .RN(n617), .Q(out[189])
         );
  DFFR_X1 ID_EX_REG_out_reg_188_ ( .D(n467), .CK(clk), .RN(n609), .Q(out[188])
         );
  DFFR_X1 ID_EX_REG_out_reg_187_ ( .D(n466), .CK(clk), .RN(n617), .Q(out[187])
         );
  DFFR_X1 ID_EX_REG_out_reg_186_ ( .D(n465), .CK(clk), .RN(n609), .Q(out[186])
         );
  DFFR_X1 ID_EX_REG_out_reg_185_ ( .D(n464), .CK(clk), .RN(n617), .Q(out[185])
         );
  DFFR_X1 ID_EX_REG_out_reg_184_ ( .D(n463), .CK(clk), .RN(n609), .Q(out[184])
         );
  DFFR_X1 ID_EX_REG_out_reg_183_ ( .D(n462), .CK(clk), .RN(n617), .Q(out[183])
         );
  DFFR_X1 ID_EX_REG_out_reg_182_ ( .D(n461), .CK(clk), .RN(n609), .Q(out[182])
         );
  DFFR_X1 ID_EX_REG_out_reg_181_ ( .D(n460), .CK(clk), .RN(n617), .Q(out[181])
         );
  DFFR_X1 ID_EX_REG_out_reg_180_ ( .D(n459), .CK(clk), .RN(n609), .Q(out[180])
         );
  DFFR_X1 ID_EX_REG_out_reg_179_ ( .D(n458), .CK(clk), .RN(n609), .Q(out[179])
         );
  DFFR_X1 ID_EX_REG_out_reg_178_ ( .D(n457), .CK(clk), .RN(n617), .Q(out[178])
         );
  DFFR_X1 ID_EX_REG_out_reg_177_ ( .D(n456), .CK(clk), .RN(n609), .Q(out[177])
         );
  DFFR_X1 ID_EX_REG_out_reg_176_ ( .D(n455), .CK(clk), .RN(n617), .Q(out[176])
         );
  DFFR_X1 ID_EX_REG_out_reg_175_ ( .D(n454), .CK(clk), .RN(n610), .Q(out[175])
         );
  DFFR_X1 ID_EX_REG_out_reg_174_ ( .D(n453), .CK(clk), .RN(n616), .Q(out[174])
         );
  DFFR_X1 ID_EX_REG_out_reg_173_ ( .D(n452), .CK(clk), .RN(n610), .Q(out[173])
         );
  DFFR_X1 ID_EX_REG_out_reg_172_ ( .D(n451), .CK(clk), .RN(n616), .Q(out[172])
         );
  DFFR_X1 ID_EX_REG_out_reg_171_ ( .D(n450), .CK(clk), .RN(n610), .Q(out[171])
         );
  DFFR_X1 ID_EX_REG_out_reg_170_ ( .D(n449), .CK(clk), .RN(n616), .Q(out[170])
         );
  DFFR_X1 ID_EX_REG_out_reg_169_ ( .D(n448), .CK(clk), .RN(n616), .Q(out[169])
         );
  DFFR_X1 ID_EX_REG_out_reg_168_ ( .D(n447), .CK(clk), .RN(n610), .Q(out[168])
         );
  DFFR_X1 ID_EX_REG_out_reg_167_ ( .D(n446), .CK(clk), .RN(n616), .Q(out[167])
         );
  DFFR_X1 ID_EX_REG_out_reg_166_ ( .D(n445), .CK(clk), .RN(n610), .Q(out[166])
         );
  DFFR_X1 ID_EX_REG_out_reg_165_ ( .D(n444), .CK(clk), .RN(n616), .Q(out[165])
         );
  DFFR_X1 ID_EX_REG_out_reg_164_ ( .D(n443), .CK(clk), .RN(n610), .Q(out[164])
         );
  DFFR_X1 ID_EX_REG_out_reg_163_ ( .D(n442), .CK(clk), .RN(n616), .Q(out[163])
         );
  DFFR_X1 ID_EX_REG_out_reg_162_ ( .D(n441), .CK(clk), .RN(n610), .Q(out[162])
         );
  DFFR_X1 ID_EX_REG_out_reg_161_ ( .D(n440), .CK(clk), .RN(n616), .Q(out[161])
         );
  DFFR_X1 ID_EX_REG_out_reg_160_ ( .D(n439), .CK(clk), .RN(n610), .Q(out[160])
         );
  DFFR_X1 ID_EX_REG_out_reg_159_ ( .D(n438), .CK(clk), .RN(n610), .Q(out[159])
         );
  DFFR_X1 ID_EX_REG_out_reg_158_ ( .D(n437), .CK(clk), .RN(n616), .Q(out[158])
         );
  DFFR_X1 ID_EX_REG_out_reg_157_ ( .D(n436), .CK(clk), .RN(n610), .Q(out[157])
         );
  DFFR_X1 ID_EX_REG_out_reg_156_ ( .D(n435), .CK(clk), .RN(n616), .Q(out[156])
         );
  DFFR_X1 ID_EX_REG_out_reg_155_ ( .D(n434), .CK(clk), .RN(n610), .Q(out[155])
         );
  DFFR_X1 ID_EX_REG_out_reg_154_ ( .D(n433), .CK(clk), .RN(n616), .Q(out[154])
         );
  DFFR_X1 ID_EX_REG_out_reg_153_ ( .D(n432), .CK(clk), .RN(n611), .Q(out[153])
         );
  DFFR_X1 ID_EX_REG_out_reg_152_ ( .D(n431), .CK(clk), .RN(n615), .Q(out[152])
         );
  DFFR_X1 ID_EX_REG_out_reg_151_ ( .D(n430), .CK(clk), .RN(n611), .Q(out[151])
         );
  DFFR_X1 ID_EX_REG_out_reg_150_ ( .D(n429), .CK(clk), .RN(n615), .Q(out[150])
         );
  DFFR_X1 ID_EX_REG_out_reg_149_ ( .D(n428), .CK(clk), .RN(n615), .Q(out[149])
         );
  DFFR_X1 ID_EX_REG_out_reg_148_ ( .D(n427), .CK(clk), .RN(n611), .Q(out[148])
         );
  DFFR_X1 ID_EX_REG_out_reg_147_ ( .D(n426), .CK(clk), .RN(n615), .Q(out[147])
         );
  DFFR_X1 ID_EX_REG_out_reg_146_ ( .D(n425), .CK(clk), .RN(n611), .Q(out[146])
         );
  DFFR_X1 ID_EX_REG_out_reg_145_ ( .D(n424), .CK(clk), .RN(n615), .Q(out[145])
         );
  DFFR_X1 ID_EX_REG_out_reg_144_ ( .D(n423), .CK(clk), .RN(n611), .Q(out[144])
         );
  DFFR_X1 ID_EX_REG_out_reg_143_ ( .D(n422), .CK(clk), .RN(n615), .Q(out[143])
         );
  DFFR_X1 ID_EX_REG_out_reg_142_ ( .D(n421), .CK(clk), .RN(n611), .Q(out[142])
         );
  DFFR_X1 ID_EX_REG_out_reg_141_ ( .D(n420), .CK(clk), .RN(n615), .Q(out[141])
         );
  DFFR_X1 ID_EX_REG_out_reg_140_ ( .D(n419), .CK(clk), .RN(n611), .Q(out[140])
         );
  DFFR_X1 ID_EX_REG_out_reg_139_ ( .D(n418), .CK(clk), .RN(n611), .Q(out[139])
         );
  DFFR_X1 ID_EX_REG_out_reg_138_ ( .D(n417), .CK(clk), .RN(n615), .Q(out[138])
         );
  DFFR_X1 ID_EX_REG_out_reg_137_ ( .D(n416), .CK(clk), .RN(n611), .Q(out[137])
         );
  DFFR_X1 ID_EX_REG_out_reg_136_ ( .D(n415), .CK(clk), .RN(n615), .Q(out[136])
         );
  DFFR_X1 ID_EX_REG_out_reg_135_ ( .D(n414), .CK(clk), .RN(n611), .Q(out[135])
         );
  DFFR_X1 ID_EX_REG_out_reg_134_ ( .D(n413), .CK(clk), .RN(n615), .Q(out[134])
         );
  DFFR_X1 ID_EX_REG_out_reg_133_ ( .D(n412), .CK(clk), .RN(n611), .Q(out[133])
         );
  DFFR_X1 ID_EX_REG_out_reg_132_ ( .D(n411), .CK(clk), .RN(n615), .Q(out[132])
         );
  DFFR_X1 ID_EX_REG_out_reg_131_ ( .D(n410), .CK(clk), .RN(n612), .Q(out[131])
         );
  DFFR_X1 ID_EX_REG_out_reg_130_ ( .D(n409), .CK(clk), .RN(n614), .Q(out[130])
         );
  DFFR_X1 ID_EX_REG_out_reg_129_ ( .D(n408), .CK(clk), .RN(n614), .Q(out[129])
         );
  DFFR_X1 ID_EX_REG_out_reg_128_ ( .D(n407), .CK(clk), .RN(n612), .Q(out[128])
         );
  DFFR_X1 ID_EX_REG_out_reg_127_ ( .D(n406), .CK(clk), .RN(n614), .Q(out[127])
         );
  DFFR_X1 ID_EX_REG_out_reg_126_ ( .D(n405), .CK(clk), .RN(n612), .Q(out[126])
         );
  DFFR_X1 ID_EX_REG_out_reg_125_ ( .D(n404), .CK(clk), .RN(n614), .Q(out[125])
         );
  DFFR_X1 ID_EX_REG_out_reg_124_ ( .D(n403), .CK(clk), .RN(n612), .Q(out[124])
         );
  DFFR_X1 ID_EX_REG_out_reg_123_ ( .D(n402), .CK(clk), .RN(n614), .Q(out[123])
         );
  DFFR_X1 ID_EX_REG_out_reg_122_ ( .D(n401), .CK(clk), .RN(n612), .Q(out[122])
         );
  DFFR_X1 ID_EX_REG_out_reg_121_ ( .D(n400), .CK(clk), .RN(n614), .Q(out[121])
         );
  DFFR_X1 ID_EX_REG_out_reg_120_ ( .D(n399), .CK(clk), .RN(n612), .Q(out[120])
         );
  DFFR_X1 ID_EX_REG_out_reg_119_ ( .D(n398), .CK(clk), .RN(n612), .Q(out[119])
         );
  DFFR_X1 ID_EX_REG_out_reg_118_ ( .D(n397), .CK(clk), .RN(n614), .Q(out[118])
         );
  DFFR_X1 ID_EX_REG_out_reg_117_ ( .D(n396), .CK(clk), .RN(n612), .Q(out[117])
         );
  DFFR_X1 ID_EX_REG_out_reg_116_ ( .D(n395), .CK(clk), .RN(n614), .Q(out[116])
         );
  DFFR_X1 ID_EX_REG_out_reg_115_ ( .D(n394), .CK(clk), .RN(n612), .Q(out[115])
         );
  DFFR_X1 ID_EX_REG_out_reg_114_ ( .D(n393), .CK(clk), .RN(n614), .Q(out[114])
         );
  DFFR_X1 ID_EX_REG_out_reg_113_ ( .D(n392), .CK(clk), .RN(n612), .Q(out[113])
         );
  DFFR_X1 ID_EX_REG_out_reg_112_ ( .D(n391), .CK(clk), .RN(n614), .Q(out[112])
         );
  DFFR_X1 ID_EX_REG_out_reg_111_ ( .D(n390), .CK(clk), .RN(n612), .Q(out[111])
         );
  DFFR_X1 ID_EX_REG_out_reg_110_ ( .D(n389), .CK(clk), .RN(n614), .Q(out[110])
         );
  DFFR_X1 ID_EX_REG_out_reg_109_ ( .D(n388), .CK(clk), .RN(n613), .Q(out[109])
         );
  DFFR_X1 ID_EX_REG_out_reg_108_ ( .D(n387), .CK(clk), .RN(n613), .Q(out[108])
         );
  DFFR_X1 ID_EX_REG_out_reg_107_ ( .D(n386), .CK(clk), .RN(n613), .Q(out[107])
         );
  DFFR_X1 ID_EX_REG_out_reg_106_ ( .D(n385), .CK(clk), .RN(n613), .Q(out[106])
         );
  DFFR_X1 ID_EX_REG_out_reg_105_ ( .D(n384), .CK(clk), .RN(n613), .Q(out[105])
         );
  DFFR_X1 ID_EX_REG_out_reg_104_ ( .D(n383), .CK(clk), .RN(n613), .Q(out[104])
         );
  DFFR_X1 ID_EX_REG_out_reg_103_ ( .D(n382), .CK(clk), .RN(n613), .Q(out[103])
         );
  DFFR_X1 ID_EX_REG_out_reg_102_ ( .D(n381), .CK(clk), .RN(n613), .Q(out[102])
         );
  DFFR_X1 ID_EX_REG_out_reg_101_ ( .D(n380), .CK(clk), .RN(n613), .Q(out[101])
         );
  DFFR_X1 ID_EX_REG_out_reg_100_ ( .D(n379), .CK(clk), .RN(n613), .Q(out[100])
         );
  DFFR_X1 ID_EX_REG_out_reg_99_ ( .D(n378), .CK(clk), .RN(n605), .Q(out[99])
         );
  DFFR_X1 ID_EX_REG_out_reg_98_ ( .D(n377), .CK(clk), .RN(n623), .Q(out[98])
         );
  DFFR_X1 ID_EX_REG_out_reg_97_ ( .D(n376), .CK(clk), .RN(n605), .Q(out[97])
         );
  DFFR_X1 ID_EX_REG_out_reg_96_ ( .D(n375), .CK(clk), .RN(n623), .Q(out[96])
         );
  DFFR_X1 ID_EX_REG_out_reg_95_ ( .D(n374), .CK(clk), .RN(n605), .Q(out[95])
         );
  DFFR_X1 ID_EX_REG_out_reg_94_ ( .D(n373), .CK(clk), .RN(n623), .Q(out[94])
         );
  DFFR_X1 ID_EX_REG_out_reg_93_ ( .D(n372), .CK(clk), .RN(n605), .Q(out[93])
         );
  DFFR_X1 ID_EX_REG_out_reg_92_ ( .D(n371), .CK(clk), .RN(n623), .Q(out[92])
         );
  DFFR_X1 ID_EX_REG_out_reg_91_ ( .D(n370), .CK(clk), .RN(n605), .Q(out[91])
         );
  DFFR_X1 ID_EX_REG_out_reg_90_ ( .D(n369), .CK(clk), .RN(n623), .Q(out[90])
         );
  DFFR_X1 ID_EX_REG_out_reg_89_ ( .D(n368), .CK(clk), .RN(n623), .Q(out[89])
         );
  DFFR_X1 ID_EX_REG_out_reg_88_ ( .D(n367), .CK(clk), .RN(n605), .Q(out[88])
         );
  DFFR_X1 ID_EX_REG_out_reg_87_ ( .D(n366), .CK(clk), .RN(n623), .Q(out[87])
         );
  DFFR_X1 ID_EX_REG_out_reg_86_ ( .D(n365), .CK(clk), .RN(n605), .Q(out[86])
         );
  DFFR_X1 ID_EX_REG_out_reg_85_ ( .D(n364), .CK(clk), .RN(n623), .Q(out[85])
         );
  DFFR_X1 ID_EX_REG_out_reg_84_ ( .D(n363), .CK(clk), .RN(n605), .Q(out[84])
         );
  DFFR_X1 ID_EX_REG_out_reg_83_ ( .D(n362), .CK(clk), .RN(n623), .Q(out[83])
         );
  DFFR_X1 ID_EX_REG_out_reg_82_ ( .D(n361), .CK(clk), .RN(n605), .Q(out[82])
         );
  DFFR_X1 ID_EX_REG_out_reg_81_ ( .D(n360), .CK(clk), .RN(n623), .Q(out[81])
         );
  DFFR_X1 ID_EX_REG_out_reg_80_ ( .D(n359), .CK(clk), .RN(n605), .Q(out[80])
         );
  DFFR_X1 ID_EX_REG_out_reg_79_ ( .D(n358), .CK(clk), .RN(n605), .Q(out[79])
         );
  DFFR_X1 ID_EX_REG_out_reg_78_ ( .D(n357), .CK(clk), .RN(n623), .Q(out[78])
         );
  DFFR_X1 ID_EX_REG_out_reg_77_ ( .D(n356), .CK(clk), .RN(n606), .Q(out[77])
         );
  DFFR_X1 ID_EX_REG_out_reg_76_ ( .D(n355), .CK(clk), .RN(n622), .Q(out[76])
         );
  DFFR_X1 ID_EX_REG_out_reg_75_ ( .D(n354), .CK(clk), .RN(n606), .Q(out[75])
         );
  DFFR_X1 ID_EX_REG_out_reg_74_ ( .D(n353), .CK(clk), .RN(n622), .Q(out[74])
         );
  DFFR_X1 ID_EX_REG_out_reg_73_ ( .D(n352), .CK(clk), .RN(n606), .Q(out[73])
         );
  DFFR_X1 ID_EX_REG_out_reg_72_ ( .D(n351), .CK(clk), .RN(n622), .Q(out[72])
         );
  DFFR_X1 ID_EX_REG_out_reg_71_ ( .D(n350), .CK(clk), .RN(n606), .Q(out[71])
         );
  DFFR_X1 ID_EX_REG_out_reg_70_ ( .D(n349), .CK(clk), .RN(n622), .Q(out[70])
         );
  DFFR_X1 ID_EX_REG_out_reg_69_ ( .D(n348), .CK(clk), .RN(n622), .Q(out[69])
         );
  DFFR_X1 ID_EX_REG_out_reg_68_ ( .D(n347), .CK(clk), .RN(n606), .Q(out[68])
         );
  DFFR_X1 ID_EX_REG_out_reg_67_ ( .D(n346), .CK(clk), .RN(n622), .Q(out[67])
         );
  DFFR_X1 ID_EX_REG_out_reg_66_ ( .D(n345), .CK(clk), .RN(n606), .Q(out[66])
         );
  DFFR_X1 ID_EX_REG_out_reg_65_ ( .D(n344), .CK(clk), .RN(n622), .Q(out[65])
         );
  DFFR_X1 ID_EX_REG_out_reg_64_ ( .D(n343), .CK(clk), .RN(n606), .Q(out[64])
         );
  DFFR_X1 ID_EX_REG_out_reg_63_ ( .D(n342), .CK(clk), .RN(n622), .Q(out[63])
         );
  DFFR_X1 ID_EX_REG_out_reg_62_ ( .D(n341), .CK(clk), .RN(n606), .Q(out[62])
         );
  DFFR_X1 ID_EX_REG_out_reg_61_ ( .D(n340), .CK(clk), .RN(n622), .Q(out[61])
         );
  DFFR_X1 ID_EX_REG_out_reg_60_ ( .D(n339), .CK(clk), .RN(n606), .Q(out[60])
         );
  DFFR_X1 ID_EX_REG_out_reg_59_ ( .D(n338), .CK(clk), .RN(n606), .Q(out[59])
         );
  DFFR_X1 ID_EX_REG_out_reg_58_ ( .D(n337), .CK(clk), .RN(n622), .Q(out[58])
         );
  DFFR_X1 ID_EX_REG_out_reg_57_ ( .D(n336), .CK(clk), .RN(n606), .Q(out[57])
         );
  DFFR_X1 ID_EX_REG_out_reg_56_ ( .D(n335), .CK(clk), .RN(n622), .Q(out[56])
         );
  DFFR_X1 ID_EX_REG_out_reg_55_ ( .D(n334), .CK(clk), .RN(n607), .Q(out[55])
         );
  DFFR_X1 ID_EX_REG_out_reg_54_ ( .D(n333), .CK(clk), .RN(n621), .Q(out[54])
         );
  DFFR_X1 ID_EX_REG_out_reg_53_ ( .D(n332), .CK(clk), .RN(n607), .Q(out[53])
         );
  DFFR_X1 ID_EX_REG_out_reg_52_ ( .D(n331), .CK(clk), .RN(n621), .Q(out[52])
         );
  DFFR_X1 ID_EX_REG_out_reg_51_ ( .D(n330), .CK(clk), .RN(n607), .Q(out[51])
         );
  DFFR_X1 ID_EX_REG_out_reg_50_ ( .D(n329), .CK(clk), .RN(n621), .Q(out[50])
         );
  DFFR_X1 ID_EX_REG_out_reg_49_ ( .D(n328), .CK(clk), .RN(n621), .Q(out[49])
         );
  DFFR_X1 ID_EX_REG_out_reg_48_ ( .D(n327), .CK(clk), .RN(n607), .Q(out[48])
         );
  DFFR_X1 ID_EX_REG_out_reg_47_ ( .D(n326), .CK(clk), .RN(n621), .Q(out[47])
         );
  DFFR_X1 ID_EX_REG_out_reg_46_ ( .D(n325), .CK(clk), .RN(n607), .Q(out[46])
         );
  DFFR_X1 ID_EX_REG_out_reg_45_ ( .D(n324), .CK(clk), .RN(n621), .Q(out[45])
         );
  DFFR_X1 ID_EX_REG_out_reg_44_ ( .D(n323), .CK(clk), .RN(n607), .Q(out[44])
         );
  DFFR_X1 ID_EX_REG_out_reg_43_ ( .D(n322), .CK(clk), .RN(n621), .Q(out[43])
         );
  DFFR_X1 ID_EX_REG_out_reg_42_ ( .D(n321), .CK(clk), .RN(n607), .Q(out[42])
         );
  DFFR_X1 ID_EX_REG_out_reg_41_ ( .D(n320), .CK(clk), .RN(n621), .Q(out[41])
         );
  DFFR_X1 ID_EX_REG_out_reg_40_ ( .D(n319), .CK(clk), .RN(n607), .Q(out[40])
         );
  DFFR_X1 ID_EX_REG_out_reg_39_ ( .D(n318), .CK(clk), .RN(n607), .Q(out[39])
         );
  DFFR_X1 ID_EX_REG_out_reg_38_ ( .D(n317), .CK(clk), .RN(n621), .Q(out[38])
         );
  DFFR_X1 ID_EX_REG_out_reg_37_ ( .D(n316), .CK(clk), .RN(n607), .Q(out[37])
         );
  DFFR_X1 ID_EX_REG_out_reg_36_ ( .D(n315), .CK(clk), .RN(n621), .Q(out[36])
         );
  DFFR_X1 ID_EX_REG_out_reg_35_ ( .D(n314), .CK(clk), .RN(n607), .Q(out[35])
         );
  DFFR_X1 ID_EX_REG_out_reg_34_ ( .D(n313), .CK(clk), .RN(n621), .Q(out[34])
         );
  DFFR_X1 ID_EX_REG_out_reg_33_ ( .D(n312), .CK(clk), .RN(n617), .Q(out[33])
         );
  DFFR_X1 ID_EX_REG_out_reg_32_ ( .D(n311), .CK(clk), .RN(n620), .Q(out[32])
         );
  DFFR_X1 ID_EX_REG_out_reg_31_ ( .D(n310), .CK(clk), .RN(n616), .Q(out[31])
         );
  DFFR_X1 ID_EX_REG_out_reg_30_ ( .D(n309), .CK(clk), .RN(n620), .Q(out[30])
         );
  DFFR_X1 ID_EX_REG_out_reg_29_ ( .D(n308), .CK(clk), .RN(n620), .Q(out[29])
         );
  DFFR_X1 ID_EX_REG_out_reg_28_ ( .D(n307), .CK(clk), .RN(n615), .Q(out[28])
         );
  DFFR_X1 ID_EX_REG_out_reg_27_ ( .D(n306), .CK(clk), .RN(n620), .Q(out[27])
         );
  DFFR_X1 ID_EX_REG_out_reg_26_ ( .D(n305), .CK(clk), .RN(n620), .Q(out[26])
         );
  DFFR_X1 ID_EX_REG_out_reg_25_ ( .D(n304), .CK(clk), .RN(n620), .Q(out[25])
         );
  DFFR_X1 ID_EX_REG_out_reg_24_ ( .D(n303), .CK(clk), .RN(n614), .Q(out[24])
         );
  DFFR_X1 ID_EX_REG_out_reg_23_ ( .D(n302), .CK(clk), .RN(n621), .Q(out[23])
         );
  DFFR_X1 ID_EX_REG_out_reg_22_ ( .D(n301), .CK(clk), .RN(n619), .Q(out[22])
         );
  DFFR_X1 ID_EX_REG_out_reg_21_ ( .D(n300), .CK(clk), .RN(n622), .Q(out[21])
         );
  DFFR_X1 ID_EX_REG_out_reg_20_ ( .D(n299), .CK(clk), .RN(n618), .Q(out[20])
         );
  DFFR_X1 ID_EX_REG_out_reg_19_ ( .D(n298), .CK(clk), .RN(n618), .Q(out[19])
         );
  DFFR_X1 ID_EX_REG_out_reg_18_ ( .D(n297), .CK(clk), .RN(n609), .Q(out[18])
         );
  DFFR_X1 ID_EX_REG_out_reg_17_ ( .D(n296), .CK(clk), .RN(n617), .Q(out[17])
         );
  DFFR_X1 ID_EX_REG_out_reg_16_ ( .D(n295), .CK(clk), .RN(n610), .Q(out[16])
         );
  DFFR_X1 ID_EX_REG_out_reg_15_ ( .D(n294), .CK(clk), .RN(n616), .Q(out[15])
         );
  DFFR_X1 ID_EX_REG_out_reg_14_ ( .D(n293), .CK(clk), .RN(n611), .Q(out[14])
         );
  DFFR_X1 ID_EX_REG_out_reg_13_ ( .D(n292), .CK(clk), .RN(n615), .Q(out[13])
         );
  DFFR_X1 ID_EX_REG_out_reg_12_ ( .D(n291), .CK(clk), .RN(n612), .Q(out[12])
         );
  DFFR_X1 ID_EX_REG_out_reg_11_ ( .D(n290), .CK(clk), .RN(n614), .Q(out[11])
         );
  DFFR_X1 ID_EX_REG_out_reg_10_ ( .D(n289), .CK(clk), .RN(n613), .Q(out[10])
         );
  DFFR_X1 ID_EX_REG_out_reg_9_ ( .D(n288), .CK(clk), .RN(reset), .Q(out[9]) );
  DFFR_X1 ID_EX_REG_out_reg_8_ ( .D(n287), .CK(clk), .RN(n605), .Q(out[8]) );
  DFFR_X1 ID_EX_REG_out_reg_7_ ( .D(n286), .CK(clk), .RN(n623), .Q(out[7]) );
  DFFR_X1 ID_EX_REG_out_reg_6_ ( .D(n285), .CK(clk), .RN(n606), .Q(out[6]) );
  DFFR_X1 ID_EX_REG_out_reg_5_ ( .D(n284), .CK(clk), .RN(n622), .Q(out[5]) );
  DFFR_X1 ID_EX_REG_out_reg_4_ ( .D(n283), .CK(clk), .RN(n607), .Q(out[4]) );
  DFFR_X1 ID_EX_REG_out_reg_3_ ( .D(n282), .CK(clk), .RN(n621), .Q(out[3]) );
  DFFR_X1 ID_EX_REG_out_reg_2_ ( .D(n281), .CK(clk), .RN(n614), .Q(out[2]) );
  DFFR_X1 ID_EX_REG_out_reg_1_ ( .D(n280), .CK(clk), .RN(n608), .Q(out[1]) );
  DFFR_X1 ID_EX_REG_out_reg_0_ ( .D(n279), .CK(clk), .RN(n613), .Q(out[0]) );
  INV_X1 U1 ( .A(n1), .ZN(n288) );
  AOI22_X1 U2 ( .A1(in[9]), .A2(n557), .B1(n586), .B2(out[9]), .ZN(n1) );
  INV_X1 U3 ( .A(n3), .ZN(n378) );
  AOI22_X1 U4 ( .A1(in[99]), .A2(n556), .B1(out[99]), .B2(n586), .ZN(n3) );
  INV_X1 U5 ( .A(n4), .ZN(n377) );
  AOI22_X1 U6 ( .A1(in[98]), .A2(n580), .B1(out[98]), .B2(n586), .ZN(n4) );
  INV_X1 U7 ( .A(n5), .ZN(n376) );
  AOI22_X1 U8 ( .A1(in[97]), .A2(n580), .B1(out[97]), .B2(n586), .ZN(n5) );
  INV_X1 U9 ( .A(n6), .ZN(n375) );
  AOI22_X1 U10 ( .A1(in[96]), .A2(n580), .B1(out[96]), .B2(n586), .ZN(n6) );
  INV_X1 U11 ( .A(n7), .ZN(n374) );
  AOI22_X1 U12 ( .A1(in[95]), .A2(n580), .B1(out[95]), .B2(n586), .ZN(n7) );
  INV_X1 U13 ( .A(n8), .ZN(n373) );
  AOI22_X1 U14 ( .A1(in[94]), .A2(n580), .B1(out[94]), .B2(n586), .ZN(n8) );
  INV_X1 U15 ( .A(n9), .ZN(n372) );
  AOI22_X1 U16 ( .A1(in[93]), .A2(n580), .B1(out[93]), .B2(n586), .ZN(n9) );
  INV_X1 U17 ( .A(n10), .ZN(n371) );
  AOI22_X1 U18 ( .A1(in[92]), .A2(n580), .B1(out[92]), .B2(n586), .ZN(n10) );
  INV_X1 U19 ( .A(n11), .ZN(n370) );
  AOI22_X1 U20 ( .A1(in[91]), .A2(n580), .B1(out[91]), .B2(n586), .ZN(n11) );
  INV_X1 U21 ( .A(n12), .ZN(n369) );
  AOI22_X1 U22 ( .A1(in[90]), .A2(n580), .B1(out[90]), .B2(n586), .ZN(n12) );
  INV_X1 U23 ( .A(n13), .ZN(n287) );
  AOI22_X1 U24 ( .A1(in[8]), .A2(n580), .B1(out[8]), .B2(n586), .ZN(n13) );
  INV_X1 U25 ( .A(n14), .ZN(n368) );
  AOI22_X1 U26 ( .A1(in[89]), .A2(n580), .B1(out[89]), .B2(n604), .ZN(n14) );
  INV_X1 U27 ( .A(n15), .ZN(n367) );
  AOI22_X1 U28 ( .A1(in[88]), .A2(n579), .B1(out[88]), .B2(n603), .ZN(n15) );
  INV_X1 U29 ( .A(n16), .ZN(n366) );
  AOI22_X1 U30 ( .A1(in[87]), .A2(n579), .B1(out[87]), .B2(n602), .ZN(n16) );
  INV_X1 U31 ( .A(n17), .ZN(n365) );
  AOI22_X1 U32 ( .A1(in[86]), .A2(n579), .B1(out[86]), .B2(n601), .ZN(n17) );
  INV_X1 U33 ( .A(n18), .ZN(n364) );
  AOI22_X1 U34 ( .A1(in[85]), .A2(n579), .B1(out[85]), .B2(n604), .ZN(n18) );
  INV_X1 U35 ( .A(n19), .ZN(n363) );
  AOI22_X1 U36 ( .A1(in[84]), .A2(n579), .B1(out[84]), .B2(n603), .ZN(n19) );
  INV_X1 U37 ( .A(n20), .ZN(n362) );
  AOI22_X1 U38 ( .A1(in[83]), .A2(n579), .B1(out[83]), .B2(n602), .ZN(n20) );
  INV_X1 U39 ( .A(n21), .ZN(n361) );
  AOI22_X1 U40 ( .A1(in[82]), .A2(n579), .B1(out[82]), .B2(n601), .ZN(n21) );
  INV_X1 U41 ( .A(n22), .ZN(n360) );
  AOI22_X1 U42 ( .A1(in[81]), .A2(n579), .B1(out[81]), .B2(n604), .ZN(n22) );
  INV_X1 U43 ( .A(n23), .ZN(n359) );
  AOI22_X1 U44 ( .A1(in[80]), .A2(n579), .B1(out[80]), .B2(n603), .ZN(n23) );
  INV_X1 U45 ( .A(n24), .ZN(n286) );
  AOI22_X1 U46 ( .A1(in[7]), .A2(n579), .B1(out[7]), .B2(n602), .ZN(n24) );
  INV_X1 U47 ( .A(n25), .ZN(n358) );
  AOI22_X1 U48 ( .A1(in[79]), .A2(n579), .B1(out[79]), .B2(n601), .ZN(n25) );
  INV_X1 U49 ( .A(n26), .ZN(n357) );
  AOI22_X1 U50 ( .A1(in[78]), .A2(n578), .B1(out[78]), .B2(n604), .ZN(n26) );
  INV_X1 U51 ( .A(n27), .ZN(n356) );
  AOI22_X1 U52 ( .A1(in[77]), .A2(n578), .B1(out[77]), .B2(n603), .ZN(n27) );
  INV_X1 U53 ( .A(n28), .ZN(n355) );
  AOI22_X1 U54 ( .A1(in[76]), .A2(n578), .B1(out[76]), .B2(n602), .ZN(n28) );
  INV_X1 U55 ( .A(n29), .ZN(n354) );
  AOI22_X1 U56 ( .A1(in[75]), .A2(n578), .B1(out[75]), .B2(n601), .ZN(n29) );
  INV_X1 U57 ( .A(n30), .ZN(n353) );
  AOI22_X1 U58 ( .A1(in[74]), .A2(n578), .B1(out[74]), .B2(n604), .ZN(n30) );
  INV_X1 U59 ( .A(n31), .ZN(n352) );
  AOI22_X1 U60 ( .A1(in[73]), .A2(n578), .B1(out[73]), .B2(n603), .ZN(n31) );
  INV_X1 U61 ( .A(n32), .ZN(n351) );
  AOI22_X1 U62 ( .A1(in[72]), .A2(n578), .B1(out[72]), .B2(n602), .ZN(n32) );
  INV_X1 U63 ( .A(n33), .ZN(n350) );
  AOI22_X1 U64 ( .A1(in[71]), .A2(n578), .B1(out[71]), .B2(n601), .ZN(n33) );
  INV_X1 U65 ( .A(n34), .ZN(n349) );
  AOI22_X1 U66 ( .A1(in[70]), .A2(n578), .B1(out[70]), .B2(n604), .ZN(n34) );
  INV_X1 U67 ( .A(n35), .ZN(n285) );
  AOI22_X1 U68 ( .A1(in[6]), .A2(n578), .B1(out[6]), .B2(n603), .ZN(n35) );
  INV_X1 U69 ( .A(n36), .ZN(n348) );
  AOI22_X1 U70 ( .A1(in[69]), .A2(n578), .B1(out[69]), .B2(n602), .ZN(n36) );
  INV_X1 U71 ( .A(n37), .ZN(n347) );
  AOI22_X1 U72 ( .A1(in[68]), .A2(n577), .B1(out[68]), .B2(n601), .ZN(n37) );
  INV_X1 U73 ( .A(n38), .ZN(n346) );
  AOI22_X1 U74 ( .A1(in[67]), .A2(n577), .B1(out[67]), .B2(n604), .ZN(n38) );
  INV_X1 U75 ( .A(n39), .ZN(n345) );
  AOI22_X1 U76 ( .A1(in[66]), .A2(n577), .B1(out[66]), .B2(n603), .ZN(n39) );
  INV_X1 U77 ( .A(n40), .ZN(n344) );
  AOI22_X1 U78 ( .A1(in[65]), .A2(n577), .B1(out[65]), .B2(n602), .ZN(n40) );
  INV_X1 U79 ( .A(n41), .ZN(n343) );
  AOI22_X1 U80 ( .A1(in[64]), .A2(n577), .B1(out[64]), .B2(n601), .ZN(n41) );
  INV_X1 U81 ( .A(n42), .ZN(n342) );
  AOI22_X1 U82 ( .A1(in[63]), .A2(n577), .B1(out[63]), .B2(n604), .ZN(n42) );
  INV_X1 U83 ( .A(n43), .ZN(n341) );
  AOI22_X1 U84 ( .A1(in[62]), .A2(n577), .B1(out[62]), .B2(n603), .ZN(n43) );
  INV_X1 U85 ( .A(n44), .ZN(n340) );
  AOI22_X1 U86 ( .A1(in[61]), .A2(n577), .B1(out[61]), .B2(n602), .ZN(n44) );
  INV_X1 U87 ( .A(n45), .ZN(n339) );
  AOI22_X1 U88 ( .A1(in[60]), .A2(n577), .B1(out[60]), .B2(n601), .ZN(n45) );
  INV_X1 U89 ( .A(n46), .ZN(n284) );
  AOI22_X1 U90 ( .A1(in[5]), .A2(n577), .B1(out[5]), .B2(n604), .ZN(n46) );
  INV_X1 U91 ( .A(n47), .ZN(n338) );
  AOI22_X1 U92 ( .A1(in[59]), .A2(n577), .B1(out[59]), .B2(n603), .ZN(n47) );
  INV_X1 U93 ( .A(n48), .ZN(n337) );
  AOI22_X1 U94 ( .A1(in[58]), .A2(n576), .B1(out[58]), .B2(n602), .ZN(n48) );
  INV_X1 U95 ( .A(n49), .ZN(n336) );
  AOI22_X1 U96 ( .A1(in[57]), .A2(n576), .B1(out[57]), .B2(n601), .ZN(n49) );
  INV_X1 U97 ( .A(n50), .ZN(n335) );
  AOI22_X1 U98 ( .A1(in[56]), .A2(n576), .B1(out[56]), .B2(n587), .ZN(n50) );
  INV_X1 U99 ( .A(n51), .ZN(n334) );
  AOI22_X1 U100 ( .A1(in[55]), .A2(n576), .B1(out[55]), .B2(n587), .ZN(n51) );
  INV_X1 U101 ( .A(n52), .ZN(n333) );
  AOI22_X1 U102 ( .A1(in[54]), .A2(n576), .B1(out[54]), .B2(n587), .ZN(n52) );
  INV_X1 U103 ( .A(n53), .ZN(n332) );
  AOI22_X1 U104 ( .A1(in[53]), .A2(n576), .B1(out[53]), .B2(n587), .ZN(n53) );
  INV_X1 U105 ( .A(n54), .ZN(n331) );
  AOI22_X1 U106 ( .A1(in[52]), .A2(n576), .B1(out[52]), .B2(n587), .ZN(n54) );
  INV_X1 U107 ( .A(n55), .ZN(n330) );
  AOI22_X1 U108 ( .A1(in[51]), .A2(n576), .B1(out[51]), .B2(n587), .ZN(n55) );
  INV_X1 U109 ( .A(n56), .ZN(n329) );
  AOI22_X1 U110 ( .A1(in[50]), .A2(n576), .B1(out[50]), .B2(n587), .ZN(n56) );
  INV_X1 U111 ( .A(n57), .ZN(n283) );
  AOI22_X1 U112 ( .A1(in[4]), .A2(n576), .B1(out[4]), .B2(n587), .ZN(n57) );
  INV_X1 U113 ( .A(n58), .ZN(n328) );
  AOI22_X1 U114 ( .A1(in[49]), .A2(n576), .B1(out[49]), .B2(n587), .ZN(n58) );
  INV_X1 U115 ( .A(n59), .ZN(n327) );
  AOI22_X1 U116 ( .A1(in[48]), .A2(n575), .B1(out[48]), .B2(n587), .ZN(n59) );
  INV_X1 U117 ( .A(n60), .ZN(n326) );
  AOI22_X1 U118 ( .A1(in[47]), .A2(n575), .B1(out[47]), .B2(n587), .ZN(n60) );
  INV_X1 U119 ( .A(n61), .ZN(n325) );
  AOI22_X1 U120 ( .A1(in[46]), .A2(n575), .B1(out[46]), .B2(n587), .ZN(n61) );
  INV_X1 U121 ( .A(n62), .ZN(n324) );
  AOI22_X1 U122 ( .A1(in[45]), .A2(n575), .B1(out[45]), .B2(n588), .ZN(n62) );
  INV_X1 U123 ( .A(n63), .ZN(n323) );
  AOI22_X1 U124 ( .A1(in[44]), .A2(n575), .B1(out[44]), .B2(n588), .ZN(n63) );
  INV_X1 U125 ( .A(n64), .ZN(n322) );
  AOI22_X1 U126 ( .A1(in[43]), .A2(n575), .B1(out[43]), .B2(n588), .ZN(n64) );
  INV_X1 U127 ( .A(n65), .ZN(n321) );
  AOI22_X1 U128 ( .A1(in[42]), .A2(n575), .B1(out[42]), .B2(n588), .ZN(n65) );
  INV_X1 U129 ( .A(n66), .ZN(n320) );
  AOI22_X1 U130 ( .A1(in[41]), .A2(n575), .B1(out[41]), .B2(n588), .ZN(n66) );
  INV_X1 U131 ( .A(n67), .ZN(n319) );
  AOI22_X1 U132 ( .A1(in[40]), .A2(n575), .B1(out[40]), .B2(n588), .ZN(n67) );
  INV_X1 U133 ( .A(n68), .ZN(n282) );
  AOI22_X1 U134 ( .A1(in[3]), .A2(n575), .B1(out[3]), .B2(n588), .ZN(n68) );
  INV_X1 U135 ( .A(n69), .ZN(n318) );
  AOI22_X1 U136 ( .A1(in[39]), .A2(n575), .B1(out[39]), .B2(n588), .ZN(n69) );
  INV_X1 U137 ( .A(n70), .ZN(n317) );
  AOI22_X1 U138 ( .A1(in[38]), .A2(n574), .B1(out[38]), .B2(n588), .ZN(n70) );
  INV_X1 U139 ( .A(n71), .ZN(n316) );
  AOI22_X1 U140 ( .A1(in[37]), .A2(n574), .B1(out[37]), .B2(n588), .ZN(n71) );
  INV_X1 U141 ( .A(n72), .ZN(n315) );
  AOI22_X1 U142 ( .A1(in[36]), .A2(n574), .B1(out[36]), .B2(n588), .ZN(n72) );
  INV_X1 U143 ( .A(n73), .ZN(n314) );
  AOI22_X1 U144 ( .A1(in[35]), .A2(n574), .B1(out[35]), .B2(n588), .ZN(n73) );
  INV_X1 U145 ( .A(n74), .ZN(n313) );
  AOI22_X1 U146 ( .A1(in[34]), .A2(n574), .B1(out[34]), .B2(n589), .ZN(n74) );
  INV_X1 U147 ( .A(n75), .ZN(n312) );
  AOI22_X1 U148 ( .A1(in[33]), .A2(n574), .B1(out[33]), .B2(n589), .ZN(n75) );
  INV_X1 U149 ( .A(n76), .ZN(n311) );
  AOI22_X1 U150 ( .A1(in[32]), .A2(n574), .B1(out[32]), .B2(n589), .ZN(n76) );
  INV_X1 U151 ( .A(n77), .ZN(n310) );
  AOI22_X1 U152 ( .A1(in[31]), .A2(n574), .B1(out[31]), .B2(n589), .ZN(n77) );
  INV_X1 U153 ( .A(n78), .ZN(n309) );
  AOI22_X1 U154 ( .A1(in[30]), .A2(n574), .B1(out[30]), .B2(n589), .ZN(n78) );
  INV_X1 U155 ( .A(n79), .ZN(n281) );
  AOI22_X1 U156 ( .A1(in[2]), .A2(n574), .B1(out[2]), .B2(n589), .ZN(n79) );
  INV_X1 U157 ( .A(n80), .ZN(n308) );
  AOI22_X1 U158 ( .A1(in[29]), .A2(n574), .B1(out[29]), .B2(n589), .ZN(n80) );
  INV_X1 U159 ( .A(n81), .ZN(n307) );
  AOI22_X1 U160 ( .A1(in[28]), .A2(n573), .B1(out[28]), .B2(n589), .ZN(n81) );
  INV_X1 U161 ( .A(n82), .ZN(n306) );
  AOI22_X1 U162 ( .A1(in[27]), .A2(n573), .B1(out[27]), .B2(n589), .ZN(n82) );
  INV_X1 U163 ( .A(n83), .ZN(n555) );
  AOI22_X1 U164 ( .A1(in[276]), .A2(n573), .B1(out[276]), .B2(n589), .ZN(n83)
         );
  INV_X1 U165 ( .A(n84), .ZN(n554) );
  AOI22_X1 U166 ( .A1(in[275]), .A2(n573), .B1(out[275]), .B2(n589), .ZN(n84)
         );
  INV_X1 U167 ( .A(n85), .ZN(n553) );
  AOI22_X1 U168 ( .A1(in[274]), .A2(n573), .B1(out[274]), .B2(n589), .ZN(n85)
         );
  INV_X1 U169 ( .A(n86), .ZN(n552) );
  AOI22_X1 U170 ( .A1(in[273]), .A2(n573), .B1(out[273]), .B2(n590), .ZN(n86)
         );
  INV_X1 U171 ( .A(n87), .ZN(n551) );
  AOI22_X1 U172 ( .A1(in[272]), .A2(n573), .B1(out[272]), .B2(n590), .ZN(n87)
         );
  INV_X1 U173 ( .A(n88), .ZN(n550) );
  AOI22_X1 U174 ( .A1(in[271]), .A2(n573), .B1(out[271]), .B2(n590), .ZN(n88)
         );
  INV_X1 U175 ( .A(n89), .ZN(n549) );
  AOI22_X1 U176 ( .A1(in[270]), .A2(n573), .B1(out[270]), .B2(n590), .ZN(n89)
         );
  INV_X1 U177 ( .A(n90), .ZN(n305) );
  AOI22_X1 U178 ( .A1(in[26]), .A2(n573), .B1(out[26]), .B2(n590), .ZN(n90) );
  INV_X1 U179 ( .A(n91), .ZN(n548) );
  AOI22_X1 U180 ( .A1(in[269]), .A2(n573), .B1(out[269]), .B2(n590), .ZN(n91)
         );
  INV_X1 U181 ( .A(n92), .ZN(n547) );
  AOI22_X1 U182 ( .A1(in[268]), .A2(n572), .B1(out[268]), .B2(n590), .ZN(n92)
         );
  INV_X1 U183 ( .A(n93), .ZN(n546) );
  AOI22_X1 U184 ( .A1(in[267]), .A2(n572), .B1(out[267]), .B2(n590), .ZN(n93)
         );
  INV_X1 U185 ( .A(n94), .ZN(n545) );
  AOI22_X1 U186 ( .A1(in[266]), .A2(n572), .B1(out[266]), .B2(n590), .ZN(n94)
         );
  INV_X1 U187 ( .A(n95), .ZN(n544) );
  AOI22_X1 U188 ( .A1(in[265]), .A2(n572), .B1(out[265]), .B2(n590), .ZN(n95)
         );
  INV_X1 U189 ( .A(n96), .ZN(n543) );
  AOI22_X1 U190 ( .A1(in[264]), .A2(n572), .B1(out[264]), .B2(n590), .ZN(n96)
         );
  INV_X1 U191 ( .A(n97), .ZN(n542) );
  AOI22_X1 U192 ( .A1(in[263]), .A2(n572), .B1(out[263]), .B2(n590), .ZN(n97)
         );
  INV_X1 U193 ( .A(n98), .ZN(n541) );
  AOI22_X1 U194 ( .A1(in[262]), .A2(n572), .B1(out[262]), .B2(n591), .ZN(n98)
         );
  INV_X1 U195 ( .A(n99), .ZN(n540) );
  AOI22_X1 U196 ( .A1(in[261]), .A2(n572), .B1(out[261]), .B2(n591), .ZN(n99)
         );
  INV_X1 U197 ( .A(n100), .ZN(n539) );
  AOI22_X1 U198 ( .A1(in[260]), .A2(n572), .B1(out[260]), .B2(n591), .ZN(n100)
         );
  INV_X1 U199 ( .A(n101), .ZN(n304) );
  AOI22_X1 U200 ( .A1(in[25]), .A2(n572), .B1(out[25]), .B2(n591), .ZN(n101)
         );
  INV_X1 U201 ( .A(n102), .ZN(n538) );
  AOI22_X1 U202 ( .A1(in[259]), .A2(n572), .B1(out[259]), .B2(n591), .ZN(n102)
         );
  INV_X1 U203 ( .A(n103), .ZN(n537) );
  AOI22_X1 U204 ( .A1(in[258]), .A2(n571), .B1(out[258]), .B2(n591), .ZN(n103)
         );
  INV_X1 U205 ( .A(n104), .ZN(n536) );
  AOI22_X1 U206 ( .A1(in[257]), .A2(n571), .B1(out[257]), .B2(n591), .ZN(n104)
         );
  INV_X1 U207 ( .A(n105), .ZN(n535) );
  AOI22_X1 U208 ( .A1(in[256]), .A2(n571), .B1(out[256]), .B2(n591), .ZN(n105)
         );
  INV_X1 U209 ( .A(n106), .ZN(n534) );
  AOI22_X1 U210 ( .A1(in[255]), .A2(n571), .B1(out[255]), .B2(n591), .ZN(n106)
         );
  INV_X1 U211 ( .A(n107), .ZN(n533) );
  AOI22_X1 U212 ( .A1(in[254]), .A2(n571), .B1(out[254]), .B2(n591), .ZN(n107)
         );
  INV_X1 U213 ( .A(n108), .ZN(n532) );
  AOI22_X1 U214 ( .A1(in[253]), .A2(n571), .B1(out[253]), .B2(n591), .ZN(n108)
         );
  INV_X1 U215 ( .A(n109), .ZN(n531) );
  AOI22_X1 U216 ( .A1(in[252]), .A2(n571), .B1(out[252]), .B2(n591), .ZN(n109)
         );
  INV_X1 U217 ( .A(n110), .ZN(n530) );
  AOI22_X1 U218 ( .A1(in[251]), .A2(n571), .B1(out[251]), .B2(n592), .ZN(n110)
         );
  INV_X1 U219 ( .A(n111), .ZN(n529) );
  AOI22_X1 U220 ( .A1(in[250]), .A2(n571), .B1(out[250]), .B2(n592), .ZN(n111)
         );
  INV_X1 U221 ( .A(n112), .ZN(n303) );
  AOI22_X1 U222 ( .A1(in[24]), .A2(n571), .B1(out[24]), .B2(n592), .ZN(n112)
         );
  INV_X1 U223 ( .A(n113), .ZN(n528) );
  AOI22_X1 U224 ( .A1(in[249]), .A2(n571), .B1(out[249]), .B2(n592), .ZN(n113)
         );
  INV_X1 U225 ( .A(n114), .ZN(n527) );
  AOI22_X1 U226 ( .A1(in[248]), .A2(n570), .B1(out[248]), .B2(n592), .ZN(n114)
         );
  INV_X1 U227 ( .A(n115), .ZN(n526) );
  AOI22_X1 U228 ( .A1(in[247]), .A2(n570), .B1(out[247]), .B2(n592), .ZN(n115)
         );
  INV_X1 U229 ( .A(n116), .ZN(n525) );
  AOI22_X1 U230 ( .A1(in[246]), .A2(n570), .B1(out[246]), .B2(n592), .ZN(n116)
         );
  INV_X1 U231 ( .A(n117), .ZN(n524) );
  AOI22_X1 U232 ( .A1(in[245]), .A2(n570), .B1(out[245]), .B2(n592), .ZN(n117)
         );
  INV_X1 U233 ( .A(n118), .ZN(n523) );
  AOI22_X1 U234 ( .A1(in[244]), .A2(n570), .B1(out[244]), .B2(n592), .ZN(n118)
         );
  INV_X1 U235 ( .A(n119), .ZN(n522) );
  AOI22_X1 U236 ( .A1(in[243]), .A2(n570), .B1(out[243]), .B2(n592), .ZN(n119)
         );
  INV_X1 U237 ( .A(n120), .ZN(n521) );
  AOI22_X1 U238 ( .A1(in[242]), .A2(n570), .B1(out[242]), .B2(n592), .ZN(n120)
         );
  INV_X1 U239 ( .A(n121), .ZN(n520) );
  AOI22_X1 U240 ( .A1(in[241]), .A2(n570), .B1(out[241]), .B2(n592), .ZN(n121)
         );
  INV_X1 U241 ( .A(n122), .ZN(n519) );
  AOI22_X1 U242 ( .A1(in[240]), .A2(n570), .B1(out[240]), .B2(n593), .ZN(n122)
         );
  INV_X1 U243 ( .A(n123), .ZN(n302) );
  AOI22_X1 U244 ( .A1(in[23]), .A2(n570), .B1(out[23]), .B2(n593), .ZN(n123)
         );
  INV_X1 U245 ( .A(n124), .ZN(n518) );
  AOI22_X1 U246 ( .A1(in[239]), .A2(n570), .B1(out[239]), .B2(n593), .ZN(n124)
         );
  INV_X1 U247 ( .A(n125), .ZN(n517) );
  AOI22_X1 U248 ( .A1(in[238]), .A2(n569), .B1(out[238]), .B2(n593), .ZN(n125)
         );
  INV_X1 U249 ( .A(n126), .ZN(n516) );
  AOI22_X1 U250 ( .A1(in[237]), .A2(n569), .B1(out[237]), .B2(n593), .ZN(n126)
         );
  INV_X1 U251 ( .A(n127), .ZN(n515) );
  AOI22_X1 U252 ( .A1(in[236]), .A2(n569), .B1(out[236]), .B2(n593), .ZN(n127)
         );
  INV_X1 U253 ( .A(n128), .ZN(n514) );
  AOI22_X1 U254 ( .A1(in[235]), .A2(n569), .B1(out[235]), .B2(n593), .ZN(n128)
         );
  INV_X1 U255 ( .A(n129), .ZN(n513) );
  AOI22_X1 U256 ( .A1(in[234]), .A2(n569), .B1(out[234]), .B2(n593), .ZN(n129)
         );
  INV_X1 U257 ( .A(n130), .ZN(n512) );
  AOI22_X1 U258 ( .A1(in[233]), .A2(n569), .B1(out[233]), .B2(n593), .ZN(n130)
         );
  INV_X1 U259 ( .A(n131), .ZN(n511) );
  AOI22_X1 U260 ( .A1(in[232]), .A2(n569), .B1(out[232]), .B2(n593), .ZN(n131)
         );
  INV_X1 U261 ( .A(n132), .ZN(n510) );
  AOI22_X1 U262 ( .A1(in[231]), .A2(n569), .B1(out[231]), .B2(n593), .ZN(n132)
         );
  INV_X1 U263 ( .A(n133), .ZN(n509) );
  AOI22_X1 U264 ( .A1(in[230]), .A2(n569), .B1(out[230]), .B2(n593), .ZN(n133)
         );
  INV_X1 U265 ( .A(n134), .ZN(n301) );
  AOI22_X1 U266 ( .A1(in[22]), .A2(n569), .B1(out[22]), .B2(n594), .ZN(n134)
         );
  INV_X1 U267 ( .A(n135), .ZN(n508) );
  AOI22_X1 U268 ( .A1(in[229]), .A2(n569), .B1(out[229]), .B2(n594), .ZN(n135)
         );
  INV_X1 U269 ( .A(n136), .ZN(n507) );
  AOI22_X1 U270 ( .A1(in[228]), .A2(n568), .B1(out[228]), .B2(n594), .ZN(n136)
         );
  INV_X1 U271 ( .A(n137), .ZN(n506) );
  AOI22_X1 U272 ( .A1(in[227]), .A2(n568), .B1(out[227]), .B2(n594), .ZN(n137)
         );
  INV_X1 U273 ( .A(n138), .ZN(n505) );
  AOI22_X1 U274 ( .A1(in[226]), .A2(n568), .B1(out[226]), .B2(n594), .ZN(n138)
         );
  INV_X1 U275 ( .A(n139), .ZN(n504) );
  AOI22_X1 U276 ( .A1(in[225]), .A2(n568), .B1(out[225]), .B2(n594), .ZN(n139)
         );
  INV_X1 U277 ( .A(n140), .ZN(n503) );
  AOI22_X1 U278 ( .A1(in[224]), .A2(n568), .B1(out[224]), .B2(n594), .ZN(n140)
         );
  INV_X1 U279 ( .A(n141), .ZN(n502) );
  AOI22_X1 U280 ( .A1(in[223]), .A2(n568), .B1(out[223]), .B2(n594), .ZN(n141)
         );
  INV_X1 U281 ( .A(n142), .ZN(n501) );
  AOI22_X1 U282 ( .A1(in[222]), .A2(n568), .B1(out[222]), .B2(n594), .ZN(n142)
         );
  INV_X1 U283 ( .A(n143), .ZN(n500) );
  AOI22_X1 U284 ( .A1(in[221]), .A2(n568), .B1(out[221]), .B2(n594), .ZN(n143)
         );
  INV_X1 U285 ( .A(n144), .ZN(n499) );
  AOI22_X1 U286 ( .A1(in[220]), .A2(n568), .B1(out[220]), .B2(n594), .ZN(n144)
         );
  INV_X1 U287 ( .A(n145), .ZN(n300) );
  AOI22_X1 U288 ( .A1(in[21]), .A2(n568), .B1(out[21]), .B2(n594), .ZN(n145)
         );
  INV_X1 U289 ( .A(n146), .ZN(n498) );
  AOI22_X1 U290 ( .A1(in[219]), .A2(n568), .B1(out[219]), .B2(n595), .ZN(n146)
         );
  INV_X1 U291 ( .A(n147), .ZN(n497) );
  AOI22_X1 U292 ( .A1(in[218]), .A2(n567), .B1(out[218]), .B2(n595), .ZN(n147)
         );
  INV_X1 U293 ( .A(n148), .ZN(n496) );
  AOI22_X1 U294 ( .A1(in[217]), .A2(n567), .B1(out[217]), .B2(n595), .ZN(n148)
         );
  INV_X1 U295 ( .A(n149), .ZN(n495) );
  AOI22_X1 U296 ( .A1(in[216]), .A2(n567), .B1(out[216]), .B2(n595), .ZN(n149)
         );
  INV_X1 U297 ( .A(n150), .ZN(n494) );
  AOI22_X1 U298 ( .A1(in[215]), .A2(n567), .B1(out[215]), .B2(n595), .ZN(n150)
         );
  INV_X1 U299 ( .A(n151), .ZN(n493) );
  AOI22_X1 U300 ( .A1(in[214]), .A2(n567), .B1(out[214]), .B2(n595), .ZN(n151)
         );
  INV_X1 U301 ( .A(n152), .ZN(n492) );
  AOI22_X1 U302 ( .A1(in[213]), .A2(n567), .B1(out[213]), .B2(n595), .ZN(n152)
         );
  INV_X1 U303 ( .A(n153), .ZN(n491) );
  AOI22_X1 U304 ( .A1(in[212]), .A2(n567), .B1(out[212]), .B2(n595), .ZN(n153)
         );
  INV_X1 U305 ( .A(n154), .ZN(n490) );
  AOI22_X1 U306 ( .A1(in[211]), .A2(n567), .B1(out[211]), .B2(n595), .ZN(n154)
         );
  INV_X1 U307 ( .A(n155), .ZN(n489) );
  AOI22_X1 U308 ( .A1(in[210]), .A2(n567), .B1(out[210]), .B2(n595), .ZN(n155)
         );
  INV_X1 U309 ( .A(n156), .ZN(n299) );
  AOI22_X1 U310 ( .A1(in[20]), .A2(n567), .B1(out[20]), .B2(n595), .ZN(n156)
         );
  INV_X1 U311 ( .A(n157), .ZN(n488) );
  AOI22_X1 U312 ( .A1(in[209]), .A2(n567), .B1(out[209]), .B2(n595), .ZN(n157)
         );
  INV_X1 U313 ( .A(n158), .ZN(n487) );
  AOI22_X1 U314 ( .A1(in[208]), .A2(n566), .B1(out[208]), .B2(n596), .ZN(n158)
         );
  INV_X1 U315 ( .A(n159), .ZN(n486) );
  AOI22_X1 U316 ( .A1(in[207]), .A2(n566), .B1(out[207]), .B2(n596), .ZN(n159)
         );
  INV_X1 U317 ( .A(n160), .ZN(n485) );
  AOI22_X1 U318 ( .A1(in[206]), .A2(n566), .B1(out[206]), .B2(n596), .ZN(n160)
         );
  INV_X1 U319 ( .A(n161), .ZN(n484) );
  AOI22_X1 U320 ( .A1(in[205]), .A2(n566), .B1(out[205]), .B2(n596), .ZN(n161)
         );
  INV_X1 U321 ( .A(n162), .ZN(n483) );
  AOI22_X1 U322 ( .A1(in[204]), .A2(n566), .B1(out[204]), .B2(n596), .ZN(n162)
         );
  INV_X1 U323 ( .A(n163), .ZN(n482) );
  AOI22_X1 U324 ( .A1(in[203]), .A2(n566), .B1(out[203]), .B2(n596), .ZN(n163)
         );
  INV_X1 U325 ( .A(n164), .ZN(n481) );
  AOI22_X1 U326 ( .A1(in[202]), .A2(n566), .B1(out[202]), .B2(n596), .ZN(n164)
         );
  INV_X1 U327 ( .A(n165), .ZN(n480) );
  AOI22_X1 U328 ( .A1(in[201]), .A2(n566), .B1(out[201]), .B2(n596), .ZN(n165)
         );
  INV_X1 U329 ( .A(n166), .ZN(n479) );
  AOI22_X1 U330 ( .A1(in[200]), .A2(n566), .B1(out[200]), .B2(n596), .ZN(n166)
         );
  INV_X1 U331 ( .A(n167), .ZN(n280) );
  AOI22_X1 U332 ( .A1(in[1]), .A2(n566), .B1(out[1]), .B2(n596), .ZN(n167) );
  INV_X1 U333 ( .A(n168), .ZN(n298) );
  AOI22_X1 U334 ( .A1(in[19]), .A2(n566), .B1(out[19]), .B2(n596), .ZN(n168)
         );
  INV_X1 U335 ( .A(n169), .ZN(n478) );
  AOI22_X1 U336 ( .A1(in[199]), .A2(n565), .B1(out[199]), .B2(n596), .ZN(n169)
         );
  INV_X1 U337 ( .A(n170), .ZN(n477) );
  AOI22_X1 U338 ( .A1(in[198]), .A2(n565), .B1(out[198]), .B2(n597), .ZN(n170)
         );
  INV_X1 U339 ( .A(n171), .ZN(n476) );
  AOI22_X1 U340 ( .A1(in[197]), .A2(n565), .B1(out[197]), .B2(n597), .ZN(n171)
         );
  INV_X1 U341 ( .A(n172), .ZN(n475) );
  AOI22_X1 U342 ( .A1(in[196]), .A2(n565), .B1(out[196]), .B2(n597), .ZN(n172)
         );
  INV_X1 U343 ( .A(n173), .ZN(n474) );
  AOI22_X1 U344 ( .A1(in[195]), .A2(n565), .B1(out[195]), .B2(n597), .ZN(n173)
         );
  INV_X1 U345 ( .A(n174), .ZN(n473) );
  AOI22_X1 U346 ( .A1(in[194]), .A2(n565), .B1(out[194]), .B2(n597), .ZN(n174)
         );
  INV_X1 U347 ( .A(n175), .ZN(n472) );
  AOI22_X1 U348 ( .A1(in[193]), .A2(n565), .B1(out[193]), .B2(n597), .ZN(n175)
         );
  INV_X1 U349 ( .A(n176), .ZN(n471) );
  AOI22_X1 U350 ( .A1(in[192]), .A2(n565), .B1(out[192]), .B2(n597), .ZN(n176)
         );
  INV_X1 U351 ( .A(n177), .ZN(n470) );
  AOI22_X1 U352 ( .A1(in[191]), .A2(n565), .B1(out[191]), .B2(n597), .ZN(n177)
         );
  INV_X1 U353 ( .A(n178), .ZN(n469) );
  AOI22_X1 U354 ( .A1(in[190]), .A2(n565), .B1(out[190]), .B2(n597), .ZN(n178)
         );
  INV_X1 U355 ( .A(n179), .ZN(n297) );
  AOI22_X1 U356 ( .A1(in[18]), .A2(n565), .B1(out[18]), .B2(n597), .ZN(n179)
         );
  INV_X1 U357 ( .A(n180), .ZN(n468) );
  AOI22_X1 U358 ( .A1(in[189]), .A2(n564), .B1(out[189]), .B2(n597), .ZN(n180)
         );
  INV_X1 U359 ( .A(n181), .ZN(n467) );
  AOI22_X1 U360 ( .A1(in[188]), .A2(n564), .B1(out[188]), .B2(n597), .ZN(n181)
         );
  INV_X1 U361 ( .A(n182), .ZN(n466) );
  AOI22_X1 U362 ( .A1(in[187]), .A2(n564), .B1(out[187]), .B2(n598), .ZN(n182)
         );
  INV_X1 U363 ( .A(n183), .ZN(n465) );
  AOI22_X1 U364 ( .A1(in[186]), .A2(n564), .B1(out[186]), .B2(n598), .ZN(n183)
         );
  INV_X1 U365 ( .A(n184), .ZN(n464) );
  AOI22_X1 U366 ( .A1(in[185]), .A2(n564), .B1(out[185]), .B2(n598), .ZN(n184)
         );
  INV_X1 U367 ( .A(n185), .ZN(n463) );
  AOI22_X1 U368 ( .A1(in[184]), .A2(n564), .B1(out[184]), .B2(n598), .ZN(n185)
         );
  INV_X1 U369 ( .A(n186), .ZN(n462) );
  AOI22_X1 U370 ( .A1(in[183]), .A2(n564), .B1(out[183]), .B2(n598), .ZN(n186)
         );
  INV_X1 U371 ( .A(n187), .ZN(n461) );
  AOI22_X1 U372 ( .A1(in[182]), .A2(n564), .B1(out[182]), .B2(n598), .ZN(n187)
         );
  INV_X1 U373 ( .A(n188), .ZN(n460) );
  AOI22_X1 U374 ( .A1(in[181]), .A2(n564), .B1(out[181]), .B2(n598), .ZN(n188)
         );
  INV_X1 U375 ( .A(n189), .ZN(n459) );
  AOI22_X1 U376 ( .A1(in[180]), .A2(n564), .B1(out[180]), .B2(n598), .ZN(n189)
         );
  INV_X1 U377 ( .A(n190), .ZN(n296) );
  AOI22_X1 U378 ( .A1(in[17]), .A2(n564), .B1(out[17]), .B2(n598), .ZN(n190)
         );
  INV_X1 U379 ( .A(n191), .ZN(n458) );
  AOI22_X1 U380 ( .A1(in[179]), .A2(n563), .B1(out[179]), .B2(n598), .ZN(n191)
         );
  INV_X1 U381 ( .A(n192), .ZN(n457) );
  AOI22_X1 U382 ( .A1(in[178]), .A2(n563), .B1(out[178]), .B2(n598), .ZN(n192)
         );
  INV_X1 U383 ( .A(n193), .ZN(n456) );
  AOI22_X1 U384 ( .A1(in[177]), .A2(n563), .B1(out[177]), .B2(n598), .ZN(n193)
         );
  INV_X1 U385 ( .A(n194), .ZN(n455) );
  AOI22_X1 U386 ( .A1(in[176]), .A2(n563), .B1(out[176]), .B2(n599), .ZN(n194)
         );
  INV_X1 U387 ( .A(n195), .ZN(n454) );
  AOI22_X1 U388 ( .A1(in[175]), .A2(n563), .B1(out[175]), .B2(n599), .ZN(n195)
         );
  INV_X1 U389 ( .A(n196), .ZN(n453) );
  AOI22_X1 U390 ( .A1(in[174]), .A2(n563), .B1(out[174]), .B2(n599), .ZN(n196)
         );
  INV_X1 U391 ( .A(n197), .ZN(n452) );
  AOI22_X1 U392 ( .A1(in[173]), .A2(n563), .B1(out[173]), .B2(n599), .ZN(n197)
         );
  INV_X1 U393 ( .A(n198), .ZN(n451) );
  AOI22_X1 U394 ( .A1(in[172]), .A2(n563), .B1(out[172]), .B2(n599), .ZN(n198)
         );
  INV_X1 U395 ( .A(n199), .ZN(n450) );
  AOI22_X1 U396 ( .A1(in[171]), .A2(n563), .B1(out[171]), .B2(n599), .ZN(n199)
         );
  INV_X1 U397 ( .A(n200), .ZN(n449) );
  AOI22_X1 U398 ( .A1(in[170]), .A2(n563), .B1(out[170]), .B2(n599), .ZN(n200)
         );
  INV_X1 U399 ( .A(n201), .ZN(n295) );
  AOI22_X1 U400 ( .A1(in[16]), .A2(n563), .B1(out[16]), .B2(n599), .ZN(n201)
         );
  INV_X1 U401 ( .A(n202), .ZN(n448) );
  AOI22_X1 U402 ( .A1(in[169]), .A2(n562), .B1(out[169]), .B2(n599), .ZN(n202)
         );
  INV_X1 U403 ( .A(n203), .ZN(n447) );
  AOI22_X1 U404 ( .A1(in[168]), .A2(n562), .B1(out[168]), .B2(n599), .ZN(n203)
         );
  INV_X1 U405 ( .A(n204), .ZN(n446) );
  AOI22_X1 U406 ( .A1(in[167]), .A2(n562), .B1(out[167]), .B2(n599), .ZN(n204)
         );
  INV_X1 U407 ( .A(n205), .ZN(n445) );
  AOI22_X1 U408 ( .A1(in[166]), .A2(n562), .B1(out[166]), .B2(n599), .ZN(n205)
         );
  INV_X1 U409 ( .A(n206), .ZN(n444) );
  AOI22_X1 U410 ( .A1(in[165]), .A2(n562), .B1(out[165]), .B2(n600), .ZN(n206)
         );
  INV_X1 U411 ( .A(n207), .ZN(n443) );
  AOI22_X1 U412 ( .A1(in[164]), .A2(n562), .B1(out[164]), .B2(n600), .ZN(n207)
         );
  INV_X1 U413 ( .A(n208), .ZN(n442) );
  AOI22_X1 U414 ( .A1(in[163]), .A2(n562), .B1(out[163]), .B2(n600), .ZN(n208)
         );
  INV_X1 U415 ( .A(n209), .ZN(n441) );
  AOI22_X1 U416 ( .A1(in[162]), .A2(n562), .B1(out[162]), .B2(n600), .ZN(n209)
         );
  INV_X1 U417 ( .A(n210), .ZN(n440) );
  AOI22_X1 U418 ( .A1(in[161]), .A2(n562), .B1(out[161]), .B2(n600), .ZN(n210)
         );
  INV_X1 U419 ( .A(n211), .ZN(n439) );
  AOI22_X1 U420 ( .A1(in[160]), .A2(n562), .B1(out[160]), .B2(n600), .ZN(n211)
         );
  INV_X1 U421 ( .A(n212), .ZN(n294) );
  AOI22_X1 U422 ( .A1(in[15]), .A2(n562), .B1(out[15]), .B2(n600), .ZN(n212)
         );
  INV_X1 U423 ( .A(n213), .ZN(n438) );
  AOI22_X1 U424 ( .A1(in[159]), .A2(n561), .B1(out[159]), .B2(n600), .ZN(n213)
         );
  INV_X1 U425 ( .A(n214), .ZN(n437) );
  AOI22_X1 U426 ( .A1(in[158]), .A2(n561), .B1(out[158]), .B2(n600), .ZN(n214)
         );
  INV_X1 U427 ( .A(n215), .ZN(n436) );
  AOI22_X1 U428 ( .A1(in[157]), .A2(n561), .B1(out[157]), .B2(n600), .ZN(n215)
         );
  INV_X1 U429 ( .A(n216), .ZN(n435) );
  AOI22_X1 U430 ( .A1(in[156]), .A2(n561), .B1(out[156]), .B2(n600), .ZN(n216)
         );
  INV_X1 U431 ( .A(n217), .ZN(n434) );
  AOI22_X1 U432 ( .A1(in[155]), .A2(n561), .B1(out[155]), .B2(n600), .ZN(n217)
         );
  INV_X1 U433 ( .A(n218), .ZN(n433) );
  AOI22_X1 U434 ( .A1(in[154]), .A2(n561), .B1(out[154]), .B2(n601), .ZN(n218)
         );
  INV_X1 U435 ( .A(n219), .ZN(n432) );
  AOI22_X1 U436 ( .A1(in[153]), .A2(n561), .B1(out[153]), .B2(n601), .ZN(n219)
         );
  INV_X1 U437 ( .A(n220), .ZN(n431) );
  AOI22_X1 U438 ( .A1(in[152]), .A2(n561), .B1(out[152]), .B2(n601), .ZN(n220)
         );
  INV_X1 U439 ( .A(n221), .ZN(n430) );
  AOI22_X1 U440 ( .A1(in[151]), .A2(n561), .B1(out[151]), .B2(n601), .ZN(n221)
         );
  INV_X1 U441 ( .A(n222), .ZN(n429) );
  AOI22_X1 U442 ( .A1(in[150]), .A2(n561), .B1(out[150]), .B2(n601), .ZN(n222)
         );
  INV_X1 U443 ( .A(n223), .ZN(n293) );
  AOI22_X1 U444 ( .A1(in[14]), .A2(n561), .B1(out[14]), .B2(n601), .ZN(n223)
         );
  INV_X1 U445 ( .A(n224), .ZN(n428) );
  AOI22_X1 U446 ( .A1(in[149]), .A2(n560), .B1(out[149]), .B2(n601), .ZN(n224)
         );
  INV_X1 U447 ( .A(n225), .ZN(n427) );
  AOI22_X1 U448 ( .A1(in[148]), .A2(n560), .B1(out[148]), .B2(n601), .ZN(n225)
         );
  INV_X1 U449 ( .A(n226), .ZN(n426) );
  AOI22_X1 U450 ( .A1(in[147]), .A2(n560), .B1(out[147]), .B2(n601), .ZN(n226)
         );
  INV_X1 U451 ( .A(n227), .ZN(n425) );
  AOI22_X1 U452 ( .A1(in[146]), .A2(n560), .B1(out[146]), .B2(n601), .ZN(n227)
         );
  INV_X1 U453 ( .A(n228), .ZN(n424) );
  AOI22_X1 U454 ( .A1(in[145]), .A2(n560), .B1(out[145]), .B2(n601), .ZN(n228)
         );
  INV_X1 U455 ( .A(n229), .ZN(n423) );
  AOI22_X1 U456 ( .A1(in[144]), .A2(n560), .B1(out[144]), .B2(n601), .ZN(n229)
         );
  INV_X1 U457 ( .A(n230), .ZN(n422) );
  AOI22_X1 U458 ( .A1(in[143]), .A2(n560), .B1(out[143]), .B2(n602), .ZN(n230)
         );
  INV_X1 U459 ( .A(n231), .ZN(n421) );
  AOI22_X1 U460 ( .A1(in[142]), .A2(n560), .B1(out[142]), .B2(n602), .ZN(n231)
         );
  INV_X1 U461 ( .A(n232), .ZN(n420) );
  AOI22_X1 U462 ( .A1(in[141]), .A2(n560), .B1(out[141]), .B2(n602), .ZN(n232)
         );
  INV_X1 U463 ( .A(n233), .ZN(n419) );
  AOI22_X1 U464 ( .A1(in[140]), .A2(n560), .B1(out[140]), .B2(n602), .ZN(n233)
         );
  INV_X1 U465 ( .A(n234), .ZN(n292) );
  AOI22_X1 U466 ( .A1(in[13]), .A2(n560), .B1(out[13]), .B2(n602), .ZN(n234)
         );
  INV_X1 U467 ( .A(n235), .ZN(n418) );
  AOI22_X1 U468 ( .A1(in[139]), .A2(n559), .B1(out[139]), .B2(n602), .ZN(n235)
         );
  INV_X1 U469 ( .A(n236), .ZN(n417) );
  AOI22_X1 U470 ( .A1(in[138]), .A2(n559), .B1(out[138]), .B2(n602), .ZN(n236)
         );
  INV_X1 U471 ( .A(n237), .ZN(n416) );
  AOI22_X1 U472 ( .A1(in[137]), .A2(n559), .B1(out[137]), .B2(n602), .ZN(n237)
         );
  INV_X1 U473 ( .A(n238), .ZN(n415) );
  AOI22_X1 U474 ( .A1(in[136]), .A2(n559), .B1(out[136]), .B2(n602), .ZN(n238)
         );
  INV_X1 U475 ( .A(n239), .ZN(n414) );
  AOI22_X1 U476 ( .A1(in[135]), .A2(n559), .B1(out[135]), .B2(n602), .ZN(n239)
         );
  INV_X1 U477 ( .A(n240), .ZN(n413) );
  AOI22_X1 U478 ( .A1(in[134]), .A2(n559), .B1(out[134]), .B2(n602), .ZN(n240)
         );
  INV_X1 U479 ( .A(n241), .ZN(n412) );
  AOI22_X1 U480 ( .A1(in[133]), .A2(n559), .B1(out[133]), .B2(n602), .ZN(n241)
         );
  INV_X1 U481 ( .A(n242), .ZN(n411) );
  AOI22_X1 U482 ( .A1(in[132]), .A2(n559), .B1(out[132]), .B2(n603), .ZN(n242)
         );
  INV_X1 U483 ( .A(n243), .ZN(n410) );
  AOI22_X1 U484 ( .A1(in[131]), .A2(n559), .B1(out[131]), .B2(n603), .ZN(n243)
         );
  INV_X1 U485 ( .A(n244), .ZN(n409) );
  AOI22_X1 U486 ( .A1(in[130]), .A2(n559), .B1(out[130]), .B2(n603), .ZN(n244)
         );
  INV_X1 U487 ( .A(n245), .ZN(n291) );
  AOI22_X1 U488 ( .A1(in[12]), .A2(n559), .B1(out[12]), .B2(n603), .ZN(n245)
         );
  INV_X1 U489 ( .A(n246), .ZN(n408) );
  AOI22_X1 U490 ( .A1(in[129]), .A2(n558), .B1(out[129]), .B2(n603), .ZN(n246)
         );
  INV_X1 U491 ( .A(n247), .ZN(n407) );
  AOI22_X1 U492 ( .A1(in[128]), .A2(n558), .B1(out[128]), .B2(n603), .ZN(n247)
         );
  INV_X1 U493 ( .A(n248), .ZN(n406) );
  AOI22_X1 U494 ( .A1(in[127]), .A2(n558), .B1(out[127]), .B2(n603), .ZN(n248)
         );
  INV_X1 U495 ( .A(n249), .ZN(n405) );
  AOI22_X1 U496 ( .A1(in[126]), .A2(n558), .B1(out[126]), .B2(n603), .ZN(n249)
         );
  INV_X1 U497 ( .A(n250), .ZN(n404) );
  AOI22_X1 U498 ( .A1(in[125]), .A2(n558), .B1(out[125]), .B2(n603), .ZN(n250)
         );
  INV_X1 U499 ( .A(n251), .ZN(n403) );
  AOI22_X1 U500 ( .A1(in[124]), .A2(n558), .B1(out[124]), .B2(n603), .ZN(n251)
         );
  INV_X1 U501 ( .A(n252), .ZN(n402) );
  AOI22_X1 U502 ( .A1(in[123]), .A2(n558), .B1(out[123]), .B2(n603), .ZN(n252)
         );
  INV_X1 U503 ( .A(n253), .ZN(n401) );
  AOI22_X1 U504 ( .A1(in[122]), .A2(n558), .B1(out[122]), .B2(n603), .ZN(n253)
         );
  INV_X1 U505 ( .A(n254), .ZN(n400) );
  AOI22_X1 U506 ( .A1(in[121]), .A2(n558), .B1(out[121]), .B2(n604), .ZN(n254)
         );
  INV_X1 U507 ( .A(n255), .ZN(n399) );
  AOI22_X1 U508 ( .A1(in[120]), .A2(n558), .B1(out[120]), .B2(n604), .ZN(n255)
         );
  INV_X1 U509 ( .A(n256), .ZN(n290) );
  AOI22_X1 U510 ( .A1(in[11]), .A2(n558), .B1(out[11]), .B2(n604), .ZN(n256)
         );
  INV_X1 U511 ( .A(n257), .ZN(n398) );
  AOI22_X1 U512 ( .A1(in[119]), .A2(n557), .B1(out[119]), .B2(n604), .ZN(n257)
         );
  INV_X1 U513 ( .A(n258), .ZN(n397) );
  AOI22_X1 U514 ( .A1(in[118]), .A2(n557), .B1(out[118]), .B2(n604), .ZN(n258)
         );
  INV_X1 U515 ( .A(n259), .ZN(n396) );
  AOI22_X1 U516 ( .A1(in[117]), .A2(n557), .B1(out[117]), .B2(n604), .ZN(n259)
         );
  INV_X1 U517 ( .A(n260), .ZN(n395) );
  AOI22_X1 U518 ( .A1(in[116]), .A2(n557), .B1(out[116]), .B2(n604), .ZN(n260)
         );
  INV_X1 U519 ( .A(n261), .ZN(n394) );
  AOI22_X1 U520 ( .A1(in[115]), .A2(n557), .B1(out[115]), .B2(n604), .ZN(n261)
         );
  INV_X1 U521 ( .A(n262), .ZN(n393) );
  AOI22_X1 U522 ( .A1(in[114]), .A2(n557), .B1(out[114]), .B2(n604), .ZN(n262)
         );
  INV_X1 U523 ( .A(n263), .ZN(n392) );
  AOI22_X1 U524 ( .A1(in[113]), .A2(n557), .B1(out[113]), .B2(n604), .ZN(n263)
         );
  INV_X1 U525 ( .A(n264), .ZN(n391) );
  AOI22_X1 U526 ( .A1(in[112]), .A2(n557), .B1(out[112]), .B2(n604), .ZN(n264)
         );
  INV_X1 U527 ( .A(n265), .ZN(n390) );
  AOI22_X1 U528 ( .A1(in[111]), .A2(n557), .B1(out[111]), .B2(n604), .ZN(n265)
         );
  INV_X1 U529 ( .A(n266), .ZN(n389) );
  AOI22_X1 U530 ( .A1(in[110]), .A2(n557), .B1(out[110]), .B2(n592), .ZN(n266)
         );
  INV_X1 U531 ( .A(n267), .ZN(n289) );
  AOI22_X1 U532 ( .A1(in[10]), .A2(n557), .B1(out[10]), .B2(n593), .ZN(n267)
         );
  INV_X1 U533 ( .A(n268), .ZN(n388) );
  AOI22_X1 U534 ( .A1(in[109]), .A2(n556), .B1(out[109]), .B2(n594), .ZN(n268)
         );
  INV_X1 U535 ( .A(n269), .ZN(n387) );
  AOI22_X1 U536 ( .A1(in[108]), .A2(n556), .B1(out[108]), .B2(n595), .ZN(n269)
         );
  INV_X1 U537 ( .A(n270), .ZN(n386) );
  AOI22_X1 U538 ( .A1(in[107]), .A2(n556), .B1(out[107]), .B2(n596), .ZN(n270)
         );
  INV_X1 U539 ( .A(n271), .ZN(n385) );
  AOI22_X1 U540 ( .A1(in[106]), .A2(n556), .B1(out[106]), .B2(n597), .ZN(n271)
         );
  INV_X1 U541 ( .A(n272), .ZN(n384) );
  AOI22_X1 U542 ( .A1(in[105]), .A2(n556), .B1(out[105]), .B2(n598), .ZN(n272)
         );
  INV_X1 U543 ( .A(n273), .ZN(n383) );
  AOI22_X1 U544 ( .A1(in[104]), .A2(n556), .B1(out[104]), .B2(n599), .ZN(n273)
         );
  INV_X1 U545 ( .A(n274), .ZN(n382) );
  AOI22_X1 U546 ( .A1(in[103]), .A2(n556), .B1(out[103]), .B2(n600), .ZN(n274)
         );
  INV_X1 U547 ( .A(n275), .ZN(n381) );
  AOI22_X1 U548 ( .A1(in[102]), .A2(n556), .B1(out[102]), .B2(n601), .ZN(n275)
         );
  INV_X1 U549 ( .A(n276), .ZN(n380) );
  AOI22_X1 U550 ( .A1(in[101]), .A2(n556), .B1(out[101]), .B2(n602), .ZN(n276)
         );
  INV_X1 U551 ( .A(n277), .ZN(n379) );
  AOI22_X1 U552 ( .A1(in[100]), .A2(n556), .B1(out[100]), .B2(n603), .ZN(n277)
         );
  INV_X1 U553 ( .A(n278), .ZN(n279) );
  AOI22_X1 U554 ( .A1(in[0]), .A2(n556), .B1(out[0]), .B2(n604), .ZN(n278) );
  BUF_X4 U556 ( .A(n2), .Z(n583) );
  BUF_X4 U557 ( .A(n2), .Z(n582) );
  BUF_X4 U558 ( .A(n585), .Z(n574) );
  BUF_X4 U559 ( .A(we), .Z(n588) );
  BUF_X4 U560 ( .A(n581), .Z(n575) );
  BUF_X4 U561 ( .A(we), .Z(n587) );
  BUF_X4 U562 ( .A(n581), .Z(n576) );
  BUF_X4 U563 ( .A(n581), .Z(n577) );
  BUF_X4 U564 ( .A(n581), .Z(n578) );
  BUF_X4 U565 ( .A(n581), .Z(n579) );
  BUF_X4 U566 ( .A(n581), .Z(n580) );
  BUF_X4 U567 ( .A(we), .Z(n586) );
  BUF_X4 U568 ( .A(n585), .Z(n558) );
  BUF_X4 U569 ( .A(n585), .Z(n559) );
  BUF_X4 U570 ( .A(n585), .Z(n560) );
  BUF_X4 U571 ( .A(n584), .Z(n561) );
  BUF_X4 U572 ( .A(we), .Z(n600) );
  BUF_X4 U573 ( .A(n584), .Z(n562) );
  BUF_X4 U574 ( .A(we), .Z(n599) );
  BUF_X4 U575 ( .A(n584), .Z(n563) );
  BUF_X4 U576 ( .A(we), .Z(n598) );
  BUF_X4 U577 ( .A(n583), .Z(n564) );
  BUF_X4 U578 ( .A(we), .Z(n597) );
  BUF_X4 U579 ( .A(n583), .Z(n565) );
  BUF_X4 U580 ( .A(n583), .Z(n566) );
  BUF_X4 U581 ( .A(we), .Z(n596) );
  BUF_X4 U582 ( .A(n582), .Z(n567) );
  BUF_X4 U583 ( .A(we), .Z(n595) );
  BUF_X4 U584 ( .A(n582), .Z(n568) );
  BUF_X4 U585 ( .A(we), .Z(n594) );
  BUF_X4 U586 ( .A(n582), .Z(n569) );
  BUF_X4 U587 ( .A(we), .Z(n593) );
  BUF_X4 U588 ( .A(n584), .Z(n570) );
  BUF_X4 U589 ( .A(we), .Z(n592) );
  BUF_X4 U590 ( .A(n585), .Z(n571) );
  BUF_X4 U591 ( .A(we), .Z(n591) );
  BUF_X4 U592 ( .A(n581), .Z(n572) );
  BUF_X4 U593 ( .A(we), .Z(n590) );
  BUF_X4 U594 ( .A(n584), .Z(n573) );
  BUF_X4 U595 ( .A(we), .Z(n589) );
  BUF_X4 U596 ( .A(reset), .Z(n614) );
  BUF_X4 U597 ( .A(reset), .Z(n615) );
  BUF_X4 U598 ( .A(reset), .Z(n616) );
  BUF_X4 U599 ( .A(reset), .Z(n605) );
  BUF_X4 U600 ( .A(reset), .Z(n617) );
  BUF_X4 U601 ( .A(reset), .Z(n606) );
  BUF_X4 U602 ( .A(reset), .Z(n607) );
  BUF_X4 U603 ( .A(reset), .Z(n608) );
  BUF_X4 U604 ( .A(reset), .Z(n609) );
  BUF_X4 U605 ( .A(reset), .Z(n610) );
  BUF_X4 U606 ( .A(reset), .Z(n618) );
  BUF_X4 U607 ( .A(reset), .Z(n619) );
  BUF_X4 U608 ( .A(reset), .Z(n613) );
  BUF_X4 U609 ( .A(reset), .Z(n612) );
  BUF_X4 U610 ( .A(reset), .Z(n611) );
  BUF_X4 U611 ( .A(n2), .Z(n581) );
  BUF_X4 U612 ( .A(n585), .Z(n556) );
  BUF_X4 U613 ( .A(n584), .Z(n557) );
  BUF_X4 U614 ( .A(we), .Z(n604) );
  BUF_X4 U615 ( .A(we), .Z(n603) );
  BUF_X4 U616 ( .A(we), .Z(n602) );
  BUF_X4 U617 ( .A(we), .Z(n601) );
  BUF_X4 U618 ( .A(reset), .Z(n623) );
  BUF_X4 U619 ( .A(reset), .Z(n622) );
  BUF_X4 U620 ( .A(reset), .Z(n621) );
  BUF_X4 U621 ( .A(reset), .Z(n620) );
  NOR2_X2 U622 ( .A1(we), .A2(flush), .ZN(n2) );
  BUF_X4 U623 ( .A(n2), .Z(n585) );
  BUF_X4 U624 ( .A(n2), .Z(n584) );
endmodule

