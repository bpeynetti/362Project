
module register_file ( rd, ra, rb, busW, clk, writeEnable, reset, busA, busB
 );
  input [0:4] rd;
  input [0:4] ra;
  input [0:4] rb;
  input [0:31] busW;
  output [0:31] busA;
  output [0:31] busB;
  input clk, writeEnable, reset;
  wire   \reg_out[1][0] , \reg_out[1][1] , \reg_out[1][2] , \reg_out[1][3] ,
         \reg_out[1][4] , \reg_out[1][5] , \reg_out[1][6] , \reg_out[1][7] ,
         \reg_out[1][8] , \reg_out[1][9] , \reg_out[1][10] , \reg_out[1][11] ,
         \reg_out[1][12] , \reg_out[1][13] , \reg_out[1][14] ,
         \reg_out[1][15] , \reg_out[1][16] , \reg_out[1][17] ,
         \reg_out[1][18] , \reg_out[1][19] , \reg_out[1][20] ,
         \reg_out[1][21] , \reg_out[1][22] , \reg_out[1][23] ,
         \reg_out[1][24] , \reg_out[1][25] , \reg_out[1][26] ,
         \reg_out[1][27] , \reg_out[1][28] , \reg_out[1][29] ,
         \reg_out[1][30] , \reg_out[1][31] , \reg_out[3][0] , \reg_out[3][1] ,
         \reg_out[3][2] , \reg_out[3][3] , \reg_out[3][4] , \reg_out[3][5] ,
         \reg_out[3][6] , \reg_out[3][7] , \reg_out[3][8] , \reg_out[3][9] ,
         \reg_out[3][10] , \reg_out[3][11] , \reg_out[3][12] ,
         \reg_out[3][13] , \reg_out[3][14] , \reg_out[3][15] ,
         \reg_out[3][16] , \reg_out[3][17] , \reg_out[3][18] ,
         \reg_out[3][19] , \reg_out[3][20] , \reg_out[3][21] ,
         \reg_out[3][22] , \reg_out[3][23] , \reg_out[3][24] ,
         \reg_out[3][25] , \reg_out[3][26] , \reg_out[3][27] ,
         \reg_out[3][28] , \reg_out[3][29] , \reg_out[3][30] ,
         \reg_out[3][31] , \reg_out[5][0] , \reg_out[5][1] , \reg_out[5][2] ,
         \reg_out[5][3] , \reg_out[5][4] , \reg_out[5][5] , \reg_out[5][6] ,
         \reg_out[5][7] , \reg_out[5][8] , \reg_out[5][9] , \reg_out[5][10] ,
         \reg_out[5][11] , \reg_out[5][12] , \reg_out[5][13] ,
         \reg_out[5][14] , \reg_out[5][15] , \reg_out[5][16] ,
         \reg_out[5][17] , \reg_out[5][18] , \reg_out[5][19] ,
         \reg_out[5][20] , \reg_out[5][21] , \reg_out[5][22] ,
         \reg_out[5][23] , \reg_out[5][24] , \reg_out[5][25] ,
         \reg_out[5][26] , \reg_out[5][27] , \reg_out[5][28] ,
         \reg_out[5][29] , \reg_out[5][30] , \reg_out[5][31] , \reg_out[7][0] ,
         \reg_out[7][1] , \reg_out[7][2] , \reg_out[7][3] , \reg_out[7][4] ,
         \reg_out[7][5] , \reg_out[7][6] , \reg_out[7][7] , \reg_out[7][8] ,
         \reg_out[7][9] , \reg_out[7][10] , \reg_out[7][11] , \reg_out[7][12] ,
         \reg_out[7][13] , \reg_out[7][14] , \reg_out[7][15] ,
         \reg_out[7][16] , \reg_out[7][17] , \reg_out[7][18] ,
         \reg_out[7][19] , \reg_out[7][20] , \reg_out[7][21] ,
         \reg_out[7][22] , \reg_out[7][23] , \reg_out[7][24] ,
         \reg_out[7][25] , \reg_out[7][26] , \reg_out[7][27] ,
         \reg_out[7][28] , \reg_out[7][29] , \reg_out[7][30] ,
         \reg_out[7][31] , \reg_out[9][0] , \reg_out[9][1] , \reg_out[9][2] ,
         \reg_out[9][3] , \reg_out[9][4] , \reg_out[9][5] , \reg_out[9][6] ,
         \reg_out[9][7] , \reg_out[9][8] , \reg_out[9][9] , \reg_out[9][10] ,
         \reg_out[9][11] , \reg_out[9][12] , \reg_out[9][13] ,
         \reg_out[9][14] , \reg_out[9][15] , \reg_out[9][16] ,
         \reg_out[9][17] , \reg_out[9][18] , \reg_out[9][19] ,
         \reg_out[9][20] , \reg_out[9][21] , \reg_out[9][22] ,
         \reg_out[9][23] , \reg_out[9][24] , \reg_out[9][25] ,
         \reg_out[9][26] , \reg_out[9][27] , \reg_out[9][28] ,
         \reg_out[9][29] , \reg_out[9][30] , \reg_out[9][31] ,
         \reg_out[11][0] , \reg_out[11][1] , \reg_out[11][2] ,
         \reg_out[11][3] , \reg_out[11][4] , \reg_out[11][5] ,
         \reg_out[11][6] , \reg_out[11][7] , \reg_out[11][8] ,
         \reg_out[11][9] , \reg_out[11][10] , \reg_out[11][11] ,
         \reg_out[11][12] , \reg_out[11][13] , \reg_out[11][14] ,
         \reg_out[11][15] , \reg_out[11][16] , \reg_out[11][17] ,
         \reg_out[11][18] , \reg_out[11][19] , \reg_out[11][20] ,
         \reg_out[11][21] , \reg_out[11][22] , \reg_out[11][23] ,
         \reg_out[11][24] , \reg_out[11][25] , \reg_out[11][26] ,
         \reg_out[11][27] , \reg_out[11][28] , \reg_out[11][29] ,
         \reg_out[11][30] , \reg_out[11][31] , \reg_out[13][0] ,
         \reg_out[13][1] , \reg_out[13][2] , \reg_out[13][3] ,
         \reg_out[13][4] , \reg_out[13][5] , \reg_out[13][6] ,
         \reg_out[13][7] , \reg_out[13][8] , \reg_out[13][9] ,
         \reg_out[13][10] , \reg_out[13][11] , \reg_out[13][12] ,
         \reg_out[13][13] , \reg_out[13][14] , \reg_out[13][15] ,
         \reg_out[13][16] , \reg_out[13][17] , \reg_out[13][18] ,
         \reg_out[13][19] , \reg_out[13][20] , \reg_out[13][21] ,
         \reg_out[13][22] , \reg_out[13][23] , \reg_out[13][24] ,
         \reg_out[13][25] , \reg_out[13][26] , \reg_out[13][27] ,
         \reg_out[13][28] , \reg_out[13][29] , \reg_out[13][30] ,
         \reg_out[13][31] , \reg_out[15][0] , \reg_out[15][1] ,
         \reg_out[15][2] , \reg_out[15][3] , \reg_out[15][4] ,
         \reg_out[15][5] , \reg_out[15][6] , \reg_out[15][7] ,
         \reg_out[15][8] , \reg_out[15][9] , \reg_out[15][10] ,
         \reg_out[15][11] , \reg_out[15][12] , \reg_out[15][13] ,
         \reg_out[15][14] , \reg_out[15][15] , \reg_out[15][16] ,
         \reg_out[15][17] , \reg_out[15][18] , \reg_out[15][19] ,
         \reg_out[15][20] , \reg_out[15][21] , \reg_out[15][22] ,
         \reg_out[15][23] , \reg_out[15][24] , \reg_out[15][25] ,
         \reg_out[15][26] , \reg_out[15][27] , \reg_out[15][28] ,
         \reg_out[15][29] , \reg_out[15][30] , \reg_out[15][31] ,
         \reg_out[17][0] , \reg_out[17][1] , \reg_out[17][2] ,
         \reg_out[17][3] , \reg_out[17][4] , \reg_out[17][5] ,
         \reg_out[17][6] , \reg_out[17][7] , \reg_out[17][8] ,
         \reg_out[17][9] , \reg_out[17][10] , \reg_out[17][11] ,
         \reg_out[17][12] , \reg_out[17][13] , \reg_out[17][14] ,
         \reg_out[17][15] , \reg_out[17][16] , \reg_out[17][17] ,
         \reg_out[17][18] , \reg_out[17][19] , \reg_out[17][20] ,
         \reg_out[17][21] , \reg_out[17][22] , \reg_out[17][23] ,
         \reg_out[17][24] , \reg_out[17][25] , \reg_out[17][26] ,
         \reg_out[17][27] , \reg_out[17][28] , \reg_out[17][29] ,
         \reg_out[17][30] , \reg_out[17][31] , \reg_out[19][0] ,
         \reg_out[19][1] , \reg_out[19][2] , \reg_out[19][3] ,
         \reg_out[19][4] , \reg_out[19][5] , \reg_out[19][6] ,
         \reg_out[19][7] , \reg_out[19][8] , \reg_out[19][9] ,
         \reg_out[19][10] , \reg_out[19][11] , \reg_out[19][12] ,
         \reg_out[19][13] , \reg_out[19][14] , \reg_out[19][15] ,
         \reg_out[19][16] , \reg_out[19][17] , \reg_out[19][18] ,
         \reg_out[19][19] , \reg_out[19][20] , \reg_out[19][21] ,
         \reg_out[19][22] , \reg_out[19][23] , \reg_out[19][24] ,
         \reg_out[19][25] , \reg_out[19][26] , \reg_out[19][27] ,
         \reg_out[19][28] , \reg_out[19][29] , \reg_out[19][30] ,
         \reg_out[19][31] , \reg_out[21][0] , \reg_out[21][1] ,
         \reg_out[21][2] , \reg_out[21][3] , \reg_out[21][4] ,
         \reg_out[21][5] , \reg_out[21][6] , \reg_out[21][7] ,
         \reg_out[21][8] , \reg_out[21][9] , \reg_out[21][10] ,
         \reg_out[21][11] , \reg_out[21][12] , \reg_out[21][13] ,
         \reg_out[21][14] , \reg_out[21][15] , \reg_out[21][16] ,
         \reg_out[21][17] , \reg_out[21][18] , \reg_out[21][19] ,
         \reg_out[21][20] , \reg_out[21][21] , \reg_out[21][22] ,
         \reg_out[21][23] , \reg_out[21][24] , \reg_out[21][25] ,
         \reg_out[21][26] , \reg_out[21][27] , \reg_out[21][28] ,
         \reg_out[21][29] , \reg_out[21][30] , \reg_out[21][31] ,
         \reg_out[23][0] , \reg_out[23][1] , \reg_out[23][2] ,
         \reg_out[23][3] , \reg_out[23][4] , \reg_out[23][5] ,
         \reg_out[23][6] , \reg_out[23][7] , \reg_out[23][8] ,
         \reg_out[23][9] , \reg_out[23][10] , \reg_out[23][11] ,
         \reg_out[23][12] , \reg_out[23][13] , \reg_out[23][14] ,
         \reg_out[23][15] , \reg_out[23][16] , \reg_out[23][17] ,
         \reg_out[23][18] , \reg_out[23][19] , \reg_out[23][20] ,
         \reg_out[23][21] , \reg_out[23][22] , \reg_out[23][23] ,
         \reg_out[23][24] , \reg_out[23][25] , \reg_out[23][26] ,
         \reg_out[23][27] , \reg_out[23][28] , \reg_out[23][29] ,
         \reg_out[23][30] , \reg_out[23][31] , \reg_out[25][0] ,
         \reg_out[25][1] , \reg_out[25][2] , \reg_out[25][3] ,
         \reg_out[25][4] , \reg_out[25][5] , \reg_out[25][6] ,
         \reg_out[25][7] , \reg_out[25][8] , \reg_out[25][9] ,
         \reg_out[25][10] , \reg_out[25][11] , \reg_out[25][12] ,
         \reg_out[25][13] , \reg_out[25][14] , \reg_out[25][15] ,
         \reg_out[25][16] , \reg_out[25][17] , \reg_out[25][18] ,
         \reg_out[25][19] , \reg_out[25][20] , \reg_out[25][21] ,
         \reg_out[25][22] , \reg_out[25][23] , \reg_out[25][24] ,
         \reg_out[25][25] , \reg_out[25][26] , \reg_out[25][27] ,
         \reg_out[25][28] , \reg_out[25][29] , \reg_out[25][30] ,
         \reg_out[25][31] , \reg_out[27][0] , \reg_out[27][1] ,
         \reg_out[27][2] , \reg_out[27][3] , \reg_out[27][4] ,
         \reg_out[27][5] , \reg_out[27][6] , \reg_out[27][7] ,
         \reg_out[27][8] , \reg_out[27][9] , \reg_out[27][10] ,
         \reg_out[27][11] , \reg_out[27][12] , \reg_out[27][13] ,
         \reg_out[27][14] , \reg_out[27][15] , \reg_out[27][16] ,
         \reg_out[27][17] , \reg_out[27][18] , \reg_out[27][19] ,
         \reg_out[27][20] , \reg_out[27][21] , \reg_out[27][22] ,
         \reg_out[27][23] , \reg_out[27][24] , \reg_out[27][25] ,
         \reg_out[27][26] , \reg_out[27][27] , \reg_out[27][28] ,
         \reg_out[27][29] , \reg_out[27][30] , \reg_out[27][31] ,
         \reg_out[29][0] , \reg_out[29][1] , \reg_out[29][2] ,
         \reg_out[29][3] , \reg_out[29][4] , \reg_out[29][5] ,
         \reg_out[29][6] , \reg_out[29][7] , \reg_out[29][8] ,
         \reg_out[29][9] , \reg_out[29][10] , \reg_out[29][11] ,
         \reg_out[29][12] , \reg_out[29][13] , \reg_out[29][14] ,
         \reg_out[29][15] , \reg_out[29][16] , \reg_out[29][17] ,
         \reg_out[29][18] , \reg_out[29][19] , \reg_out[29][20] ,
         \reg_out[29][21] , \reg_out[29][22] , \reg_out[29][23] ,
         \reg_out[29][24] , \reg_out[29][25] , \reg_out[29][26] ,
         \reg_out[29][27] , \reg_out[29][28] , \reg_out[29][29] ,
         \reg_out[29][30] , \reg_out[29][31] , \reg_out[31][0] ,
         \reg_out[31][1] , \reg_out[31][2] , \reg_out[31][3] ,
         \reg_out[31][4] , \reg_out[31][5] , \reg_out[31][6] ,
         \reg_out[31][7] , \reg_out[31][8] , \reg_out[31][9] ,
         \reg_out[31][10] , \reg_out[31][11] , \reg_out[31][12] ,
         \reg_out[31][13] , \reg_out[31][14] , \reg_out[31][15] ,
         \reg_out[31][16] , \reg_out[31][17] , \reg_out[31][18] ,
         \reg_out[31][19] , \reg_out[31][20] , \reg_out[31][21] ,
         \reg_out[31][22] , \reg_out[31][23] , \reg_out[31][24] ,
         \reg_out[31][25] , \reg_out[31][26] , \reg_out[31][27] ,
         \reg_out[31][28] , \reg_out[31][29] , \reg_out[31][30] ,
         \reg_out[31][31] ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n2061, n2062, n2063, n2064, n2065, n2066, n2070, n2075,
         n2078, n2079, n2081, n2082, n2083, n2084, n2086, n2087, n2088, n2089,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2726, n2731, n2734, n2735, n2737, n2738, n2739, n2740,
         n2742, n2743, n2744, n2745, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3407, n3408, n3411,
         n3414, n3415, n3418, n3423, n3426, n3429, n3434, n3436, n3438, n3440,
         n3441, n3443, n3445, n3447, n3448, n3450, n3451, n3453, n3455, n3457,
         n3459, n3461, n3470, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912;

  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n4443) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3911) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3602) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3993) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3999) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n4005) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n4011) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n4017) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3769) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3777) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4449) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4455) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4461) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4467) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3881) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3886) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3891) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4474) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4480) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3903) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3919) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3927) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3935) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3943) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3951) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3959) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3967) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3975) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3983) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4486) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3610) );
  DFF_X1 \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3987) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[1][0] ), .QN(n4509) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[1][1] ), .QN(n4085) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[1][2] ), .QN(n4095) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[1][3] ), .QN(n4098) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[1][4] ), .QN(n4099) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[1][5] ), .QN(n4100) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[1][6] ), .QN(n4101) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[1][7] ), .QN(n4102) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[1][8] ), .QN(n4103) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[1][9] ), .QN(n4104) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][10] ), .QN(n4510) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][11] ), .QN(n4511) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][12] ), .QN(n4512) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][13] ), .QN(n4513) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][14] ), .QN(n4514) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][15] ), .QN(n4515) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][16] ), .QN(n4516) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][17] ), .QN(n4517) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][18] ), .QN(n4518) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][19] ), .QN(n4084) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][20] ), .QN(n4086) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][21] ), .QN(n4087) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][22] ), .QN(n4088) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][23] ), .QN(n4089) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][24] ), .QN(n4090) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][25] ), .QN(n4091) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][26] ), .QN(n4092) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][27] ), .QN(n4093) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][28] ), .QN(n4094) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][29] ), .QN(n4519) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][30] ), .QN(n4096) );
  DFF_X1 \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[1][31] ), .QN(n4097) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3829) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3659) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3525) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3718) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3724) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3730) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3736) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3742) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3586) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3594) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3833) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3837) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3841) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3845) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3634) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3636) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3638) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3853) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3857) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3651) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3667) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3497) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3505) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3513) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3677) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3685) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3693) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3701) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3709) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3863) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3533) );
  DFF_X1 \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3712) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[3][0] ), .QN(n4348) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[3][1] ), .QN(n4359) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[3][2] ), .QN(n4370) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[3][3] ), .QN(n3813) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[3][4] ), .QN(n3814) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[3][5] ), .QN(n3815) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[3][6] ), .QN(n3816) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[3][7] ), .QN(n3817) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[3][8] ), .QN(n3818) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[3][9] ), .QN(n4372) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][10] ), .QN(n4349) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][11] ), .QN(n4350) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][12] ), .QN(n4351) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][13] ), .QN(n4352) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][14] ), .QN(n4353) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][15] ), .QN(n4354) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][16] ), .QN(n4355) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][17] ), .QN(n4356) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][18] ), .QN(n4357) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][19] ), .QN(n4358) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][20] ), .QN(n4360) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][21] ), .QN(n4361) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][22] ), .QN(n4362) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][23] ), .QN(n4363) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][24] ), .QN(n4364) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][25] ), .QN(n4365) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][26] ), .QN(n4366) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][27] ), .QN(n4367) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][28] ), .QN(n4368) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][29] ), .QN(n4369) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][30] ), .QN(n4371) );
  DFF_X1 \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[3][31] ), .QN(n3812) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3870) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3912) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3603) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3756) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3758) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3760) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3762) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3764) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3770) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3778) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3872) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3874) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3876) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3878) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3882) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3887) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3892) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3894) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3896) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3904) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3920) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3928) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3936) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3944) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3952) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3960) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3968) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3976) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3984) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3986) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3611) );
  DFF_X1 \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3754) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[5][0] ), .QN(n4168) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[5][1] ), .QN(n4179) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[5][2] ), .QN(n4190) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[5][3] ), .QN(n3792) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[5][4] ), .QN(n3793) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[5][5] ), .QN(n3794) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[5][6] ), .QN(n3795) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[5][7] ), .QN(n3796) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[5][8] ), .QN(n3797) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[5][9] ), .QN(n4192) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][10] ), .QN(n4169) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][11] ), .QN(n4170) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][12] ), .QN(n4171) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][13] ), .QN(n4172) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][14] ), .QN(n4173) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][15] ), .QN(n4174) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][16] ), .QN(n4175) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][17] ), .QN(n4176) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][18] ), .QN(n4177) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][19] ), .QN(n4178) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][20] ), .QN(n4180) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][21] ), .QN(n4181) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][22] ), .QN(n4182) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][23] ), .QN(n4183) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][24] ), .QN(n4184) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][25] ), .QN(n4185) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][26] ), .QN(n4186) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][27] ), .QN(n4187) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][28] ), .QN(n4188) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][29] ), .QN(n4189) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][30] ), .QN(n4191) );
  DFF_X1 \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[5][31] ), .QN(n3791) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3620) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3660) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3526) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3577) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3578) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3579) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3580) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3581) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3587) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3595) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3623) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3626) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3629) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3632) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3635) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3637) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3639) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3641) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3644) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3652) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3668) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3498) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3506) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3514) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3678) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3686) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3694) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3702) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3710) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3711) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3534) );
  DFF_X1 \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3576) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[7][0] ), .QN(n4373) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[7][1] ), .QN(n4384) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[7][2] ), .QN(n4395) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[7][3] ), .QN(n3820) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[7][4] ), .QN(n3821) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[7][5] ), .QN(n3822) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[7][6] ), .QN(n3823) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[7][7] ), .QN(n3824) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[7][8] ), .QN(n3825) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[7][9] ), .QN(n4397) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][10] ), .QN(n4374) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][11] ), .QN(n4375) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][12] ), .QN(n4376) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][13] ), .QN(n4377) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][14] ), .QN(n4378) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][15] ), .QN(n4379) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][16] ), .QN(n4380) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][17] ), .QN(n4381) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][18] ), .QN(n4382) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][19] ), .QN(n4383) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][20] ), .QN(n4385) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][21] ), .QN(n4386) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][22] ), .QN(n4387) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][23] ), .QN(n4388) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][24] ), .QN(n4389) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][25] ), .QN(n4390) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][26] ), .QN(n4391) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][27] ), .QN(n4392) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][28] ), .QN(n4393) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][29] ), .QN(n4394) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][30] ), .QN(n4396) );
  DFF_X1 \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[7][31] ), .QN(n3819) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3869) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3907) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3598) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3755) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3757) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3759) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3761) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3763) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3765) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .QN(n3773) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3871) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3873) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3875) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3877) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3879) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3883) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3888) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3893) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3895) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3899) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3915) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3923) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3931) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3939) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3947) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3955) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3963) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3971) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3979) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3985) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3606) );
  DFF_X1 \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3614) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[9][0] ), .QN(n4193) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[9][1] ), .QN(n4204) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[9][2] ), .QN(n4215) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[9][3] ), .QN(n3799) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[9][4] ), .QN(n3800) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[9][5] ), .QN(n3801) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[9][6] ), .QN(n3802) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[9][7] ), .QN(n3803) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[9][8] ), .QN(n3804) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), 
        .CK(clk), .Q(\reg_out[9][9] ), .QN(n4217) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][10] ), .QN(n4194) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][11] ), .QN(n4195) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][12] ), .QN(n4196) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][13] ), .QN(n4197) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][14] ), .QN(n4198) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][15] ), .QN(n4199) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][16] ), .QN(n4200) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][17] ), .QN(n4201) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][18] ), .QN(n4202) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][19] ), .QN(n4203) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][20] ), .QN(n4205) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][21] ), .QN(n4206) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][22] ), .QN(n4207) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][23] ), .QN(n4208) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][24] ), .QN(n4209) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][25] ), .QN(n4210) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][26] ), .QN(n4211) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][27] ), .QN(n4212) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][28] ), .QN(n4213) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][29] ), .QN(n4214) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][30] ), .QN(n4216) );
  DFF_X1 \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[9][31] ), .QN(n3798) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4429) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3655) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3521) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3864) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3865) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3866) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3867) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3868) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3582) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3590) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4430) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4431) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4432) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4433) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4434) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3566) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3571) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4435) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4436) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3647) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3663) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3671) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3501) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3509) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3517) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3681) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3689) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3697) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3705) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4437) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3529) );
  DFF_X1 \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3537) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][0] ), .QN(n4553) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][1] ), .QN(n4219) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][2] ), .QN(n4229) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][3] ), .QN(n4232) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][4] ), .QN(n4233) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][5] ), .QN(n4234) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][6] ), .QN(n4235) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][7] ), .QN(n4236) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][8] ), .QN(n4237) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][9] ), .QN(n4238) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][10] ), .QN(n4554) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][11] ), .QN(n4555) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][12] ), .QN(n4556) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][13] ), .QN(n4557) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][14] ), .QN(n4558) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][15] ), .QN(n4559) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][16] ), .QN(n4560) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][17] ), .QN(n4561) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][18] ), .QN(n4562) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][19] ), .QN(n4218) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][20] ), .QN(n4220) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][21] ), .QN(n4221) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][22] ), .QN(n4222) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][23] ), .QN(n4223) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][24] ), .QN(n4224) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][25] ), .QN(n4225) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][26] ), .QN(n4226) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][27] ), .QN(n4227) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][28] ), .QN(n4228) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][29] ), .QN(n4563) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][30] ), .QN(n4230) );
  DFF_X1 \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[11][31] ), .QN(n4231) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4440) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3908) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3599) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3990) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3996) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4002) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4008) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4014) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3766) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3774) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4446) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4452) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4458) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4464) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4470) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3884) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3889) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4471) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4477) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3900) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3916) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3924) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3932) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3940) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3948) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3956) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3964) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3972) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3980) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4483) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3607) );
  DFF_X1 \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3615) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][0] ), .QN(n4487) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][1] ), .QN(n4043) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][2] ), .QN(n4053) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][3] ), .QN(n4056) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][4] ), .QN(n4057) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][5] ), .QN(n4058) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][6] ), .QN(n4059) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][7] ), .QN(n4060) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][8] ), .QN(n4061) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][9] ), .QN(n4062) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][10] ), .QN(n4488) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][11] ), .QN(n4489) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][12] ), .QN(n4490) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][13] ), .QN(n4491) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][14] ), .QN(n4492) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][15] ), .QN(n4493) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][16] ), .QN(n4494) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][17] ), .QN(n4495) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][18] ), .QN(n4496) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][19] ), .QN(n4042) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][20] ), .QN(n4044) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][21] ), .QN(n4045) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][22] ), .QN(n4046) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][23] ), .QN(n4047) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][24] ), .QN(n4048) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][25] ), .QN(n4049) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][26] ), .QN(n4050) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][27] ), .QN(n4051) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][28] ), .QN(n4052) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][29] ), .QN(n4497) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][30] ), .QN(n4054) );
  DFF_X1 \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[13][31] ), .QN(n4055) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3827) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3656) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3522) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3715) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3721) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3727) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3733) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3739) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3583) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3591) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3831) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3835) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3839) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3843) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3847) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3567) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3572) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3851) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3855) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3648) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3664) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3672) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3502) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3510) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3518) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3682) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3690) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3698) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3706) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3860) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3530) );
  DFF_X1 \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3538) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][0] ), .QN(n4564) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][1] ), .QN(n4240) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][2] ), .QN(n4250) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][3] ), .QN(n4253) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][4] ), .QN(n4254) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][5] ), .QN(n4255) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][6] ), .QN(n4256) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][7] ), .QN(n4257) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][8] ), .QN(n4258) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][9] ), .QN(n4259) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][10] ), .QN(n4565) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][11] ), .QN(n4566) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][12] ), .QN(n4567) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][13] ), .QN(n4568) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][14] ), .QN(n4569) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][15] ), .QN(n4570) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][16] ), .QN(n4571) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][17] ), .QN(n4572) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][18] ), .QN(n4573) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][19] ), .QN(n4239) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][20] ), .QN(n4241) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][21] ), .QN(n4242) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][22] ), .QN(n4243) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][23] ), .QN(n4244) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][24] ), .QN(n4245) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][25] ), .QN(n4246) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][26] ), .QN(n4247) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][27] ), .QN(n4248) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][28] ), .QN(n4249) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][29] ), .QN(n4574) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][30] ), .QN(n4251) );
  DFF_X1 \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[15][31] ), .QN(n4252) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4441) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3909) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3600) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3991) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3997) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4003) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4009) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4015) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3767) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3775) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4447) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4453) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4459) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4465) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3880) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3885) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3890) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4472) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4478) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3901) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3917) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3925) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3933) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3941) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3949) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3957) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3965) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3973) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3981) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4484) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3608) );
  DFF_X1 \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3616) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][0] ), .QN(n4498) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][1] ), .QN(n4064) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][2] ), .QN(n4074) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][3] ), .QN(n4077) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][4] ), .QN(n4078) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][5] ), .QN(n4079) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][6] ), .QN(n4080) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][7] ), .QN(n4081) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][8] ), .QN(n4082) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][9] ), .QN(n4083) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][10] ), .QN(n4499) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][11] ), .QN(n4500) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][12] ), .QN(n4501) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][13] ), .QN(n4502) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][14] ), .QN(n4503) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][15] ), .QN(n4504) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][16] ), .QN(n4505) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][17] ), .QN(n4506) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][18] ), .QN(n4507) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][19] ), .QN(n4063) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][20] ), .QN(n4065) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][21] ), .QN(n4066) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][22] ), .QN(n4067) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][23] ), .QN(n4068) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][24] ), .QN(n4069) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][25] ), .QN(n4070) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][26] ), .QN(n4071) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][27] ), .QN(n4072) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][28] ), .QN(n4073) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][29] ), .QN(n4508) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][30] ), .QN(n4075) );
  DFF_X1 \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[17][31] ), .QN(n4076) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3828) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3657) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3523) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3716) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3722) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3728) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3734) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3740) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3584) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3592) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3832) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3836) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3840) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3844) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3563) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3568) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3573) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3852) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3856) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3649) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3665) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3673) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3503) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3511) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3675) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3683) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3691) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3699) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3707) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3861) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3531) );
  DFF_X1 \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3539) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][0] ), .QN(n4575) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][1] ), .QN(n4261) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][2] ), .QN(n4271) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][3] ), .QN(n4274) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][4] ), .QN(n4275) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][5] ), .QN(n4276) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][6] ), .QN(n4277) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][7] ), .QN(n4278) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][8] ), .QN(n4279) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][9] ), .QN(n4280) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][10] ), .QN(n4576) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][11] ), .QN(n4577) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][12] ), .QN(n4578) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][13] ), .QN(n4579) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][14] ), .QN(n4580) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][15] ), .QN(n4581) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][16] ), .QN(n4582) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][17] ), .QN(n4583) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][18] ), .QN(n4584) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][19] ), .QN(n4260) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][20] ), .QN(n4262) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][21] ), .QN(n4263) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][22] ), .QN(n4264) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][23] ), .QN(n4265) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][24] ), .QN(n4266) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][25] ), .QN(n4267) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][26] ), .QN(n4268) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][27] ), .QN(n4269) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][28] ), .QN(n4270) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][29] ), .QN(n4585) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][30] ), .QN(n4272) );
  DFF_X1 \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[19][31] ), .QN(n4273) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4442) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3910) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3601) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3992) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3998) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4004) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4010) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4016) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3768) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3776) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4448) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4454) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4460) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4466) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3745) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3748) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3751) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4473) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4479) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3902) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3918) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3926) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3934) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3942) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3950) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3958) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3966) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3974) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3982) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4485) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3609) );
  DFF_X1 \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3617) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][0] ), .QN(n4520) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][1] ), .QN(n4106) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][2] ), .QN(n4116) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][3] ), .QN(n4119) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][4] ), .QN(n4120) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][5] ), .QN(n4121) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][6] ), .QN(n4122) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][7] ), .QN(n4123) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][8] ), .QN(n4124) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][9] ), .QN(n4125) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][10] ), .QN(n4521) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][11] ), .QN(n4522) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][12] ), .QN(n4523) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][13] ), .QN(n4524) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][14] ), .QN(n4525) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][15] ), .QN(n4526) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][16] ), .QN(n4527) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][17] ), .QN(n4528) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][18] ), .QN(n4529) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][19] ), .QN(n4105) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][20] ), .QN(n4107) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][21] ), .QN(n4108) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][22] ), .QN(n4109) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][23] ), .QN(n4110) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][24] ), .QN(n4111) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][25] ), .QN(n4112) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][26] ), .QN(n4113) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][27] ), .QN(n4114) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][28] ), .QN(n4115) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][29] ), .QN(n4530) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][30] ), .QN(n4117) );
  DFF_X1 \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[21][31] ), .QN(n4118) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3619) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3658) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3524) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3717) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3723) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3729) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3735) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3741) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3585) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3593) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3622) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3625) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3628) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3631) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3564) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3569) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3574) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3640) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3643) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3650) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3666) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3674) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3504) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3512) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3676) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3684) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3692) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3700) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3708) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3862) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3532) );
  DFF_X1 \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3540) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][0] ), .QN(n4586) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][1] ), .QN(n4282) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][2] ), .QN(n4292) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][3] ), .QN(n4295) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][4] ), .QN(n4296) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][5] ), .QN(n4297) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][6] ), .QN(n4298) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][7] ), .QN(n4299) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][8] ), .QN(n4300) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][9] ), .QN(n4301) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][10] ), .QN(n4587) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][11] ), .QN(n4588) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][12] ), .QN(n4589) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][13] ), .QN(n4590) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][14] ), .QN(n4591) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][15] ), .QN(n4592) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][16] ), .QN(n4593) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][17] ), .QN(n4594) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][18] ), .QN(n4595) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][19] ), .QN(n4281) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][20] ), .QN(n4283) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][21] ), .QN(n4284) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][22] ), .QN(n4285) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][23] ), .QN(n4286) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][24] ), .QN(n4287) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][25] ), .QN(n4288) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][26] ), .QN(n4289) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][27] ), .QN(n4290) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][28] ), .QN(n4291) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][29] ), .QN(n4596) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][30] ), .QN(n4293) );
  DFF_X1 \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[23][31] ), .QN(n4294) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4438) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3905) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3596) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3988) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3994) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4000) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4006) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4012) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4018) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3771) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4444) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4450) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4456) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4462) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4468) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3746) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3749) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3752) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4475) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3897) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3913) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3921) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3929) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3937) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3945) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3953) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3961) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3969) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3977) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4481) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3604) );
  DFF_X1 \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3612) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][0] ), .QN(n4531) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][1] ), .QN(n4127) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][2] ), .QN(n4137) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][3] ), .QN(n4140) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][4] ), .QN(n4141) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][5] ), .QN(n4142) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][6] ), .QN(n4143) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][7] ), .QN(n4144) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][8] ), .QN(n4145) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][9] ), .QN(n4146) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][10] ), .QN(n4532) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][11] ), .QN(n4533) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][12] ), .QN(n4534) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][13] ), .QN(n4535) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][14] ), .QN(n4536) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][15] ), .QN(n4537) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][16] ), .QN(n4538) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][17] ), .QN(n4539) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][18] ), .QN(n4540) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][19] ), .QN(n4126) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][20] ), .QN(n4128) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][21] ), .QN(n4129) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][22] ), .QN(n4130) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][23] ), .QN(n4131) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][24] ), .QN(n4132) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][25] ), .QN(n4133) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][26] ), .QN(n4134) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][27] ), .QN(n4135) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][28] ), .QN(n4136) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][29] ), .QN(n4541) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][30] ), .QN(n4138) );
  DFF_X1 \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[25][31] ), .QN(n4139) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3618) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3653) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3519) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3713) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3719) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3725) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3731) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3737) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3743) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3588) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3621) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3624) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3627) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3630) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3633) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3565) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3570) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3575) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3642) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3645) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3661) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3669) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3499) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3507) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3515) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3679) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3687) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3695) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3703) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3858) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3527) );
  DFF_X1 \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3535) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][0] ), .QN(n4597) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][1] ), .QN(n4303) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][2] ), .QN(n4313) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][3] ), .QN(n4316) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][4] ), .QN(n4317) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][5] ), .QN(n4318) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][6] ), .QN(n4319) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][7] ), .QN(n4320) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][8] ), .QN(n4321) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][9] ), .QN(n4322) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][10] ), .QN(n4598) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][11] ), .QN(n4599) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][12] ), .QN(n4600) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][13] ), .QN(n4601) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][14] ), .QN(n4602) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][15] ), .QN(n4603) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][16] ), .QN(n4604) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][17] ), .QN(n4605) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][18] ), .QN(n4606) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][19] ), .QN(n4302) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][20] ), .QN(n4304) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][21] ), .QN(n4305) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][22] ), .QN(n4306) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][23] ), .QN(n4307) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][24] ), .QN(n4308) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][25] ), .QN(n4309) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][26] ), .QN(n4310) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][27] ), .QN(n4311) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][28] ), .QN(n4312) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][29] ), .QN(n4607) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][30] ), .QN(n4314) );
  DFF_X1 \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[27][31] ), .QN(n4315) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4439) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3906) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3597) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3989) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3995) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4001) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4007) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4013) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4019) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3772) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4445) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4451) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4457) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4463) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4469) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3747) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3750) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3753) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4476) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3898) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3914) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3922) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3930) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3938) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3946) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3954) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3962) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3970) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3978) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n4482) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3605) );
  DFF_X1 \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3613) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][0] ), .QN(n4542) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][1] ), .QN(n4148) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][2] ), .QN(n4158) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][3] ), .QN(n4161) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][4] ), .QN(n4162) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][5] ), .QN(n4163) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][6] ), .QN(n4164) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][7] ), .QN(n4165) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][8] ), .QN(n4166) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][9] ), .QN(n4167) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][10] ), .QN(n4543) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][11] ), .QN(n4544) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][12] ), .QN(n4545) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][13] ), .QN(n4546) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][14] ), .QN(n4547) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][15] ), .QN(n4548) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][16] ), .QN(n4549) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][17] ), .QN(n4550) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][18] ), .QN(n4551) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][19] ), .QN(n4147) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][20] ), .QN(n4149) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][21] ), .QN(n4150) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][22] ), .QN(n4151) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][23] ), .QN(n4152) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][24] ), .QN(n4153) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][25] ), .QN(n4154) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][26] ), .QN(n4155) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][27] ), .QN(n4156) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][28] ), .QN(n4157) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][29] ), .QN(n4552) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][30] ), .QN(n4159) );
  DFF_X1 \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[29][31] ), .QN(n4160) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3826) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3654) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3520) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3714) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3720) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3726) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3732) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3738) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3744) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3589) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3830) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3834) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3838) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3842) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3846) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3848) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3849) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3850) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3854) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3646) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3662) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3670) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3500) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3508) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3516) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3680) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3688) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3696) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3704) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3859) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3528) );
  DFF_X1 \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n3536) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][0] ), .QN(n4323) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][1] ), .QN(n4334) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][2] ), .QN(n4345) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][3] ), .QN(n3806) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][4] ), .QN(n3807) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][5] ), .QN(n3808) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][6] ), .QN(n3809) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][7] ), .QN(n3810) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][8] ), .QN(n3811) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][9] ), .QN(n4347) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][10] ), .QN(n4324) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][11] ), .QN(n4325) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][12] ), .QN(n4326) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][13] ), .QN(n4327) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][14] ), .QN(n4328) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][15] ), .QN(n4329) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][16] ), .QN(n4330) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][17] ), .QN(n4331) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][18] ), .QN(n4332) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][19] ), .QN(n4333) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][20] ), .QN(n4335) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][21] ), .QN(n4336) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][22] ), .QN(n4337) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][23] ), .QN(n4338) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][24] ), .QN(n4339) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][25] ), .QN(n4340) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][26] ), .QN(n4341) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][27] ), .QN(n4342) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][28] ), .QN(n4343) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][29] ), .QN(n4344) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][30] ), .QN(n4346) );
  DFF_X1 \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\reg_out[31][31] ), .QN(n3805) );
  NAND4_X2 U1 ( .A1(n2061), .A2(n2062), .A3(n2063), .A4(n2064), .ZN(busB[9])
         );
  OAI221_X2 U3 ( .B1(n4905), .B2(n3778), .C1(n4892), .C2(n3595), .A(n2070), 
        .ZN(n2066) );
  AOI22_X2 U4 ( .A1(\reg_out[5][9] ), .A2(n4887), .B1(\reg_out[7][9] ), .B2(
        n4885), .ZN(n2070) );
  OAI221_X2 U5 ( .B1(n4878), .B2(n3777), .C1(n4866), .C2(n3594), .A(n2075), 
        .ZN(n2065) );
  AOI22_X2 U6 ( .A1(\reg_out[1][9] ), .A2(n4859), .B1(\reg_out[3][9] ), .B2(
        n4857), .ZN(n2075) );
  OAI221_X2 U8 ( .B1(n4905), .B2(n3776), .C1(n4892), .C2(n3593), .A(n2081), 
        .ZN(n2079) );
  AOI22_X2 U9 ( .A1(\reg_out[21][9] ), .A2(n4887), .B1(\reg_out[23][9] ), .B2(
        n4885), .ZN(n2081) );
  OAI221_X2 U10 ( .B1(n4878), .B2(n3775), .C1(n4866), .C2(n3592), .A(n2082), 
        .ZN(n2078) );
  AOI22_X2 U11 ( .A1(\reg_out[17][9] ), .A2(n4859), .B1(\reg_out[19][9] ), 
        .B2(n4857), .ZN(n2082) );
  OAI221_X2 U13 ( .B1(n4905), .B2(n3774), .C1(n4892), .C2(n3591), .A(n2086), 
        .ZN(n2084) );
  AOI22_X2 U14 ( .A1(\reg_out[13][9] ), .A2(n4887), .B1(\reg_out[15][9] ), 
        .B2(n4885), .ZN(n2086) );
  OAI221_X2 U15 ( .B1(n4878), .B2(n3773), .C1(n4866), .C2(n3590), .A(n2087), 
        .ZN(n2083) );
  AOI22_X2 U16 ( .A1(\reg_out[9][9] ), .A2(n4859), .B1(\reg_out[11][9] ), .B2(
        n4857), .ZN(n2087) );
  OAI221_X2 U18 ( .B1(n4905), .B2(n3772), .C1(n4898), .C2(n3589), .A(n2091), 
        .ZN(n2089) );
  AOI22_X2 U19 ( .A1(\reg_out[29][9] ), .A2(n4887), .B1(\reg_out[31][9] ), 
        .B2(n4885), .ZN(n2091) );
  OAI221_X2 U20 ( .B1(n4878), .B2(n3771), .C1(n4871), .C2(n3588), .A(n2092), 
        .ZN(n2088) );
  AOI22_X2 U21 ( .A1(\reg_out[25][9] ), .A2(n4859), .B1(\reg_out[27][9] ), 
        .B2(n4857), .ZN(n2092) );
  NAND4_X2 U22 ( .A1(n2093), .A2(n2094), .A3(n2095), .A4(n2096), .ZN(busB[8])
         );
  OAI221_X2 U24 ( .B1(n4906), .B2(n3770), .C1(n4892), .C2(n3587), .A(n2099), 
        .ZN(n2098) );
  AOI22_X2 U25 ( .A1(\reg_out[5][8] ), .A2(n4887), .B1(\reg_out[7][8] ), .B2(
        n4886), .ZN(n2099) );
  OAI221_X2 U26 ( .B1(n4879), .B2(n3769), .C1(n4866), .C2(n3586), .A(n2100), 
        .ZN(n2097) );
  AOI22_X2 U27 ( .A1(\reg_out[1][8] ), .A2(n4859), .B1(\reg_out[3][8] ), .B2(
        n4858), .ZN(n2100) );
  OAI221_X2 U29 ( .B1(n4906), .B2(n3768), .C1(n4892), .C2(n3585), .A(n2103), 
        .ZN(n2102) );
  AOI22_X2 U30 ( .A1(\reg_out[21][8] ), .A2(n4887), .B1(\reg_out[23][8] ), 
        .B2(n4886), .ZN(n2103) );
  OAI221_X2 U31 ( .B1(n4879), .B2(n3767), .C1(n4866), .C2(n3584), .A(n2104), 
        .ZN(n2101) );
  AOI22_X2 U32 ( .A1(\reg_out[17][8] ), .A2(n4859), .B1(\reg_out[19][8] ), 
        .B2(n4858), .ZN(n2104) );
  OAI221_X2 U34 ( .B1(n4906), .B2(n3766), .C1(n4892), .C2(n3583), .A(n2107), 
        .ZN(n2106) );
  AOI22_X2 U35 ( .A1(\reg_out[13][8] ), .A2(n4887), .B1(\reg_out[15][8] ), 
        .B2(n4886), .ZN(n2107) );
  OAI221_X2 U36 ( .B1(n4879), .B2(n3765), .C1(n4866), .C2(n3582), .A(n2108), 
        .ZN(n2105) );
  AOI22_X2 U37 ( .A1(\reg_out[9][8] ), .A2(n4859), .B1(\reg_out[11][8] ), .B2(
        n4858), .ZN(n2108) );
  OAI221_X2 U39 ( .B1(n4906), .B2(n4019), .C1(n4899), .C2(n3744), .A(n2111), 
        .ZN(n2110) );
  AOI22_X2 U40 ( .A1(\reg_out[29][8] ), .A2(n4888), .B1(\reg_out[31][8] ), 
        .B2(n4886), .ZN(n2111) );
  OAI221_X2 U41 ( .B1(n4879), .B2(n4018), .C1(n4872), .C2(n3743), .A(n2112), 
        .ZN(n2109) );
  AOI22_X2 U42 ( .A1(\reg_out[25][8] ), .A2(n4863), .B1(\reg_out[27][8] ), 
        .B2(n4858), .ZN(n2112) );
  NAND4_X2 U43 ( .A1(n2113), .A2(n2114), .A3(n2115), .A4(n2116), .ZN(busB[7])
         );
  OAI221_X2 U45 ( .B1(n4906), .B2(n3764), .C1(n4899), .C2(n3581), .A(n2119), 
        .ZN(n2118) );
  AOI22_X2 U46 ( .A1(\reg_out[5][7] ), .A2(n4888), .B1(\reg_out[7][7] ), .B2(
        n4886), .ZN(n2119) );
  OAI221_X2 U47 ( .B1(n4879), .B2(n4017), .C1(n4872), .C2(n3742), .A(n2120), 
        .ZN(n2117) );
  AOI22_X2 U48 ( .A1(\reg_out[1][7] ), .A2(n4863), .B1(\reg_out[3][7] ), .B2(
        n4858), .ZN(n2120) );
  OAI221_X2 U50 ( .B1(n4906), .B2(n4016), .C1(n4899), .C2(n3741), .A(n2123), 
        .ZN(n2122) );
  AOI22_X2 U51 ( .A1(\reg_out[21][7] ), .A2(n4890), .B1(\reg_out[23][7] ), 
        .B2(n4886), .ZN(n2123) );
  OAI221_X2 U52 ( .B1(n4879), .B2(n4015), .C1(n4872), .C2(n3740), .A(n2124), 
        .ZN(n2121) );
  AOI22_X2 U53 ( .A1(\reg_out[17][7] ), .A2(n4864), .B1(\reg_out[19][7] ), 
        .B2(n4858), .ZN(n2124) );
  OAI221_X2 U55 ( .B1(n4906), .B2(n4014), .C1(n4899), .C2(n3739), .A(n2127), 
        .ZN(n2126) );
  AOI22_X2 U56 ( .A1(\reg_out[13][7] ), .A2(n4890), .B1(\reg_out[15][7] ), 
        .B2(n4886), .ZN(n2127) );
  OAI221_X2 U57 ( .B1(n4879), .B2(n3763), .C1(n4872), .C2(n3868), .A(n2128), 
        .ZN(n2125) );
  AOI22_X2 U58 ( .A1(\reg_out[9][7] ), .A2(n4864), .B1(\reg_out[11][7] ), .B2(
        n4858), .ZN(n2128) );
  OAI221_X2 U60 ( .B1(n4906), .B2(n4013), .C1(n4899), .C2(n3738), .A(n2131), 
        .ZN(n2130) );
  AOI22_X2 U61 ( .A1(\reg_out[29][7] ), .A2(n4890), .B1(\reg_out[31][7] ), 
        .B2(n4886), .ZN(n2131) );
  OAI221_X2 U62 ( .B1(n4879), .B2(n4012), .C1(n4872), .C2(n3737), .A(n2132), 
        .ZN(n2129) );
  AOI22_X2 U63 ( .A1(\reg_out[25][7] ), .A2(n4864), .B1(\reg_out[27][7] ), 
        .B2(n4858), .ZN(n2132) );
  NAND4_X2 U64 ( .A1(n2133), .A2(n2134), .A3(n2135), .A4(n2136), .ZN(busB[6])
         );
  OAI221_X2 U66 ( .B1(n4906), .B2(n3762), .C1(n4899), .C2(n3580), .A(n2139), 
        .ZN(n2138) );
  AOI22_X2 U67 ( .A1(\reg_out[5][6] ), .A2(n4891), .B1(\reg_out[7][6] ), .B2(
        n4886), .ZN(n2139) );
  OAI221_X2 U68 ( .B1(n4879), .B2(n4011), .C1(n4872), .C2(n3736), .A(n2140), 
        .ZN(n2137) );
  AOI22_X2 U69 ( .A1(\reg_out[1][6] ), .A2(n4861), .B1(\reg_out[3][6] ), .B2(
        n4858), .ZN(n2140) );
  OAI221_X2 U71 ( .B1(n4906), .B2(n4010), .C1(n4899), .C2(n3735), .A(n2143), 
        .ZN(n2142) );
  AOI22_X2 U72 ( .A1(\reg_out[21][6] ), .A2(n4891), .B1(\reg_out[23][6] ), 
        .B2(n4886), .ZN(n2143) );
  OAI221_X2 U73 ( .B1(n4879), .B2(n4009), .C1(n4872), .C2(n3734), .A(n2144), 
        .ZN(n2141) );
  AOI22_X2 U74 ( .A1(\reg_out[17][6] ), .A2(n4861), .B1(\reg_out[19][6] ), 
        .B2(n4858), .ZN(n2144) );
  OAI221_X2 U76 ( .B1(n4906), .B2(n4008), .C1(n4899), .C2(n3733), .A(n2147), 
        .ZN(n2146) );
  AOI22_X2 U77 ( .A1(\reg_out[13][6] ), .A2(n4891), .B1(\reg_out[15][6] ), 
        .B2(n4886), .ZN(n2147) );
  OAI221_X2 U78 ( .B1(n4879), .B2(n3761), .C1(n4872), .C2(n3867), .A(n2148), 
        .ZN(n2145) );
  AOI22_X2 U79 ( .A1(\reg_out[9][6] ), .A2(n4861), .B1(\reg_out[11][6] ), .B2(
        n4858), .ZN(n2148) );
  OAI221_X2 U81 ( .B1(n4906), .B2(n4007), .C1(n4899), .C2(n3732), .A(n2151), 
        .ZN(n2150) );
  AOI22_X2 U82 ( .A1(\reg_out[29][6] ), .A2(n4891), .B1(\reg_out[31][6] ), 
        .B2(n4886), .ZN(n2151) );
  OAI221_X2 U83 ( .B1(n4879), .B2(n4006), .C1(n4872), .C2(n3731), .A(n2152), 
        .ZN(n2149) );
  AOI22_X2 U84 ( .A1(\reg_out[25][6] ), .A2(n4865), .B1(\reg_out[27][6] ), 
        .B2(n4858), .ZN(n2152) );
  NAND4_X2 U85 ( .A1(n2153), .A2(n2154), .A3(n2155), .A4(n2156), .ZN(busB[5])
         );
  OAI221_X2 U87 ( .B1(n4906), .B2(n3760), .C1(n4899), .C2(n3579), .A(n2159), 
        .ZN(n2158) );
  AOI22_X2 U88 ( .A1(\reg_out[5][5] ), .A2(n4888), .B1(\reg_out[7][5] ), .B2(
        n4886), .ZN(n2159) );
  OAI221_X2 U89 ( .B1(n4879), .B2(n4005), .C1(n4872), .C2(n3730), .A(n2160), 
        .ZN(n2157) );
  AOI22_X2 U90 ( .A1(\reg_out[1][5] ), .A2(n4863), .B1(\reg_out[3][5] ), .B2(
        n4858), .ZN(n2160) );
  OAI221_X2 U92 ( .B1(n4906), .B2(n4004), .C1(n4899), .C2(n3729), .A(n2163), 
        .ZN(n2162) );
  AOI22_X2 U93 ( .A1(\reg_out[21][5] ), .A2(n4888), .B1(\reg_out[23][5] ), 
        .B2(n4886), .ZN(n2163) );
  OAI221_X2 U94 ( .B1(n4879), .B2(n4003), .C1(n4872), .C2(n3728), .A(n2164), 
        .ZN(n2161) );
  AOI22_X2 U95 ( .A1(\reg_out[17][5] ), .A2(n4863), .B1(\reg_out[19][5] ), 
        .B2(n4858), .ZN(n2164) );
  OAI221_X2 U97 ( .B1(n4905), .B2(n4002), .C1(n4898), .C2(n3727), .A(n2167), 
        .ZN(n2166) );
  AOI22_X2 U98 ( .A1(\reg_out[13][5] ), .A2(n4889), .B1(\reg_out[15][5] ), 
        .B2(n4885), .ZN(n2167) );
  OAI221_X2 U99 ( .B1(n4878), .B2(n3759), .C1(n4871), .C2(n3866), .A(n2168), 
        .ZN(n2165) );
  AOI22_X2 U100 ( .A1(\reg_out[9][5] ), .A2(n4865), .B1(\reg_out[11][5] ), 
        .B2(n4857), .ZN(n2168) );
  OAI221_X2 U102 ( .B1(n4905), .B2(n4001), .C1(n4898), .C2(n3726), .A(n2171), 
        .ZN(n2170) );
  AOI22_X2 U103 ( .A1(\reg_out[29][5] ), .A2(n4890), .B1(\reg_out[31][5] ), 
        .B2(n4885), .ZN(n2171) );
  OAI221_X2 U104 ( .B1(n4878), .B2(n4000), .C1(n4871), .C2(n3725), .A(n2172), 
        .ZN(n2169) );
  AOI22_X2 U105 ( .A1(\reg_out[25][5] ), .A2(n4865), .B1(\reg_out[27][5] ), 
        .B2(n4857), .ZN(n2172) );
  NAND4_X2 U106 ( .A1(n2173), .A2(n2174), .A3(n2175), .A4(n2176), .ZN(busB[4])
         );
  OAI221_X2 U108 ( .B1(n4905), .B2(n3758), .C1(n4898), .C2(n3578), .A(n2179), 
        .ZN(n2178) );
  AOI22_X2 U109 ( .A1(\reg_out[5][4] ), .A2(n4890), .B1(\reg_out[7][4] ), .B2(
        n4885), .ZN(n2179) );
  OAI221_X2 U110 ( .B1(n4878), .B2(n3999), .C1(n4871), .C2(n3724), .A(n2180), 
        .ZN(n2177) );
  AOI22_X2 U111 ( .A1(\reg_out[1][4] ), .A2(n4865), .B1(\reg_out[3][4] ), .B2(
        n4857), .ZN(n2180) );
  OAI221_X2 U113 ( .B1(n4905), .B2(n3998), .C1(n4898), .C2(n3723), .A(n2183), 
        .ZN(n2182) );
  AOI22_X2 U114 ( .A1(\reg_out[21][4] ), .A2(n4888), .B1(\reg_out[23][4] ), 
        .B2(n4885), .ZN(n2183) );
  OAI221_X2 U115 ( .B1(n4878), .B2(n3997), .C1(n4871), .C2(n3722), .A(n2184), 
        .ZN(n2181) );
  AOI22_X2 U116 ( .A1(\reg_out[17][4] ), .A2(n4865), .B1(\reg_out[19][4] ), 
        .B2(n4857), .ZN(n2184) );
  OAI221_X2 U118 ( .B1(n4905), .B2(n3996), .C1(n4898), .C2(n3721), .A(n2187), 
        .ZN(n2186) );
  AOI22_X2 U119 ( .A1(\reg_out[13][4] ), .A2(n4891), .B1(\reg_out[15][4] ), 
        .B2(n4885), .ZN(n2187) );
  OAI221_X2 U120 ( .B1(n4878), .B2(n3757), .C1(n4871), .C2(n3865), .A(n2188), 
        .ZN(n2185) );
  AOI22_X2 U121 ( .A1(\reg_out[9][4] ), .A2(n4865), .B1(\reg_out[11][4] ), 
        .B2(n4857), .ZN(n2188) );
  OAI221_X2 U123 ( .B1(n4905), .B2(n3995), .C1(n4898), .C2(n3720), .A(n2191), 
        .ZN(n2190) );
  AOI22_X2 U124 ( .A1(\reg_out[29][4] ), .A2(n4889), .B1(\reg_out[31][4] ), 
        .B2(n4885), .ZN(n2191) );
  OAI221_X2 U125 ( .B1(n4878), .B2(n3994), .C1(n4871), .C2(n3719), .A(n2192), 
        .ZN(n2189) );
  AOI22_X2 U126 ( .A1(\reg_out[25][4] ), .A2(n4865), .B1(\reg_out[27][4] ), 
        .B2(n4857), .ZN(n2192) );
  NAND4_X2 U127 ( .A1(n2193), .A2(n2194), .A3(n2195), .A4(n2196), .ZN(busB[3])
         );
  OAI221_X2 U129 ( .B1(n4905), .B2(n3756), .C1(n4898), .C2(n3577), .A(n2199), 
        .ZN(n2198) );
  AOI22_X2 U130 ( .A1(\reg_out[5][3] ), .A2(n4889), .B1(\reg_out[7][3] ), .B2(
        n4885), .ZN(n2199) );
  OAI221_X2 U131 ( .B1(n4878), .B2(n3993), .C1(n4871), .C2(n3718), .A(n2200), 
        .ZN(n2197) );
  AOI22_X2 U132 ( .A1(\reg_out[1][3] ), .A2(n4865), .B1(\reg_out[3][3] ), .B2(
        n4857), .ZN(n2200) );
  OAI221_X2 U134 ( .B1(n4905), .B2(n3992), .C1(n4898), .C2(n3717), .A(n2203), 
        .ZN(n2202) );
  AOI22_X2 U135 ( .A1(\reg_out[21][3] ), .A2(n4890), .B1(\reg_out[23][3] ), 
        .B2(n4885), .ZN(n2203) );
  OAI221_X2 U136 ( .B1(n4878), .B2(n3991), .C1(n4871), .C2(n3716), .A(n2204), 
        .ZN(n2201) );
  AOI22_X2 U137 ( .A1(\reg_out[17][3] ), .A2(n4865), .B1(\reg_out[19][3] ), 
        .B2(n4857), .ZN(n2204) );
  OAI221_X2 U139 ( .B1(n4905), .B2(n3990), .C1(n4898), .C2(n3715), .A(n2207), 
        .ZN(n2206) );
  AOI22_X2 U140 ( .A1(\reg_out[13][3] ), .A2(n4888), .B1(\reg_out[15][3] ), 
        .B2(n4885), .ZN(n2207) );
  OAI221_X2 U141 ( .B1(n4878), .B2(n3755), .C1(n4871), .C2(n3864), .A(n2208), 
        .ZN(n2205) );
  AOI22_X2 U142 ( .A1(\reg_out[9][3] ), .A2(n4865), .B1(\reg_out[11][3] ), 
        .B2(n4857), .ZN(n2208) );
  OAI221_X2 U144 ( .B1(n4905), .B2(n3989), .C1(n4898), .C2(n3714), .A(n2211), 
        .ZN(n2210) );
  AOI22_X2 U145 ( .A1(\reg_out[29][3] ), .A2(n4891), .B1(\reg_out[31][3] ), 
        .B2(n4885), .ZN(n2211) );
  OAI221_X2 U146 ( .B1(n4878), .B2(n3988), .C1(n4871), .C2(n3713), .A(n2212), 
        .ZN(n2209) );
  AOI22_X2 U147 ( .A1(\reg_out[25][3] ), .A2(n4865), .B1(\reg_out[27][3] ), 
        .B2(n4857), .ZN(n2212) );
  NAND4_X2 U148 ( .A1(n2213), .A2(n2214), .A3(n2215), .A4(n2216), .ZN(busB[31]) );
  OAI221_X2 U150 ( .B1(n4905), .B2(n3754), .C1(n4898), .C2(n3576), .A(n2219), 
        .ZN(n2218) );
  AOI22_X2 U151 ( .A1(\reg_out[5][31] ), .A2(n4891), .B1(\reg_out[7][31] ), 
        .B2(n4885), .ZN(n2219) );
  OAI221_X2 U152 ( .B1(n4878), .B2(n3987), .C1(n4871), .C2(n3712), .A(n2220), 
        .ZN(n2217) );
  AOI22_X2 U153 ( .A1(\reg_out[1][31] ), .A2(n4865), .B1(\reg_out[3][31] ), 
        .B2(n4857), .ZN(n2220) );
  OAI221_X2 U155 ( .B1(n4903), .B2(n3617), .C1(n4896), .C2(n3540), .A(n2223), 
        .ZN(n2222) );
  AOI22_X2 U156 ( .A1(\reg_out[21][31] ), .A2(n4890), .B1(\reg_out[23][31] ), 
        .B2(n4884), .ZN(n2223) );
  OAI221_X2 U157 ( .B1(n4877), .B2(n3616), .C1(n4870), .C2(n3539), .A(n2224), 
        .ZN(n2221) );
  AOI22_X2 U158 ( .A1(\reg_out[17][31] ), .A2(n4863), .B1(\reg_out[19][31] ), 
        .B2(n4855), .ZN(n2224) );
  OAI221_X2 U160 ( .B1(n4904), .B2(n3615), .C1(n4897), .C2(n3538), .A(n2227), 
        .ZN(n2226) );
  AOI22_X2 U161 ( .A1(\reg_out[13][31] ), .A2(n4891), .B1(\reg_out[15][31] ), 
        .B2(n4884), .ZN(n2227) );
  OAI221_X2 U162 ( .B1(n4876), .B2(n3614), .C1(n4869), .C2(n3537), .A(n2228), 
        .ZN(n2225) );
  AOI22_X2 U163 ( .A1(\reg_out[9][31] ), .A2(n4864), .B1(\reg_out[11][31] ), 
        .B2(n4853), .ZN(n2228) );
  OAI221_X2 U165 ( .B1(n4903), .B2(n3613), .C1(n4896), .C2(n3536), .A(n2231), 
        .ZN(n2230) );
  AOI22_X2 U166 ( .A1(\reg_out[29][31] ), .A2(n4890), .B1(\reg_out[31][31] ), 
        .B2(n4884), .ZN(n2231) );
  OAI221_X2 U167 ( .B1(n4877), .B2(n3612), .C1(n4870), .C2(n3535), .A(n2232), 
        .ZN(n2229) );
  AOI22_X2 U168 ( .A1(\reg_out[25][31] ), .A2(n4863), .B1(\reg_out[27][31] ), 
        .B2(n4855), .ZN(n2232) );
  NAND4_X2 U169 ( .A1(n2233), .A2(n2234), .A3(n2235), .A4(n2236), .ZN(busB[30]) );
  OAI221_X2 U171 ( .B1(n4903), .B2(n3611), .C1(n4896), .C2(n3534), .A(n2239), 
        .ZN(n2238) );
  AOI22_X2 U172 ( .A1(\reg_out[5][30] ), .A2(n4890), .B1(\reg_out[7][30] ), 
        .B2(n4883), .ZN(n2239) );
  OAI221_X2 U173 ( .B1(n4877), .B2(n3610), .C1(n4870), .C2(n3533), .A(n2240), 
        .ZN(n2237) );
  AOI22_X2 U174 ( .A1(\reg_out[1][30] ), .A2(n4863), .B1(\reg_out[3][30] ), 
        .B2(n4855), .ZN(n2240) );
  OAI221_X2 U176 ( .B1(n4904), .B2(n3609), .C1(n4897), .C2(n3532), .A(n2243), 
        .ZN(n2242) );
  AOI22_X2 U177 ( .A1(\reg_out[21][30] ), .A2(n4891), .B1(\reg_out[23][30] ), 
        .B2(n4884), .ZN(n2243) );
  OAI221_X2 U178 ( .B1(n4876), .B2(n3608), .C1(n4869), .C2(n3531), .A(n2244), 
        .ZN(n2241) );
  AOI22_X2 U179 ( .A1(\reg_out[17][30] ), .A2(n4864), .B1(\reg_out[19][30] ), 
        .B2(n4855), .ZN(n2244) );
  OAI221_X2 U181 ( .B1(n4903), .B2(n3607), .C1(n4896), .C2(n3530), .A(n2247), 
        .ZN(n2246) );
  AOI22_X2 U182 ( .A1(\reg_out[13][30] ), .A2(n4890), .B1(\reg_out[15][30] ), 
        .B2(n4883), .ZN(n2247) );
  OAI221_X2 U183 ( .B1(n4877), .B2(n3606), .C1(n4870), .C2(n3529), .A(n2248), 
        .ZN(n2245) );
  AOI22_X2 U184 ( .A1(\reg_out[9][30] ), .A2(n4863), .B1(\reg_out[11][30] ), 
        .B2(n4856), .ZN(n2248) );
  OAI221_X2 U186 ( .B1(n4904), .B2(n3605), .C1(n4897), .C2(n3528), .A(n2251), 
        .ZN(n2250) );
  AOI22_X2 U187 ( .A1(\reg_out[29][30] ), .A2(n4891), .B1(\reg_out[31][30] ), 
        .B2(n4883), .ZN(n2251) );
  OAI221_X2 U188 ( .B1(n4876), .B2(n3604), .C1(n4869), .C2(n3527), .A(n2252), 
        .ZN(n2249) );
  AOI22_X2 U189 ( .A1(\reg_out[25][30] ), .A2(n4864), .B1(\reg_out[27][30] ), 
        .B2(n4853), .ZN(n2252) );
  NAND4_X2 U190 ( .A1(n2253), .A2(n2254), .A3(n2255), .A4(n2256), .ZN(busB[2])
         );
  OAI221_X2 U192 ( .B1(n4904), .B2(n3603), .C1(n4897), .C2(n3526), .A(n2259), 
        .ZN(n2258) );
  AOI22_X2 U193 ( .A1(\reg_out[5][2] ), .A2(n4891), .B1(\reg_out[7][2] ), .B2(
        n4884), .ZN(n2259) );
  OAI221_X2 U194 ( .B1(n4876), .B2(n3602), .C1(n4869), .C2(n3525), .A(n2260), 
        .ZN(n2257) );
  AOI22_X2 U195 ( .A1(\reg_out[1][2] ), .A2(n4864), .B1(\reg_out[3][2] ), .B2(
        n4856), .ZN(n2260) );
  OAI221_X2 U197 ( .B1(n4903), .B2(n3601), .C1(n4896), .C2(n3524), .A(n2263), 
        .ZN(n2262) );
  AOI22_X2 U198 ( .A1(\reg_out[21][2] ), .A2(n4890), .B1(\reg_out[23][2] ), 
        .B2(n4883), .ZN(n2263) );
  OAI221_X2 U199 ( .B1(n4877), .B2(n3600), .C1(n4870), .C2(n3523), .A(n2264), 
        .ZN(n2261) );
  AOI22_X2 U200 ( .A1(\reg_out[17][2] ), .A2(n4863), .B1(\reg_out[19][2] ), 
        .B2(n4856), .ZN(n2264) );
  OAI221_X2 U202 ( .B1(n4904), .B2(n3599), .C1(n4897), .C2(n3522), .A(n2267), 
        .ZN(n2266) );
  AOI22_X2 U203 ( .A1(\reg_out[13][2] ), .A2(n4891), .B1(\reg_out[15][2] ), 
        .B2(n4883), .ZN(n2267) );
  OAI221_X2 U204 ( .B1(n4876), .B2(n3598), .C1(n4869), .C2(n3521), .A(n2268), 
        .ZN(n2265) );
  AOI22_X2 U205 ( .A1(\reg_out[9][2] ), .A2(n4864), .B1(\reg_out[11][2] ), 
        .B2(n4854), .ZN(n2268) );
  OAI221_X2 U207 ( .B1(n4903), .B2(n3597), .C1(n4896), .C2(n3520), .A(n2271), 
        .ZN(n2270) );
  AOI22_X2 U208 ( .A1(\reg_out[29][2] ), .A2(n4888), .B1(\reg_out[31][2] ), 
        .B2(n4884), .ZN(n2271) );
  OAI221_X2 U209 ( .B1(n4877), .B2(n3596), .C1(n4870), .C2(n3519), .A(n2272), 
        .ZN(n2269) );
  AOI22_X2 U210 ( .A1(\reg_out[25][2] ), .A2(n4861), .B1(\reg_out[27][2] ), 
        .B2(n4856), .ZN(n2272) );
  NAND4_X2 U211 ( .A1(n2273), .A2(n2274), .A3(n2275), .A4(n2276), .ZN(busB[29]) );
  OAI221_X2 U213 ( .B1(n4904), .B2(n3986), .C1(n4897), .C2(n3711), .A(n2279), 
        .ZN(n2278) );
  AOI22_X2 U214 ( .A1(\reg_out[5][29] ), .A2(n4891), .B1(\reg_out[7][29] ), 
        .B2(n4884), .ZN(n2279) );
  OAI221_X2 U215 ( .B1(n4877), .B2(n4486), .C1(n4870), .C2(n3863), .A(n2280), 
        .ZN(n2277) );
  AOI22_X2 U216 ( .A1(\reg_out[1][29] ), .A2(n4864), .B1(\reg_out[3][29] ), 
        .B2(n4856), .ZN(n2280) );
  OAI221_X2 U218 ( .B1(n4904), .B2(n4485), .C1(n4897), .C2(n3862), .A(n2283), 
        .ZN(n2282) );
  AOI22_X2 U219 ( .A1(\reg_out[21][29] ), .A2(n4891), .B1(\reg_out[23][29] ), 
        .B2(n4884), .ZN(n2283) );
  OAI221_X2 U220 ( .B1(n4877), .B2(n4484), .C1(n4870), .C2(n3861), .A(n2284), 
        .ZN(n2281) );
  AOI22_X2 U221 ( .A1(\reg_out[17][29] ), .A2(n4864), .B1(\reg_out[19][29] ), 
        .B2(n4856), .ZN(n2284) );
  OAI221_X2 U223 ( .B1(n4904), .B2(n4483), .C1(n4897), .C2(n3860), .A(n2287), 
        .ZN(n2286) );
  AOI22_X2 U224 ( .A1(\reg_out[13][29] ), .A2(n4891), .B1(\reg_out[15][29] ), 
        .B2(n4884), .ZN(n2287) );
  OAI221_X2 U225 ( .B1(n4877), .B2(n3985), .C1(n4870), .C2(n4437), .A(n2288), 
        .ZN(n2285) );
  AOI22_X2 U226 ( .A1(\reg_out[9][29] ), .A2(n4864), .B1(\reg_out[11][29] ), 
        .B2(n4856), .ZN(n2288) );
  OAI221_X2 U228 ( .B1(n4904), .B2(n4482), .C1(n4897), .C2(n3859), .A(n2291), 
        .ZN(n2290) );
  AOI22_X2 U229 ( .A1(\reg_out[29][29] ), .A2(n4891), .B1(\reg_out[31][29] ), 
        .B2(n4884), .ZN(n2291) );
  OAI221_X2 U230 ( .B1(n4877), .B2(n4481), .C1(n4870), .C2(n3858), .A(n2292), 
        .ZN(n2289) );
  AOI22_X2 U231 ( .A1(\reg_out[25][29] ), .A2(n4864), .B1(\reg_out[27][29] ), 
        .B2(n4856), .ZN(n2292) );
  NAND4_X2 U232 ( .A1(n2293), .A2(n2294), .A3(n2295), .A4(n2296), .ZN(busB[28]) );
  OAI221_X2 U234 ( .B1(n4904), .B2(n3984), .C1(n4897), .C2(n3710), .A(n2299), 
        .ZN(n2298) );
  AOI22_X2 U235 ( .A1(\reg_out[5][28] ), .A2(n4891), .B1(\reg_out[7][28] ), 
        .B2(n4884), .ZN(n2299) );
  OAI221_X2 U236 ( .B1(n4877), .B2(n3983), .C1(n4870), .C2(n3709), .A(n2300), 
        .ZN(n2297) );
  AOI22_X2 U237 ( .A1(\reg_out[1][28] ), .A2(n4864), .B1(\reg_out[3][28] ), 
        .B2(n4856), .ZN(n2300) );
  OAI221_X2 U239 ( .B1(n4904), .B2(n3982), .C1(n4897), .C2(n3708), .A(n2303), 
        .ZN(n2302) );
  AOI22_X2 U240 ( .A1(\reg_out[21][28] ), .A2(n4891), .B1(\reg_out[23][28] ), 
        .B2(n4884), .ZN(n2303) );
  OAI221_X2 U241 ( .B1(n4877), .B2(n3981), .C1(n4870), .C2(n3707), .A(n2304), 
        .ZN(n2301) );
  AOI22_X2 U242 ( .A1(\reg_out[17][28] ), .A2(n4864), .B1(\reg_out[19][28] ), 
        .B2(n4856), .ZN(n2304) );
  OAI221_X2 U244 ( .B1(n4904), .B2(n3980), .C1(n4897), .C2(n3706), .A(n2307), 
        .ZN(n2306) );
  AOI22_X2 U245 ( .A1(\reg_out[13][28] ), .A2(n4891), .B1(\reg_out[15][28] ), 
        .B2(n4884), .ZN(n2307) );
  OAI221_X2 U246 ( .B1(n4877), .B2(n3979), .C1(n4870), .C2(n3705), .A(n2308), 
        .ZN(n2305) );
  AOI22_X2 U247 ( .A1(\reg_out[9][28] ), .A2(n4864), .B1(\reg_out[11][28] ), 
        .B2(n4856), .ZN(n2308) );
  OAI221_X2 U249 ( .B1(n4904), .B2(n3978), .C1(n4897), .C2(n3704), .A(n2311), 
        .ZN(n2310) );
  AOI22_X2 U250 ( .A1(\reg_out[29][28] ), .A2(n4891), .B1(\reg_out[31][28] ), 
        .B2(n4884), .ZN(n2311) );
  OAI221_X2 U251 ( .B1(n4877), .B2(n3977), .C1(n4870), .C2(n3703), .A(n2312), 
        .ZN(n2309) );
  AOI22_X2 U252 ( .A1(\reg_out[25][28] ), .A2(n4864), .B1(\reg_out[27][28] ), 
        .B2(n4856), .ZN(n2312) );
  NAND4_X2 U253 ( .A1(n2313), .A2(n2314), .A3(n2315), .A4(n2316), .ZN(busB[27]) );
  OAI221_X2 U255 ( .B1(n4904), .B2(n3976), .C1(n4897), .C2(n3702), .A(n2319), 
        .ZN(n2318) );
  AOI22_X2 U256 ( .A1(\reg_out[5][27] ), .A2(n4891), .B1(\reg_out[7][27] ), 
        .B2(n4884), .ZN(n2319) );
  OAI221_X2 U257 ( .B1(n4877), .B2(n3975), .C1(n4870), .C2(n3701), .A(n2320), 
        .ZN(n2317) );
  AOI22_X2 U258 ( .A1(\reg_out[1][27] ), .A2(n4864), .B1(\reg_out[3][27] ), 
        .B2(n4856), .ZN(n2320) );
  OAI221_X2 U260 ( .B1(n4904), .B2(n3974), .C1(n4897), .C2(n3700), .A(n2323), 
        .ZN(n2322) );
  AOI22_X2 U261 ( .A1(\reg_out[21][27] ), .A2(n4891), .B1(\reg_out[23][27] ), 
        .B2(n4884), .ZN(n2323) );
  OAI221_X2 U262 ( .B1(n4877), .B2(n3973), .C1(n4870), .C2(n3699), .A(n2324), 
        .ZN(n2321) );
  AOI22_X2 U263 ( .A1(\reg_out[17][27] ), .A2(n4864), .B1(\reg_out[19][27] ), 
        .B2(n4856), .ZN(n2324) );
  OAI221_X2 U265 ( .B1(n4904), .B2(n3972), .C1(n4897), .C2(n3698), .A(n2327), 
        .ZN(n2326) );
  AOI22_X2 U266 ( .A1(\reg_out[13][27] ), .A2(n4891), .B1(\reg_out[15][27] ), 
        .B2(n4884), .ZN(n2327) );
  OAI221_X2 U267 ( .B1(n4877), .B2(n3971), .C1(n4870), .C2(n3697), .A(n2328), 
        .ZN(n2325) );
  AOI22_X2 U268 ( .A1(\reg_out[9][27] ), .A2(n4864), .B1(\reg_out[11][27] ), 
        .B2(n4856), .ZN(n2328) );
  OAI221_X2 U270 ( .B1(n4903), .B2(n3970), .C1(n4896), .C2(n3696), .A(n2331), 
        .ZN(n2330) );
  AOI22_X2 U271 ( .A1(\reg_out[29][27] ), .A2(n4890), .B1(\reg_out[31][27] ), 
        .B2(n4883), .ZN(n2331) );
  OAI221_X2 U272 ( .B1(n4876), .B2(n3969), .C1(n4869), .C2(n3695), .A(n2332), 
        .ZN(n2329) );
  AOI22_X2 U273 ( .A1(\reg_out[25][27] ), .A2(n4863), .B1(\reg_out[27][27] ), 
        .B2(n4855), .ZN(n2332) );
  NAND4_X2 U274 ( .A1(n2333), .A2(n2334), .A3(n2335), .A4(n2336), .ZN(busB[26]) );
  OAI221_X2 U276 ( .B1(n4903), .B2(n3968), .C1(n4896), .C2(n3694), .A(n2339), 
        .ZN(n2338) );
  AOI22_X2 U277 ( .A1(\reg_out[5][26] ), .A2(n4890), .B1(\reg_out[7][26] ), 
        .B2(n4883), .ZN(n2339) );
  OAI221_X2 U278 ( .B1(n4876), .B2(n3967), .C1(n4869), .C2(n3693), .A(n2340), 
        .ZN(n2337) );
  AOI22_X2 U279 ( .A1(\reg_out[1][26] ), .A2(n4863), .B1(\reg_out[3][26] ), 
        .B2(n4855), .ZN(n2340) );
  OAI221_X2 U281 ( .B1(n4903), .B2(n3966), .C1(n4896), .C2(n3692), .A(n2343), 
        .ZN(n2342) );
  AOI22_X2 U282 ( .A1(\reg_out[21][26] ), .A2(n4890), .B1(\reg_out[23][26] ), 
        .B2(n4883), .ZN(n2343) );
  OAI221_X2 U283 ( .B1(n4876), .B2(n3965), .C1(n4869), .C2(n3691), .A(n2344), 
        .ZN(n2341) );
  AOI22_X2 U284 ( .A1(\reg_out[17][26] ), .A2(n4863), .B1(\reg_out[19][26] ), 
        .B2(n4855), .ZN(n2344) );
  OAI221_X2 U286 ( .B1(n4903), .B2(n3964), .C1(n4896), .C2(n3690), .A(n2347), 
        .ZN(n2346) );
  AOI22_X2 U287 ( .A1(\reg_out[13][26] ), .A2(n4890), .B1(\reg_out[15][26] ), 
        .B2(n4883), .ZN(n2347) );
  OAI221_X2 U288 ( .B1(n4876), .B2(n3963), .C1(n4869), .C2(n3689), .A(n2348), 
        .ZN(n2345) );
  AOI22_X2 U289 ( .A1(\reg_out[9][26] ), .A2(n4863), .B1(\reg_out[11][26] ), 
        .B2(n4855), .ZN(n2348) );
  OAI221_X2 U291 ( .B1(n4903), .B2(n3962), .C1(n4896), .C2(n3688), .A(n2351), 
        .ZN(n2350) );
  AOI22_X2 U292 ( .A1(\reg_out[29][26] ), .A2(n4890), .B1(\reg_out[31][26] ), 
        .B2(n4883), .ZN(n2351) );
  OAI221_X2 U293 ( .B1(n4876), .B2(n3961), .C1(n4869), .C2(n3687), .A(n2352), 
        .ZN(n2349) );
  AOI22_X2 U294 ( .A1(\reg_out[25][26] ), .A2(n4863), .B1(\reg_out[27][26] ), 
        .B2(n4855), .ZN(n2352) );
  NAND4_X2 U295 ( .A1(n2353), .A2(n2354), .A3(n2355), .A4(n2356), .ZN(busB[25]) );
  OAI221_X2 U297 ( .B1(n4903), .B2(n3960), .C1(n4896), .C2(n3686), .A(n2359), 
        .ZN(n2358) );
  AOI22_X2 U298 ( .A1(\reg_out[5][25] ), .A2(n4890), .B1(\reg_out[7][25] ), 
        .B2(n4883), .ZN(n2359) );
  OAI221_X2 U299 ( .B1(n4876), .B2(n3959), .C1(n4869), .C2(n3685), .A(n2360), 
        .ZN(n2357) );
  AOI22_X2 U300 ( .A1(\reg_out[1][25] ), .A2(n4863), .B1(\reg_out[3][25] ), 
        .B2(n4855), .ZN(n2360) );
  OAI221_X2 U302 ( .B1(n4903), .B2(n3958), .C1(n4896), .C2(n3684), .A(n2363), 
        .ZN(n2362) );
  AOI22_X2 U303 ( .A1(\reg_out[21][25] ), .A2(n4890), .B1(\reg_out[23][25] ), 
        .B2(n4883), .ZN(n2363) );
  OAI221_X2 U304 ( .B1(n4876), .B2(n3957), .C1(n4869), .C2(n3683), .A(n2364), 
        .ZN(n2361) );
  AOI22_X2 U305 ( .A1(\reg_out[17][25] ), .A2(n4863), .B1(\reg_out[19][25] ), 
        .B2(n4855), .ZN(n2364) );
  OAI221_X2 U307 ( .B1(n4903), .B2(n3956), .C1(n4896), .C2(n3682), .A(n2367), 
        .ZN(n2366) );
  AOI22_X2 U308 ( .A1(\reg_out[13][25] ), .A2(n4890), .B1(\reg_out[15][25] ), 
        .B2(n4883), .ZN(n2367) );
  OAI221_X2 U309 ( .B1(n4876), .B2(n3955), .C1(n4869), .C2(n3681), .A(n2368), 
        .ZN(n2365) );
  AOI22_X2 U310 ( .A1(\reg_out[9][25] ), .A2(n4863), .B1(\reg_out[11][25] ), 
        .B2(n4855), .ZN(n2368) );
  OAI221_X2 U312 ( .B1(n4903), .B2(n3954), .C1(n4896), .C2(n3680), .A(n2371), 
        .ZN(n2370) );
  AOI22_X2 U313 ( .A1(\reg_out[29][25] ), .A2(n4890), .B1(\reg_out[31][25] ), 
        .B2(n4883), .ZN(n2371) );
  OAI221_X2 U314 ( .B1(n4876), .B2(n3953), .C1(n4869), .C2(n3679), .A(n2372), 
        .ZN(n2369) );
  AOI22_X2 U315 ( .A1(\reg_out[25][25] ), .A2(n4863), .B1(\reg_out[27][25] ), 
        .B2(n4855), .ZN(n2372) );
  NAND4_X2 U316 ( .A1(n2373), .A2(n2374), .A3(n2375), .A4(n2376), .ZN(busB[24]) );
  OAI221_X2 U318 ( .B1(n4903), .B2(n3952), .C1(n4896), .C2(n3678), .A(n2379), 
        .ZN(n2378) );
  AOI22_X2 U319 ( .A1(\reg_out[5][24] ), .A2(n4890), .B1(\reg_out[7][24] ), 
        .B2(n4883), .ZN(n2379) );
  OAI221_X2 U320 ( .B1(n4876), .B2(n3951), .C1(n4869), .C2(n3677), .A(n2380), 
        .ZN(n2377) );
  AOI22_X2 U321 ( .A1(\reg_out[1][24] ), .A2(n4863), .B1(\reg_out[3][24] ), 
        .B2(n4855), .ZN(n2380) );
  OAI221_X2 U323 ( .B1(n4903), .B2(n3950), .C1(n4896), .C2(n3676), .A(n2383), 
        .ZN(n2382) );
  AOI22_X2 U324 ( .A1(\reg_out[21][24] ), .A2(n4890), .B1(\reg_out[23][24] ), 
        .B2(n4883), .ZN(n2383) );
  OAI221_X2 U325 ( .B1(n4876), .B2(n3949), .C1(n4869), .C2(n3675), .A(n2384), 
        .ZN(n2381) );
  AOI22_X2 U326 ( .A1(\reg_out[17][24] ), .A2(n4863), .B1(\reg_out[19][24] ), 
        .B2(n4855), .ZN(n2384) );
  OAI221_X2 U328 ( .B1(n4902), .B2(n3948), .C1(n4895), .C2(n3518), .A(n2387), 
        .ZN(n2386) );
  AOI22_X2 U329 ( .A1(\reg_out[13][24] ), .A2(n4889), .B1(\reg_out[15][24] ), 
        .B2(n4882), .ZN(n2387) );
  OAI221_X2 U330 ( .B1(n4875), .B2(n3947), .C1(n4868), .C2(n3517), .A(n2388), 
        .ZN(n2385) );
  AOI22_X2 U331 ( .A1(\reg_out[9][24] ), .A2(n4862), .B1(\reg_out[11][24] ), 
        .B2(n4854), .ZN(n2388) );
  OAI221_X2 U333 ( .B1(n4901), .B2(n3946), .C1(n4894), .C2(n3516), .A(n2391), 
        .ZN(n2390) );
  AOI22_X2 U334 ( .A1(\reg_out[29][24] ), .A2(n4889), .B1(\reg_out[31][24] ), 
        .B2(n4882), .ZN(n2391) );
  OAI221_X2 U335 ( .B1(n4874), .B2(n3945), .C1(n4867), .C2(n3515), .A(n2392), 
        .ZN(n2389) );
  AOI22_X2 U336 ( .A1(\reg_out[25][24] ), .A2(n4862), .B1(\reg_out[27][24] ), 
        .B2(n4854), .ZN(n2392) );
  NAND4_X2 U337 ( .A1(n2393), .A2(n2394), .A3(n2395), .A4(n2396), .ZN(busB[23]) );
  OAI221_X2 U339 ( .B1(n4901), .B2(n3944), .C1(n4894), .C2(n3514), .A(n2399), 
        .ZN(n2398) );
  AOI22_X2 U340 ( .A1(\reg_out[5][23] ), .A2(n4889), .B1(\reg_out[7][23] ), 
        .B2(n4882), .ZN(n2399) );
  OAI221_X2 U341 ( .B1(n4874), .B2(n3943), .C1(n4867), .C2(n3513), .A(n2400), 
        .ZN(n2397) );
  AOI22_X2 U342 ( .A1(\reg_out[1][23] ), .A2(n4862), .B1(\reg_out[3][23] ), 
        .B2(n4854), .ZN(n2400) );
  OAI221_X2 U344 ( .B1(n4902), .B2(n3942), .C1(n4895), .C2(n3512), .A(n2403), 
        .ZN(n2402) );
  AOI22_X2 U345 ( .A1(\reg_out[21][23] ), .A2(n4889), .B1(\reg_out[23][23] ), 
        .B2(n4882), .ZN(n2403) );
  OAI221_X2 U346 ( .B1(n4875), .B2(n3941), .C1(n4868), .C2(n3511), .A(n2404), 
        .ZN(n2401) );
  AOI22_X2 U347 ( .A1(\reg_out[17][23] ), .A2(n4862), .B1(\reg_out[19][23] ), 
        .B2(n4854), .ZN(n2404) );
  OAI221_X2 U349 ( .B1(n4901), .B2(n3940), .C1(n4894), .C2(n3510), .A(n2407), 
        .ZN(n2406) );
  AOI22_X2 U350 ( .A1(\reg_out[13][23] ), .A2(n4889), .B1(\reg_out[15][23] ), 
        .B2(n4881), .ZN(n2407) );
  OAI221_X2 U351 ( .B1(n4874), .B2(n3939), .C1(n4867), .C2(n3509), .A(n2408), 
        .ZN(n2405) );
  AOI22_X2 U352 ( .A1(\reg_out[9][23] ), .A2(n4862), .B1(\reg_out[11][23] ), 
        .B2(n4854), .ZN(n2408) );
  OAI221_X2 U354 ( .B1(n4902), .B2(n3938), .C1(n4895), .C2(n3508), .A(n2411), 
        .ZN(n2410) );
  AOI22_X2 U355 ( .A1(\reg_out[29][23] ), .A2(n4889), .B1(\reg_out[31][23] ), 
        .B2(n4882), .ZN(n2411) );
  OAI221_X2 U356 ( .B1(n4875), .B2(n3937), .C1(n4868), .C2(n3507), .A(n2412), 
        .ZN(n2409) );
  AOI22_X2 U357 ( .A1(\reg_out[25][23] ), .A2(n4862), .B1(\reg_out[27][23] ), 
        .B2(n4854), .ZN(n2412) );
  NAND4_X2 U358 ( .A1(n2413), .A2(n2414), .A3(n2415), .A4(n2416), .ZN(busB[22]) );
  OAI221_X2 U360 ( .B1(n4902), .B2(n3936), .C1(n4895), .C2(n3506), .A(n2419), 
        .ZN(n2418) );
  AOI22_X2 U361 ( .A1(\reg_out[5][22] ), .A2(n4889), .B1(\reg_out[7][22] ), 
        .B2(n4882), .ZN(n2419) );
  OAI221_X2 U362 ( .B1(n4875), .B2(n3935), .C1(n4868), .C2(n3505), .A(n2420), 
        .ZN(n2417) );
  AOI22_X2 U363 ( .A1(\reg_out[1][22] ), .A2(n4862), .B1(\reg_out[3][22] ), 
        .B2(n4854), .ZN(n2420) );
  OAI221_X2 U365 ( .B1(n4901), .B2(n3934), .C1(n4894), .C2(n3504), .A(n2423), 
        .ZN(n2422) );
  AOI22_X2 U366 ( .A1(\reg_out[21][22] ), .A2(n4889), .B1(\reg_out[23][22] ), 
        .B2(n4881), .ZN(n2423) );
  OAI221_X2 U367 ( .B1(n4874), .B2(n3933), .C1(n4867), .C2(n3503), .A(n2424), 
        .ZN(n2421) );
  AOI22_X2 U368 ( .A1(\reg_out[17][22] ), .A2(n4862), .B1(\reg_out[19][22] ), 
        .B2(n4854), .ZN(n2424) );
  OAI221_X2 U370 ( .B1(n4902), .B2(n3932), .C1(n4895), .C2(n3502), .A(n2427), 
        .ZN(n2426) );
  AOI22_X2 U371 ( .A1(\reg_out[13][22] ), .A2(n4889), .B1(\reg_out[15][22] ), 
        .B2(n4881), .ZN(n2427) );
  OAI221_X2 U372 ( .B1(n4875), .B2(n3931), .C1(n4868), .C2(n3501), .A(n2428), 
        .ZN(n2425) );
  AOI22_X2 U373 ( .A1(\reg_out[9][22] ), .A2(n4862), .B1(\reg_out[11][22] ), 
        .B2(n4854), .ZN(n2428) );
  OAI221_X2 U375 ( .B1(n4901), .B2(n3930), .C1(n4894), .C2(n3500), .A(n2431), 
        .ZN(n2430) );
  AOI22_X2 U376 ( .A1(\reg_out[29][22] ), .A2(n4889), .B1(\reg_out[31][22] ), 
        .B2(n4881), .ZN(n2431) );
  OAI221_X2 U377 ( .B1(n4874), .B2(n3929), .C1(n4867), .C2(n3499), .A(n2432), 
        .ZN(n2429) );
  AOI22_X2 U378 ( .A1(\reg_out[25][22] ), .A2(n4862), .B1(\reg_out[27][22] ), 
        .B2(n4854), .ZN(n2432) );
  NAND4_X2 U379 ( .A1(n2433), .A2(n2434), .A3(n2435), .A4(n2436), .ZN(busB[21]) );
  OAI221_X2 U381 ( .B1(n4901), .B2(n3928), .C1(n4894), .C2(n3498), .A(n2439), 
        .ZN(n2438) );
  AOI22_X2 U382 ( .A1(\reg_out[5][21] ), .A2(n4889), .B1(\reg_out[7][21] ), 
        .B2(n4881), .ZN(n2439) );
  OAI221_X2 U383 ( .B1(n4874), .B2(n3927), .C1(n4867), .C2(n3497), .A(n2440), 
        .ZN(n2437) );
  AOI22_X2 U384 ( .A1(\reg_out[1][21] ), .A2(n4862), .B1(\reg_out[3][21] ), 
        .B2(n4854), .ZN(n2440) );
  OAI221_X2 U386 ( .B1(n4902), .B2(n3926), .C1(n4895), .C2(n3674), .A(n2443), 
        .ZN(n2442) );
  AOI22_X2 U387 ( .A1(\reg_out[21][21] ), .A2(n4889), .B1(\reg_out[23][21] ), 
        .B2(n4882), .ZN(n2443) );
  OAI221_X2 U388 ( .B1(n4875), .B2(n3925), .C1(n4868), .C2(n3673), .A(n2444), 
        .ZN(n2441) );
  AOI22_X2 U389 ( .A1(\reg_out[17][21] ), .A2(n4862), .B1(\reg_out[19][21] ), 
        .B2(n4853), .ZN(n2444) );
  OAI221_X2 U391 ( .B1(n4902), .B2(n3924), .C1(n4895), .C2(n3672), .A(n2447), 
        .ZN(n2446) );
  AOI22_X2 U392 ( .A1(\reg_out[13][21] ), .A2(n4889), .B1(\reg_out[15][21] ), 
        .B2(n4882), .ZN(n2447) );
  OAI221_X2 U393 ( .B1(n4875), .B2(n3923), .C1(n4868), .C2(n3671), .A(n2448), 
        .ZN(n2445) );
  AOI22_X2 U394 ( .A1(\reg_out[9][21] ), .A2(n4862), .B1(\reg_out[11][21] ), 
        .B2(n4853), .ZN(n2448) );
  OAI221_X2 U396 ( .B1(n4902), .B2(n3922), .C1(n4895), .C2(n3670), .A(n2451), 
        .ZN(n2450) );
  AOI22_X2 U397 ( .A1(\reg_out[29][21] ), .A2(n4889), .B1(\reg_out[31][21] ), 
        .B2(n4882), .ZN(n2451) );
  OAI221_X2 U398 ( .B1(n4875), .B2(n3921), .C1(n4868), .C2(n3669), .A(n2452), 
        .ZN(n2449) );
  AOI22_X2 U399 ( .A1(\reg_out[25][21] ), .A2(n4862), .B1(\reg_out[27][21] ), 
        .B2(n4853), .ZN(n2452) );
  NAND4_X2 U400 ( .A1(n2453), .A2(n2454), .A3(n2455), .A4(n2456), .ZN(busB[20]) );
  OAI221_X2 U402 ( .B1(n4902), .B2(n3920), .C1(n4895), .C2(n3668), .A(n2459), 
        .ZN(n2458) );
  AOI22_X2 U403 ( .A1(\reg_out[5][20] ), .A2(n4889), .B1(\reg_out[7][20] ), 
        .B2(n4882), .ZN(n2459) );
  OAI221_X2 U404 ( .B1(n4875), .B2(n3919), .C1(n4868), .C2(n3667), .A(n2460), 
        .ZN(n2457) );
  AOI22_X2 U405 ( .A1(\reg_out[1][20] ), .A2(n4862), .B1(\reg_out[3][20] ), 
        .B2(n4853), .ZN(n2460) );
  OAI221_X2 U407 ( .B1(n4902), .B2(n3918), .C1(n4895), .C2(n3666), .A(n2463), 
        .ZN(n2462) );
  AOI22_X2 U408 ( .A1(\reg_out[21][20] ), .A2(n4889), .B1(\reg_out[23][20] ), 
        .B2(n4882), .ZN(n2463) );
  OAI221_X2 U409 ( .B1(n4875), .B2(n3917), .C1(n4868), .C2(n3665), .A(n2464), 
        .ZN(n2461) );
  AOI22_X2 U410 ( .A1(\reg_out[17][20] ), .A2(n4862), .B1(\reg_out[19][20] ), 
        .B2(n4853), .ZN(n2464) );
  OAI221_X2 U412 ( .B1(n4902), .B2(n3916), .C1(n4895), .C2(n3664), .A(n2467), 
        .ZN(n2466) );
  AOI22_X2 U413 ( .A1(\reg_out[13][20] ), .A2(n4889), .B1(\reg_out[15][20] ), 
        .B2(n4882), .ZN(n2467) );
  OAI221_X2 U414 ( .B1(n4875), .B2(n3915), .C1(n4868), .C2(n3663), .A(n2468), 
        .ZN(n2465) );
  AOI22_X2 U415 ( .A1(\reg_out[9][20] ), .A2(n4862), .B1(\reg_out[11][20] ), 
        .B2(n4853), .ZN(n2468) );
  OAI221_X2 U417 ( .B1(n4902), .B2(n3914), .C1(n4895), .C2(n3662), .A(n2471), 
        .ZN(n2470) );
  AOI22_X2 U418 ( .A1(\reg_out[29][20] ), .A2(n4889), .B1(\reg_out[31][20] ), 
        .B2(n4882), .ZN(n2471) );
  OAI221_X2 U419 ( .B1(n4875), .B2(n3913), .C1(n4868), .C2(n3661), .A(n2472), 
        .ZN(n2469) );
  AOI22_X2 U420 ( .A1(\reg_out[25][20] ), .A2(n4862), .B1(\reg_out[27][20] ), 
        .B2(n4853), .ZN(n2472) );
  NAND4_X2 U421 ( .A1(n2473), .A2(n2474), .A3(n2475), .A4(n2476), .ZN(busB[1])
         );
  OAI221_X2 U423 ( .B1(n4902), .B2(n3912), .C1(n4895), .C2(n3660), .A(n2479), 
        .ZN(n2478) );
  AOI22_X2 U424 ( .A1(\reg_out[5][1] ), .A2(n4889), .B1(\reg_out[7][1] ), .B2(
        n4882), .ZN(n2479) );
  OAI221_X2 U425 ( .B1(n4875), .B2(n3911), .C1(n4868), .C2(n3659), .A(n2480), 
        .ZN(n2477) );
  AOI22_X2 U426 ( .A1(\reg_out[1][1] ), .A2(n4862), .B1(\reg_out[3][1] ), .B2(
        n4853), .ZN(n2480) );
  OAI221_X2 U428 ( .B1(n4902), .B2(n3910), .C1(n4895), .C2(n3658), .A(n2483), 
        .ZN(n2482) );
  AOI22_X2 U429 ( .A1(\reg_out[21][1] ), .A2(n4889), .B1(\reg_out[23][1] ), 
        .B2(n4882), .ZN(n2483) );
  OAI221_X2 U430 ( .B1(n4875), .B2(n3909), .C1(n4868), .C2(n3657), .A(n2484), 
        .ZN(n2481) );
  AOI22_X2 U431 ( .A1(\reg_out[17][1] ), .A2(n4862), .B1(\reg_out[19][1] ), 
        .B2(n4853), .ZN(n2484) );
  OAI221_X2 U433 ( .B1(n4902), .B2(n3908), .C1(n4895), .C2(n3656), .A(n2487), 
        .ZN(n2486) );
  AOI22_X2 U434 ( .A1(\reg_out[13][1] ), .A2(n4889), .B1(\reg_out[15][1] ), 
        .B2(n4882), .ZN(n2487) );
  OAI221_X2 U435 ( .B1(n4875), .B2(n3907), .C1(n4868), .C2(n3655), .A(n2488), 
        .ZN(n2485) );
  AOI22_X2 U436 ( .A1(\reg_out[9][1] ), .A2(n4862), .B1(\reg_out[11][1] ), 
        .B2(n4853), .ZN(n2488) );
  OAI221_X2 U438 ( .B1(n4902), .B2(n3906), .C1(n4895), .C2(n3654), .A(n2491), 
        .ZN(n2490) );
  AOI22_X2 U439 ( .A1(\reg_out[29][1] ), .A2(n4889), .B1(\reg_out[31][1] ), 
        .B2(n4882), .ZN(n2491) );
  OAI221_X2 U440 ( .B1(n4875), .B2(n3905), .C1(n4868), .C2(n3653), .A(n2492), 
        .ZN(n2489) );
  AOI22_X2 U441 ( .A1(\reg_out[25][1] ), .A2(n4862), .B1(\reg_out[27][1] ), 
        .B2(n4853), .ZN(n2492) );
  NAND4_X2 U442 ( .A1(n2493), .A2(n2494), .A3(n2495), .A4(n2496), .ZN(busB[19]) );
  OAI221_X2 U444 ( .B1(n4901), .B2(n3904), .C1(n4894), .C2(n3652), .A(n2499), 
        .ZN(n2498) );
  AOI22_X2 U445 ( .A1(\reg_out[5][19] ), .A2(n4888), .B1(\reg_out[7][19] ), 
        .B2(n4881), .ZN(n2499) );
  OAI221_X2 U446 ( .B1(n4874), .B2(n3903), .C1(n4867), .C2(n3651), .A(n2500), 
        .ZN(n2497) );
  AOI22_X2 U447 ( .A1(\reg_out[1][19] ), .A2(n4861), .B1(\reg_out[3][19] ), 
        .B2(n4854), .ZN(n2500) );
  OAI221_X2 U449 ( .B1(n4901), .B2(n3902), .C1(n4894), .C2(n3650), .A(n2503), 
        .ZN(n2502) );
  AOI22_X2 U450 ( .A1(\reg_out[21][19] ), .A2(n4888), .B1(\reg_out[23][19] ), 
        .B2(n4881), .ZN(n2503) );
  OAI221_X2 U451 ( .B1(n4874), .B2(n3901), .C1(n4867), .C2(n3649), .A(n2504), 
        .ZN(n2501) );
  AOI22_X2 U452 ( .A1(\reg_out[17][19] ), .A2(n4861), .B1(\reg_out[19][19] ), 
        .B2(n4854), .ZN(n2504) );
  OAI221_X2 U454 ( .B1(n4901), .B2(n3900), .C1(n4894), .C2(n3648), .A(n2507), 
        .ZN(n2506) );
  AOI22_X2 U455 ( .A1(\reg_out[13][19] ), .A2(n4888), .B1(\reg_out[15][19] ), 
        .B2(n4881), .ZN(n2507) );
  OAI221_X2 U456 ( .B1(n4874), .B2(n3899), .C1(n4867), .C2(n3647), .A(n2508), 
        .ZN(n2505) );
  AOI22_X2 U457 ( .A1(\reg_out[9][19] ), .A2(n4861), .B1(\reg_out[11][19] ), 
        .B2(n4854), .ZN(n2508) );
  OAI221_X2 U459 ( .B1(n4901), .B2(n3898), .C1(n4894), .C2(n3646), .A(n2511), 
        .ZN(n2510) );
  AOI22_X2 U460 ( .A1(\reg_out[29][19] ), .A2(n4888), .B1(\reg_out[31][19] ), 
        .B2(n4881), .ZN(n2511) );
  OAI221_X2 U461 ( .B1(n4874), .B2(n3897), .C1(n4867), .C2(n3645), .A(n2512), 
        .ZN(n2509) );
  AOI22_X2 U462 ( .A1(\reg_out[25][19] ), .A2(n4861), .B1(\reg_out[27][19] ), 
        .B2(n4854), .ZN(n2512) );
  NAND4_X2 U463 ( .A1(n2513), .A2(n2514), .A3(n2515), .A4(n2516), .ZN(busB[18]) );
  OAI221_X2 U465 ( .B1(n4901), .B2(n3896), .C1(n4894), .C2(n3644), .A(n2519), 
        .ZN(n2518) );
  AOI22_X2 U466 ( .A1(\reg_out[5][18] ), .A2(n4888), .B1(\reg_out[7][18] ), 
        .B2(n4881), .ZN(n2519) );
  OAI221_X2 U467 ( .B1(n4874), .B2(n4480), .C1(n4867), .C2(n3857), .A(n2520), 
        .ZN(n2517) );
  AOI22_X2 U468 ( .A1(\reg_out[1][18] ), .A2(n4861), .B1(\reg_out[3][18] ), 
        .B2(n4854), .ZN(n2520) );
  OAI221_X2 U470 ( .B1(n4901), .B2(n4479), .C1(n4894), .C2(n3643), .A(n2523), 
        .ZN(n2522) );
  AOI22_X2 U471 ( .A1(\reg_out[21][18] ), .A2(n4888), .B1(\reg_out[23][18] ), 
        .B2(n4881), .ZN(n2523) );
  OAI221_X2 U472 ( .B1(n4874), .B2(n4478), .C1(n4867), .C2(n3856), .A(n2524), 
        .ZN(n2521) );
  AOI22_X2 U473 ( .A1(\reg_out[17][18] ), .A2(n4861), .B1(\reg_out[19][18] ), 
        .B2(n4854), .ZN(n2524) );
  OAI221_X2 U475 ( .B1(n4901), .B2(n4477), .C1(n4894), .C2(n3855), .A(n2527), 
        .ZN(n2526) );
  AOI22_X2 U476 ( .A1(\reg_out[13][18] ), .A2(n4888), .B1(\reg_out[15][18] ), 
        .B2(n4881), .ZN(n2527) );
  OAI221_X2 U477 ( .B1(n4874), .B2(n3895), .C1(n4867), .C2(n4436), .A(n2528), 
        .ZN(n2525) );
  AOI22_X2 U478 ( .A1(\reg_out[9][18] ), .A2(n4861), .B1(\reg_out[11][18] ), 
        .B2(n4854), .ZN(n2528) );
  OAI221_X2 U480 ( .B1(n4901), .B2(n4476), .C1(n4894), .C2(n3854), .A(n2531), 
        .ZN(n2530) );
  AOI22_X2 U481 ( .A1(\reg_out[29][18] ), .A2(n4888), .B1(\reg_out[31][18] ), 
        .B2(n4881), .ZN(n2531) );
  OAI221_X2 U482 ( .B1(n4874), .B2(n4475), .C1(n4867), .C2(n3642), .A(n2532), 
        .ZN(n2529) );
  AOI22_X2 U483 ( .A1(\reg_out[25][18] ), .A2(n4861), .B1(\reg_out[27][18] ), 
        .B2(n4854), .ZN(n2532) );
  NAND4_X2 U484 ( .A1(n2533), .A2(n2534), .A3(n2535), .A4(n2536), .ZN(busB[17]) );
  OAI221_X2 U486 ( .B1(n4901), .B2(n3894), .C1(n4894), .C2(n3641), .A(n2539), 
        .ZN(n2538) );
  AOI22_X2 U487 ( .A1(\reg_out[5][17] ), .A2(n4888), .B1(\reg_out[7][17] ), 
        .B2(n4881), .ZN(n2539) );
  OAI221_X2 U488 ( .B1(n4874), .B2(n4474), .C1(n4867), .C2(n3853), .A(n2540), 
        .ZN(n2537) );
  AOI22_X2 U489 ( .A1(\reg_out[1][17] ), .A2(n4861), .B1(\reg_out[3][17] ), 
        .B2(n4854), .ZN(n2540) );
  OAI221_X2 U491 ( .B1(n4901), .B2(n4473), .C1(n4894), .C2(n3640), .A(n2543), 
        .ZN(n2542) );
  AOI22_X2 U492 ( .A1(\reg_out[21][17] ), .A2(n4888), .B1(\reg_out[23][17] ), 
        .B2(n4881), .ZN(n2543) );
  OAI221_X2 U493 ( .B1(n4874), .B2(n4472), .C1(n4867), .C2(n3852), .A(n2544), 
        .ZN(n2541) );
  AOI22_X2 U494 ( .A1(\reg_out[17][17] ), .A2(n4861), .B1(\reg_out[19][17] ), 
        .B2(n4854), .ZN(n2544) );
  OAI221_X2 U496 ( .B1(n4901), .B2(n4471), .C1(n4894), .C2(n3851), .A(n2547), 
        .ZN(n2546) );
  AOI22_X2 U497 ( .A1(\reg_out[13][17] ), .A2(n4888), .B1(\reg_out[15][17] ), 
        .B2(n4881), .ZN(n2547) );
  OAI221_X2 U498 ( .B1(n4874), .B2(n3893), .C1(n4867), .C2(n4435), .A(n2548), 
        .ZN(n2545) );
  AOI22_X2 U499 ( .A1(\reg_out[9][17] ), .A2(n4861), .B1(\reg_out[11][17] ), 
        .B2(n4854), .ZN(n2548) );
  OAI221_X2 U501 ( .B1(n4900), .B2(n3753), .C1(n4899), .C2(n3850), .A(n2551), 
        .ZN(n2550) );
  AOI22_X2 U502 ( .A1(\reg_out[29][17] ), .A2(n4891), .B1(\reg_out[31][17] ), 
        .B2(n4880), .ZN(n2551) );
  OAI221_X2 U503 ( .B1(n4873), .B2(n3752), .C1(n4872), .C2(n3575), .A(n2552), 
        .ZN(n2549) );
  AOI22_X2 U504 ( .A1(\reg_out[25][17] ), .A2(n4863), .B1(\reg_out[27][17] ), 
        .B2(n4852), .ZN(n2552) );
  NAND4_X2 U505 ( .A1(n2553), .A2(n2554), .A3(n2555), .A4(n2556), .ZN(busB[16]) );
  OAI221_X2 U507 ( .B1(n4900), .B2(n3892), .C1(n4899), .C2(n3639), .A(n2559), 
        .ZN(n2558) );
  AOI22_X2 U508 ( .A1(\reg_out[5][16] ), .A2(n4888), .B1(\reg_out[7][16] ), 
        .B2(n4880), .ZN(n2559) );
  OAI221_X2 U509 ( .B1(n4873), .B2(n3891), .C1(n4872), .C2(n3638), .A(n2560), 
        .ZN(n2557) );
  AOI22_X2 U510 ( .A1(\reg_out[1][16] ), .A2(n4861), .B1(\reg_out[3][16] ), 
        .B2(n4852), .ZN(n2560) );
  OAI221_X2 U512 ( .B1(n4900), .B2(n3751), .C1(n4899), .C2(n3574), .A(n2563), 
        .ZN(n2562) );
  AOI22_X2 U513 ( .A1(\reg_out[21][16] ), .A2(n4888), .B1(\reg_out[23][16] ), 
        .B2(n4880), .ZN(n2563) );
  OAI221_X2 U514 ( .B1(n4873), .B2(n3890), .C1(n4872), .C2(n3573), .A(n2564), 
        .ZN(n2561) );
  AOI22_X2 U515 ( .A1(\reg_out[17][16] ), .A2(n4861), .B1(\reg_out[19][16] ), 
        .B2(n4852), .ZN(n2564) );
  OAI221_X2 U517 ( .B1(n4900), .B2(n3889), .C1(n4899), .C2(n3572), .A(n2567), 
        .ZN(n2566) );
  AOI22_X2 U518 ( .A1(\reg_out[13][16] ), .A2(n4888), .B1(\reg_out[15][16] ), 
        .B2(n4880), .ZN(n2567) );
  OAI221_X2 U519 ( .B1(n4873), .B2(n3888), .C1(n4872), .C2(n3571), .A(n2568), 
        .ZN(n2565) );
  AOI22_X2 U520 ( .A1(\reg_out[9][16] ), .A2(n4861), .B1(\reg_out[11][16] ), 
        .B2(n4852), .ZN(n2568) );
  OAI221_X2 U522 ( .B1(n4900), .B2(n3750), .C1(n4899), .C2(n3849), .A(n2571), 
        .ZN(n2570) );
  AOI22_X2 U523 ( .A1(\reg_out[29][16] ), .A2(n4888), .B1(\reg_out[31][16] ), 
        .B2(n4880), .ZN(n2571) );
  OAI221_X2 U524 ( .B1(n4873), .B2(n3749), .C1(n4872), .C2(n3570), .A(n2572), 
        .ZN(n2569) );
  AOI22_X2 U525 ( .A1(\reg_out[25][16] ), .A2(n4861), .B1(\reg_out[27][16] ), 
        .B2(n4852), .ZN(n2572) );
  NAND4_X2 U526 ( .A1(n2573), .A2(n2574), .A3(n2575), .A4(n2576), .ZN(busB[15]) );
  OAI221_X2 U528 ( .B1(n4900), .B2(n3887), .C1(n4899), .C2(n3637), .A(n2579), 
        .ZN(n2578) );
  AOI22_X2 U529 ( .A1(\reg_out[5][15] ), .A2(n4888), .B1(\reg_out[7][15] ), 
        .B2(n4880), .ZN(n2579) );
  OAI221_X2 U530 ( .B1(n4873), .B2(n3886), .C1(n4872), .C2(n3636), .A(n2580), 
        .ZN(n2577) );
  AOI22_X2 U531 ( .A1(\reg_out[1][15] ), .A2(n4861), .B1(\reg_out[3][15] ), 
        .B2(n4852), .ZN(n2580) );
  OAI221_X2 U533 ( .B1(n4900), .B2(n3748), .C1(n4899), .C2(n3569), .A(n2583), 
        .ZN(n2582) );
  AOI22_X2 U534 ( .A1(\reg_out[21][15] ), .A2(n4890), .B1(\reg_out[23][15] ), 
        .B2(n4880), .ZN(n2583) );
  OAI221_X2 U535 ( .B1(n4873), .B2(n3885), .C1(n4872), .C2(n3568), .A(n2584), 
        .ZN(n2581) );
  AOI22_X2 U536 ( .A1(\reg_out[17][15] ), .A2(n4864), .B1(\reg_out[19][15] ), 
        .B2(n4852), .ZN(n2584) );
  OAI221_X2 U538 ( .B1(n4900), .B2(n3884), .C1(n4899), .C2(n3567), .A(n2587), 
        .ZN(n2586) );
  AOI22_X2 U539 ( .A1(\reg_out[13][15] ), .A2(n4890), .B1(\reg_out[15][15] ), 
        .B2(n4880), .ZN(n2587) );
  OAI221_X2 U540 ( .B1(n4873), .B2(n3883), .C1(n4872), .C2(n3566), .A(n2588), 
        .ZN(n2585) );
  AOI22_X2 U541 ( .A1(\reg_out[9][15] ), .A2(n4864), .B1(\reg_out[11][15] ), 
        .B2(n4852), .ZN(n2588) );
  OAI221_X2 U543 ( .B1(n4900), .B2(n3747), .C1(n4899), .C2(n3848), .A(n2591), 
        .ZN(n2590) );
  AOI22_X2 U544 ( .A1(\reg_out[29][15] ), .A2(n4890), .B1(\reg_out[31][15] ), 
        .B2(n4880), .ZN(n2591) );
  OAI221_X2 U545 ( .B1(n4873), .B2(n3746), .C1(n4872), .C2(n3565), .A(n2592), 
        .ZN(n2589) );
  AOI22_X2 U546 ( .A1(\reg_out[25][15] ), .A2(n4864), .B1(\reg_out[27][15] ), 
        .B2(n4852), .ZN(n2592) );
  NAND4_X2 U547 ( .A1(n2593), .A2(n2594), .A3(n2595), .A4(n2596), .ZN(busB[14]) );
  OAI221_X2 U549 ( .B1(n4900), .B2(n3882), .C1(n4899), .C2(n3635), .A(n2599), 
        .ZN(n2598) );
  AOI22_X2 U550 ( .A1(\reg_out[5][14] ), .A2(n4888), .B1(\reg_out[7][14] ), 
        .B2(n4880), .ZN(n2599) );
  OAI221_X2 U551 ( .B1(n4873), .B2(n3881), .C1(n4872), .C2(n3634), .A(n2600), 
        .ZN(n2597) );
  AOI22_X2 U552 ( .A1(\reg_out[1][14] ), .A2(n4861), .B1(\reg_out[3][14] ), 
        .B2(n4852), .ZN(n2600) );
  OAI221_X2 U554 ( .B1(n4900), .B2(n3745), .C1(n4899), .C2(n3564), .A(n2603), 
        .ZN(n2602) );
  AOI22_X2 U555 ( .A1(\reg_out[21][14] ), .A2(n4891), .B1(\reg_out[23][14] ), 
        .B2(n4880), .ZN(n2603) );
  OAI221_X2 U556 ( .B1(n4873), .B2(n3880), .C1(n4872), .C2(n3563), .A(n2604), 
        .ZN(n2601) );
  AOI22_X2 U557 ( .A1(\reg_out[17][14] ), .A2(n4863), .B1(\reg_out[19][14] ), 
        .B2(n4852), .ZN(n2604) );
  OAI221_X2 U559 ( .B1(n4904), .B2(n4470), .C1(n4897), .C2(n3847), .A(n2607), 
        .ZN(n2606) );
  AOI22_X2 U560 ( .A1(\reg_out[13][14] ), .A2(n4887), .B1(\reg_out[15][14] ), 
        .B2(n4883), .ZN(n2607) );
  OAI221_X2 U561 ( .B1(n4876), .B2(n3879), .C1(n4871), .C2(n4434), .A(n2608), 
        .ZN(n2605) );
  AOI22_X2 U562 ( .A1(\reg_out[9][14] ), .A2(n4865), .B1(\reg_out[11][14] ), 
        .B2(n4857), .ZN(n2608) );
  OAI221_X2 U564 ( .B1(n4904), .B2(n4469), .C1(n4897), .C2(n3846), .A(n2611), 
        .ZN(n2610) );
  AOI22_X2 U565 ( .A1(\reg_out[29][14] ), .A2(n4887), .B1(\reg_out[31][14] ), 
        .B2(n4882), .ZN(n2611) );
  OAI221_X2 U566 ( .B1(n4876), .B2(n4468), .C1(n4871), .C2(n3633), .A(n2612), 
        .ZN(n2609) );
  AOI22_X2 U567 ( .A1(\reg_out[25][14] ), .A2(n4865), .B1(\reg_out[27][14] ), 
        .B2(n4858), .ZN(n2612) );
  NAND4_X2 U568 ( .A1(n2613), .A2(n2614), .A3(n2615), .A4(n2616), .ZN(busB[13]) );
  OAI221_X2 U570 ( .B1(n4904), .B2(n3878), .C1(n4898), .C2(n3632), .A(n2619), 
        .ZN(n2618) );
  AOI22_X2 U571 ( .A1(\reg_out[5][13] ), .A2(n4887), .B1(\reg_out[7][13] ), 
        .B2(n4886), .ZN(n2619) );
  OAI221_X2 U572 ( .B1(n4876), .B2(n4467), .C1(n4871), .C2(n3845), .A(n2620), 
        .ZN(n2617) );
  AOI22_X2 U573 ( .A1(\reg_out[1][13] ), .A2(n4865), .B1(\reg_out[3][13] ), 
        .B2(n4853), .ZN(n2620) );
  OAI221_X2 U575 ( .B1(n4903), .B2(n4466), .C1(n4898), .C2(n3631), .A(n2623), 
        .ZN(n2622) );
  AOI22_X2 U576 ( .A1(\reg_out[21][13] ), .A2(n4887), .B1(\reg_out[23][13] ), 
        .B2(n4886), .ZN(n2623) );
  OAI221_X2 U577 ( .B1(n4877), .B2(n4465), .C1(n4871), .C2(n3844), .A(n2624), 
        .ZN(n2621) );
  AOI22_X2 U578 ( .A1(\reg_out[17][13] ), .A2(n4865), .B1(\reg_out[19][13] ), 
        .B2(n4858), .ZN(n2624) );
  OAI221_X2 U580 ( .B1(n4903), .B2(n4464), .C1(n4895), .C2(n3843), .A(n2627), 
        .ZN(n2626) );
  AOI22_X2 U581 ( .A1(\reg_out[13][13] ), .A2(n4888), .B1(\reg_out[15][13] ), 
        .B2(n4886), .ZN(n2627) );
  OAI221_X2 U582 ( .B1(n4877), .B2(n3877), .C1(n4868), .C2(n4433), .A(n2628), 
        .ZN(n2625) );
  AOI22_X2 U583 ( .A1(\reg_out[9][13] ), .A2(n4865), .B1(\reg_out[11][13] ), 
        .B2(n4856), .ZN(n2628) );
  OAI221_X2 U585 ( .B1(n4903), .B2(n4463), .C1(n4896), .C2(n3842), .A(n2631), 
        .ZN(n2630) );
  AOI22_X2 U586 ( .A1(\reg_out[29][13] ), .A2(n4887), .B1(\reg_out[31][13] ), 
        .B2(n4885), .ZN(n2631) );
  OAI221_X2 U587 ( .B1(n4877), .B2(n4462), .C1(n4868), .C2(n3630), .A(n2632), 
        .ZN(n2629) );
  AOI22_X2 U588 ( .A1(\reg_out[25][13] ), .A2(n4865), .B1(\reg_out[27][13] ), 
        .B2(n4858), .ZN(n2632) );
  NAND4_X2 U589 ( .A1(n2633), .A2(n2634), .A3(n2635), .A4(n2636), .ZN(busB[12]) );
  OAI221_X2 U591 ( .B1(n4903), .B2(n3876), .C1(n4898), .C2(n3629), .A(n2639), 
        .ZN(n2638) );
  AOI22_X2 U592 ( .A1(\reg_out[5][12] ), .A2(n4887), .B1(\reg_out[7][12] ), 
        .B2(n4885), .ZN(n2639) );
  OAI221_X2 U593 ( .B1(n4877), .B2(n4461), .C1(n4871), .C2(n3841), .A(n2640), 
        .ZN(n2637) );
  AOI22_X2 U594 ( .A1(\reg_out[1][12] ), .A2(n4865), .B1(\reg_out[3][12] ), 
        .B2(n4853), .ZN(n2640) );
  OAI221_X2 U596 ( .B1(n4906), .B2(n4460), .C1(n4898), .C2(n3628), .A(n2643), 
        .ZN(n2642) );
  AOI22_X2 U597 ( .A1(\reg_out[21][12] ), .A2(n4887), .B1(\reg_out[23][12] ), 
        .B2(n4885), .ZN(n2643) );
  OAI221_X2 U598 ( .B1(n4879), .B2(n4459), .C1(n4871), .C2(n3840), .A(n2644), 
        .ZN(n2641) );
  AOI22_X2 U599 ( .A1(\reg_out[17][12] ), .A2(n4865), .B1(\reg_out[19][12] ), 
        .B2(n4855), .ZN(n2644) );
  OAI221_X2 U601 ( .B1(n4906), .B2(n4458), .C1(n4898), .C2(n3839), .A(n2647), 
        .ZN(n2646) );
  AOI22_X2 U602 ( .A1(\reg_out[13][12] ), .A2(n4887), .B1(\reg_out[15][12] ), 
        .B2(n4881), .ZN(n2647) );
  OAI221_X2 U603 ( .B1(n4879), .B2(n3875), .C1(n4869), .C2(n4432), .A(n2648), 
        .ZN(n2645) );
  AOI22_X2 U604 ( .A1(\reg_out[9][12] ), .A2(n4865), .B1(\reg_out[11][12] ), 
        .B2(n4853), .ZN(n2648) );
  OAI221_X2 U606 ( .B1(n4906), .B2(n4457), .C1(n4893), .C2(n3838), .A(n2651), 
        .ZN(n2650) );
  AOI22_X2 U607 ( .A1(\reg_out[29][12] ), .A2(n4888), .B1(\reg_out[31][12] ), 
        .B2(n4886), .ZN(n2651) );
  OAI221_X2 U608 ( .B1(n4879), .B2(n4456), .C1(n4869), .C2(n3627), .A(n2652), 
        .ZN(n2649) );
  AOI22_X2 U609 ( .A1(\reg_out[25][12] ), .A2(n4860), .B1(\reg_out[27][12] ), 
        .B2(n4855), .ZN(n2652) );
  NAND4_X2 U610 ( .A1(n2653), .A2(n2654), .A3(n2655), .A4(n2656), .ZN(busB[11]) );
  OAI221_X2 U612 ( .B1(n4904), .B2(n3874), .C1(n4898), .C2(n3626), .A(n2659), 
        .ZN(n2658) );
  AOI22_X2 U613 ( .A1(\reg_out[5][11] ), .A2(n4887), .B1(\reg_out[7][11] ), 
        .B2(n4881), .ZN(n2659) );
  OAI221_X2 U614 ( .B1(n4876), .B2(n4455), .C1(n4871), .C2(n3837), .A(n2660), 
        .ZN(n2657) );
  AOI22_X2 U615 ( .A1(\reg_out[1][11] ), .A2(n4865), .B1(\reg_out[3][11] ), 
        .B2(n4853), .ZN(n2660) );
  OAI221_X2 U617 ( .B1(n4906), .B2(n4454), .C1(n4893), .C2(n3625), .A(n2663), 
        .ZN(n2662) );
  AOI22_X2 U618 ( .A1(\reg_out[21][11] ), .A2(n4887), .B1(\reg_out[23][11] ), 
        .B2(n4880), .ZN(n2663) );
  OAI221_X2 U619 ( .B1(n4879), .B2(n4453), .C1(n4866), .C2(n3836), .A(n2664), 
        .ZN(n2661) );
  AOI22_X2 U620 ( .A1(\reg_out[17][11] ), .A2(n4860), .B1(\reg_out[19][11] ), 
        .B2(n4852), .ZN(n2664) );
  OAI221_X2 U622 ( .B1(n4904), .B2(n4452), .C1(n4893), .C2(n3835), .A(n2667), 
        .ZN(n2666) );
  AOI22_X2 U623 ( .A1(\reg_out[13][11] ), .A2(n4887), .B1(\reg_out[15][11] ), 
        .B2(n4880), .ZN(n2667) );
  OAI221_X2 U624 ( .B1(n4876), .B2(n3873), .C1(n4866), .C2(n4431), .A(n2668), 
        .ZN(n2665) );
  AOI22_X2 U625 ( .A1(\reg_out[9][11] ), .A2(n4860), .B1(\reg_out[11][11] ), 
        .B2(n4852), .ZN(n2668) );
  OAI221_X2 U627 ( .B1(n4904), .B2(n4451), .C1(n4893), .C2(n3834), .A(n2671), 
        .ZN(n2670) );
  AOI22_X2 U628 ( .A1(\reg_out[29][11] ), .A2(n4887), .B1(\reg_out[31][11] ), 
        .B2(n4884), .ZN(n2671) );
  OAI221_X2 U629 ( .B1(n4876), .B2(n4450), .C1(n4866), .C2(n3624), .A(n2672), 
        .ZN(n2669) );
  AOI22_X2 U630 ( .A1(\reg_out[25][11] ), .A2(n4860), .B1(\reg_out[27][11] ), 
        .B2(n4856), .ZN(n2672) );
  NAND4_X2 U631 ( .A1(n2673), .A2(n2674), .A3(n2675), .A4(n2676), .ZN(busB[10]) );
  OAI221_X2 U633 ( .B1(n4906), .B2(n3872), .C1(n4893), .C2(n3623), .A(n2679), 
        .ZN(n2678) );
  AOI22_X2 U634 ( .A1(\reg_out[5][10] ), .A2(n4887), .B1(\reg_out[7][10] ), 
        .B2(n4880), .ZN(n2679) );
  OAI221_X2 U635 ( .B1(n4879), .B2(n4449), .C1(n4866), .C2(n3833), .A(n2680), 
        .ZN(n2677) );
  AOI22_X2 U636 ( .A1(\reg_out[1][10] ), .A2(n4860), .B1(\reg_out[3][10] ), 
        .B2(n4852), .ZN(n2680) );
  OAI221_X2 U638 ( .B1(n4904), .B2(n4448), .C1(n4893), .C2(n3622), .A(n2683), 
        .ZN(n2682) );
  AOI22_X2 U639 ( .A1(\reg_out[21][10] ), .A2(n4887), .B1(\reg_out[23][10] ), 
        .B2(n4880), .ZN(n2683) );
  OAI221_X2 U640 ( .B1(n4876), .B2(n4447), .C1(n4866), .C2(n3832), .A(n2684), 
        .ZN(n2681) );
  AOI22_X2 U641 ( .A1(\reg_out[17][10] ), .A2(n4860), .B1(\reg_out[19][10] ), 
        .B2(n4852), .ZN(n2684) );
  OAI221_X2 U643 ( .B1(n4906), .B2(n4446), .C1(n4893), .C2(n3831), .A(n2687), 
        .ZN(n2686) );
  AOI22_X2 U644 ( .A1(\reg_out[13][10] ), .A2(n4887), .B1(\reg_out[15][10] ), 
        .B2(n4880), .ZN(n2687) );
  OAI221_X2 U645 ( .B1(n4879), .B2(n3871), .C1(n4866), .C2(n4430), .A(n2688), 
        .ZN(n2685) );
  AOI22_X2 U646 ( .A1(\reg_out[9][10] ), .A2(n4860), .B1(\reg_out[11][10] ), 
        .B2(n4857), .ZN(n2688) );
  OAI221_X2 U648 ( .B1(n4906), .B2(n4445), .C1(n4893), .C2(n3830), .A(n2691), 
        .ZN(n2690) );
  AOI22_X2 U649 ( .A1(\reg_out[29][10] ), .A2(n4887), .B1(\reg_out[31][10] ), 
        .B2(n4881), .ZN(n2691) );
  OAI221_X2 U650 ( .B1(n4879), .B2(n4444), .C1(n4866), .C2(n3621), .A(n2692), 
        .ZN(n2689) );
  AOI22_X2 U651 ( .A1(\reg_out[25][10] ), .A2(n4860), .B1(\reg_out[27][10] ), 
        .B2(n4852), .ZN(n2692) );
  NAND4_X2 U652 ( .A1(n2693), .A2(n2694), .A3(n2695), .A4(n2696), .ZN(busB[0])
         );
  OAI221_X2 U655 ( .B1(n4906), .B2(n3870), .C1(n4893), .C2(n3620), .A(n2699), 
        .ZN(n2698) );
  AOI22_X2 U656 ( .A1(\reg_out[5][0] ), .A2(n4887), .B1(\reg_out[7][0] ), .B2(
        n4880), .ZN(n2699) );
  OAI221_X2 U657 ( .B1(n4879), .B2(n4443), .C1(n4866), .C2(n3829), .A(n2700), 
        .ZN(n2697) );
  AOI22_X2 U658 ( .A1(\reg_out[1][0] ), .A2(n4860), .B1(\reg_out[3][0] ), .B2(
        n4852), .ZN(n2700) );
  OAI221_X2 U661 ( .B1(n4906), .B2(n4442), .C1(n4893), .C2(n3619), .A(n2703), 
        .ZN(n2702) );
  AOI22_X2 U662 ( .A1(\reg_out[21][0] ), .A2(n4887), .B1(\reg_out[23][0] ), 
        .B2(n4880), .ZN(n2703) );
  OAI221_X2 U663 ( .B1(n4879), .B2(n4441), .C1(n4866), .C2(n3828), .A(n2704), 
        .ZN(n2701) );
  AOI22_X2 U664 ( .A1(\reg_out[17][0] ), .A2(n4860), .B1(\reg_out[19][0] ), 
        .B2(n4852), .ZN(n2704) );
  OAI221_X2 U667 ( .B1(n4903), .B2(n4440), .C1(n4893), .C2(n3827), .A(n2707), 
        .ZN(n2706) );
  AOI22_X2 U668 ( .A1(\reg_out[13][0] ), .A2(n4887), .B1(\reg_out[15][0] ), 
        .B2(n4880), .ZN(n2707) );
  OAI221_X2 U669 ( .B1(n4877), .B2(n3869), .C1(n4866), .C2(n4429), .A(n2708), 
        .ZN(n2705) );
  AOI22_X2 U670 ( .A1(\reg_out[9][0] ), .A2(n4860), .B1(\reg_out[11][0] ), 
        .B2(n4852), .ZN(n2708) );
  OAI221_X2 U673 ( .B1(n4903), .B2(n4439), .C1(n4893), .C2(n3826), .A(n2711), 
        .ZN(n2710) );
  AOI22_X2 U674 ( .A1(\reg_out[29][0] ), .A2(n4889), .B1(\reg_out[31][0] ), 
        .B2(n4883), .ZN(n2711) );
  OAI221_X2 U679 ( .B1(n4877), .B2(n4438), .C1(n4866), .C2(n3618), .A(n2716), 
        .ZN(n2709) );
  AOI22_X2 U680 ( .A1(\reg_out[25][0] ), .A2(n4860), .B1(\reg_out[27][0] ), 
        .B2(n4853), .ZN(n2716) );
  AND2_X2 U682 ( .A1(rb[4]), .A2(rb[3]), .ZN(n2712) );
  AND2_X2 U684 ( .A1(rb[4]), .A2(n1035), .ZN(n2713) );
  NAND4_X2 U689 ( .A1(n2717), .A2(n2718), .A3(n2719), .A4(n2720), .ZN(busA[9])
         );
  OAI221_X2 U691 ( .B1(n3778), .B2(n4837), .C1(n3595), .C2(n4835), .A(n2726), 
        .ZN(n2722) );
  AOI22_X2 U692 ( .A1(n4829), .A2(\reg_out[5][9] ), .B1(n4815), .B2(
        \reg_out[7][9] ), .ZN(n2726) );
  OAI221_X2 U693 ( .B1(n3777), .B2(n4808), .C1(n3594), .C2(n4806), .A(n2731), 
        .ZN(n2721) );
  AOI22_X2 U694 ( .A1(n4800), .A2(\reg_out[1][9] ), .B1(n4786), .B2(
        \reg_out[3][9] ), .ZN(n2731) );
  OAI221_X2 U696 ( .B1(n3776), .B2(n4837), .C1(n3593), .C2(n4835), .A(n2737), 
        .ZN(n2735) );
  AOI22_X2 U697 ( .A1(n4829), .A2(\reg_out[21][9] ), .B1(n4815), .B2(
        \reg_out[23][9] ), .ZN(n2737) );
  OAI221_X2 U698 ( .B1(n3775), .B2(n4808), .C1(n3592), .C2(n4806), .A(n2738), 
        .ZN(n2734) );
  AOI22_X2 U699 ( .A1(n4800), .A2(\reg_out[17][9] ), .B1(n4786), .B2(
        \reg_out[19][9] ), .ZN(n2738) );
  OAI221_X2 U701 ( .B1(n3774), .B2(n4837), .C1(n3591), .C2(n4835), .A(n2742), 
        .ZN(n2740) );
  AOI22_X2 U702 ( .A1(n4829), .A2(\reg_out[13][9] ), .B1(n4815), .B2(
        \reg_out[15][9] ), .ZN(n2742) );
  OAI221_X2 U703 ( .B1(n3773), .B2(n4808), .C1(n3590), .C2(n4806), .A(n2743), 
        .ZN(n2739) );
  AOI22_X2 U704 ( .A1(n4800), .A2(\reg_out[9][9] ), .B1(n4786), .B2(
        \reg_out[11][9] ), .ZN(n2743) );
  OAI221_X2 U706 ( .B1(n3772), .B2(n4842), .C1(n3589), .C2(n4835), .A(n2747), 
        .ZN(n2745) );
  AOI22_X2 U707 ( .A1(n4826), .A2(\reg_out[29][9] ), .B1(n4820), .B2(
        \reg_out[31][9] ), .ZN(n2747) );
  OAI221_X2 U708 ( .B1(n3771), .B2(n4813), .C1(n3588), .C2(n4806), .A(n2748), 
        .ZN(n2744) );
  AOI22_X2 U709 ( .A1(n4797), .A2(\reg_out[25][9] ), .B1(n4791), .B2(
        \reg_out[27][9] ), .ZN(n2748) );
  NAND4_X2 U710 ( .A1(n2749), .A2(n2750), .A3(n2751), .A4(n2752), .ZN(busA[8])
         );
  OAI221_X2 U712 ( .B1(n3770), .B2(n4837), .C1(n3587), .C2(n4836), .A(n2755), 
        .ZN(n2754) );
  AOI22_X2 U713 ( .A1(n4828), .A2(\reg_out[5][8] ), .B1(n4815), .B2(
        \reg_out[7][8] ), .ZN(n2755) );
  OAI221_X2 U714 ( .B1(n3769), .B2(n4808), .C1(n3586), .C2(n4807), .A(n2756), 
        .ZN(n2753) );
  AOI22_X2 U715 ( .A1(n4799), .A2(\reg_out[1][8] ), .B1(n4786), .B2(
        \reg_out[3][8] ), .ZN(n2756) );
  OAI221_X2 U717 ( .B1(n3768), .B2(n4837), .C1(n3585), .C2(n4836), .A(n2759), 
        .ZN(n2758) );
  AOI22_X2 U718 ( .A1(n4828), .A2(\reg_out[21][8] ), .B1(n4815), .B2(
        \reg_out[23][8] ), .ZN(n2759) );
  OAI221_X2 U719 ( .B1(n3767), .B2(n4808), .C1(n3584), .C2(n4807), .A(n2760), 
        .ZN(n2757) );
  AOI22_X2 U720 ( .A1(n4799), .A2(\reg_out[17][8] ), .B1(n4786), .B2(
        \reg_out[19][8] ), .ZN(n2760) );
  OAI221_X2 U722 ( .B1(n3766), .B2(n4837), .C1(n3583), .C2(n4836), .A(n2763), 
        .ZN(n2762) );
  AOI22_X2 U723 ( .A1(n4826), .A2(\reg_out[13][8] ), .B1(n4815), .B2(
        \reg_out[15][8] ), .ZN(n2763) );
  OAI221_X2 U724 ( .B1(n3765), .B2(n4808), .C1(n3582), .C2(n4807), .A(n2764), 
        .ZN(n2761) );
  AOI22_X2 U725 ( .A1(n4797), .A2(\reg_out[9][8] ), .B1(n4786), .B2(
        \reg_out[11][8] ), .ZN(n2764) );
  OAI221_X2 U727 ( .B1(n4019), .B2(n4843), .C1(n3744), .C2(n4836), .A(n2767), 
        .ZN(n2766) );
  AOI22_X2 U728 ( .A1(n4829), .A2(\reg_out[29][8] ), .B1(n4821), .B2(
        \reg_out[31][8] ), .ZN(n2767) );
  OAI221_X2 U729 ( .B1(n4018), .B2(n4814), .C1(n3743), .C2(n4807), .A(n2768), 
        .ZN(n2765) );
  AOI22_X2 U730 ( .A1(n4800), .A2(\reg_out[25][8] ), .B1(n4792), .B2(
        \reg_out[27][8] ), .ZN(n2768) );
  NAND4_X2 U731 ( .A1(n2769), .A2(n2770), .A3(n2771), .A4(n2772), .ZN(busA[7])
         );
  OAI221_X2 U733 ( .B1(n3764), .B2(n4843), .C1(n3581), .C2(n4836), .A(n2775), 
        .ZN(n2774) );
  AOI22_X2 U734 ( .A1(n4829), .A2(\reg_out[5][7] ), .B1(n4821), .B2(
        \reg_out[7][7] ), .ZN(n2775) );
  OAI221_X2 U735 ( .B1(n4017), .B2(n4814), .C1(n3742), .C2(n4807), .A(n2776), 
        .ZN(n2773) );
  AOI22_X2 U736 ( .A1(n4800), .A2(\reg_out[1][7] ), .B1(n4792), .B2(
        \reg_out[3][7] ), .ZN(n2776) );
  OAI221_X2 U738 ( .B1(n4016), .B2(n4843), .C1(n3741), .C2(n4836), .A(n2779), 
        .ZN(n2778) );
  AOI22_X2 U739 ( .A1(n4829), .A2(\reg_out[21][7] ), .B1(n4821), .B2(
        \reg_out[23][7] ), .ZN(n2779) );
  OAI221_X2 U740 ( .B1(n4015), .B2(n4814), .C1(n3740), .C2(n4807), .A(n2780), 
        .ZN(n2777) );
  AOI22_X2 U741 ( .A1(n4800), .A2(\reg_out[17][7] ), .B1(n4792), .B2(
        \reg_out[19][7] ), .ZN(n2780) );
  OAI221_X2 U743 ( .B1(n4014), .B2(n4843), .C1(n3739), .C2(n4836), .A(n2783), 
        .ZN(n2782) );
  AOI22_X2 U744 ( .A1(n4829), .A2(\reg_out[13][7] ), .B1(n4821), .B2(
        \reg_out[15][7] ), .ZN(n2783) );
  OAI221_X2 U745 ( .B1(n3763), .B2(n4814), .C1(n3868), .C2(n4807), .A(n2784), 
        .ZN(n2781) );
  AOI22_X2 U746 ( .A1(n4800), .A2(\reg_out[9][7] ), .B1(n4792), .B2(
        \reg_out[11][7] ), .ZN(n2784) );
  OAI221_X2 U748 ( .B1(n4013), .B2(n4843), .C1(n3738), .C2(n4836), .A(n2787), 
        .ZN(n2786) );
  AOI22_X2 U749 ( .A1(n4829), .A2(\reg_out[29][7] ), .B1(n4821), .B2(
        \reg_out[31][7] ), .ZN(n2787) );
  OAI221_X2 U750 ( .B1(n4012), .B2(n4814), .C1(n3737), .C2(n4807), .A(n2788), 
        .ZN(n2785) );
  AOI22_X2 U751 ( .A1(n4800), .A2(\reg_out[25][7] ), .B1(n4792), .B2(
        \reg_out[27][7] ), .ZN(n2788) );
  NAND4_X2 U752 ( .A1(n2789), .A2(n2790), .A3(n2791), .A4(n2792), .ZN(busA[6])
         );
  OAI221_X2 U754 ( .B1(n3762), .B2(n4843), .C1(n3580), .C2(n4836), .A(n2795), 
        .ZN(n2794) );
  AOI22_X2 U755 ( .A1(n4829), .A2(\reg_out[5][6] ), .B1(n4821), .B2(
        \reg_out[7][6] ), .ZN(n2795) );
  OAI221_X2 U756 ( .B1(n4011), .B2(n4814), .C1(n3736), .C2(n4807), .A(n2796), 
        .ZN(n2793) );
  AOI22_X2 U757 ( .A1(n4800), .A2(\reg_out[1][6] ), .B1(n4792), .B2(
        \reg_out[3][6] ), .ZN(n2796) );
  OAI221_X2 U759 ( .B1(n4010), .B2(n4843), .C1(n3735), .C2(n4836), .A(n2799), 
        .ZN(n2798) );
  AOI22_X2 U760 ( .A1(n4829), .A2(\reg_out[21][6] ), .B1(n4821), .B2(
        \reg_out[23][6] ), .ZN(n2799) );
  OAI221_X2 U761 ( .B1(n4009), .B2(n4814), .C1(n3734), .C2(n4807), .A(n2800), 
        .ZN(n2797) );
  AOI22_X2 U762 ( .A1(n4800), .A2(\reg_out[17][6] ), .B1(n4792), .B2(
        \reg_out[19][6] ), .ZN(n2800) );
  OAI221_X2 U764 ( .B1(n4008), .B2(n4843), .C1(n3733), .C2(n4836), .A(n2803), 
        .ZN(n2802) );
  AOI22_X2 U765 ( .A1(n4829), .A2(\reg_out[13][6] ), .B1(n4821), .B2(
        \reg_out[15][6] ), .ZN(n2803) );
  OAI221_X2 U766 ( .B1(n3761), .B2(n4814), .C1(n3867), .C2(n4807), .A(n2804), 
        .ZN(n2801) );
  AOI22_X2 U767 ( .A1(n4800), .A2(\reg_out[9][6] ), .B1(n4792), .B2(
        \reg_out[11][6] ), .ZN(n2804) );
  OAI221_X2 U769 ( .B1(n4007), .B2(n4843), .C1(n3732), .C2(n4836), .A(n2807), 
        .ZN(n2806) );
  AOI22_X2 U770 ( .A1(n4829), .A2(\reg_out[29][6] ), .B1(n4821), .B2(
        \reg_out[31][6] ), .ZN(n2807) );
  OAI221_X2 U771 ( .B1(n4006), .B2(n4814), .C1(n3731), .C2(n4807), .A(n2808), 
        .ZN(n2805) );
  AOI22_X2 U772 ( .A1(n4800), .A2(\reg_out[25][6] ), .B1(n4792), .B2(
        \reg_out[27][6] ), .ZN(n2808) );
  NAND4_X2 U773 ( .A1(n2809), .A2(n2810), .A3(n2811), .A4(n2812), .ZN(busA[5])
         );
  OAI221_X2 U775 ( .B1(n3760), .B2(n4843), .C1(n3579), .C2(n4836), .A(n2815), 
        .ZN(n2814) );
  AOI22_X2 U776 ( .A1(n4829), .A2(\reg_out[5][5] ), .B1(n4821), .B2(
        \reg_out[7][5] ), .ZN(n2815) );
  OAI221_X2 U777 ( .B1(n4005), .B2(n4814), .C1(n3730), .C2(n4807), .A(n2816), 
        .ZN(n2813) );
  AOI22_X2 U778 ( .A1(n4800), .A2(\reg_out[1][5] ), .B1(n4792), .B2(
        \reg_out[3][5] ), .ZN(n2816) );
  OAI221_X2 U780 ( .B1(n4004), .B2(n4843), .C1(n3729), .C2(n4836), .A(n2819), 
        .ZN(n2818) );
  AOI22_X2 U781 ( .A1(n4829), .A2(\reg_out[21][5] ), .B1(n4821), .B2(
        \reg_out[23][5] ), .ZN(n2819) );
  OAI221_X2 U782 ( .B1(n4003), .B2(n4814), .C1(n3728), .C2(n4807), .A(n2820), 
        .ZN(n2817) );
  AOI22_X2 U783 ( .A1(n4800), .A2(\reg_out[17][5] ), .B1(n4792), .B2(
        \reg_out[19][5] ), .ZN(n2820) );
  OAI221_X2 U785 ( .B1(n4002), .B2(n4842), .C1(n3727), .C2(n4835), .A(n2823), 
        .ZN(n2822) );
  AOI22_X2 U786 ( .A1(n4828), .A2(\reg_out[13][5] ), .B1(n4820), .B2(
        \reg_out[15][5] ), .ZN(n2823) );
  OAI221_X2 U787 ( .B1(n3759), .B2(n4813), .C1(n3866), .C2(n4806), .A(n2824), 
        .ZN(n2821) );
  AOI22_X2 U788 ( .A1(n4799), .A2(\reg_out[9][5] ), .B1(n4791), .B2(
        \reg_out[11][5] ), .ZN(n2824) );
  OAI221_X2 U790 ( .B1(n4001), .B2(n4842), .C1(n3726), .C2(n4835), .A(n2827), 
        .ZN(n2826) );
  AOI22_X2 U791 ( .A1(n4828), .A2(\reg_out[29][5] ), .B1(n4820), .B2(
        \reg_out[31][5] ), .ZN(n2827) );
  OAI221_X2 U792 ( .B1(n4000), .B2(n4813), .C1(n3725), .C2(n4806), .A(n2828), 
        .ZN(n2825) );
  AOI22_X2 U793 ( .A1(n4799), .A2(\reg_out[25][5] ), .B1(n4791), .B2(
        \reg_out[27][5] ), .ZN(n2828) );
  NAND4_X2 U794 ( .A1(n2829), .A2(n2830), .A3(n2831), .A4(n2832), .ZN(busA[4])
         );
  OAI221_X2 U796 ( .B1(n3758), .B2(n4842), .C1(n3578), .C2(n4835), .A(n2835), 
        .ZN(n2834) );
  AOI22_X2 U797 ( .A1(n4828), .A2(\reg_out[5][4] ), .B1(n4820), .B2(
        \reg_out[7][4] ), .ZN(n2835) );
  OAI221_X2 U798 ( .B1(n3999), .B2(n4813), .C1(n3724), .C2(n4806), .A(n2836), 
        .ZN(n2833) );
  AOI22_X2 U799 ( .A1(n4799), .A2(\reg_out[1][4] ), .B1(n4791), .B2(
        \reg_out[3][4] ), .ZN(n2836) );
  OAI221_X2 U801 ( .B1(n3998), .B2(n4842), .C1(n3723), .C2(n4835), .A(n2839), 
        .ZN(n2838) );
  AOI22_X2 U802 ( .A1(n4828), .A2(\reg_out[21][4] ), .B1(n4820), .B2(
        \reg_out[23][4] ), .ZN(n2839) );
  OAI221_X2 U803 ( .B1(n3997), .B2(n4813), .C1(n3722), .C2(n4806), .A(n2840), 
        .ZN(n2837) );
  AOI22_X2 U804 ( .A1(n4799), .A2(\reg_out[17][4] ), .B1(n4791), .B2(
        \reg_out[19][4] ), .ZN(n2840) );
  OAI221_X2 U806 ( .B1(n3996), .B2(n4842), .C1(n3721), .C2(n4835), .A(n2843), 
        .ZN(n2842) );
  AOI22_X2 U807 ( .A1(n4828), .A2(\reg_out[13][4] ), .B1(n4820), .B2(
        \reg_out[15][4] ), .ZN(n2843) );
  OAI221_X2 U808 ( .B1(n3757), .B2(n4813), .C1(n3865), .C2(n4806), .A(n2844), 
        .ZN(n2841) );
  AOI22_X2 U809 ( .A1(n4799), .A2(\reg_out[9][4] ), .B1(n4791), .B2(
        \reg_out[11][4] ), .ZN(n2844) );
  OAI221_X2 U811 ( .B1(n3995), .B2(n4842), .C1(n3720), .C2(n4835), .A(n2847), 
        .ZN(n2846) );
  AOI22_X2 U812 ( .A1(n4828), .A2(\reg_out[29][4] ), .B1(n4820), .B2(
        \reg_out[31][4] ), .ZN(n2847) );
  OAI221_X2 U813 ( .B1(n3994), .B2(n4813), .C1(n3719), .C2(n4806), .A(n2848), 
        .ZN(n2845) );
  AOI22_X2 U814 ( .A1(n4799), .A2(\reg_out[25][4] ), .B1(n4791), .B2(
        \reg_out[27][4] ), .ZN(n2848) );
  NAND4_X2 U815 ( .A1(n2849), .A2(n2850), .A3(n2851), .A4(n2852), .ZN(busA[3])
         );
  OAI221_X2 U817 ( .B1(n3756), .B2(n4842), .C1(n3577), .C2(n4835), .A(n2855), 
        .ZN(n2854) );
  AOI22_X2 U818 ( .A1(n4828), .A2(\reg_out[5][3] ), .B1(n4820), .B2(
        \reg_out[7][3] ), .ZN(n2855) );
  OAI221_X2 U819 ( .B1(n3993), .B2(n4813), .C1(n3718), .C2(n4806), .A(n2856), 
        .ZN(n2853) );
  AOI22_X2 U820 ( .A1(n4799), .A2(\reg_out[1][3] ), .B1(n4791), .B2(
        \reg_out[3][3] ), .ZN(n2856) );
  OAI221_X2 U822 ( .B1(n3992), .B2(n4842), .C1(n3717), .C2(n4835), .A(n2859), 
        .ZN(n2858) );
  AOI22_X2 U823 ( .A1(n4828), .A2(\reg_out[21][3] ), .B1(n4820), .B2(
        \reg_out[23][3] ), .ZN(n2859) );
  OAI221_X2 U824 ( .B1(n3991), .B2(n4813), .C1(n3716), .C2(n4806), .A(n2860), 
        .ZN(n2857) );
  AOI22_X2 U825 ( .A1(n4799), .A2(\reg_out[17][3] ), .B1(n4791), .B2(
        \reg_out[19][3] ), .ZN(n2860) );
  OAI221_X2 U827 ( .B1(n3990), .B2(n4842), .C1(n3715), .C2(n4835), .A(n2863), 
        .ZN(n2862) );
  AOI22_X2 U828 ( .A1(n4828), .A2(\reg_out[13][3] ), .B1(n4820), .B2(
        \reg_out[15][3] ), .ZN(n2863) );
  OAI221_X2 U829 ( .B1(n3755), .B2(n4813), .C1(n3864), .C2(n4806), .A(n2864), 
        .ZN(n2861) );
  AOI22_X2 U830 ( .A1(n4799), .A2(\reg_out[9][3] ), .B1(n4791), .B2(
        \reg_out[11][3] ), .ZN(n2864) );
  OAI221_X2 U832 ( .B1(n3989), .B2(n4842), .C1(n3714), .C2(n4835), .A(n2867), 
        .ZN(n2866) );
  AOI22_X2 U833 ( .A1(n4828), .A2(\reg_out[29][3] ), .B1(n4820), .B2(
        \reg_out[31][3] ), .ZN(n2867) );
  OAI221_X2 U834 ( .B1(n3988), .B2(n4813), .C1(n3713), .C2(n4806), .A(n2868), 
        .ZN(n2865) );
  AOI22_X2 U835 ( .A1(n4799), .A2(\reg_out[25][3] ), .B1(n4791), .B2(
        \reg_out[27][3] ), .ZN(n2868) );
  NAND4_X2 U836 ( .A1(n2869), .A2(n2870), .A3(n2871), .A4(n2872), .ZN(busA[31]) );
  OAI221_X2 U838 ( .B1(n3754), .B2(n4842), .C1(n3576), .C2(n4835), .A(n2875), 
        .ZN(n2874) );
  AOI22_X2 U839 ( .A1(n4828), .A2(\reg_out[5][31] ), .B1(n4820), .B2(
        \reg_out[7][31] ), .ZN(n2875) );
  OAI221_X2 U840 ( .B1(n3987), .B2(n4813), .C1(n3712), .C2(n4806), .A(n2876), 
        .ZN(n2873) );
  AOI22_X2 U841 ( .A1(n4799), .A2(\reg_out[1][31] ), .B1(n4791), .B2(
        \reg_out[3][31] ), .ZN(n2876) );
  OAI221_X2 U843 ( .B1(n3617), .B2(n4840), .C1(n3540), .C2(n4833), .A(n2879), 
        .ZN(n2878) );
  AOI22_X2 U844 ( .A1(n4824), .A2(\reg_out[21][31] ), .B1(n4818), .B2(
        \reg_out[23][31] ), .ZN(n2879) );
  OAI221_X2 U845 ( .B1(n3616), .B2(n4811), .C1(n3539), .C2(n4805), .A(n2880), 
        .ZN(n2877) );
  AOI22_X2 U846 ( .A1(n4795), .A2(\reg_out[17][31] ), .B1(n4789), .B2(
        \reg_out[19][31] ), .ZN(n2880) );
  OAI221_X2 U848 ( .B1(n3615), .B2(n4841), .C1(n3538), .C2(n4834), .A(n2883), 
        .ZN(n2882) );
  AOI22_X2 U849 ( .A1(n4827), .A2(\reg_out[13][31] ), .B1(n4819), .B2(
        \reg_out[15][31] ), .ZN(n2883) );
  OAI221_X2 U850 ( .B1(n3614), .B2(n4812), .C1(n3537), .C2(n4804), .A(n2884), 
        .ZN(n2881) );
  AOI22_X2 U851 ( .A1(n4798), .A2(\reg_out[9][31] ), .B1(n4790), .B2(
        \reg_out[11][31] ), .ZN(n2884) );
  OAI221_X2 U853 ( .B1(n3613), .B2(n4840), .C1(n3536), .C2(n4833), .A(n2887), 
        .ZN(n2886) );
  AOI22_X2 U854 ( .A1(n4825), .A2(\reg_out[29][31] ), .B1(n4818), .B2(
        \reg_out[31][31] ), .ZN(n2887) );
  OAI221_X2 U855 ( .B1(n3612), .B2(n4811), .C1(n3535), .C2(n4805), .A(n2888), 
        .ZN(n2885) );
  AOI22_X2 U856 ( .A1(n4796), .A2(\reg_out[25][31] ), .B1(n4789), .B2(
        \reg_out[27][31] ), .ZN(n2888) );
  NAND4_X2 U857 ( .A1(n2889), .A2(n2890), .A3(n2891), .A4(n2892), .ZN(busA[30]) );
  OAI221_X2 U859 ( .B1(n3611), .B2(n4840), .C1(n3534), .C2(n4833), .A(n2895), 
        .ZN(n2894) );
  AOI22_X2 U860 ( .A1(n4826), .A2(\reg_out[5][30] ), .B1(n4818), .B2(
        \reg_out[7][30] ), .ZN(n2895) );
  OAI221_X2 U861 ( .B1(n3610), .B2(n4811), .C1(n3533), .C2(n4805), .A(n2896), 
        .ZN(n2893) );
  AOI22_X2 U862 ( .A1(n4797), .A2(\reg_out[1][30] ), .B1(n4789), .B2(
        \reg_out[3][30] ), .ZN(n2896) );
  OAI221_X2 U864 ( .B1(n3609), .B2(n4841), .C1(n3532), .C2(n4834), .A(n2899), 
        .ZN(n2898) );
  AOI22_X2 U865 ( .A1(n4826), .A2(\reg_out[21][30] ), .B1(n4819), .B2(
        \reg_out[23][30] ), .ZN(n2899) );
  OAI221_X2 U866 ( .B1(n3608), .B2(n4812), .C1(n3531), .C2(n4804), .A(n2900), 
        .ZN(n2897) );
  AOI22_X2 U867 ( .A1(n4797), .A2(\reg_out[17][30] ), .B1(n4790), .B2(
        \reg_out[19][30] ), .ZN(n2900) );
  OAI221_X2 U869 ( .B1(n3607), .B2(n4840), .C1(n3530), .C2(n4833), .A(n2903), 
        .ZN(n2902) );
  AOI22_X2 U870 ( .A1(n4826), .A2(\reg_out[13][30] ), .B1(n4818), .B2(
        \reg_out[15][30] ), .ZN(n2903) );
  OAI221_X2 U871 ( .B1(n3606), .B2(n4811), .C1(n3529), .C2(n4805), .A(n2904), 
        .ZN(n2901) );
  AOI22_X2 U872 ( .A1(n4797), .A2(\reg_out[9][30] ), .B1(n4789), .B2(
        \reg_out[11][30] ), .ZN(n2904) );
  OAI221_X2 U874 ( .B1(n3605), .B2(n4841), .C1(n3528), .C2(n4834), .A(n2907), 
        .ZN(n2906) );
  AOI22_X2 U875 ( .A1(n4827), .A2(\reg_out[29][30] ), .B1(n4819), .B2(
        \reg_out[31][30] ), .ZN(n2907) );
  OAI221_X2 U876 ( .B1(n3604), .B2(n4812), .C1(n3527), .C2(n4804), .A(n2908), 
        .ZN(n2905) );
  AOI22_X2 U877 ( .A1(n4798), .A2(\reg_out[25][30] ), .B1(n4790), .B2(
        \reg_out[27][30] ), .ZN(n2908) );
  NAND4_X2 U878 ( .A1(n2909), .A2(n2910), .A3(n2911), .A4(n2912), .ZN(busA[2])
         );
  OAI221_X2 U880 ( .B1(n3603), .B2(n4841), .C1(n3526), .C2(n4834), .A(n2915), 
        .ZN(n2914) );
  AOI22_X2 U881 ( .A1(n4827), .A2(\reg_out[5][2] ), .B1(n4819), .B2(
        \reg_out[7][2] ), .ZN(n2915) );
  OAI221_X2 U882 ( .B1(n3602), .B2(n4812), .C1(n3525), .C2(n4804), .A(n2916), 
        .ZN(n2913) );
  AOI22_X2 U883 ( .A1(n4798), .A2(\reg_out[1][2] ), .B1(n4790), .B2(
        \reg_out[3][2] ), .ZN(n2916) );
  OAI221_X2 U885 ( .B1(n3601), .B2(n4840), .C1(n3524), .C2(n4833), .A(n2919), 
        .ZN(n2918) );
  AOI22_X2 U886 ( .A1(n4825), .A2(\reg_out[21][2] ), .B1(n4818), .B2(
        \reg_out[23][2] ), .ZN(n2919) );
  OAI221_X2 U887 ( .B1(n3600), .B2(n4811), .C1(n3523), .C2(n4805), .A(n2920), 
        .ZN(n2917) );
  AOI22_X2 U888 ( .A1(n4796), .A2(\reg_out[17][2] ), .B1(n4789), .B2(
        \reg_out[19][2] ), .ZN(n2920) );
  OAI221_X2 U890 ( .B1(n3599), .B2(n4841), .C1(n3522), .C2(n4834), .A(n2923), 
        .ZN(n2922) );
  AOI22_X2 U891 ( .A1(n4824), .A2(\reg_out[13][2] ), .B1(n4819), .B2(
        \reg_out[15][2] ), .ZN(n2923) );
  OAI221_X2 U892 ( .B1(n3598), .B2(n4812), .C1(n3521), .C2(n4804), .A(n2924), 
        .ZN(n2921) );
  AOI22_X2 U893 ( .A1(n4795), .A2(\reg_out[9][2] ), .B1(n4790), .B2(
        \reg_out[11][2] ), .ZN(n2924) );
  OAI221_X2 U895 ( .B1(n3597), .B2(n4840), .C1(n3520), .C2(n4833), .A(n2927), 
        .ZN(n2926) );
  AOI22_X2 U896 ( .A1(n4826), .A2(\reg_out[29][2] ), .B1(n4818), .B2(
        \reg_out[31][2] ), .ZN(n2927) );
  OAI221_X2 U897 ( .B1(n3596), .B2(n4811), .C1(n3519), .C2(n4805), .A(n2928), 
        .ZN(n2925) );
  AOI22_X2 U898 ( .A1(n4797), .A2(\reg_out[25][2] ), .B1(n4789), .B2(
        \reg_out[27][2] ), .ZN(n2928) );
  NAND4_X2 U899 ( .A1(n2929), .A2(n2930), .A3(n2931), .A4(n2932), .ZN(busA[29]) );
  OAI221_X2 U901 ( .B1(n3986), .B2(n4841), .C1(n3711), .C2(n4834), .A(n2935), 
        .ZN(n2934) );
  AOI22_X2 U902 ( .A1(n4827), .A2(\reg_out[5][29] ), .B1(n4819), .B2(
        \reg_out[7][29] ), .ZN(n2935) );
  OAI221_X2 U903 ( .B1(n4486), .B2(n4812), .C1(n3863), .C2(n4805), .A(n2936), 
        .ZN(n2933) );
  AOI22_X2 U904 ( .A1(n4798), .A2(\reg_out[1][29] ), .B1(n4790), .B2(
        \reg_out[3][29] ), .ZN(n2936) );
  OAI221_X2 U906 ( .B1(n4485), .B2(n4841), .C1(n3862), .C2(n4834), .A(n2939), 
        .ZN(n2938) );
  AOI22_X2 U907 ( .A1(n4827), .A2(\reg_out[21][29] ), .B1(n4819), .B2(
        \reg_out[23][29] ), .ZN(n2939) );
  OAI221_X2 U908 ( .B1(n4484), .B2(n4812), .C1(n3861), .C2(n4805), .A(n2940), 
        .ZN(n2937) );
  AOI22_X2 U909 ( .A1(n4798), .A2(\reg_out[17][29] ), .B1(n4790), .B2(
        \reg_out[19][29] ), .ZN(n2940) );
  OAI221_X2 U911 ( .B1(n4483), .B2(n4841), .C1(n3860), .C2(n4834), .A(n2943), 
        .ZN(n2942) );
  AOI22_X2 U912 ( .A1(n4827), .A2(\reg_out[13][29] ), .B1(n4819), .B2(
        \reg_out[15][29] ), .ZN(n2943) );
  OAI221_X2 U913 ( .B1(n3985), .B2(n4812), .C1(n4437), .C2(n4805), .A(n2944), 
        .ZN(n2941) );
  AOI22_X2 U914 ( .A1(n4798), .A2(\reg_out[9][29] ), .B1(n4790), .B2(
        \reg_out[11][29] ), .ZN(n2944) );
  OAI221_X2 U916 ( .B1(n4482), .B2(n4841), .C1(n3859), .C2(n4834), .A(n2947), 
        .ZN(n2946) );
  AOI22_X2 U917 ( .A1(n4827), .A2(\reg_out[29][29] ), .B1(n4819), .B2(
        \reg_out[31][29] ), .ZN(n2947) );
  OAI221_X2 U918 ( .B1(n4481), .B2(n4812), .C1(n3858), .C2(n4805), .A(n2948), 
        .ZN(n2945) );
  AOI22_X2 U919 ( .A1(n4798), .A2(\reg_out[25][29] ), .B1(n4790), .B2(
        \reg_out[27][29] ), .ZN(n2948) );
  NAND4_X2 U920 ( .A1(n2949), .A2(n2950), .A3(n2951), .A4(n2952), .ZN(busA[28]) );
  OAI221_X2 U922 ( .B1(n3984), .B2(n4841), .C1(n3710), .C2(n4834), .A(n2955), 
        .ZN(n2954) );
  AOI22_X2 U923 ( .A1(n4827), .A2(\reg_out[5][28] ), .B1(n4819), .B2(
        \reg_out[7][28] ), .ZN(n2955) );
  OAI221_X2 U924 ( .B1(n3983), .B2(n4812), .C1(n3709), .C2(n4805), .A(n2956), 
        .ZN(n2953) );
  AOI22_X2 U925 ( .A1(n4798), .A2(\reg_out[1][28] ), .B1(n4790), .B2(
        \reg_out[3][28] ), .ZN(n2956) );
  OAI221_X2 U927 ( .B1(n3982), .B2(n4841), .C1(n3708), .C2(n4834), .A(n2959), 
        .ZN(n2958) );
  AOI22_X2 U928 ( .A1(n4827), .A2(\reg_out[21][28] ), .B1(n4819), .B2(
        \reg_out[23][28] ), .ZN(n2959) );
  OAI221_X2 U929 ( .B1(n3981), .B2(n4812), .C1(n3707), .C2(n4805), .A(n2960), 
        .ZN(n2957) );
  AOI22_X2 U930 ( .A1(n4798), .A2(\reg_out[17][28] ), .B1(n4790), .B2(
        \reg_out[19][28] ), .ZN(n2960) );
  OAI221_X2 U932 ( .B1(n3980), .B2(n4841), .C1(n3706), .C2(n4834), .A(n2963), 
        .ZN(n2962) );
  AOI22_X2 U933 ( .A1(n4827), .A2(\reg_out[13][28] ), .B1(n4819), .B2(
        \reg_out[15][28] ), .ZN(n2963) );
  OAI221_X2 U934 ( .B1(n3979), .B2(n4812), .C1(n3705), .C2(n4805), .A(n2964), 
        .ZN(n2961) );
  AOI22_X2 U935 ( .A1(n4798), .A2(\reg_out[9][28] ), .B1(n4790), .B2(
        \reg_out[11][28] ), .ZN(n2964) );
  OAI221_X2 U937 ( .B1(n3978), .B2(n4841), .C1(n3704), .C2(n4834), .A(n2967), 
        .ZN(n2966) );
  AOI22_X2 U938 ( .A1(n4827), .A2(\reg_out[29][28] ), .B1(n4819), .B2(
        \reg_out[31][28] ), .ZN(n2967) );
  OAI221_X2 U939 ( .B1(n3977), .B2(n4812), .C1(n3703), .C2(n4805), .A(n2968), 
        .ZN(n2965) );
  AOI22_X2 U940 ( .A1(n4798), .A2(\reg_out[25][28] ), .B1(n4790), .B2(
        \reg_out[27][28] ), .ZN(n2968) );
  NAND4_X2 U941 ( .A1(n2969), .A2(n2970), .A3(n2971), .A4(n2972), .ZN(busA[27]) );
  OAI221_X2 U943 ( .B1(n3976), .B2(n4841), .C1(n3702), .C2(n4834), .A(n2975), 
        .ZN(n2974) );
  AOI22_X2 U944 ( .A1(n4827), .A2(\reg_out[5][27] ), .B1(n4819), .B2(
        \reg_out[7][27] ), .ZN(n2975) );
  OAI221_X2 U945 ( .B1(n3975), .B2(n4812), .C1(n3701), .C2(n4805), .A(n2976), 
        .ZN(n2973) );
  AOI22_X2 U946 ( .A1(n4798), .A2(\reg_out[1][27] ), .B1(n4790), .B2(
        \reg_out[3][27] ), .ZN(n2976) );
  OAI221_X2 U948 ( .B1(n3974), .B2(n4841), .C1(n3700), .C2(n4834), .A(n2979), 
        .ZN(n2978) );
  AOI22_X2 U949 ( .A1(n4827), .A2(\reg_out[21][27] ), .B1(n4819), .B2(
        \reg_out[23][27] ), .ZN(n2979) );
  OAI221_X2 U950 ( .B1(n3973), .B2(n4812), .C1(n3699), .C2(n4805), .A(n2980), 
        .ZN(n2977) );
  AOI22_X2 U951 ( .A1(n4798), .A2(\reg_out[17][27] ), .B1(n4790), .B2(
        \reg_out[19][27] ), .ZN(n2980) );
  OAI221_X2 U953 ( .B1(n3972), .B2(n4841), .C1(n3698), .C2(n4834), .A(n2983), 
        .ZN(n2982) );
  AOI22_X2 U954 ( .A1(n4827), .A2(\reg_out[13][27] ), .B1(n4819), .B2(
        \reg_out[15][27] ), .ZN(n2983) );
  OAI221_X2 U955 ( .B1(n3971), .B2(n4812), .C1(n3697), .C2(n4805), .A(n2984), 
        .ZN(n2981) );
  AOI22_X2 U956 ( .A1(n4798), .A2(\reg_out[9][27] ), .B1(n4790), .B2(
        \reg_out[11][27] ), .ZN(n2984) );
  OAI221_X2 U958 ( .B1(n3970), .B2(n4840), .C1(n3696), .C2(n4833), .A(n2987), 
        .ZN(n2986) );
  AOI22_X2 U959 ( .A1(n4826), .A2(\reg_out[29][27] ), .B1(n4818), .B2(
        \reg_out[31][27] ), .ZN(n2987) );
  OAI221_X2 U960 ( .B1(n3969), .B2(n4811), .C1(n3695), .C2(n4804), .A(n2988), 
        .ZN(n2985) );
  AOI22_X2 U961 ( .A1(n4797), .A2(\reg_out[25][27] ), .B1(n4789), .B2(
        \reg_out[27][27] ), .ZN(n2988) );
  NAND4_X2 U962 ( .A1(n2989), .A2(n2990), .A3(n2991), .A4(n2992), .ZN(busA[26]) );
  OAI221_X2 U964 ( .B1(n3968), .B2(n4840), .C1(n3694), .C2(n4833), .A(n2995), 
        .ZN(n2994) );
  AOI22_X2 U965 ( .A1(n4826), .A2(\reg_out[5][26] ), .B1(n4818), .B2(
        \reg_out[7][26] ), .ZN(n2995) );
  OAI221_X2 U966 ( .B1(n3967), .B2(n4811), .C1(n3693), .C2(n4804), .A(n2996), 
        .ZN(n2993) );
  AOI22_X2 U967 ( .A1(n4797), .A2(\reg_out[1][26] ), .B1(n4789), .B2(
        \reg_out[3][26] ), .ZN(n2996) );
  OAI221_X2 U969 ( .B1(n3966), .B2(n4840), .C1(n3692), .C2(n4833), .A(n2999), 
        .ZN(n2998) );
  AOI22_X2 U970 ( .A1(n4826), .A2(\reg_out[21][26] ), .B1(n4818), .B2(
        \reg_out[23][26] ), .ZN(n2999) );
  OAI221_X2 U971 ( .B1(n3965), .B2(n4811), .C1(n3691), .C2(n4804), .A(n3000), 
        .ZN(n2997) );
  AOI22_X2 U972 ( .A1(n4797), .A2(\reg_out[17][26] ), .B1(n4789), .B2(
        \reg_out[19][26] ), .ZN(n3000) );
  OAI221_X2 U974 ( .B1(n3964), .B2(n4840), .C1(n3690), .C2(n4833), .A(n3003), 
        .ZN(n3002) );
  AOI22_X2 U975 ( .A1(n4826), .A2(\reg_out[13][26] ), .B1(n4818), .B2(
        \reg_out[15][26] ), .ZN(n3003) );
  OAI221_X2 U976 ( .B1(n3963), .B2(n4811), .C1(n3689), .C2(n4804), .A(n3004), 
        .ZN(n3001) );
  AOI22_X2 U977 ( .A1(n4797), .A2(\reg_out[9][26] ), .B1(n4789), .B2(
        \reg_out[11][26] ), .ZN(n3004) );
  OAI221_X2 U979 ( .B1(n3962), .B2(n4840), .C1(n3688), .C2(n4833), .A(n3007), 
        .ZN(n3006) );
  AOI22_X2 U980 ( .A1(n4826), .A2(\reg_out[29][26] ), .B1(n4818), .B2(
        \reg_out[31][26] ), .ZN(n3007) );
  OAI221_X2 U981 ( .B1(n3961), .B2(n4811), .C1(n3687), .C2(n4804), .A(n3008), 
        .ZN(n3005) );
  AOI22_X2 U982 ( .A1(n4797), .A2(\reg_out[25][26] ), .B1(n4789), .B2(
        \reg_out[27][26] ), .ZN(n3008) );
  NAND4_X2 U983 ( .A1(n3009), .A2(n3010), .A3(n3011), .A4(n3012), .ZN(busA[25]) );
  OAI221_X2 U985 ( .B1(n3960), .B2(n4840), .C1(n3686), .C2(n4833), .A(n3015), 
        .ZN(n3014) );
  AOI22_X2 U986 ( .A1(n4826), .A2(\reg_out[5][25] ), .B1(n4818), .B2(
        \reg_out[7][25] ), .ZN(n3015) );
  OAI221_X2 U987 ( .B1(n3959), .B2(n4811), .C1(n3685), .C2(n4804), .A(n3016), 
        .ZN(n3013) );
  AOI22_X2 U988 ( .A1(n4797), .A2(\reg_out[1][25] ), .B1(n4789), .B2(
        \reg_out[3][25] ), .ZN(n3016) );
  OAI221_X2 U990 ( .B1(n3958), .B2(n4840), .C1(n3684), .C2(n4833), .A(n3019), 
        .ZN(n3018) );
  AOI22_X2 U991 ( .A1(n4826), .A2(\reg_out[21][25] ), .B1(n4818), .B2(
        \reg_out[23][25] ), .ZN(n3019) );
  OAI221_X2 U992 ( .B1(n3957), .B2(n4811), .C1(n3683), .C2(n4804), .A(n3020), 
        .ZN(n3017) );
  AOI22_X2 U993 ( .A1(n4797), .A2(\reg_out[17][25] ), .B1(n4789), .B2(
        \reg_out[19][25] ), .ZN(n3020) );
  OAI221_X2 U995 ( .B1(n3956), .B2(n4840), .C1(n3682), .C2(n4833), .A(n3023), 
        .ZN(n3022) );
  AOI22_X2 U996 ( .A1(n4826), .A2(\reg_out[13][25] ), .B1(n4818), .B2(
        \reg_out[15][25] ), .ZN(n3023) );
  OAI221_X2 U997 ( .B1(n3955), .B2(n4811), .C1(n3681), .C2(n4804), .A(n3024), 
        .ZN(n3021) );
  AOI22_X2 U998 ( .A1(n4797), .A2(\reg_out[9][25] ), .B1(n4789), .B2(
        \reg_out[11][25] ), .ZN(n3024) );
  OAI221_X2 U1000 ( .B1(n3954), .B2(n4840), .C1(n3680), .C2(n4833), .A(n3027), 
        .ZN(n3026) );
  AOI22_X2 U1001 ( .A1(n4826), .A2(\reg_out[29][25] ), .B1(n4818), .B2(
        \reg_out[31][25] ), .ZN(n3027) );
  OAI221_X2 U1002 ( .B1(n3953), .B2(n4811), .C1(n3679), .C2(n4804), .A(n3028), 
        .ZN(n3025) );
  AOI22_X2 U1003 ( .A1(n4797), .A2(\reg_out[25][25] ), .B1(n4789), .B2(
        \reg_out[27][25] ), .ZN(n3028) );
  NAND4_X2 U1004 ( .A1(n3029), .A2(n3030), .A3(n3031), .A4(n3032), .ZN(
        busA[24]) );
  OAI221_X2 U1006 ( .B1(n3952), .B2(n4840), .C1(n3678), .C2(n4833), .A(n3035), 
        .ZN(n3034) );
  AOI22_X2 U1007 ( .A1(n4826), .A2(\reg_out[5][24] ), .B1(n4818), .B2(
        \reg_out[7][24] ), .ZN(n3035) );
  OAI221_X2 U1008 ( .B1(n3951), .B2(n4811), .C1(n3677), .C2(n4804), .A(n3036), 
        .ZN(n3033) );
  AOI22_X2 U1009 ( .A1(n4797), .A2(\reg_out[1][24] ), .B1(n4789), .B2(
        \reg_out[3][24] ), .ZN(n3036) );
  OAI221_X2 U1011 ( .B1(n3950), .B2(n4840), .C1(n3676), .C2(n4833), .A(n3039), 
        .ZN(n3038) );
  AOI22_X2 U1012 ( .A1(n4826), .A2(\reg_out[21][24] ), .B1(n4818), .B2(
        \reg_out[23][24] ), .ZN(n3039) );
  OAI221_X2 U1013 ( .B1(n3949), .B2(n4811), .C1(n3675), .C2(n4804), .A(n3040), 
        .ZN(n3037) );
  AOI22_X2 U1014 ( .A1(n4797), .A2(\reg_out[17][24] ), .B1(n4789), .B2(
        \reg_out[19][24] ), .ZN(n3040) );
  OAI221_X2 U1016 ( .B1(n3948), .B2(n4839), .C1(n3518), .C2(n4831), .A(n3043), 
        .ZN(n3042) );
  AOI22_X2 U1017 ( .A1(n4826), .A2(\reg_out[13][24] ), .B1(n4817), .B2(
        \reg_out[15][24] ), .ZN(n3043) );
  OAI221_X2 U1018 ( .B1(n3947), .B2(n4810), .C1(n3517), .C2(n4802), .A(n3044), 
        .ZN(n3041) );
  AOI22_X2 U1019 ( .A1(n4797), .A2(\reg_out[9][24] ), .B1(n4787), .B2(
        \reg_out[11][24] ), .ZN(n3044) );
  OAI221_X2 U1021 ( .B1(n3946), .B2(n4838), .C1(n3516), .C2(n4831), .A(n3047), 
        .ZN(n3046) );
  AOI22_X2 U1022 ( .A1(n4826), .A2(\reg_out[29][24] ), .B1(n4816), .B2(
        \reg_out[31][24] ), .ZN(n3047) );
  OAI221_X2 U1023 ( .B1(n3945), .B2(n4809), .C1(n3515), .C2(n4802), .A(n3048), 
        .ZN(n3045) );
  AOI22_X2 U1024 ( .A1(n4797), .A2(\reg_out[25][24] ), .B1(n4788), .B2(
        \reg_out[27][24] ), .ZN(n3048) );
  NAND4_X2 U1025 ( .A1(n3049), .A2(n3050), .A3(n3051), .A4(n3052), .ZN(
        busA[23]) );
  OAI221_X2 U1027 ( .B1(n3944), .B2(n4838), .C1(n3514), .C2(n4831), .A(n3055), 
        .ZN(n3054) );
  AOI22_X2 U1028 ( .A1(n4826), .A2(\reg_out[5][23] ), .B1(n4816), .B2(
        \reg_out[7][23] ), .ZN(n3055) );
  OAI221_X2 U1029 ( .B1(n3943), .B2(n4809), .C1(n3513), .C2(n4802), .A(n3056), 
        .ZN(n3053) );
  AOI22_X2 U1030 ( .A1(n4797), .A2(\reg_out[1][23] ), .B1(n4788), .B2(
        \reg_out[3][23] ), .ZN(n3056) );
  OAI221_X2 U1032 ( .B1(n3942), .B2(n4839), .C1(n3512), .C2(n4831), .A(n3059), 
        .ZN(n3058) );
  AOI22_X2 U1033 ( .A1(n4826), .A2(\reg_out[21][23] ), .B1(n4817), .B2(
        \reg_out[23][23] ), .ZN(n3059) );
  OAI221_X2 U1034 ( .B1(n3941), .B2(n4810), .C1(n3511), .C2(n4802), .A(n3060), 
        .ZN(n3057) );
  AOI22_X2 U1035 ( .A1(n4797), .A2(\reg_out[17][23] ), .B1(n4788), .B2(
        \reg_out[19][23] ), .ZN(n3060) );
  OAI221_X2 U1037 ( .B1(n3940), .B2(n4838), .C1(n3510), .C2(n4832), .A(n3063), 
        .ZN(n3062) );
  AOI22_X2 U1038 ( .A1(n4826), .A2(\reg_out[13][23] ), .B1(n4816), .B2(
        \reg_out[15][23] ), .ZN(n3063) );
  OAI221_X2 U1039 ( .B1(n3939), .B2(n4809), .C1(n3509), .C2(n4803), .A(n3064), 
        .ZN(n3061) );
  AOI22_X2 U1040 ( .A1(n4797), .A2(\reg_out[9][23] ), .B1(n4788), .B2(
        \reg_out[11][23] ), .ZN(n3064) );
  OAI221_X2 U1042 ( .B1(n3938), .B2(n4839), .C1(n3508), .C2(n4831), .A(n3067), 
        .ZN(n3066) );
  AOI22_X2 U1043 ( .A1(n4826), .A2(\reg_out[29][23] ), .B1(n4817), .B2(
        \reg_out[31][23] ), .ZN(n3067) );
  OAI221_X2 U1044 ( .B1(n3937), .B2(n4810), .C1(n3507), .C2(n4802), .A(n3068), 
        .ZN(n3065) );
  AOI22_X2 U1045 ( .A1(n4797), .A2(\reg_out[25][23] ), .B1(n4787), .B2(
        \reg_out[27][23] ), .ZN(n3068) );
  NAND4_X2 U1046 ( .A1(n3069), .A2(n3070), .A3(n3071), .A4(n3072), .ZN(
        busA[22]) );
  OAI221_X2 U1048 ( .B1(n3936), .B2(n4839), .C1(n3506), .C2(n4831), .A(n3075), 
        .ZN(n3074) );
  AOI22_X2 U1049 ( .A1(n4826), .A2(\reg_out[5][22] ), .B1(n4817), .B2(
        \reg_out[7][22] ), .ZN(n3075) );
  OAI221_X2 U1050 ( .B1(n3935), .B2(n4810), .C1(n3505), .C2(n4802), .A(n3076), 
        .ZN(n3073) );
  AOI22_X2 U1051 ( .A1(n4797), .A2(\reg_out[1][22] ), .B1(n4788), .B2(
        \reg_out[3][22] ), .ZN(n3076) );
  OAI221_X2 U1053 ( .B1(n3934), .B2(n4838), .C1(n3504), .C2(n4832), .A(n3079), 
        .ZN(n3078) );
  AOI22_X2 U1054 ( .A1(n4826), .A2(\reg_out[21][22] ), .B1(n4816), .B2(
        \reg_out[23][22] ), .ZN(n3079) );
  OAI221_X2 U1055 ( .B1(n3933), .B2(n4809), .C1(n3503), .C2(n4803), .A(n3080), 
        .ZN(n3077) );
  AOI22_X2 U1056 ( .A1(n4797), .A2(\reg_out[17][22] ), .B1(n4788), .B2(
        \reg_out[19][22] ), .ZN(n3080) );
  OAI221_X2 U1058 ( .B1(n3932), .B2(n4839), .C1(n3502), .C2(n4832), .A(n3083), 
        .ZN(n3082) );
  AOI22_X2 U1059 ( .A1(n4826), .A2(\reg_out[13][22] ), .B1(n4817), .B2(
        \reg_out[15][22] ), .ZN(n3083) );
  OAI221_X2 U1060 ( .B1(n3931), .B2(n4810), .C1(n3501), .C2(n4803), .A(n3084), 
        .ZN(n3081) );
  AOI22_X2 U1061 ( .A1(n4797), .A2(\reg_out[9][22] ), .B1(n4787), .B2(
        \reg_out[11][22] ), .ZN(n3084) );
  OAI221_X2 U1063 ( .B1(n3930), .B2(n4838), .C1(n3500), .C2(n4832), .A(n3087), 
        .ZN(n3086) );
  AOI22_X2 U1064 ( .A1(n4826), .A2(\reg_out[29][22] ), .B1(n4816), .B2(
        \reg_out[31][22] ), .ZN(n3087) );
  OAI221_X2 U1065 ( .B1(n3929), .B2(n4809), .C1(n3499), .C2(n4803), .A(n3088), 
        .ZN(n3085) );
  AOI22_X2 U1066 ( .A1(n4797), .A2(\reg_out[25][22] ), .B1(n4788), .B2(
        \reg_out[27][22] ), .ZN(n3088) );
  NAND4_X2 U1067 ( .A1(n3089), .A2(n3090), .A3(n3091), .A4(n3092), .ZN(
        busA[21]) );
  OAI221_X2 U1069 ( .B1(n3928), .B2(n4838), .C1(n3498), .C2(n4832), .A(n3095), 
        .ZN(n3094) );
  AOI22_X2 U1070 ( .A1(n4826), .A2(\reg_out[5][21] ), .B1(n4816), .B2(
        \reg_out[7][21] ), .ZN(n3095) );
  OAI221_X2 U1071 ( .B1(n3927), .B2(n4809), .C1(n3497), .C2(n4803), .A(n3096), 
        .ZN(n3093) );
  AOI22_X2 U1072 ( .A1(n4797), .A2(\reg_out[1][21] ), .B1(n4788), .B2(
        \reg_out[3][21] ), .ZN(n3096) );
  OAI221_X2 U1074 ( .B1(n3926), .B2(n4839), .C1(n3674), .C2(n4832), .A(n3099), 
        .ZN(n3098) );
  AOI22_X2 U1075 ( .A1(n4825), .A2(\reg_out[21][21] ), .B1(n4817), .B2(
        \reg_out[23][21] ), .ZN(n3099) );
  OAI221_X2 U1076 ( .B1(n3925), .B2(n4810), .C1(n3673), .C2(n4803), .A(n3100), 
        .ZN(n3097) );
  AOI22_X2 U1077 ( .A1(n4796), .A2(\reg_out[17][21] ), .B1(n4788), .B2(
        \reg_out[19][21] ), .ZN(n3100) );
  OAI221_X2 U1079 ( .B1(n3924), .B2(n4839), .C1(n3672), .C2(n4832), .A(n3103), 
        .ZN(n3102) );
  AOI22_X2 U1080 ( .A1(n4825), .A2(\reg_out[13][21] ), .B1(n4817), .B2(
        \reg_out[15][21] ), .ZN(n3103) );
  OAI221_X2 U1081 ( .B1(n3923), .B2(n4810), .C1(n3671), .C2(n4803), .A(n3104), 
        .ZN(n3101) );
  AOI22_X2 U1082 ( .A1(n4796), .A2(\reg_out[9][21] ), .B1(n4788), .B2(
        \reg_out[11][21] ), .ZN(n3104) );
  OAI221_X2 U1084 ( .B1(n3922), .B2(n4839), .C1(n3670), .C2(n4832), .A(n3107), 
        .ZN(n3106) );
  AOI22_X2 U1085 ( .A1(n4825), .A2(\reg_out[29][21] ), .B1(n4817), .B2(
        \reg_out[31][21] ), .ZN(n3107) );
  OAI221_X2 U1086 ( .B1(n3921), .B2(n4810), .C1(n3669), .C2(n4803), .A(n3108), 
        .ZN(n3105) );
  AOI22_X2 U1087 ( .A1(n4796), .A2(\reg_out[25][21] ), .B1(n4788), .B2(
        \reg_out[27][21] ), .ZN(n3108) );
  NAND4_X2 U1088 ( .A1(n3109), .A2(n3110), .A3(n3111), .A4(n3112), .ZN(
        busA[20]) );
  OAI221_X2 U1090 ( .B1(n3920), .B2(n4839), .C1(n3668), .C2(n4832), .A(n3115), 
        .ZN(n3114) );
  AOI22_X2 U1091 ( .A1(n4825), .A2(\reg_out[5][20] ), .B1(n4817), .B2(
        \reg_out[7][20] ), .ZN(n3115) );
  OAI221_X2 U1092 ( .B1(n3919), .B2(n4810), .C1(n3667), .C2(n4803), .A(n3116), 
        .ZN(n3113) );
  AOI22_X2 U1093 ( .A1(n4796), .A2(\reg_out[1][20] ), .B1(n4788), .B2(
        \reg_out[3][20] ), .ZN(n3116) );
  OAI221_X2 U1095 ( .B1(n3918), .B2(n4839), .C1(n3666), .C2(n4832), .A(n3119), 
        .ZN(n3118) );
  AOI22_X2 U1096 ( .A1(n4825), .A2(\reg_out[21][20] ), .B1(n4817), .B2(
        \reg_out[23][20] ), .ZN(n3119) );
  OAI221_X2 U1097 ( .B1(n3917), .B2(n4810), .C1(n3665), .C2(n4803), .A(n3120), 
        .ZN(n3117) );
  AOI22_X2 U1098 ( .A1(n4796), .A2(\reg_out[17][20] ), .B1(n4788), .B2(
        \reg_out[19][20] ), .ZN(n3120) );
  OAI221_X2 U1100 ( .B1(n3916), .B2(n4839), .C1(n3664), .C2(n4832), .A(n3123), 
        .ZN(n3122) );
  AOI22_X2 U1101 ( .A1(n4825), .A2(\reg_out[13][20] ), .B1(n4817), .B2(
        \reg_out[15][20] ), .ZN(n3123) );
  OAI221_X2 U1102 ( .B1(n3915), .B2(n4810), .C1(n3663), .C2(n4803), .A(n3124), 
        .ZN(n3121) );
  AOI22_X2 U1103 ( .A1(n4796), .A2(\reg_out[9][20] ), .B1(n4788), .B2(
        \reg_out[11][20] ), .ZN(n3124) );
  OAI221_X2 U1105 ( .B1(n3914), .B2(n4839), .C1(n3662), .C2(n4832), .A(n3127), 
        .ZN(n3126) );
  AOI22_X2 U1106 ( .A1(n4825), .A2(\reg_out[29][20] ), .B1(n4817), .B2(
        \reg_out[31][20] ), .ZN(n3127) );
  OAI221_X2 U1107 ( .B1(n3913), .B2(n4810), .C1(n3661), .C2(n4803), .A(n3128), 
        .ZN(n3125) );
  AOI22_X2 U1108 ( .A1(n4796), .A2(\reg_out[25][20] ), .B1(n4788), .B2(
        \reg_out[27][20] ), .ZN(n3128) );
  NAND4_X2 U1109 ( .A1(n3129), .A2(n3130), .A3(n3131), .A4(n3132), .ZN(busA[1]) );
  OAI221_X2 U1111 ( .B1(n3912), .B2(n4839), .C1(n3660), .C2(n4832), .A(n3135), 
        .ZN(n3134) );
  AOI22_X2 U1112 ( .A1(n4825), .A2(\reg_out[5][1] ), .B1(n4817), .B2(
        \reg_out[7][1] ), .ZN(n3135) );
  OAI221_X2 U1113 ( .B1(n3911), .B2(n4810), .C1(n3659), .C2(n4803), .A(n3136), 
        .ZN(n3133) );
  AOI22_X2 U1114 ( .A1(n4796), .A2(\reg_out[1][1] ), .B1(n4788), .B2(
        \reg_out[3][1] ), .ZN(n3136) );
  OAI221_X2 U1116 ( .B1(n3910), .B2(n4839), .C1(n3658), .C2(n4832), .A(n3139), 
        .ZN(n3138) );
  AOI22_X2 U1117 ( .A1(n4825), .A2(\reg_out[21][1] ), .B1(n4817), .B2(
        \reg_out[23][1] ), .ZN(n3139) );
  OAI221_X2 U1118 ( .B1(n3909), .B2(n4810), .C1(n3657), .C2(n4803), .A(n3140), 
        .ZN(n3137) );
  AOI22_X2 U1119 ( .A1(n4796), .A2(\reg_out[17][1] ), .B1(n4788), .B2(
        \reg_out[19][1] ), .ZN(n3140) );
  OAI221_X2 U1121 ( .B1(n3908), .B2(n4839), .C1(n3656), .C2(n4832), .A(n3143), 
        .ZN(n3142) );
  AOI22_X2 U1122 ( .A1(n4825), .A2(\reg_out[13][1] ), .B1(n4817), .B2(
        \reg_out[15][1] ), .ZN(n3143) );
  OAI221_X2 U1123 ( .B1(n3907), .B2(n4810), .C1(n3655), .C2(n4803), .A(n3144), 
        .ZN(n3141) );
  AOI22_X2 U1124 ( .A1(n4796), .A2(\reg_out[9][1] ), .B1(n4788), .B2(
        \reg_out[11][1] ), .ZN(n3144) );
  OAI221_X2 U1126 ( .B1(n3906), .B2(n4839), .C1(n3654), .C2(n4832), .A(n3147), 
        .ZN(n3146) );
  AOI22_X2 U1127 ( .A1(n4825), .A2(\reg_out[29][1] ), .B1(n4817), .B2(
        \reg_out[31][1] ), .ZN(n3147) );
  OAI221_X2 U1128 ( .B1(n3905), .B2(n4810), .C1(n3653), .C2(n4803), .A(n3148), 
        .ZN(n3145) );
  AOI22_X2 U1129 ( .A1(n4796), .A2(\reg_out[25][1] ), .B1(n4788), .B2(
        \reg_out[27][1] ), .ZN(n3148) );
  NAND4_X2 U1130 ( .A1(n3149), .A2(n3150), .A3(n3151), .A4(n3152), .ZN(
        busA[19]) );
  OAI221_X2 U1132 ( .B1(n3904), .B2(n4838), .C1(n3652), .C2(n4831), .A(n3155), 
        .ZN(n3154) );
  AOI22_X2 U1133 ( .A1(n4824), .A2(\reg_out[5][19] ), .B1(n4816), .B2(
        \reg_out[7][19] ), .ZN(n3155) );
  OAI221_X2 U1134 ( .B1(n3903), .B2(n4809), .C1(n3651), .C2(n4802), .A(n3156), 
        .ZN(n3153) );
  AOI22_X2 U1135 ( .A1(n4795), .A2(\reg_out[1][19] ), .B1(n4787), .B2(
        \reg_out[3][19] ), .ZN(n3156) );
  OAI221_X2 U1137 ( .B1(n3902), .B2(n4838), .C1(n3650), .C2(n4831), .A(n3159), 
        .ZN(n3158) );
  AOI22_X2 U1138 ( .A1(n4824), .A2(\reg_out[21][19] ), .B1(n4816), .B2(
        \reg_out[23][19] ), .ZN(n3159) );
  OAI221_X2 U1139 ( .B1(n3901), .B2(n4809), .C1(n3649), .C2(n4802), .A(n3160), 
        .ZN(n3157) );
  AOI22_X2 U1140 ( .A1(n4795), .A2(\reg_out[17][19] ), .B1(n4787), .B2(
        \reg_out[19][19] ), .ZN(n3160) );
  OAI221_X2 U1142 ( .B1(n3900), .B2(n4838), .C1(n3648), .C2(n4831), .A(n3163), 
        .ZN(n3162) );
  AOI22_X2 U1143 ( .A1(n4824), .A2(\reg_out[13][19] ), .B1(n4816), .B2(
        \reg_out[15][19] ), .ZN(n3163) );
  OAI221_X2 U1144 ( .B1(n3899), .B2(n4809), .C1(n3647), .C2(n4802), .A(n3164), 
        .ZN(n3161) );
  AOI22_X2 U1145 ( .A1(n4795), .A2(\reg_out[9][19] ), .B1(n4787), .B2(
        \reg_out[11][19] ), .ZN(n3164) );
  OAI221_X2 U1147 ( .B1(n3898), .B2(n4838), .C1(n3646), .C2(n4831), .A(n3167), 
        .ZN(n3166) );
  AOI22_X2 U1148 ( .A1(n4824), .A2(\reg_out[29][19] ), .B1(n4816), .B2(
        \reg_out[31][19] ), .ZN(n3167) );
  OAI221_X2 U1149 ( .B1(n3897), .B2(n4809), .C1(n3645), .C2(n4802), .A(n3168), 
        .ZN(n3165) );
  AOI22_X2 U1150 ( .A1(n4795), .A2(\reg_out[25][19] ), .B1(n4787), .B2(
        \reg_out[27][19] ), .ZN(n3168) );
  NAND4_X2 U1151 ( .A1(n3169), .A2(n3170), .A3(n3171), .A4(n3172), .ZN(
        busA[18]) );
  OAI221_X2 U1153 ( .B1(n3896), .B2(n4838), .C1(n3644), .C2(n4831), .A(n3175), 
        .ZN(n3174) );
  AOI22_X2 U1154 ( .A1(n4824), .A2(\reg_out[5][18] ), .B1(n4816), .B2(
        \reg_out[7][18] ), .ZN(n3175) );
  OAI221_X2 U1155 ( .B1(n4480), .B2(n4809), .C1(n3857), .C2(n4802), .A(n3176), 
        .ZN(n3173) );
  AOI22_X2 U1156 ( .A1(n4795), .A2(\reg_out[1][18] ), .B1(n4787), .B2(
        \reg_out[3][18] ), .ZN(n3176) );
  OAI221_X2 U1158 ( .B1(n4479), .B2(n4838), .C1(n3643), .C2(n4831), .A(n3179), 
        .ZN(n3178) );
  AOI22_X2 U1159 ( .A1(n4824), .A2(\reg_out[21][18] ), .B1(n4816), .B2(
        \reg_out[23][18] ), .ZN(n3179) );
  OAI221_X2 U1160 ( .B1(n4478), .B2(n4809), .C1(n3856), .C2(n4802), .A(n3180), 
        .ZN(n3177) );
  AOI22_X2 U1161 ( .A1(n4795), .A2(\reg_out[17][18] ), .B1(n4787), .B2(
        \reg_out[19][18] ), .ZN(n3180) );
  OAI221_X2 U1163 ( .B1(n4477), .B2(n4838), .C1(n3855), .C2(n4831), .A(n3183), 
        .ZN(n3182) );
  AOI22_X2 U1164 ( .A1(n4824), .A2(\reg_out[13][18] ), .B1(n4816), .B2(
        \reg_out[15][18] ), .ZN(n3183) );
  OAI221_X2 U1165 ( .B1(n3895), .B2(n4809), .C1(n4436), .C2(n4802), .A(n3184), 
        .ZN(n3181) );
  AOI22_X2 U1166 ( .A1(n4795), .A2(\reg_out[9][18] ), .B1(n4787), .B2(
        \reg_out[11][18] ), .ZN(n3184) );
  OAI221_X2 U1168 ( .B1(n4476), .B2(n4838), .C1(n3854), .C2(n4831), .A(n3187), 
        .ZN(n3186) );
  AOI22_X2 U1169 ( .A1(n4824), .A2(\reg_out[29][18] ), .B1(n4816), .B2(
        \reg_out[31][18] ), .ZN(n3187) );
  OAI221_X2 U1170 ( .B1(n4475), .B2(n4809), .C1(n3642), .C2(n4802), .A(n3188), 
        .ZN(n3185) );
  AOI22_X2 U1171 ( .A1(n4795), .A2(\reg_out[25][18] ), .B1(n4787), .B2(
        \reg_out[27][18] ), .ZN(n3188) );
  NAND4_X2 U1172 ( .A1(n3189), .A2(n3190), .A3(n3191), .A4(n3192), .ZN(
        busA[17]) );
  OAI221_X2 U1174 ( .B1(n3894), .B2(n4838), .C1(n3641), .C2(n4831), .A(n3195), 
        .ZN(n3194) );
  AOI22_X2 U1175 ( .A1(n4824), .A2(\reg_out[5][17] ), .B1(n4816), .B2(
        \reg_out[7][17] ), .ZN(n3195) );
  OAI221_X2 U1176 ( .B1(n4474), .B2(n4809), .C1(n3853), .C2(n4802), .A(n3196), 
        .ZN(n3193) );
  AOI22_X2 U1177 ( .A1(n4795), .A2(\reg_out[1][17] ), .B1(n4787), .B2(
        \reg_out[3][17] ), .ZN(n3196) );
  OAI221_X2 U1179 ( .B1(n4473), .B2(n4838), .C1(n3640), .C2(n4831), .A(n3199), 
        .ZN(n3198) );
  AOI22_X2 U1180 ( .A1(n4824), .A2(\reg_out[21][17] ), .B1(n4816), .B2(
        \reg_out[23][17] ), .ZN(n3199) );
  OAI221_X2 U1181 ( .B1(n4472), .B2(n4809), .C1(n3852), .C2(n4802), .A(n3200), 
        .ZN(n3197) );
  AOI22_X2 U1182 ( .A1(n4795), .A2(\reg_out[17][17] ), .B1(n4787), .B2(
        \reg_out[19][17] ), .ZN(n3200) );
  OAI221_X2 U1184 ( .B1(n4471), .B2(n4838), .C1(n3851), .C2(n4831), .A(n3203), 
        .ZN(n3202) );
  AOI22_X2 U1185 ( .A1(n4824), .A2(\reg_out[13][17] ), .B1(n4816), .B2(
        \reg_out[15][17] ), .ZN(n3203) );
  OAI221_X2 U1186 ( .B1(n3893), .B2(n4809), .C1(n4435), .C2(n4802), .A(n3204), 
        .ZN(n3201) );
  AOI22_X2 U1187 ( .A1(n4795), .A2(\reg_out[9][17] ), .B1(n4787), .B2(
        \reg_out[11][17] ), .ZN(n3204) );
  OAI221_X2 U1189 ( .B1(n3753), .B2(n4843), .C1(n3850), .C2(n4830), .A(n3207), 
        .ZN(n3206) );
  AOI22_X2 U1190 ( .A1(n4822), .A2(\reg_out[29][17] ), .B1(n4821), .B2(
        \reg_out[31][17] ), .ZN(n3207) );
  OAI221_X2 U1191 ( .B1(n3752), .B2(n4814), .C1(n3575), .C2(n4801), .A(n3208), 
        .ZN(n3205) );
  AOI22_X2 U1192 ( .A1(n4793), .A2(\reg_out[25][17] ), .B1(n4792), .B2(
        \reg_out[27][17] ), .ZN(n3208) );
  NAND4_X2 U1193 ( .A1(n3209), .A2(n3210), .A3(n3211), .A4(n3212), .ZN(
        busA[16]) );
  OAI221_X2 U1195 ( .B1(n3892), .B2(n4843), .C1(n3639), .C2(n4830), .A(n3215), 
        .ZN(n3214) );
  AOI22_X2 U1196 ( .A1(n4822), .A2(\reg_out[5][16] ), .B1(n4821), .B2(
        \reg_out[7][16] ), .ZN(n3215) );
  OAI221_X2 U1197 ( .B1(n3891), .B2(n4814), .C1(n3638), .C2(n4801), .A(n3216), 
        .ZN(n3213) );
  AOI22_X2 U1198 ( .A1(n4793), .A2(\reg_out[1][16] ), .B1(n4792), .B2(
        \reg_out[3][16] ), .ZN(n3216) );
  OAI221_X2 U1200 ( .B1(n3751), .B2(n4843), .C1(n3574), .C2(n4830), .A(n3219), 
        .ZN(n3218) );
  AOI22_X2 U1201 ( .A1(n4822), .A2(\reg_out[21][16] ), .B1(n4821), .B2(
        \reg_out[23][16] ), .ZN(n3219) );
  OAI221_X2 U1202 ( .B1(n3890), .B2(n4814), .C1(n3573), .C2(n4801), .A(n3220), 
        .ZN(n3217) );
  AOI22_X2 U1203 ( .A1(n4793), .A2(\reg_out[17][16] ), .B1(n4792), .B2(
        \reg_out[19][16] ), .ZN(n3220) );
  OAI221_X2 U1205 ( .B1(n3889), .B2(n4843), .C1(n3572), .C2(n4830), .A(n3223), 
        .ZN(n3222) );
  AOI22_X2 U1206 ( .A1(n4822), .A2(\reg_out[13][16] ), .B1(n4821), .B2(
        \reg_out[15][16] ), .ZN(n3223) );
  OAI221_X2 U1207 ( .B1(n3888), .B2(n4814), .C1(n3571), .C2(n4801), .A(n3224), 
        .ZN(n3221) );
  AOI22_X2 U1208 ( .A1(n4793), .A2(\reg_out[9][16] ), .B1(n4792), .B2(
        \reg_out[11][16] ), .ZN(n3224) );
  OAI221_X2 U1210 ( .B1(n3750), .B2(n4843), .C1(n3849), .C2(n4830), .A(n3227), 
        .ZN(n3226) );
  AOI22_X2 U1211 ( .A1(n4822), .A2(\reg_out[29][16] ), .B1(n4821), .B2(
        \reg_out[31][16] ), .ZN(n3227) );
  OAI221_X2 U1212 ( .B1(n3749), .B2(n4814), .C1(n3570), .C2(n4801), .A(n3228), 
        .ZN(n3225) );
  AOI22_X2 U1213 ( .A1(n4793), .A2(\reg_out[25][16] ), .B1(n4792), .B2(
        \reg_out[27][16] ), .ZN(n3228) );
  NAND4_X2 U1214 ( .A1(n3229), .A2(n3230), .A3(n3231), .A4(n3232), .ZN(
        busA[15]) );
  OAI221_X2 U1216 ( .B1(n3887), .B2(n4843), .C1(n3637), .C2(n4830), .A(n3235), 
        .ZN(n3234) );
  AOI22_X2 U1217 ( .A1(n4822), .A2(\reg_out[5][15] ), .B1(n4821), .B2(
        \reg_out[7][15] ), .ZN(n3235) );
  OAI221_X2 U1218 ( .B1(n3886), .B2(n4814), .C1(n3636), .C2(n4801), .A(n3236), 
        .ZN(n3233) );
  AOI22_X2 U1219 ( .A1(n4793), .A2(\reg_out[1][15] ), .B1(n4792), .B2(
        \reg_out[3][15] ), .ZN(n3236) );
  OAI221_X2 U1221 ( .B1(n3748), .B2(n4843), .C1(n3569), .C2(n4830), .A(n3239), 
        .ZN(n3238) );
  AOI22_X2 U1222 ( .A1(n4822), .A2(\reg_out[21][15] ), .B1(n4821), .B2(
        \reg_out[23][15] ), .ZN(n3239) );
  OAI221_X2 U1223 ( .B1(n3885), .B2(n4814), .C1(n3568), .C2(n4801), .A(n3240), 
        .ZN(n3237) );
  AOI22_X2 U1224 ( .A1(n4793), .A2(\reg_out[17][15] ), .B1(n4792), .B2(
        \reg_out[19][15] ), .ZN(n3240) );
  OAI221_X2 U1226 ( .B1(n3884), .B2(n4843), .C1(n3567), .C2(n4830), .A(n3243), 
        .ZN(n3242) );
  AOI22_X2 U1227 ( .A1(n4822), .A2(\reg_out[13][15] ), .B1(n4821), .B2(
        \reg_out[15][15] ), .ZN(n3243) );
  OAI221_X2 U1228 ( .B1(n3883), .B2(n4814), .C1(n3566), .C2(n4801), .A(n3244), 
        .ZN(n3241) );
  AOI22_X2 U1229 ( .A1(n4793), .A2(\reg_out[9][15] ), .B1(n4792), .B2(
        \reg_out[11][15] ), .ZN(n3244) );
  OAI221_X2 U1231 ( .B1(n3747), .B2(n4843), .C1(n3848), .C2(n4830), .A(n3247), 
        .ZN(n3246) );
  AOI22_X2 U1232 ( .A1(n4822), .A2(\reg_out[29][15] ), .B1(n4821), .B2(
        \reg_out[31][15] ), .ZN(n3247) );
  OAI221_X2 U1233 ( .B1(n3746), .B2(n4814), .C1(n3565), .C2(n4801), .A(n3248), 
        .ZN(n3245) );
  AOI22_X2 U1234 ( .A1(n4793), .A2(\reg_out[25][15] ), .B1(n4792), .B2(
        \reg_out[27][15] ), .ZN(n3248) );
  NAND4_X2 U1235 ( .A1(n3249), .A2(n3250), .A3(n3251), .A4(n3252), .ZN(
        busA[14]) );
  OAI221_X2 U1237 ( .B1(n3882), .B2(n4843), .C1(n3635), .C2(n4830), .A(n3255), 
        .ZN(n3254) );
  AOI22_X2 U1238 ( .A1(n4822), .A2(\reg_out[5][14] ), .B1(n4821), .B2(
        \reg_out[7][14] ), .ZN(n3255) );
  OAI221_X2 U1239 ( .B1(n3881), .B2(n4814), .C1(n3634), .C2(n4801), .A(n3256), 
        .ZN(n3253) );
  AOI22_X2 U1240 ( .A1(n4793), .A2(\reg_out[1][14] ), .B1(n4792), .B2(
        \reg_out[3][14] ), .ZN(n3256) );
  OAI221_X2 U1242 ( .B1(n3745), .B2(n4843), .C1(n3564), .C2(n4830), .A(n3259), 
        .ZN(n3258) );
  AOI22_X2 U1243 ( .A1(n4822), .A2(\reg_out[21][14] ), .B1(n4821), .B2(
        \reg_out[23][14] ), .ZN(n3259) );
  OAI221_X2 U1244 ( .B1(n3880), .B2(n4814), .C1(n3563), .C2(n4801), .A(n3260), 
        .ZN(n3257) );
  AOI22_X2 U1245 ( .A1(n4793), .A2(\reg_out[17][14] ), .B1(n4792), .B2(
        \reg_out[19][14] ), .ZN(n3260) );
  OAI221_X2 U1247 ( .B1(n4470), .B2(n4842), .C1(n3847), .C2(n4830), .A(n3263), 
        .ZN(n3262) );
  AOI22_X2 U1248 ( .A1(n4823), .A2(\reg_out[13][14] ), .B1(n4820), .B2(
        \reg_out[15][14] ), .ZN(n3263) );
  OAI221_X2 U1249 ( .B1(n3879), .B2(n4813), .C1(n4434), .C2(n4801), .A(n3264), 
        .ZN(n3261) );
  AOI22_X2 U1250 ( .A1(n4794), .A2(\reg_out[9][14] ), .B1(n4791), .B2(
        \reg_out[11][14] ), .ZN(n3264) );
  OAI221_X2 U1252 ( .B1(n4469), .B2(n4842), .C1(n3846), .C2(n4830), .A(n3267), 
        .ZN(n3266) );
  AOI22_X2 U1253 ( .A1(n4823), .A2(\reg_out[29][14] ), .B1(n4820), .B2(
        \reg_out[31][14] ), .ZN(n3267) );
  OAI221_X2 U1254 ( .B1(n4468), .B2(n4813), .C1(n3633), .C2(n4801), .A(n3268), 
        .ZN(n3265) );
  AOI22_X2 U1255 ( .A1(n4794), .A2(\reg_out[25][14] ), .B1(n4787), .B2(
        \reg_out[27][14] ), .ZN(n3268) );
  NAND4_X2 U1256 ( .A1(n3269), .A2(n3270), .A3(n3271), .A4(n3272), .ZN(
        busA[13]) );
  OAI221_X2 U1258 ( .B1(n3878), .B2(n4842), .C1(n3632), .C2(n4830), .A(n3275), 
        .ZN(n3274) );
  AOI22_X2 U1259 ( .A1(n4823), .A2(\reg_out[5][13] ), .B1(n4820), .B2(
        \reg_out[7][13] ), .ZN(n3275) );
  OAI221_X2 U1260 ( .B1(n4467), .B2(n4813), .C1(n3845), .C2(n4801), .A(n3276), 
        .ZN(n3273) );
  AOI22_X2 U1261 ( .A1(n4794), .A2(\reg_out[1][13] ), .B1(n4791), .B2(
        \reg_out[3][13] ), .ZN(n3276) );
  OAI221_X2 U1263 ( .B1(n4466), .B2(n4842), .C1(n3631), .C2(n4830), .A(n3279), 
        .ZN(n3278) );
  AOI22_X2 U1264 ( .A1(n4823), .A2(\reg_out[21][13] ), .B1(n4820), .B2(
        \reg_out[23][13] ), .ZN(n3279) );
  OAI221_X2 U1265 ( .B1(n4465), .B2(n4813), .C1(n3844), .C2(n4801), .A(n3280), 
        .ZN(n3277) );
  AOI22_X2 U1266 ( .A1(n4794), .A2(\reg_out[17][13] ), .B1(n4791), .B2(
        \reg_out[19][13] ), .ZN(n3280) );
  OAI221_X2 U1268 ( .B1(n4464), .B2(n4842), .C1(n3843), .C2(n4830), .A(n3283), 
        .ZN(n3282) );
  AOI22_X2 U1269 ( .A1(n4823), .A2(\reg_out[13][13] ), .B1(n4819), .B2(
        \reg_out[15][13] ), .ZN(n3283) );
  OAI221_X2 U1270 ( .B1(n3877), .B2(n4813), .C1(n4433), .C2(n4801), .A(n3284), 
        .ZN(n3281) );
  AOI22_X2 U1271 ( .A1(n4794), .A2(\reg_out[9][13] ), .B1(n4787), .B2(
        \reg_out[11][13] ), .ZN(n3284) );
  OAI221_X2 U1273 ( .B1(n4463), .B2(n4839), .C1(n3842), .C2(n4831), .A(n3287), 
        .ZN(n3286) );
  AOI22_X2 U1274 ( .A1(n4823), .A2(\reg_out[29][13] ), .B1(n4819), .B2(
        \reg_out[31][13] ), .ZN(n3287) );
  OAI221_X2 U1275 ( .B1(n4462), .B2(n4810), .C1(n3630), .C2(n4802), .A(n3288), 
        .ZN(n3285) );
  AOI22_X2 U1276 ( .A1(n4794), .A2(\reg_out[25][13] ), .B1(n4791), .B2(
        \reg_out[27][13] ), .ZN(n3288) );
  NAND4_X2 U1277 ( .A1(n3289), .A2(n3290), .A3(n3291), .A4(n3292), .ZN(
        busA[12]) );
  OAI221_X2 U1279 ( .B1(n3876), .B2(n4842), .C1(n3629), .C2(n4830), .A(n3295), 
        .ZN(n3294) );
  AOI22_X2 U1280 ( .A1(n4823), .A2(\reg_out[5][12] ), .B1(n4820), .B2(
        \reg_out[7][12] ), .ZN(n3295) );
  OAI221_X2 U1281 ( .B1(n4461), .B2(n4813), .C1(n3841), .C2(n4801), .A(n3296), 
        .ZN(n3293) );
  AOI22_X2 U1282 ( .A1(n4794), .A2(\reg_out[1][12] ), .B1(n4791), .B2(
        \reg_out[3][12] ), .ZN(n3296) );
  OAI221_X2 U1284 ( .B1(n4460), .B2(n4842), .C1(n3628), .C2(n4830), .A(n3299), 
        .ZN(n3298) );
  AOI22_X2 U1285 ( .A1(n4823), .A2(\reg_out[21][12] ), .B1(n4820), .B2(
        \reg_out[23][12] ), .ZN(n3299) );
  OAI221_X2 U1286 ( .B1(n4459), .B2(n4813), .C1(n3840), .C2(n4801), .A(n3300), 
        .ZN(n3297) );
  AOI22_X2 U1287 ( .A1(n4794), .A2(\reg_out[17][12] ), .B1(n4787), .B2(
        \reg_out[19][12] ), .ZN(n3300) );
  OAI221_X2 U1289 ( .B1(n4458), .B2(n4842), .C1(n3839), .C2(n4830), .A(n3303), 
        .ZN(n3302) );
  AOI22_X2 U1290 ( .A1(n4823), .A2(\reg_out[13][12] ), .B1(n4817), .B2(
        \reg_out[15][12] ), .ZN(n3303) );
  OAI221_X2 U1291 ( .B1(n3875), .B2(n4813), .C1(n4432), .C2(n4801), .A(n3304), 
        .ZN(n3301) );
  AOI22_X2 U1292 ( .A1(n4794), .A2(\reg_out[9][12] ), .B1(n4791), .B2(
        \reg_out[11][12] ), .ZN(n3304) );
  OAI221_X2 U1294 ( .B1(n4457), .B2(n4841), .C1(n3838), .C2(n4832), .A(n3307), 
        .ZN(n3306) );
  AOI22_X2 U1295 ( .A1(n4823), .A2(\reg_out[29][12] ), .B1(n4817), .B2(
        \reg_out[31][12] ), .ZN(n3307) );
  OAI221_X2 U1296 ( .B1(n4456), .B2(n4812), .C1(n3627), .C2(n4803), .A(n3308), 
        .ZN(n3305) );
  AOI22_X2 U1297 ( .A1(n4794), .A2(\reg_out[25][12] ), .B1(n4790), .B2(
        \reg_out[27][12] ), .ZN(n3308) );
  NAND4_X2 U1298 ( .A1(n3309), .A2(n3310), .A3(n3311), .A4(n3312), .ZN(
        busA[11]) );
  OAI221_X2 U1300 ( .B1(n3874), .B2(n4842), .C1(n3626), .C2(n4830), .A(n3315), 
        .ZN(n3314) );
  AOI22_X2 U1301 ( .A1(n4823), .A2(\reg_out[5][11] ), .B1(n4820), .B2(
        \reg_out[7][11] ), .ZN(n3315) );
  OAI221_X2 U1302 ( .B1(n4455), .B2(n4813), .C1(n3837), .C2(n4801), .A(n3316), 
        .ZN(n3313) );
  AOI22_X2 U1303 ( .A1(n4794), .A2(\reg_out[1][11] ), .B1(n4787), .B2(
        \reg_out[3][11] ), .ZN(n3316) );
  OAI221_X2 U1305 ( .B1(n4454), .B2(n4837), .C1(n3625), .C2(n4835), .A(n3319), 
        .ZN(n3318) );
  AOI22_X2 U1306 ( .A1(n4823), .A2(\reg_out[21][11] ), .B1(n4815), .B2(
        \reg_out[23][11] ), .ZN(n3319) );
  OAI221_X2 U1307 ( .B1(n4453), .B2(n4808), .C1(n3836), .C2(n4806), .A(n3320), 
        .ZN(n3317) );
  AOI22_X2 U1308 ( .A1(n4794), .A2(\reg_out[17][11] ), .B1(n4786), .B2(
        \reg_out[19][11] ), .ZN(n3320) );
  OAI221_X2 U1310 ( .B1(n4452), .B2(n4837), .C1(n3835), .C2(n4835), .A(n3323), 
        .ZN(n3322) );
  AOI22_X2 U1311 ( .A1(n4825), .A2(\reg_out[13][11] ), .B1(n4815), .B2(
        \reg_out[15][11] ), .ZN(n3323) );
  OAI221_X2 U1312 ( .B1(n3873), .B2(n4808), .C1(n4431), .C2(n4806), .A(n3324), 
        .ZN(n3321) );
  AOI22_X2 U1313 ( .A1(n4799), .A2(\reg_out[9][11] ), .B1(n4786), .B2(
        \reg_out[11][11] ), .ZN(n3324) );
  OAI221_X2 U1315 ( .B1(n4451), .B2(n4837), .C1(n3834), .C2(n4833), .A(n3327), 
        .ZN(n3326) );
  AOI22_X2 U1316 ( .A1(n4828), .A2(\reg_out[29][11] ), .B1(n4815), .B2(
        \reg_out[31][11] ), .ZN(n3327) );
  OAI221_X2 U1317 ( .B1(n4450), .B2(n4808), .C1(n3624), .C2(n4805), .A(n3328), 
        .ZN(n3325) );
  AOI22_X2 U1318 ( .A1(n4796), .A2(\reg_out[25][11] ), .B1(n4786), .B2(
        \reg_out[27][11] ), .ZN(n3328) );
  NAND4_X2 U1319 ( .A1(n3329), .A2(n3330), .A3(n3331), .A4(n3332), .ZN(
        busA[10]) );
  OAI221_X2 U1321 ( .B1(n3872), .B2(n4837), .C1(n3623), .C2(n4836), .A(n3335), 
        .ZN(n3334) );
  AOI22_X2 U1322 ( .A1(n4823), .A2(\reg_out[5][10] ), .B1(n4815), .B2(
        \reg_out[7][10] ), .ZN(n3335) );
  OAI221_X2 U1323 ( .B1(n4449), .B2(n4808), .C1(n3833), .C2(n4807), .A(n3336), 
        .ZN(n3333) );
  AOI22_X2 U1324 ( .A1(n4794), .A2(\reg_out[1][10] ), .B1(n4786), .B2(
        \reg_out[3][10] ), .ZN(n3336) );
  OAI221_X2 U1326 ( .B1(n4448), .B2(n4837), .C1(n3622), .C2(n4834), .A(n3339), 
        .ZN(n3338) );
  AOI22_X2 U1327 ( .A1(n4822), .A2(\reg_out[21][10] ), .B1(n4815), .B2(
        \reg_out[23][10] ), .ZN(n3339) );
  OAI221_X2 U1328 ( .B1(n4447), .B2(n4808), .C1(n3832), .C2(n4804), .A(n3340), 
        .ZN(n3337) );
  AOI22_X2 U1329 ( .A1(n4793), .A2(\reg_out[17][10] ), .B1(n4786), .B2(
        \reg_out[19][10] ), .ZN(n3340) );
  OAI221_X2 U1331 ( .B1(n4446), .B2(n4837), .C1(n3831), .C2(n4832), .A(n3343), 
        .ZN(n3342) );
  AOI22_X2 U1332 ( .A1(n4824), .A2(\reg_out[13][10] ), .B1(n4815), .B2(
        \reg_out[15][10] ), .ZN(n3343) );
  OAI221_X2 U1333 ( .B1(n3871), .B2(n4808), .C1(n4430), .C2(n4803), .A(n3344), 
        .ZN(n3341) );
  AOI22_X2 U1334 ( .A1(n4795), .A2(\reg_out[9][10] ), .B1(n4786), .B2(
        \reg_out[11][10] ), .ZN(n3344) );
  OAI221_X2 U1336 ( .B1(n4445), .B2(n4837), .C1(n3830), .C2(n4836), .A(n3347), 
        .ZN(n3346) );
  AOI22_X2 U1337 ( .A1(n4822), .A2(\reg_out[29][10] ), .B1(n4815), .B2(
        \reg_out[31][10] ), .ZN(n3347) );
  OAI221_X2 U1338 ( .B1(n4444), .B2(n4808), .C1(n3621), .C2(n4807), .A(n3348), 
        .ZN(n3345) );
  AOI22_X2 U1339 ( .A1(n4799), .A2(\reg_out[25][10] ), .B1(n4786), .B2(
        \reg_out[27][10] ), .ZN(n3348) );
  NAND4_X2 U1340 ( .A1(n3349), .A2(n3350), .A3(n3351), .A4(n3352), .ZN(busA[0]) );
  OAI221_X2 U1343 ( .B1(n3870), .B2(n4837), .C1(n3620), .C2(n4836), .A(n3355), 
        .ZN(n3354) );
  AOI22_X2 U1344 ( .A1(n4823), .A2(\reg_out[5][0] ), .B1(n4815), .B2(
        \reg_out[7][0] ), .ZN(n3355) );
  OAI221_X2 U1345 ( .B1(n4443), .B2(n4808), .C1(n3829), .C2(n4807), .A(n3356), 
        .ZN(n3353) );
  AOI22_X2 U1346 ( .A1(n4794), .A2(\reg_out[1][0] ), .B1(n4786), .B2(
        \reg_out[3][0] ), .ZN(n3356) );
  OAI221_X2 U1349 ( .B1(n4442), .B2(n4837), .C1(n3619), .C2(n4836), .A(n3359), 
        .ZN(n3358) );
  AOI22_X2 U1350 ( .A1(n4828), .A2(\reg_out[21][0] ), .B1(n4815), .B2(
        \reg_out[23][0] ), .ZN(n3359) );
  OAI221_X2 U1351 ( .B1(n4441), .B2(n4808), .C1(n3828), .C2(n4807), .A(n3360), 
        .ZN(n3357) );
  AOI22_X2 U1352 ( .A1(n4793), .A2(\reg_out[17][0] ), .B1(n4786), .B2(
        \reg_out[19][0] ), .ZN(n3360) );
  OAI221_X2 U1355 ( .B1(n4440), .B2(n4837), .C1(n3827), .C2(n4834), .A(n3363), 
        .ZN(n3362) );
  AOI22_X2 U1356 ( .A1(n4822), .A2(\reg_out[13][0] ), .B1(n4815), .B2(
        \reg_out[15][0] ), .ZN(n3363) );
  OAI221_X2 U1357 ( .B1(n3869), .B2(n4808), .C1(n4429), .C2(n4804), .A(n3364), 
        .ZN(n3361) );
  AOI22_X2 U1358 ( .A1(n4793), .A2(\reg_out[9][0] ), .B1(n4786), .B2(
        \reg_out[11][0] ), .ZN(n3364) );
  OAI221_X2 U1361 ( .B1(n4439), .B2(n4837), .C1(n3826), .C2(n4835), .A(n3367), 
        .ZN(n3366) );
  AOI22_X2 U1362 ( .A1(n4825), .A2(\reg_out[29][0] ), .B1(n4815), .B2(
        \reg_out[31][0] ), .ZN(n3367) );
  OAI221_X2 U1367 ( .B1(n4438), .B2(n4808), .C1(n3618), .C2(n4806), .A(n3372), 
        .ZN(n3365) );
  AOI22_X2 U1368 ( .A1(n4795), .A2(\reg_out[25][0] ), .B1(n4786), .B2(
        \reg_out[27][0] ), .ZN(n3372) );
  AND2_X2 U1370 ( .A1(ra[4]), .A2(ra[3]), .ZN(n3368) );
  AND2_X2 U1372 ( .A1(ra[4]), .A2(n1031), .ZN(n3369) );
  OAI22_X2 U1377 ( .A1(n4779), .A2(n4777), .B1(n4217), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1378 ( .A1(n4776), .A2(n3376), .B1(n3804), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1379 ( .A1(n4776), .A2(n3377), .B1(n3803), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1380 ( .A1(n4776), .A2(n3378), .B1(n3802), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1381 ( .A1(n4776), .A2(n3379), .B1(n3801), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1382 ( .A1(n4776), .A2(n3380), .B1(n3800), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1383 ( .A1(n4776), .A2(n3381), .B1(n3799), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1384 ( .A1(n4776), .A2(n3382), .B1(n3798), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1385 ( .A1(n4777), .A2(n4758), .B1(n4216), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1386 ( .A1(n4776), .A2(n4756), .B1(n4215), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1387 ( .A1(n4776), .A2(n4754), .B1(n4214), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1388 ( .A1(n4776), .A2(n4752), .B1(n4213), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1389 ( .A1(n4776), .A2(n4750), .B1(n4212), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1390 ( .A1(n4777), .A2(n4748), .B1(n4211), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1391 ( .A1(n4777), .A2(n4746), .B1(n4210), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1392 ( .A1(n4777), .A2(n4744), .B1(n4209), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1393 ( .A1(n4777), .A2(n4742), .B1(n4208), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1394 ( .A1(n4777), .A2(n4740), .B1(n4207), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1395 ( .A1(n4777), .A2(n4738), .B1(n4206), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1396 ( .A1(n4777), .A2(n4736), .B1(n4205), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1397 ( .A1(n4777), .A2(n4734), .B1(n4204), .B2(n4775), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1398 ( .A1(n4777), .A2(n4732), .B1(n4203), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1399 ( .A1(n4777), .A2(n4730), .B1(n4202), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1400 ( .A1(n4777), .A2(n4728), .B1(n4201), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1401 ( .A1(n4777), .A2(n4726), .B1(n4200), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1402 ( .A1(n4777), .A2(n4724), .B1(n4199), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1403 ( .A1(n4777), .A2(n4722), .B1(n4198), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1404 ( .A1(n4777), .A2(n4720), .B1(n4197), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1405 ( .A1(n4777), .A2(n4718), .B1(n4196), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1406 ( .A1(n4777), .A2(n4716), .B1(n4195), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1407 ( .A1(n4777), .A2(n4714), .B1(n4194), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1408 ( .A1(n4777), .A2(n4712), .B1(n4193), .B2(n4774), .ZN(
        \REGISTER_FILE_32[9].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1411 ( .A1(n4778), .A2(n4710), .B1(n3773), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1412 ( .A1(n4772), .A2(n4710), .B1(n3765), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1413 ( .A1(n4770), .A2(n4710), .B1(n3763), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1414 ( .A1(n4768), .A2(n4710), .B1(n3761), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1415 ( .A1(n4766), .A2(n4710), .B1(n3759), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1416 ( .A1(n4764), .A2(n4710), .B1(n3757), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1417 ( .A1(n4762), .A2(n4710), .B1(n3755), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1418 ( .A1(n4760), .A2(n4710), .B1(n3614), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1419 ( .A1(n4759), .A2(n4710), .B1(n3606), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1420 ( .A1(n4757), .A2(n4710), .B1(n3598), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1421 ( .A1(n4755), .A2(n4710), .B1(n3985), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1422 ( .A1(n4753), .A2(n4711), .B1(n3979), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1423 ( .A1(n4751), .A2(n4711), .B1(n3971), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1424 ( .A1(n4749), .A2(n4711), .B1(n3963), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1425 ( .A1(n4747), .A2(n4711), .B1(n3955), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1426 ( .A1(n4745), .A2(n4711), .B1(n3947), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1427 ( .A1(n4743), .A2(n4711), .B1(n3939), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1428 ( .A1(n4741), .A2(n4711), .B1(n3931), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1429 ( .A1(n4739), .A2(n4711), .B1(n3923), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1430 ( .A1(n4737), .A2(n4711), .B1(n3915), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1431 ( .A1(n4735), .A2(n4711), .B1(n3907), .B2(n4709), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1432 ( .A1(n4733), .A2(n4711), .B1(n3899), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1433 ( .A1(n4731), .A2(n4711), .B1(n3895), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1434 ( .A1(n4729), .A2(n4711), .B1(n3893), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1435 ( .A1(n4727), .A2(n4711), .B1(n3888), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1436 ( .A1(n4725), .A2(n4711), .B1(n3883), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1437 ( .A1(n4723), .A2(n4711), .B1(n3879), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1438 ( .A1(n4721), .A2(n4711), .B1(n3877), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1439 ( .A1(n4719), .A2(n4711), .B1(n3875), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1440 ( .A1(n4717), .A2(n4711), .B1(n3873), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1441 ( .A1(n4715), .A2(n4711), .B1(n3871), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1442 ( .A1(n4713), .A2(n4711), .B1(n3869), .B2(n4708), .ZN(
        \REGISTER_FILE_32[8].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1445 ( .A1(n4778), .A2(n4706), .B1(n4397), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1446 ( .A1(n3376), .A2(n4706), .B1(n3825), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1447 ( .A1(n3377), .A2(n4706), .B1(n3824), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1448 ( .A1(n3378), .A2(n4706), .B1(n3823), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1449 ( .A1(n3379), .A2(n4706), .B1(n3822), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1450 ( .A1(n3380), .A2(n4706), .B1(n3821), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1451 ( .A1(n3381), .A2(n4706), .B1(n3820), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1452 ( .A1(n3382), .A2(n4706), .B1(n3819), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1453 ( .A1(n4759), .A2(n4706), .B1(n4396), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1454 ( .A1(n4757), .A2(n4706), .B1(n4395), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1455 ( .A1(n4755), .A2(n4706), .B1(n4394), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1456 ( .A1(n4753), .A2(n4707), .B1(n4393), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1457 ( .A1(n4751), .A2(n4707), .B1(n4392), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1458 ( .A1(n4749), .A2(n4707), .B1(n4391), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1459 ( .A1(n4747), .A2(n4707), .B1(n4390), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1460 ( .A1(n4745), .A2(n4707), .B1(n4389), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1461 ( .A1(n4743), .A2(n4707), .B1(n4388), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1462 ( .A1(n4741), .A2(n4707), .B1(n4387), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1463 ( .A1(n4739), .A2(n4707), .B1(n4386), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1464 ( .A1(n4737), .A2(n4707), .B1(n4385), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1465 ( .A1(n4735), .A2(n4707), .B1(n4384), .B2(n4705), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1466 ( .A1(n4733), .A2(n4707), .B1(n4383), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1467 ( .A1(n4731), .A2(n4707), .B1(n4382), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1468 ( .A1(n4729), .A2(n4707), .B1(n4381), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1469 ( .A1(n4727), .A2(n4707), .B1(n4380), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1470 ( .A1(n4725), .A2(n4707), .B1(n4379), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1471 ( .A1(n4723), .A2(n4707), .B1(n4378), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1472 ( .A1(n4721), .A2(n4707), .B1(n4377), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1473 ( .A1(n4719), .A2(n4707), .B1(n4376), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1474 ( .A1(n4717), .A2(n4707), .B1(n4375), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1475 ( .A1(n4715), .A2(n4707), .B1(n4374), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1476 ( .A1(n4713), .A2(n4707), .B1(n4373), .B2(n4704), .ZN(
        \REGISTER_FILE_32[7].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1479 ( .A1(n4779), .A2(n4702), .B1(n3595), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1480 ( .A1(n4772), .A2(n4702), .B1(n3587), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1481 ( .A1(n4770), .A2(n4702), .B1(n3581), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1482 ( .A1(n4768), .A2(n4702), .B1(n3580), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1483 ( .A1(n4766), .A2(n4702), .B1(n3579), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1484 ( .A1(n4764), .A2(n4702), .B1(n3578), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1485 ( .A1(n4762), .A2(n4702), .B1(n3577), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1486 ( .A1(n4760), .A2(n4702), .B1(n3576), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1487 ( .A1(n4759), .A2(n4702), .B1(n3534), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1488 ( .A1(n4757), .A2(n4702), .B1(n3526), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1489 ( .A1(n4755), .A2(n4702), .B1(n3711), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1490 ( .A1(n4753), .A2(n4703), .B1(n3710), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1491 ( .A1(n4751), .A2(n4703), .B1(n3702), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1492 ( .A1(n4749), .A2(n4703), .B1(n3694), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1493 ( .A1(n4747), .A2(n4703), .B1(n3686), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1494 ( .A1(n4745), .A2(n4703), .B1(n3678), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1495 ( .A1(n4743), .A2(n4703), .B1(n3514), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1496 ( .A1(n4741), .A2(n4703), .B1(n3506), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1497 ( .A1(n4739), .A2(n4703), .B1(n3498), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1498 ( .A1(n4737), .A2(n4703), .B1(n3668), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1499 ( .A1(n4735), .A2(n4703), .B1(n3660), .B2(n4701), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1500 ( .A1(n4733), .A2(n4703), .B1(n3652), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1501 ( .A1(n4731), .A2(n4703), .B1(n3644), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1502 ( .A1(n4729), .A2(n4703), .B1(n3641), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1503 ( .A1(n4727), .A2(n4703), .B1(n3639), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1504 ( .A1(n4725), .A2(n4703), .B1(n3637), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1505 ( .A1(n4723), .A2(n4703), .B1(n3635), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1506 ( .A1(n4721), .A2(n4703), .B1(n3632), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1507 ( .A1(n4719), .A2(n4703), .B1(n3629), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1508 ( .A1(n4717), .A2(n4703), .B1(n3626), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1509 ( .A1(n4715), .A2(n4703), .B1(n3623), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1510 ( .A1(n4713), .A2(n4703), .B1(n3620), .B2(n4700), .ZN(
        \REGISTER_FILE_32[6].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1513 ( .A1(n4779), .A2(n4698), .B1(n4192), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1514 ( .A1(n3376), .A2(n4698), .B1(n3797), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1515 ( .A1(n3377), .A2(n4698), .B1(n3796), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1516 ( .A1(n3378), .A2(n4698), .B1(n3795), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1517 ( .A1(n3379), .A2(n4698), .B1(n3794), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1518 ( .A1(n3380), .A2(n4698), .B1(n3793), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1519 ( .A1(n3381), .A2(n4698), .B1(n3792), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1520 ( .A1(n3382), .A2(n4698), .B1(n3791), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1521 ( .A1(n4759), .A2(n4698), .B1(n4191), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1522 ( .A1(n4757), .A2(n4698), .B1(n4190), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1523 ( .A1(n4755), .A2(n4698), .B1(n4189), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1524 ( .A1(n4753), .A2(n4699), .B1(n4188), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1525 ( .A1(n4751), .A2(n4699), .B1(n4187), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1526 ( .A1(n4749), .A2(n4699), .B1(n4186), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1527 ( .A1(n4747), .A2(n4699), .B1(n4185), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1528 ( .A1(n4745), .A2(n4699), .B1(n4184), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1529 ( .A1(n4743), .A2(n4699), .B1(n4183), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1530 ( .A1(n4741), .A2(n4699), .B1(n4182), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1531 ( .A1(n4739), .A2(n4699), .B1(n4181), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1532 ( .A1(n4737), .A2(n4699), .B1(n4180), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1533 ( .A1(n4735), .A2(n4699), .B1(n4179), .B2(n4697), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1534 ( .A1(n4733), .A2(n4699), .B1(n4178), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1535 ( .A1(n4731), .A2(n4699), .B1(n4177), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1536 ( .A1(n4729), .A2(n4699), .B1(n4176), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1537 ( .A1(n4727), .A2(n4699), .B1(n4175), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1538 ( .A1(n4725), .A2(n4699), .B1(n4174), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1539 ( .A1(n4723), .A2(n4699), .B1(n4173), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1540 ( .A1(n4721), .A2(n4699), .B1(n4172), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1541 ( .A1(n4719), .A2(n4699), .B1(n4171), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1542 ( .A1(n4717), .A2(n4699), .B1(n4170), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1543 ( .A1(n4715), .A2(n4699), .B1(n4169), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1544 ( .A1(n4713), .A2(n4699), .B1(n4168), .B2(n4696), .ZN(
        \REGISTER_FILE_32[5].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1547 ( .A1(n4778), .A2(n4694), .B1(n3778), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1548 ( .A1(n4772), .A2(n4694), .B1(n3770), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1549 ( .A1(n4770), .A2(n4694), .B1(n3764), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1550 ( .A1(n4768), .A2(n4694), .B1(n3762), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1551 ( .A1(n4766), .A2(n4694), .B1(n3760), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1552 ( .A1(n4764), .A2(n4694), .B1(n3758), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1553 ( .A1(n4762), .A2(n4694), .B1(n3756), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1554 ( .A1(n4760), .A2(n4694), .B1(n3754), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1555 ( .A1(n4759), .A2(n4694), .B1(n3611), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1556 ( .A1(n4757), .A2(n4694), .B1(n3603), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1557 ( .A1(n4755), .A2(n4694), .B1(n3986), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1558 ( .A1(n4753), .A2(n4695), .B1(n3984), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1559 ( .A1(n4751), .A2(n4695), .B1(n3976), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1560 ( .A1(n4749), .A2(n4695), .B1(n3968), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1561 ( .A1(n4747), .A2(n4695), .B1(n3960), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1562 ( .A1(n4745), .A2(n4695), .B1(n3952), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1563 ( .A1(n4743), .A2(n4695), .B1(n3944), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1564 ( .A1(n4741), .A2(n4695), .B1(n3936), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1565 ( .A1(n4739), .A2(n4695), .B1(n3928), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1566 ( .A1(n4737), .A2(n4695), .B1(n3920), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1567 ( .A1(n4735), .A2(n4695), .B1(n3912), .B2(n4693), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1568 ( .A1(n4733), .A2(n4695), .B1(n3904), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1569 ( .A1(n4731), .A2(n4695), .B1(n3896), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1570 ( .A1(n4729), .A2(n4695), .B1(n3894), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1571 ( .A1(n4727), .A2(n4695), .B1(n3892), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1572 ( .A1(n4725), .A2(n4695), .B1(n3887), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1573 ( .A1(n4723), .A2(n4695), .B1(n3882), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1574 ( .A1(n4721), .A2(n4695), .B1(n3878), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1575 ( .A1(n4719), .A2(n4695), .B1(n3876), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1576 ( .A1(n4717), .A2(n4695), .B1(n3874), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1577 ( .A1(n4715), .A2(n4695), .B1(n3872), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1578 ( .A1(n4713), .A2(n4695), .B1(n3870), .B2(n4692), .ZN(
        \REGISTER_FILE_32[4].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 )
         );
  AND3_X2 U1581 ( .A1(n1025), .A2(n1026), .A3(n3423), .ZN(n3414) );
  OAI22_X2 U1582 ( .A1(n4778), .A2(n4690), .B1(n4372), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1583 ( .A1(n3376), .A2(n4690), .B1(n3818), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1584 ( .A1(n3377), .A2(n4690), .B1(n3817), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1585 ( .A1(n3378), .A2(n4690), .B1(n3816), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1586 ( .A1(n3379), .A2(n4690), .B1(n3815), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1587 ( .A1(n3380), .A2(n4690), .B1(n3814), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1588 ( .A1(n3381), .A2(n4690), .B1(n3813), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1589 ( .A1(n3382), .A2(n4690), .B1(n3812), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1590 ( .A1(n4759), .A2(n4690), .B1(n4371), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1591 ( .A1(n4757), .A2(n4690), .B1(n4370), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1592 ( .A1(n4755), .A2(n4690), .B1(n4369), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1593 ( .A1(n4753), .A2(n4691), .B1(n4368), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1594 ( .A1(n4751), .A2(n4691), .B1(n4367), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1595 ( .A1(n4749), .A2(n4691), .B1(n4366), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1596 ( .A1(n4747), .A2(n4691), .B1(n4365), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1597 ( .A1(n4745), .A2(n4691), .B1(n4364), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1598 ( .A1(n4743), .A2(n4691), .B1(n4363), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1599 ( .A1(n4741), .A2(n4691), .B1(n4362), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1600 ( .A1(n4739), .A2(n4691), .B1(n4361), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1601 ( .A1(n4737), .A2(n4691), .B1(n4360), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1602 ( .A1(n4735), .A2(n4691), .B1(n4359), .B2(n4689), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1603 ( .A1(n4733), .A2(n4691), .B1(n4358), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1604 ( .A1(n4731), .A2(n4691), .B1(n4357), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1605 ( .A1(n4729), .A2(n4691), .B1(n4356), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1606 ( .A1(n4727), .A2(n4691), .B1(n4355), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1607 ( .A1(n4725), .A2(n4691), .B1(n4354), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1608 ( .A1(n4723), .A2(n4691), .B1(n4353), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1609 ( .A1(n4721), .A2(n4691), .B1(n4352), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1610 ( .A1(n4719), .A2(n4691), .B1(n4351), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1611 ( .A1(n4717), .A2(n4691), .B1(n4350), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1612 ( .A1(n4715), .A2(n4691), .B1(n4349), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1613 ( .A1(n4713), .A2(n4691), .B1(n4348), .B2(n4688), .ZN(
        \REGISTER_FILE_32[3].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1616 ( .A1(n4779), .A2(n4686), .B1(n4347), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1617 ( .A1(n4772), .A2(n4686), .B1(n3811), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1618 ( .A1(n4770), .A2(n4686), .B1(n3810), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1619 ( .A1(n4768), .A2(n4686), .B1(n3809), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1620 ( .A1(n4766), .A2(n4686), .B1(n3808), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1621 ( .A1(n4764), .A2(n4686), .B1(n3807), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1622 ( .A1(n4762), .A2(n4686), .B1(n3806), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1623 ( .A1(n4760), .A2(n4686), .B1(n3805), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1624 ( .A1(n4759), .A2(n4686), .B1(n4346), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1625 ( .A1(n4757), .A2(n4686), .B1(n4345), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1626 ( .A1(n4755), .A2(n4686), .B1(n4344), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1627 ( .A1(n4753), .A2(n4687), .B1(n4343), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1628 ( .A1(n4751), .A2(n4687), .B1(n4342), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1629 ( .A1(n4749), .A2(n4687), .B1(n4341), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1630 ( .A1(n4747), .A2(n4687), .B1(n4340), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1631 ( .A1(n4745), .A2(n4687), .B1(n4339), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1632 ( .A1(n4743), .A2(n4687), .B1(n4338), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1633 ( .A1(n4741), .A2(n4687), .B1(n4337), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1634 ( .A1(n4739), .A2(n4687), .B1(n4336), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1635 ( .A1(n4737), .A2(n4687), .B1(n4335), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1636 ( .A1(n4735), .A2(n4687), .B1(n4334), .B2(n4685), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1637 ( .A1(n4733), .A2(n4687), .B1(n4333), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1638 ( .A1(n4731), .A2(n4687), .B1(n4332), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1639 ( .A1(n4729), .A2(n4687), .B1(n4331), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1640 ( .A1(n4727), .A2(n4687), .B1(n4330), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1641 ( .A1(n4725), .A2(n4687), .B1(n4329), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1642 ( .A1(n4723), .A2(n4687), .B1(n4328), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1643 ( .A1(n4721), .A2(n4687), .B1(n4327), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1644 ( .A1(n4719), .A2(n4687), .B1(n4326), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1645 ( .A1(n4717), .A2(n4687), .B1(n4325), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1646 ( .A1(n4715), .A2(n4687), .B1(n4324), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1647 ( .A1(n4713), .A2(n4687), .B1(n4323), .B2(n4684), .ZN(
        \REGISTER_FILE_32[31].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1650 ( .A1(n4779), .A2(n4682), .B1(n3589), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1651 ( .A1(n4772), .A2(n4682), .B1(n3744), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1652 ( .A1(n4770), .A2(n4682), .B1(n3738), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1653 ( .A1(n4768), .A2(n4682), .B1(n3732), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1654 ( .A1(n4766), .A2(n4682), .B1(n3726), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1655 ( .A1(n4764), .A2(n4682), .B1(n3720), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1656 ( .A1(n4762), .A2(n4682), .B1(n3714), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1657 ( .A1(n4760), .A2(n4682), .B1(n3536), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1658 ( .A1(n4759), .A2(n4682), .B1(n3528), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1659 ( .A1(n4757), .A2(n4682), .B1(n3520), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1660 ( .A1(n4754), .A2(n4682), .B1(n3859), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1661 ( .A1(n4752), .A2(n4683), .B1(n3704), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1662 ( .A1(n4750), .A2(n4682), .B1(n3696), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1663 ( .A1(n4748), .A2(n4683), .B1(n3688), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1664 ( .A1(n4746), .A2(n4682), .B1(n3680), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1665 ( .A1(n4744), .A2(n4683), .B1(n3516), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1666 ( .A1(n4742), .A2(n4682), .B1(n3508), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1667 ( .A1(n4740), .A2(n4683), .B1(n3500), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1668 ( .A1(n4738), .A2(n4682), .B1(n3670), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1669 ( .A1(n4736), .A2(n4683), .B1(n3662), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1670 ( .A1(n4734), .A2(n4682), .B1(n3654), .B2(n4681), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1671 ( .A1(n4732), .A2(n4683), .B1(n3646), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1672 ( .A1(n4730), .A2(n4683), .B1(n3854), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1673 ( .A1(n4728), .A2(n4683), .B1(n3850), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1674 ( .A1(n4726), .A2(n4683), .B1(n3849), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1675 ( .A1(n4724), .A2(n4683), .B1(n3848), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1676 ( .A1(n4722), .A2(n4683), .B1(n3846), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1677 ( .A1(n4720), .A2(n4683), .B1(n3842), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1678 ( .A1(n4718), .A2(n4683), .B1(n3838), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1679 ( .A1(n4716), .A2(n4683), .B1(n3834), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1680 ( .A1(n4714), .A2(n4683), .B1(n3830), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1681 ( .A1(n4712), .A2(n4683), .B1(n3826), .B2(n4680), .ZN(
        \REGISTER_FILE_32[30].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1684 ( .A1(n4778), .A2(n4678), .B1(n3594), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1685 ( .A1(n4772), .A2(n4678), .B1(n3586), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1686 ( .A1(n4770), .A2(n4678), .B1(n3742), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1687 ( .A1(n4768), .A2(n4678), .B1(n3736), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1688 ( .A1(n4766), .A2(n4678), .B1(n3730), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1689 ( .A1(n4764), .A2(n4678), .B1(n3724), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1690 ( .A1(n4762), .A2(n4678), .B1(n3718), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1691 ( .A1(n4760), .A2(n4678), .B1(n3712), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1692 ( .A1(n4759), .A2(n4678), .B1(n3533), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1693 ( .A1(n4757), .A2(n4678), .B1(n3525), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1694 ( .A1(n4755), .A2(n4678), .B1(n3863), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1695 ( .A1(n4753), .A2(n4679), .B1(n3709), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1696 ( .A1(n4751), .A2(n4678), .B1(n3701), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1697 ( .A1(n4749), .A2(n4679), .B1(n3693), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1698 ( .A1(n4747), .A2(n4678), .B1(n3685), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1699 ( .A1(n4745), .A2(n4679), .B1(n3677), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1700 ( .A1(n4743), .A2(n4678), .B1(n3513), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1701 ( .A1(n4741), .A2(n4679), .B1(n3505), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1702 ( .A1(n4739), .A2(n4678), .B1(n3497), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1703 ( .A1(n4737), .A2(n4679), .B1(n3667), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1704 ( .A1(n4735), .A2(n4678), .B1(n3659), .B2(n4677), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1705 ( .A1(n4733), .A2(n4679), .B1(n3651), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1706 ( .A1(n4731), .A2(n4679), .B1(n3857), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1707 ( .A1(n4729), .A2(n4679), .B1(n3853), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1708 ( .A1(n4727), .A2(n4679), .B1(n3638), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1709 ( .A1(n4725), .A2(n4679), .B1(n3636), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1710 ( .A1(n4723), .A2(n4679), .B1(n3634), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1711 ( .A1(n4721), .A2(n4679), .B1(n3845), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1712 ( .A1(n4719), .A2(n4679), .B1(n3841), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1713 ( .A1(n4717), .A2(n4679), .B1(n3837), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1714 ( .A1(n4715), .A2(n4679), .B1(n3833), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1715 ( .A1(n4713), .A2(n4679), .B1(n3829), .B2(n4676), .ZN(
        \REGISTER_FILE_32[2].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U1718 ( .A1(n4779), .A2(n4674), .B1(n4167), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1719 ( .A1(n3376), .A2(n4674), .B1(n4166), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1720 ( .A1(n3377), .A2(n4674), .B1(n4165), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1721 ( .A1(n3378), .A2(n4674), .B1(n4164), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1722 ( .A1(n3379), .A2(n4674), .B1(n4163), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1723 ( .A1(n3380), .A2(n4674), .B1(n4162), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1724 ( .A1(n3381), .A2(n4674), .B1(n4161), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1725 ( .A1(n3382), .A2(n4674), .B1(n4160), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1726 ( .A1(n4759), .A2(n4674), .B1(n4159), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1727 ( .A1(n4757), .A2(n4674), .B1(n4158), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1728 ( .A1(n4755), .A2(n4674), .B1(n4552), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1729 ( .A1(n4753), .A2(n4674), .B1(n4157), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1730 ( .A1(n4751), .A2(n4674), .B1(n4156), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1731 ( .A1(n4749), .A2(n4674), .B1(n4155), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1732 ( .A1(n4747), .A2(n4674), .B1(n4154), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1733 ( .A1(n4745), .A2(n4674), .B1(n4153), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1734 ( .A1(n4743), .A2(n4674), .B1(n4152), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1735 ( .A1(n4741), .A2(n4674), .B1(n4151), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1736 ( .A1(n4739), .A2(n4674), .B1(n4150), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1737 ( .A1(n4737), .A2(n4674), .B1(n4149), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1738 ( .A1(n4735), .A2(n4674), .B1(n4148), .B2(n4673), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1739 ( .A1(n4733), .A2(n4674), .B1(n4147), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1740 ( .A1(n4731), .A2(n3434), .B1(n4551), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1741 ( .A1(n4729), .A2(n3434), .B1(n4550), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1742 ( .A1(n4727), .A2(n3434), .B1(n4549), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1743 ( .A1(n4725), .A2(n3434), .B1(n4548), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1744 ( .A1(n4723), .A2(n3434), .B1(n4547), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1745 ( .A1(n4721), .A2(n3434), .B1(n4546), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1746 ( .A1(n4719), .A2(n3434), .B1(n4545), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1747 ( .A1(n4717), .A2(n3434), .B1(n4544), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1748 ( .A1(n4715), .A2(n3434), .B1(n4543), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1749 ( .A1(n4713), .A2(n4674), .B1(n4542), .B2(n4672), .ZN(
        \REGISTER_FILE_32[29].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U1751 ( .A1(n3429), .A2(n3408), .ZN(n3434) );
  OAI22_X2 U1752 ( .A1(n4779), .A2(n4670), .B1(n3772), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1753 ( .A1(n3376), .A2(n4670), .B1(n4019), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1754 ( .A1(n3377), .A2(n4670), .B1(n4013), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1755 ( .A1(n3378), .A2(n4670), .B1(n4007), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1756 ( .A1(n3379), .A2(n4670), .B1(n4001), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1757 ( .A1(n3380), .A2(n4670), .B1(n3995), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1758 ( .A1(n3381), .A2(n4670), .B1(n3989), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1759 ( .A1(n3382), .A2(n4670), .B1(n3613), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1760 ( .A1(n4759), .A2(n4670), .B1(n3605), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1761 ( .A1(n4757), .A2(n4670), .B1(n3597), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1762 ( .A1(n4755), .A2(n4670), .B1(n4482), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1763 ( .A1(n4753), .A2(n4670), .B1(n3978), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1764 ( .A1(n4751), .A2(n4670), .B1(n3970), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1765 ( .A1(n4749), .A2(n4670), .B1(n3962), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1766 ( .A1(n4747), .A2(n4670), .B1(n3954), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1767 ( .A1(n4745), .A2(n4670), .B1(n3946), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1768 ( .A1(n4743), .A2(n4670), .B1(n3938), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1769 ( .A1(n4741), .A2(n4670), .B1(n3930), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1770 ( .A1(n4739), .A2(n4670), .B1(n3922), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1771 ( .A1(n4737), .A2(n4670), .B1(n3914), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1772 ( .A1(n4735), .A2(n4670), .B1(n3906), .B2(n4669), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1773 ( .A1(n4733), .A2(n4670), .B1(n3898), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1774 ( .A1(n4731), .A2(n3436), .B1(n4476), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1775 ( .A1(n4729), .A2(n3436), .B1(n3753), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1776 ( .A1(n4727), .A2(n3436), .B1(n3750), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1777 ( .A1(n4725), .A2(n3436), .B1(n3747), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1778 ( .A1(n4723), .A2(n3436), .B1(n4469), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1779 ( .A1(n4721), .A2(n3436), .B1(n4463), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1780 ( .A1(n4719), .A2(n3436), .B1(n4457), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1781 ( .A1(n4717), .A2(n3436), .B1(n4451), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1782 ( .A1(n4715), .A2(n3436), .B1(n4445), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1783 ( .A1(n4713), .A2(n4670), .B1(n4439), .B2(n4668), .ZN(
        \REGISTER_FILE_32[28].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U1785 ( .A1(n3429), .A2(n3411), .ZN(n3436) );
  AND3_X2 U1786 ( .A1(n3423), .A2(rd[1]), .A3(rd[0]), .ZN(n3429) );
  OAI22_X2 U1787 ( .A1(n4779), .A2(n4666), .B1(n4322), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1788 ( .A1(n3376), .A2(n4666), .B1(n4321), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1789 ( .A1(n3377), .A2(n4666), .B1(n4320), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1790 ( .A1(n3378), .A2(n4666), .B1(n4319), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1791 ( .A1(n3379), .A2(n4666), .B1(n4318), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1792 ( .A1(n3380), .A2(n4666), .B1(n4317), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1793 ( .A1(n3381), .A2(n4666), .B1(n4316), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1794 ( .A1(n3382), .A2(n4666), .B1(n4315), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1795 ( .A1(n4759), .A2(n4666), .B1(n4314), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1796 ( .A1(n4757), .A2(n4666), .B1(n4313), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1797 ( .A1(n4755), .A2(n4666), .B1(n4607), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1798 ( .A1(n4753), .A2(n4666), .B1(n4312), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1799 ( .A1(n4751), .A2(n4666), .B1(n4311), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1800 ( .A1(n4749), .A2(n4666), .B1(n4310), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1801 ( .A1(n4747), .A2(n4666), .B1(n4309), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1802 ( .A1(n4745), .A2(n4666), .B1(n4308), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1803 ( .A1(n4743), .A2(n4666), .B1(n4307), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1804 ( .A1(n4741), .A2(n4666), .B1(n4306), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1805 ( .A1(n4739), .A2(n4666), .B1(n4305), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1806 ( .A1(n4737), .A2(n4666), .B1(n4304), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1807 ( .A1(n4735), .A2(n4666), .B1(n4303), .B2(n4665), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1808 ( .A1(n4733), .A2(n4666), .B1(n4302), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1809 ( .A1(n4731), .A2(n3438), .B1(n4606), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1810 ( .A1(n4729), .A2(n3438), .B1(n4605), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1811 ( .A1(n4727), .A2(n3438), .B1(n4604), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1812 ( .A1(n4725), .A2(n3438), .B1(n4603), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1813 ( .A1(n4723), .A2(n3438), .B1(n4602), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1814 ( .A1(n4721), .A2(n3438), .B1(n4601), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1815 ( .A1(n4719), .A2(n3438), .B1(n4600), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1816 ( .A1(n4717), .A2(n3438), .B1(n4599), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1817 ( .A1(n4715), .A2(n4666), .B1(n4598), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1818 ( .A1(n4713), .A2(n4666), .B1(n4597), .B2(n4664), .ZN(
        \REGISTER_FILE_32[27].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U1820 ( .A1(n3440), .A2(n3415), .ZN(n3438) );
  OAI22_X2 U1821 ( .A1(n4779), .A2(n4662), .B1(n3588), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1822 ( .A1(n3376), .A2(n4662), .B1(n3743), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1823 ( .A1(n3377), .A2(n4662), .B1(n3737), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1824 ( .A1(n3378), .A2(n4662), .B1(n3731), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1825 ( .A1(n3379), .A2(n4662), .B1(n3725), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1826 ( .A1(n3380), .A2(n4662), .B1(n3719), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1827 ( .A1(n3381), .A2(n4662), .B1(n3713), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1828 ( .A1(n3382), .A2(n4662), .B1(n3535), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1829 ( .A1(n4759), .A2(n4662), .B1(n3527), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1830 ( .A1(n4757), .A2(n4662), .B1(n3519), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1831 ( .A1(n4755), .A2(n4662), .B1(n3858), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1832 ( .A1(n4753), .A2(n4662), .B1(n3703), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1833 ( .A1(n4751), .A2(n4662), .B1(n3695), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1834 ( .A1(n4749), .A2(n4662), .B1(n3687), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1835 ( .A1(n4747), .A2(n4662), .B1(n3679), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1836 ( .A1(n4745), .A2(n4662), .B1(n3515), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1837 ( .A1(n4743), .A2(n4662), .B1(n3507), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1838 ( .A1(n4741), .A2(n4662), .B1(n3499), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1839 ( .A1(n4739), .A2(n4662), .B1(n3669), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1840 ( .A1(n4737), .A2(n4662), .B1(n3661), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1841 ( .A1(n4735), .A2(n4662), .B1(n3653), .B2(n4661), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1842 ( .A1(n4733), .A2(n4662), .B1(n3645), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1843 ( .A1(n4731), .A2(n3441), .B1(n3642), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1844 ( .A1(n4729), .A2(n3441), .B1(n3575), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1845 ( .A1(n4727), .A2(n3441), .B1(n3570), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1846 ( .A1(n4725), .A2(n3441), .B1(n3565), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1847 ( .A1(n4723), .A2(n3441), .B1(n3633), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1848 ( .A1(n4721), .A2(n3441), .B1(n3630), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1849 ( .A1(n4719), .A2(n3441), .B1(n3627), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1850 ( .A1(n4717), .A2(n3441), .B1(n3624), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1851 ( .A1(n4715), .A2(n4662), .B1(n3621), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1852 ( .A1(n4713), .A2(n4662), .B1(n3618), .B2(n4660), .ZN(
        \REGISTER_FILE_32[26].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U1854 ( .A1(n3440), .A2(n3418), .ZN(n3441) );
  OAI22_X2 U1855 ( .A1(n4779), .A2(n4658), .B1(n4146), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1856 ( .A1(n3376), .A2(n4658), .B1(n4145), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1857 ( .A1(n3377), .A2(n4658), .B1(n4144), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1858 ( .A1(n3378), .A2(n4658), .B1(n4143), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1859 ( .A1(n3379), .A2(n4658), .B1(n4142), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1860 ( .A1(n3380), .A2(n4658), .B1(n4141), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1861 ( .A1(n3381), .A2(n4658), .B1(n4140), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1862 ( .A1(n3382), .A2(n4658), .B1(n4139), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1863 ( .A1(n4759), .A2(n4658), .B1(n4138), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1864 ( .A1(n4757), .A2(n4658), .B1(n4137), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1865 ( .A1(n4755), .A2(n4658), .B1(n4541), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1866 ( .A1(n4753), .A2(n4658), .B1(n4136), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1867 ( .A1(n4751), .A2(n4658), .B1(n4135), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1868 ( .A1(n4749), .A2(n4658), .B1(n4134), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1869 ( .A1(n4747), .A2(n4658), .B1(n4133), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1870 ( .A1(n4745), .A2(n4658), .B1(n4132), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1871 ( .A1(n4743), .A2(n4658), .B1(n4131), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1872 ( .A1(n4741), .A2(n4658), .B1(n4130), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1873 ( .A1(n4739), .A2(n4658), .B1(n4129), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1874 ( .A1(n4737), .A2(n4658), .B1(n4128), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1875 ( .A1(n4735), .A2(n4658), .B1(n4127), .B2(n4657), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1876 ( .A1(n4733), .A2(n4658), .B1(n4126), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1877 ( .A1(n4731), .A2(n3443), .B1(n4540), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1878 ( .A1(n4729), .A2(n3443), .B1(n4539), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1879 ( .A1(n4727), .A2(n3443), .B1(n4538), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1880 ( .A1(n4725), .A2(n3443), .B1(n4537), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1881 ( .A1(n4723), .A2(n3443), .B1(n4536), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1882 ( .A1(n4721), .A2(n3443), .B1(n4535), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1883 ( .A1(n4719), .A2(n3443), .B1(n4534), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1884 ( .A1(n4717), .A2(n4658), .B1(n4533), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1885 ( .A1(n4715), .A2(n4658), .B1(n4532), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1886 ( .A1(n4713), .A2(n4658), .B1(n4531), .B2(n4656), .ZN(
        \REGISTER_FILE_32[25].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U1888 ( .A1(n3440), .A2(n3408), .ZN(n3443) );
  OAI22_X2 U1889 ( .A1(n4779), .A2(n4654), .B1(n3771), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1890 ( .A1(n3376), .A2(n4654), .B1(n4018), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1891 ( .A1(n3377), .A2(n4654), .B1(n4012), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1892 ( .A1(n3378), .A2(n4654), .B1(n4006), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1893 ( .A1(n3379), .A2(n4654), .B1(n4000), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1894 ( .A1(n3380), .A2(n4654), .B1(n3994), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1895 ( .A1(n3381), .A2(n4654), .B1(n3988), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1896 ( .A1(n3382), .A2(n4654), .B1(n3612), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1897 ( .A1(n4759), .A2(n4654), .B1(n3604), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1898 ( .A1(n4757), .A2(n4654), .B1(n3596), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1899 ( .A1(n4755), .A2(n4654), .B1(n4481), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1900 ( .A1(n4753), .A2(n4654), .B1(n3977), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1901 ( .A1(n4751), .A2(n4654), .B1(n3969), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1902 ( .A1(n4749), .A2(n4654), .B1(n3961), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1903 ( .A1(n4747), .A2(n4654), .B1(n3953), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1904 ( .A1(n4745), .A2(n4654), .B1(n3945), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1905 ( .A1(n4743), .A2(n4654), .B1(n3937), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1906 ( .A1(n4741), .A2(n4654), .B1(n3929), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1907 ( .A1(n4739), .A2(n4654), .B1(n3921), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1908 ( .A1(n4737), .A2(n4654), .B1(n3913), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1909 ( .A1(n4735), .A2(n4654), .B1(n3905), .B2(n4653), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1910 ( .A1(n4733), .A2(n4654), .B1(n3897), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1911 ( .A1(n4731), .A2(n3445), .B1(n4475), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1912 ( .A1(n4729), .A2(n3445), .B1(n3752), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1913 ( .A1(n4727), .A2(n3445), .B1(n3749), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1914 ( .A1(n4725), .A2(n3445), .B1(n3746), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1915 ( .A1(n4723), .A2(n3445), .B1(n4468), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1916 ( .A1(n4721), .A2(n3445), .B1(n4462), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1917 ( .A1(n4719), .A2(n3445), .B1(n4456), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1918 ( .A1(n4717), .A2(n4654), .B1(n4450), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1919 ( .A1(n4715), .A2(n4654), .B1(n4444), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1920 ( .A1(n4713), .A2(n4654), .B1(n4438), .B2(n4652), .ZN(
        \REGISTER_FILE_32[24].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U1922 ( .A1(n3440), .A2(n3411), .ZN(n3445) );
  AND3_X2 U1923 ( .A1(rd[1]), .A2(n3447), .A3(rd[0]), .ZN(n3440) );
  OAI22_X2 U1924 ( .A1(n4779), .A2(n4650), .B1(n4301), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1925 ( .A1(n3376), .A2(n4650), .B1(n4300), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1926 ( .A1(n3377), .A2(n4650), .B1(n4299), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1927 ( .A1(n3378), .A2(n4650), .B1(n4298), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1928 ( .A1(n3379), .A2(n4650), .B1(n4297), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1929 ( .A1(n3380), .A2(n4650), .B1(n4296), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1930 ( .A1(n3381), .A2(n4650), .B1(n4295), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1931 ( .A1(n3382), .A2(n4650), .B1(n4294), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1932 ( .A1(n4759), .A2(n4650), .B1(n4293), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1933 ( .A1(n4757), .A2(n4650), .B1(n4292), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1934 ( .A1(n4755), .A2(n4650), .B1(n4596), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1935 ( .A1(n4753), .A2(n4650), .B1(n4291), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1936 ( .A1(n4751), .A2(n4650), .B1(n4290), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1937 ( .A1(n4749), .A2(n4650), .B1(n4289), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1938 ( .A1(n4747), .A2(n4650), .B1(n4288), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1939 ( .A1(n4745), .A2(n4650), .B1(n4287), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1940 ( .A1(n4743), .A2(n4650), .B1(n4286), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1941 ( .A1(n4741), .A2(n4650), .B1(n4285), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1942 ( .A1(n4739), .A2(n4650), .B1(n4284), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1943 ( .A1(n4737), .A2(n4650), .B1(n4283), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1944 ( .A1(n4735), .A2(n4650), .B1(n4282), .B2(n4649), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1945 ( .A1(n4733), .A2(n4650), .B1(n4281), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1946 ( .A1(n4731), .A2(n3448), .B1(n4595), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1947 ( .A1(n4729), .A2(n3448), .B1(n4594), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1948 ( .A1(n4727), .A2(n3448), .B1(n4593), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1949 ( .A1(n4725), .A2(n3448), .B1(n4592), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1950 ( .A1(n4723), .A2(n3448), .B1(n4591), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1951 ( .A1(n4721), .A2(n3448), .B1(n4590), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1952 ( .A1(n4719), .A2(n3448), .B1(n4589), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1953 ( .A1(n4717), .A2(n3448), .B1(n4588), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1954 ( .A1(n4715), .A2(n3448), .B1(n4587), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1955 ( .A1(n4713), .A2(n4650), .B1(n4586), .B2(n4648), .ZN(
        \REGISTER_FILE_32[23].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U1957 ( .A1(n3450), .A2(n3415), .ZN(n3448) );
  OAI22_X2 U1958 ( .A1(n4779), .A2(n4646), .B1(n3593), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1959 ( .A1(n3376), .A2(n4646), .B1(n3585), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1960 ( .A1(n3377), .A2(n4646), .B1(n3741), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1961 ( .A1(n3378), .A2(n4646), .B1(n3735), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1962 ( .A1(n3379), .A2(n4646), .B1(n3729), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1963 ( .A1(n3380), .A2(n4646), .B1(n3723), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1964 ( .A1(n3381), .A2(n4646), .B1(n3717), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1965 ( .A1(n3382), .A2(n4646), .B1(n3540), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1966 ( .A1(n4759), .A2(n4646), .B1(n3532), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1967 ( .A1(n4757), .A2(n4646), .B1(n3524), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1968 ( .A1(n4755), .A2(n4646), .B1(n3862), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1969 ( .A1(n4753), .A2(n4646), .B1(n3708), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1970 ( .A1(n4751), .A2(n4646), .B1(n3700), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1971 ( .A1(n4749), .A2(n4646), .B1(n3692), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1972 ( .A1(n4747), .A2(n4646), .B1(n3684), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1973 ( .A1(n4745), .A2(n4646), .B1(n3676), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1974 ( .A1(n4743), .A2(n4646), .B1(n3512), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1975 ( .A1(n4741), .A2(n4646), .B1(n3504), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1976 ( .A1(n4739), .A2(n4646), .B1(n3674), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1977 ( .A1(n4737), .A2(n4646), .B1(n3666), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1978 ( .A1(n4735), .A2(n4646), .B1(n3658), .B2(n4645), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1979 ( .A1(n4733), .A2(n4646), .B1(n3650), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1980 ( .A1(n4731), .A2(n3451), .B1(n3643), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1981 ( .A1(n4729), .A2(n3451), .B1(n3640), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1982 ( .A1(n4727), .A2(n3451), .B1(n3574), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1983 ( .A1(n4725), .A2(n3451), .B1(n3569), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1984 ( .A1(n4723), .A2(n3451), .B1(n3564), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1985 ( .A1(n4721), .A2(n3451), .B1(n3631), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1986 ( .A1(n4719), .A2(n3451), .B1(n3628), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1987 ( .A1(n4717), .A2(n3451), .B1(n3625), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1988 ( .A1(n4715), .A2(n3451), .B1(n3622), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1989 ( .A1(n4713), .A2(n4646), .B1(n3619), .B2(n4644), .ZN(
        \REGISTER_FILE_32[22].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U1991 ( .A1(n3450), .A2(n3418), .ZN(n3451) );
  OAI22_X2 U1992 ( .A1(n4779), .A2(n4642), .B1(n4125), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1993 ( .A1(n3376), .A2(n4642), .B1(n4124), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1994 ( .A1(n3377), .A2(n4642), .B1(n4123), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1995 ( .A1(n3378), .A2(n4642), .B1(n4122), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1996 ( .A1(n3379), .A2(n4642), .B1(n4121), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1997 ( .A1(n3380), .A2(n4642), .B1(n4120), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1998 ( .A1(n3381), .A2(n4642), .B1(n4119), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1999 ( .A1(n3382), .A2(n4642), .B1(n4118), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2000 ( .A1(n4759), .A2(n4642), .B1(n4117), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2001 ( .A1(n4757), .A2(n4642), .B1(n4116), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2002 ( .A1(n4755), .A2(n4642), .B1(n4530), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2003 ( .A1(n4753), .A2(n4642), .B1(n4115), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2004 ( .A1(n4751), .A2(n4642), .B1(n4114), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2005 ( .A1(n4749), .A2(n4642), .B1(n4113), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2006 ( .A1(n4747), .A2(n4642), .B1(n4112), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2007 ( .A1(n4745), .A2(n4642), .B1(n4111), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2008 ( .A1(n4743), .A2(n4642), .B1(n4110), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2009 ( .A1(n4741), .A2(n4642), .B1(n4109), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2010 ( .A1(n4739), .A2(n4642), .B1(n4108), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2011 ( .A1(n4737), .A2(n4642), .B1(n4107), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2012 ( .A1(n4735), .A2(n4642), .B1(n4106), .B2(n4641), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2013 ( .A1(n4733), .A2(n4642), .B1(n4105), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2014 ( .A1(n4731), .A2(n3453), .B1(n4529), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2015 ( .A1(n4729), .A2(n3453), .B1(n4528), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2016 ( .A1(n4727), .A2(n3453), .B1(n4527), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2017 ( .A1(n4725), .A2(n3453), .B1(n4526), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2018 ( .A1(n4723), .A2(n3453), .B1(n4525), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2019 ( .A1(n4721), .A2(n3453), .B1(n4524), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2020 ( .A1(n4719), .A2(n3453), .B1(n4523), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2021 ( .A1(n4717), .A2(n3453), .B1(n4522), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2022 ( .A1(n4715), .A2(n3453), .B1(n4521), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2023 ( .A1(n4713), .A2(n4642), .B1(n4520), .B2(n4640), .ZN(
        \REGISTER_FILE_32[21].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U2025 ( .A1(n3450), .A2(n3408), .ZN(n3453) );
  OAI22_X2 U2026 ( .A1(n4779), .A2(n4638), .B1(n3776), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2027 ( .A1(n3376), .A2(n4638), .B1(n3768), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2028 ( .A1(n3377), .A2(n4638), .B1(n4016), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2029 ( .A1(n3378), .A2(n4638), .B1(n4010), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2030 ( .A1(n3379), .A2(n4638), .B1(n4004), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2031 ( .A1(n3380), .A2(n4638), .B1(n3998), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2032 ( .A1(n3381), .A2(n4638), .B1(n3992), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2033 ( .A1(n3382), .A2(n4638), .B1(n3617), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2034 ( .A1(n4759), .A2(n4638), .B1(n3609), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2035 ( .A1(n4757), .A2(n4638), .B1(n3601), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2036 ( .A1(n4755), .A2(n4638), .B1(n4485), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2037 ( .A1(n4753), .A2(n4638), .B1(n3982), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2038 ( .A1(n4751), .A2(n4638), .B1(n3974), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2039 ( .A1(n4749), .A2(n4638), .B1(n3966), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2040 ( .A1(n4747), .A2(n4638), .B1(n3958), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2041 ( .A1(n4745), .A2(n4638), .B1(n3950), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2042 ( .A1(n4743), .A2(n4638), .B1(n3942), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2043 ( .A1(n4741), .A2(n4638), .B1(n3934), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2044 ( .A1(n4739), .A2(n4638), .B1(n3926), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2045 ( .A1(n4737), .A2(n4638), .B1(n3918), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2046 ( .A1(n4735), .A2(n4638), .B1(n3910), .B2(n4637), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2047 ( .A1(n4733), .A2(n4638), .B1(n3902), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2048 ( .A1(n4731), .A2(n3455), .B1(n4479), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2049 ( .A1(n4729), .A2(n3455), .B1(n4473), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2050 ( .A1(n4727), .A2(n3455), .B1(n3751), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2051 ( .A1(n4725), .A2(n3455), .B1(n3748), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2052 ( .A1(n4723), .A2(n3455), .B1(n3745), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2053 ( .A1(n4721), .A2(n3455), .B1(n4466), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2054 ( .A1(n4719), .A2(n3455), .B1(n4460), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2055 ( .A1(n4717), .A2(n3455), .B1(n4454), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2056 ( .A1(n4715), .A2(n3455), .B1(n4448), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2057 ( .A1(n4713), .A2(n4638), .B1(n4442), .B2(n4636), .ZN(
        \REGISTER_FILE_32[20].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U2059 ( .A1(n3450), .A2(n3411), .ZN(n3455) );
  AND3_X2 U2060 ( .A1(n3423), .A2(n1026), .A3(rd[0]), .ZN(n3450) );
  OAI22_X2 U2061 ( .A1(n4779), .A2(n4634), .B1(n4104), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U2062 ( .A1(n3376), .A2(n4634), .B1(n4103), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U2063 ( .A1(n3377), .A2(n4634), .B1(n4102), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U2064 ( .A1(n3378), .A2(n4634), .B1(n4101), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U2065 ( .A1(n3379), .A2(n4634), .B1(n4100), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U2066 ( .A1(n3380), .A2(n4634), .B1(n4099), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U2067 ( .A1(n3381), .A2(n4634), .B1(n4098), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U2068 ( .A1(n3382), .A2(n4634), .B1(n4097), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2069 ( .A1(n4759), .A2(n4634), .B1(n4096), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2070 ( .A1(n4757), .A2(n4634), .B1(n4095), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U2071 ( .A1(n4755), .A2(n4634), .B1(n4519), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2072 ( .A1(n4753), .A2(n4634), .B1(n4094), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2073 ( .A1(n4751), .A2(n4634), .B1(n4093), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2074 ( .A1(n4749), .A2(n4634), .B1(n4092), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2075 ( .A1(n4747), .A2(n4634), .B1(n4091), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2076 ( .A1(n4745), .A2(n4634), .B1(n4090), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2077 ( .A1(n4743), .A2(n4634), .B1(n4089), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2078 ( .A1(n4741), .A2(n4634), .B1(n4088), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2079 ( .A1(n4739), .A2(n4634), .B1(n4087), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2080 ( .A1(n4737), .A2(n4634), .B1(n4086), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2081 ( .A1(n4735), .A2(n4634), .B1(n4085), .B2(n4633), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U2082 ( .A1(n4733), .A2(n4634), .B1(n4084), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2083 ( .A1(n4731), .A2(n3457), .B1(n4518), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2084 ( .A1(n4729), .A2(n3457), .B1(n4517), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2085 ( .A1(n4727), .A2(n3457), .B1(n4516), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2086 ( .A1(n4725), .A2(n3457), .B1(n4515), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2087 ( .A1(n4723), .A2(n3457), .B1(n4514), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2088 ( .A1(n4721), .A2(n3457), .B1(n4513), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2089 ( .A1(n4719), .A2(n3457), .B1(n4512), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2090 ( .A1(n4717), .A2(n3457), .B1(n4511), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2091 ( .A1(n4715), .A2(n3457), .B1(n4510), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2092 ( .A1(n4713), .A2(n4634), .B1(n4509), .B2(n4632), .ZN(
        \REGISTER_FILE_32[1].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 )
         );
  NAND2_X2 U2094 ( .A1(n3426), .A2(n3408), .ZN(n3457) );
  OAI22_X2 U2095 ( .A1(n4778), .A2(n4630), .B1(n4280), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2096 ( .A1(n4772), .A2(n4630), .B1(n4279), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2097 ( .A1(n4770), .A2(n4630), .B1(n4278), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2098 ( .A1(n4768), .A2(n4630), .B1(n4277), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2099 ( .A1(n4766), .A2(n4630), .B1(n4276), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2100 ( .A1(n4764), .A2(n4630), .B1(n4275), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2101 ( .A1(n4762), .A2(n4630), .B1(n4274), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2102 ( .A1(n4760), .A2(n4630), .B1(n4273), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2103 ( .A1(n4758), .A2(n4630), .B1(n4272), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2104 ( .A1(n4756), .A2(n4630), .B1(n4271), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2105 ( .A1(n4754), .A2(n4630), .B1(n4585), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2106 ( .A1(n4752), .A2(n4630), .B1(n4270), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2107 ( .A1(n4750), .A2(n4630), .B1(n4269), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2108 ( .A1(n4748), .A2(n4630), .B1(n4268), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2109 ( .A1(n4746), .A2(n4630), .B1(n4267), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2110 ( .A1(n4744), .A2(n4630), .B1(n4266), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2111 ( .A1(n4742), .A2(n4630), .B1(n4265), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2112 ( .A1(n4740), .A2(n4630), .B1(n4264), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2113 ( .A1(n4738), .A2(n4630), .B1(n4263), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2114 ( .A1(n4736), .A2(n4630), .B1(n4262), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2115 ( .A1(n4734), .A2(n4630), .B1(n4261), .B2(n4629), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2116 ( .A1(n4732), .A2(n4630), .B1(n4260), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2117 ( .A1(n4730), .A2(n3459), .B1(n4584), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2118 ( .A1(n4728), .A2(n3459), .B1(n4583), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2119 ( .A1(n4726), .A2(n3459), .B1(n4582), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2120 ( .A1(n4724), .A2(n3459), .B1(n4581), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2121 ( .A1(n4722), .A2(n3459), .B1(n4580), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2122 ( .A1(n4720), .A2(n3459), .B1(n4579), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2123 ( .A1(n4718), .A2(n3459), .B1(n4578), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2124 ( .A1(n4716), .A2(n4630), .B1(n4577), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2125 ( .A1(n4714), .A2(n4630), .B1(n4576), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2126 ( .A1(n4712), .A2(n4630), .B1(n4575), .B2(n4628), .ZN(
        \REGISTER_FILE_32[19].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U2128 ( .A1(n3461), .A2(n3415), .ZN(n3459) );
  OAI22_X2 U2129 ( .A1(n4778), .A2(n3552), .B1(n3592), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2130 ( .A1(n4772), .A2(n3552), .B1(n3584), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2131 ( .A1(n4770), .A2(n3552), .B1(n3740), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2132 ( .A1(n4768), .A2(n3552), .B1(n3734), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2133 ( .A1(n4766), .A2(n3552), .B1(n3728), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2134 ( .A1(n4764), .A2(n3552), .B1(n3722), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2135 ( .A1(n4762), .A2(n3552), .B1(n3716), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2136 ( .A1(n4760), .A2(n3552), .B1(n3539), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2137 ( .A1(n4758), .A2(n3552), .B1(n3531), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2138 ( .A1(n4756), .A2(n3552), .B1(n3523), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2139 ( .A1(n4754), .A2(n3552), .B1(n3861), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2140 ( .A1(n4752), .A2(n3552), .B1(n3707), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2141 ( .A1(n4750), .A2(n3552), .B1(n3699), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2142 ( .A1(n4748), .A2(n3552), .B1(n3691), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2143 ( .A1(n4746), .A2(n3552), .B1(n3683), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2144 ( .A1(n4744), .A2(n3552), .B1(n3675), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2145 ( .A1(n4742), .A2(n3552), .B1(n3511), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2146 ( .A1(n4740), .A2(n3552), .B1(n3503), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2147 ( .A1(n4738), .A2(n3552), .B1(n3673), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2148 ( .A1(n4736), .A2(n3552), .B1(n3665), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2149 ( .A1(n4734), .A2(n3552), .B1(n3657), .B2(n4627), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2150 ( .A1(n4732), .A2(n3552), .B1(n3649), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2151 ( .A1(n4730), .A2(n3552), .B1(n3856), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2152 ( .A1(n4728), .A2(n3552), .B1(n3852), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2153 ( .A1(n4726), .A2(n3552), .B1(n3573), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2154 ( .A1(n4724), .A2(n3552), .B1(n3568), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2155 ( .A1(n4722), .A2(n3552), .B1(n3563), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2156 ( .A1(n4720), .A2(n3552), .B1(n3844), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2157 ( .A1(n4718), .A2(n3552), .B1(n3840), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2158 ( .A1(n4716), .A2(n3552), .B1(n3836), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2159 ( .A1(n4714), .A2(n3552), .B1(n3832), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2160 ( .A1(n4712), .A2(n3552), .B1(n3828), .B2(n4626), .ZN(
        \REGISTER_FILE_32[18].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2163 ( .A1(n4778), .A2(n3551), .B1(n4083), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2164 ( .A1(n4772), .A2(n3551), .B1(n4082), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2165 ( .A1(n4770), .A2(n3551), .B1(n4081), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2166 ( .A1(n4768), .A2(n3551), .B1(n4080), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2167 ( .A1(n4766), .A2(n3551), .B1(n4079), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2168 ( .A1(n4764), .A2(n3551), .B1(n4078), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2169 ( .A1(n4762), .A2(n3551), .B1(n4077), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2170 ( .A1(n4760), .A2(n3551), .B1(n4076), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2171 ( .A1(n4758), .A2(n3551), .B1(n4075), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2172 ( .A1(n4756), .A2(n3551), .B1(n4074), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2173 ( .A1(n4754), .A2(n3551), .B1(n4508), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2174 ( .A1(n4752), .A2(n3551), .B1(n4073), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2175 ( .A1(n4750), .A2(n3551), .B1(n4072), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2176 ( .A1(n4748), .A2(n3551), .B1(n4071), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2177 ( .A1(n4746), .A2(n3551), .B1(n4070), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2178 ( .A1(n4744), .A2(n3551), .B1(n4069), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2179 ( .A1(n4742), .A2(n3551), .B1(n4068), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2180 ( .A1(n4740), .A2(n3551), .B1(n4067), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2181 ( .A1(n4738), .A2(n3551), .B1(n4066), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2182 ( .A1(n4736), .A2(n3551), .B1(n4065), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2183 ( .A1(n4734), .A2(n3551), .B1(n4064), .B2(n4625), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2184 ( .A1(n4732), .A2(n3551), .B1(n4063), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2185 ( .A1(n4730), .A2(n3551), .B1(n4507), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2186 ( .A1(n4728), .A2(n3551), .B1(n4506), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2187 ( .A1(n4726), .A2(n3551), .B1(n4505), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2188 ( .A1(n4724), .A2(n3551), .B1(n4504), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2189 ( .A1(n4722), .A2(n3551), .B1(n4503), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2190 ( .A1(n4720), .A2(n3551), .B1(n4502), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2191 ( .A1(n4718), .A2(n3551), .B1(n4501), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2192 ( .A1(n4716), .A2(n3551), .B1(n4500), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2193 ( .A1(n4714), .A2(n3551), .B1(n4499), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2194 ( .A1(n4712), .A2(n3551), .B1(n4498), .B2(n4624), .ZN(
        \REGISTER_FILE_32[17].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2197 ( .A1(n4778), .A2(n3550), .B1(n3775), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2198 ( .A1(n4772), .A2(n3550), .B1(n3767), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2199 ( .A1(n4770), .A2(n3550), .B1(n4015), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2200 ( .A1(n4768), .A2(n3550), .B1(n4009), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2201 ( .A1(n4766), .A2(n3550), .B1(n4003), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2202 ( .A1(n4764), .A2(n3550), .B1(n3997), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2203 ( .A1(n4762), .A2(n3550), .B1(n3991), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2204 ( .A1(n4760), .A2(n3550), .B1(n3616), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2205 ( .A1(n4758), .A2(n3550), .B1(n3608), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2206 ( .A1(n4756), .A2(n3550), .B1(n3600), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2207 ( .A1(n4754), .A2(n3550), .B1(n4484), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2208 ( .A1(n4752), .A2(n3550), .B1(n3981), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2209 ( .A1(n4750), .A2(n3550), .B1(n3973), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2210 ( .A1(n4748), .A2(n3550), .B1(n3965), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2211 ( .A1(n4746), .A2(n3550), .B1(n3957), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2212 ( .A1(n4744), .A2(n3550), .B1(n3949), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2213 ( .A1(n4742), .A2(n3550), .B1(n3941), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2214 ( .A1(n4740), .A2(n3550), .B1(n3933), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2215 ( .A1(n4738), .A2(n3550), .B1(n3925), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2216 ( .A1(n4736), .A2(n3550), .B1(n3917), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2217 ( .A1(n4734), .A2(n3550), .B1(n3909), .B2(n4623), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2218 ( .A1(n4732), .A2(n3550), .B1(n3901), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2219 ( .A1(n4730), .A2(n3550), .B1(n4478), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2220 ( .A1(n4728), .A2(n3550), .B1(n4472), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2221 ( .A1(n4726), .A2(n3550), .B1(n3890), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2222 ( .A1(n4724), .A2(n3550), .B1(n3885), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2223 ( .A1(n4722), .A2(n3550), .B1(n3880), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2224 ( .A1(n4720), .A2(n3550), .B1(n4465), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2225 ( .A1(n4718), .A2(n3550), .B1(n4459), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2226 ( .A1(n4716), .A2(n3550), .B1(n4453), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2227 ( .A1(n4714), .A2(n3550), .B1(n4447), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2228 ( .A1(n4712), .A2(n3550), .B1(n4441), .B2(n4622), .ZN(
        \REGISTER_FILE_32[16].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  AND3_X2 U2231 ( .A1(n3447), .A2(n1026), .A3(rd[0]), .ZN(n3461) );
  OAI22_X2 U2232 ( .A1(n4778), .A2(n3549), .B1(n4259), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2233 ( .A1(n4772), .A2(n3549), .B1(n4258), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2234 ( .A1(n4770), .A2(n3549), .B1(n4257), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2235 ( .A1(n4768), .A2(n3549), .B1(n4256), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2236 ( .A1(n4766), .A2(n3549), .B1(n4255), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2237 ( .A1(n4764), .A2(n3549), .B1(n4254), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2238 ( .A1(n4762), .A2(n3549), .B1(n4253), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2239 ( .A1(n4760), .A2(n3549), .B1(n4252), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2240 ( .A1(n4758), .A2(n3549), .B1(n4251), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2241 ( .A1(n4756), .A2(n3549), .B1(n4250), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2242 ( .A1(n4754), .A2(n3549), .B1(n4574), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2243 ( .A1(n4752), .A2(n3549), .B1(n4249), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2244 ( .A1(n4750), .A2(n3549), .B1(n4248), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2245 ( .A1(n4748), .A2(n3549), .B1(n4247), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2246 ( .A1(n4746), .A2(n3549), .B1(n4246), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2247 ( .A1(n4744), .A2(n3549), .B1(n4245), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2248 ( .A1(n4742), .A2(n3549), .B1(n4244), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2249 ( .A1(n4740), .A2(n3549), .B1(n4243), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2250 ( .A1(n4738), .A2(n3549), .B1(n4242), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2251 ( .A1(n4736), .A2(n3549), .B1(n4241), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2252 ( .A1(n4734), .A2(n3549), .B1(n4240), .B2(n4621), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2253 ( .A1(n4732), .A2(n3549), .B1(n4239), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2254 ( .A1(n4730), .A2(n3549), .B1(n4573), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2255 ( .A1(n4728), .A2(n3549), .B1(n4572), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2256 ( .A1(n4726), .A2(n3549), .B1(n4571), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2257 ( .A1(n4724), .A2(n3549), .B1(n4570), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2258 ( .A1(n4722), .A2(n3549), .B1(n4569), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2259 ( .A1(n4720), .A2(n3549), .B1(n4568), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2260 ( .A1(n4718), .A2(n3549), .B1(n4567), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2261 ( .A1(n4716), .A2(n3549), .B1(n4566), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2262 ( .A1(n4714), .A2(n3549), .B1(n4565), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2263 ( .A1(n4712), .A2(n3549), .B1(n4564), .B2(n4620), .ZN(
        \REGISTER_FILE_32[15].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2266 ( .A1(n4778), .A2(n3548), .B1(n3591), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2267 ( .A1(n4772), .A2(n3548), .B1(n3583), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2268 ( .A1(n4770), .A2(n3548), .B1(n3739), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2269 ( .A1(n4768), .A2(n3548), .B1(n3733), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2270 ( .A1(n4766), .A2(n3548), .B1(n3727), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2271 ( .A1(n4764), .A2(n3548), .B1(n3721), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2272 ( .A1(n4762), .A2(n3548), .B1(n3715), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2273 ( .A1(n4760), .A2(n3548), .B1(n3538), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2274 ( .A1(n4758), .A2(n3548), .B1(n3530), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2275 ( .A1(n4756), .A2(n3548), .B1(n3522), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2276 ( .A1(n4754), .A2(n3548), .B1(n3860), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2277 ( .A1(n4752), .A2(n3548), .B1(n3706), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2278 ( .A1(n4750), .A2(n3548), .B1(n3698), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2279 ( .A1(n4748), .A2(n3548), .B1(n3690), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2280 ( .A1(n4746), .A2(n3548), .B1(n3682), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2281 ( .A1(n4744), .A2(n3548), .B1(n3518), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2282 ( .A1(n4742), .A2(n3548), .B1(n3510), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2283 ( .A1(n4740), .A2(n3548), .B1(n3502), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2284 ( .A1(n4738), .A2(n3548), .B1(n3672), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2285 ( .A1(n4736), .A2(n3548), .B1(n3664), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2286 ( .A1(n4734), .A2(n3548), .B1(n3656), .B2(n4619), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2287 ( .A1(n4732), .A2(n3548), .B1(n3648), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2288 ( .A1(n4730), .A2(n3548), .B1(n3855), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2289 ( .A1(n4728), .A2(n3548), .B1(n3851), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2290 ( .A1(n4726), .A2(n3548), .B1(n3572), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2291 ( .A1(n4724), .A2(n3548), .B1(n3567), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2292 ( .A1(n4722), .A2(n3548), .B1(n3847), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2293 ( .A1(n4720), .A2(n3548), .B1(n3843), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2294 ( .A1(n4718), .A2(n3548), .B1(n3839), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2295 ( .A1(n4716), .A2(n3548), .B1(n3835), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2296 ( .A1(n4714), .A2(n3548), .B1(n3831), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2297 ( .A1(n4712), .A2(n3548), .B1(n3827), .B2(n4618), .ZN(
        \REGISTER_FILE_32[14].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2300 ( .A1(n4778), .A2(n3547), .B1(n4062), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2301 ( .A1(n4772), .A2(n3547), .B1(n4061), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2302 ( .A1(n4770), .A2(n3547), .B1(n4060), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2303 ( .A1(n4768), .A2(n3547), .B1(n4059), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2304 ( .A1(n4766), .A2(n3547), .B1(n4058), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2305 ( .A1(n4764), .A2(n3547), .B1(n4057), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2306 ( .A1(n4762), .A2(n3547), .B1(n4056), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2307 ( .A1(n4760), .A2(n3547), .B1(n4055), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2308 ( .A1(n4758), .A2(n3547), .B1(n4054), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2309 ( .A1(n4756), .A2(n3547), .B1(n4053), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2310 ( .A1(n4754), .A2(n3547), .B1(n4497), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2311 ( .A1(n4752), .A2(n3547), .B1(n4052), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2312 ( .A1(n4750), .A2(n3547), .B1(n4051), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2313 ( .A1(n4748), .A2(n3547), .B1(n4050), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2314 ( .A1(n4746), .A2(n3547), .B1(n4049), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2315 ( .A1(n4744), .A2(n3547), .B1(n4048), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2316 ( .A1(n4742), .A2(n3547), .B1(n4047), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2317 ( .A1(n4740), .A2(n3547), .B1(n4046), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2318 ( .A1(n4738), .A2(n3547), .B1(n4045), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2319 ( .A1(n4736), .A2(n3547), .B1(n4044), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2320 ( .A1(n4734), .A2(n3547), .B1(n4043), .B2(n4617), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2321 ( .A1(n4732), .A2(n3547), .B1(n4042), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2322 ( .A1(n4730), .A2(n3547), .B1(n4496), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2323 ( .A1(n4728), .A2(n3547), .B1(n4495), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2324 ( .A1(n4726), .A2(n3547), .B1(n4494), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2325 ( .A1(n4724), .A2(n3547), .B1(n4493), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2326 ( .A1(n4722), .A2(n3547), .B1(n4492), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2327 ( .A1(n4720), .A2(n3547), .B1(n4491), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2328 ( .A1(n4718), .A2(n3547), .B1(n4490), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2329 ( .A1(n4716), .A2(n3547), .B1(n4489), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2330 ( .A1(n4714), .A2(n3547), .B1(n4488), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2331 ( .A1(n4712), .A2(n3547), .B1(n4487), .B2(n4616), .ZN(
        \REGISTER_FILE_32[13].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2335 ( .A1(n4778), .A2(n3546), .B1(n3774), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2336 ( .A1(n4772), .A2(n3546), .B1(n3766), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2337 ( .A1(n4770), .A2(n3546), .B1(n4014), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2338 ( .A1(n4768), .A2(n3546), .B1(n4008), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2339 ( .A1(n4766), .A2(n3546), .B1(n4002), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2340 ( .A1(n4764), .A2(n3546), .B1(n3996), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2341 ( .A1(n4762), .A2(n3546), .B1(n3990), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2342 ( .A1(n4760), .A2(n3546), .B1(n3615), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2343 ( .A1(n4758), .A2(n3546), .B1(n3607), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2344 ( .A1(n4756), .A2(n3546), .B1(n3599), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2345 ( .A1(n4754), .A2(n3546), .B1(n4483), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2346 ( .A1(n4752), .A2(n3546), .B1(n3980), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2347 ( .A1(n4750), .A2(n3546), .B1(n3972), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2348 ( .A1(n4748), .A2(n3546), .B1(n3964), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2349 ( .A1(n4746), .A2(n3546), .B1(n3956), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2350 ( .A1(n4744), .A2(n3546), .B1(n3948), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2351 ( .A1(n4742), .A2(n3546), .B1(n3940), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2352 ( .A1(n4740), .A2(n3546), .B1(n3932), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2353 ( .A1(n4738), .A2(n3546), .B1(n3924), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2354 ( .A1(n4736), .A2(n3546), .B1(n3916), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2355 ( .A1(n4734), .A2(n3546), .B1(n3908), .B2(n4615), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2356 ( .A1(n4732), .A2(n3546), .B1(n3900), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2357 ( .A1(n4730), .A2(n3546), .B1(n4477), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2358 ( .A1(n4728), .A2(n3546), .B1(n4471), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2359 ( .A1(n4726), .A2(n3546), .B1(n3889), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2360 ( .A1(n4724), .A2(n3546), .B1(n3884), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2361 ( .A1(n4722), .A2(n3546), .B1(n4470), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2362 ( .A1(n4720), .A2(n3546), .B1(n4464), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2363 ( .A1(n4718), .A2(n3546), .B1(n4458), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2364 ( .A1(n4716), .A2(n3546), .B1(n4452), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2365 ( .A1(n4714), .A2(n3546), .B1(n4446), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2366 ( .A1(n4712), .A2(n3546), .B1(n4440), .B2(n4614), .ZN(
        \REGISTER_FILE_32[12].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  AND3_X2 U2369 ( .A1(rd[1]), .A2(n1025), .A3(n3423), .ZN(n3470) );
  AND2_X2 U2370 ( .A1(rd[2]), .A2(writeEnable), .ZN(n3423) );
  OAI22_X2 U2371 ( .A1(n4778), .A2(n3545), .B1(n4238), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2372 ( .A1(n4772), .A2(n3545), .B1(n4237), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2373 ( .A1(n4770), .A2(n3545), .B1(n4236), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2374 ( .A1(n4768), .A2(n3545), .B1(n4235), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2375 ( .A1(n4766), .A2(n3545), .B1(n4234), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2376 ( .A1(n4764), .A2(n3545), .B1(n4233), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2377 ( .A1(n4762), .A2(n3545), .B1(n4232), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2378 ( .A1(n4760), .A2(n3545), .B1(n4231), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2379 ( .A1(n4758), .A2(n3545), .B1(n4230), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2380 ( .A1(n4756), .A2(n3545), .B1(n4229), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2381 ( .A1(n4754), .A2(n3545), .B1(n4563), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2382 ( .A1(n4752), .A2(n3545), .B1(n4228), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2383 ( .A1(n4750), .A2(n3545), .B1(n4227), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2384 ( .A1(n4748), .A2(n3545), .B1(n4226), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2385 ( .A1(n4746), .A2(n3545), .B1(n4225), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2386 ( .A1(n4744), .A2(n3545), .B1(n4224), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2387 ( .A1(n4742), .A2(n3545), .B1(n4223), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2388 ( .A1(n4740), .A2(n3545), .B1(n4222), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2389 ( .A1(n4738), .A2(n3545), .B1(n4221), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2390 ( .A1(n4736), .A2(n3545), .B1(n4220), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2391 ( .A1(n4734), .A2(n3545), .B1(n4219), .B2(n4613), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2392 ( .A1(n4732), .A2(n3545), .B1(n4218), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2393 ( .A1(n4730), .A2(n3545), .B1(n4562), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2394 ( .A1(n4728), .A2(n3545), .B1(n4561), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2395 ( .A1(n4726), .A2(n3545), .B1(n4560), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2396 ( .A1(n4724), .A2(n3545), .B1(n4559), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2397 ( .A1(n4722), .A2(n3545), .B1(n4558), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2398 ( .A1(n4720), .A2(n3545), .B1(n4557), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2399 ( .A1(n4718), .A2(n3545), .B1(n4556), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2400 ( .A1(n4716), .A2(n3545), .B1(n4555), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2401 ( .A1(n4714), .A2(n3545), .B1(n4554), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2402 ( .A1(n4712), .A2(n3545), .B1(n4553), .B2(n4612), .ZN(
        \REGISTER_FILE_32[11].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  AND2_X2 U2405 ( .A1(rd[3]), .A2(rd[4]), .ZN(n3415) );
  OAI22_X2 U2406 ( .A1(n4778), .A2(n3544), .B1(n3590), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2407 ( .A1(n4772), .A2(n3544), .B1(n3582), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2408 ( .A1(n4770), .A2(n3544), .B1(n3868), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2409 ( .A1(n4768), .A2(n3544), .B1(n3867), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2410 ( .A1(n4766), .A2(n3544), .B1(n3866), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2411 ( .A1(n4764), .A2(n3544), .B1(n3865), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2412 ( .A1(n4762), .A2(n3544), .B1(n3864), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2413 ( .A1(n4760), .A2(n3544), .B1(n3537), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2414 ( .A1(n4758), .A2(n3544), .B1(n3529), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2415 ( .A1(n4756), .A2(n3544), .B1(n3521), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2416 ( .A1(n4754), .A2(n3544), .B1(n4437), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2417 ( .A1(n4752), .A2(n3544), .B1(n3705), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2418 ( .A1(n4750), .A2(n3544), .B1(n3697), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2419 ( .A1(n4748), .A2(n3544), .B1(n3689), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2420 ( .A1(n4746), .A2(n3544), .B1(n3681), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2421 ( .A1(n4744), .A2(n3544), .B1(n3517), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2422 ( .A1(n4742), .A2(n3544), .B1(n3509), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2423 ( .A1(n4740), .A2(n3544), .B1(n3501), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2424 ( .A1(n4738), .A2(n3544), .B1(n3671), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2425 ( .A1(n4736), .A2(n3544), .B1(n3663), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2426 ( .A1(n4734), .A2(n3544), .B1(n3655), .B2(n4611), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2427 ( .A1(n4732), .A2(n3544), .B1(n3647), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2428 ( .A1(n4730), .A2(n3544), .B1(n4436), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2429 ( .A1(n4728), .A2(n3544), .B1(n4435), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2430 ( .A1(n4726), .A2(n3544), .B1(n3571), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2431 ( .A1(n4724), .A2(n3544), .B1(n3566), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2432 ( .A1(n4722), .A2(n3544), .B1(n4434), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2433 ( .A1(n4720), .A2(n3544), .B1(n4433), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2434 ( .A1(n4718), .A2(n3544), .B1(n4432), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2435 ( .A1(n4716), .A2(n3544), .B1(n4431), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2436 ( .A1(n4714), .A2(n3544), .B1(n4430), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2437 ( .A1(n4712), .A2(n3544), .B1(n4429), .B2(n4610), .ZN(
        \REGISTER_FILE_32[10].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  AND3_X2 U2440 ( .A1(n3447), .A2(n1025), .A3(rd[1]), .ZN(n3407) );
  AND2_X2 U2441 ( .A1(rd[3]), .A2(n1027), .ZN(n3418) );
  OAI22_X2 U2442 ( .A1(n4778), .A2(n3543), .B1(n3777), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U2444 ( .A1(n4772), .A2(n3543), .B1(n3769), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 )
         );
  NAND2_X2 U2445 ( .A1(busW[8]), .A2(reset), .ZN(n3376) );
  OAI22_X2 U2446 ( .A1(n4770), .A2(n3543), .B1(n4017), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 )
         );
  NAND2_X2 U2447 ( .A1(busW[7]), .A2(n4911), .ZN(n3377) );
  OAI22_X2 U2448 ( .A1(n4768), .A2(n3543), .B1(n4011), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 )
         );
  NAND2_X2 U2449 ( .A1(busW[6]), .A2(reset), .ZN(n3378) );
  OAI22_X2 U2450 ( .A1(n4766), .A2(n3543), .B1(n4005), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 )
         );
  NAND2_X2 U2451 ( .A1(busW[5]), .A2(n4911), .ZN(n3379) );
  OAI22_X2 U2452 ( .A1(n4764), .A2(n3543), .B1(n3999), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 )
         );
  NAND2_X2 U2453 ( .A1(busW[4]), .A2(reset), .ZN(n3380) );
  OAI22_X2 U2454 ( .A1(n4762), .A2(n3543), .B1(n3993), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 )
         );
  NAND2_X2 U2455 ( .A1(busW[3]), .A2(n4911), .ZN(n3381) );
  OAI22_X2 U2456 ( .A1(n4760), .A2(n3543), .B1(n3987), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U2457 ( .A1(busW[31]), .A2(reset), .ZN(n3382) );
  OAI22_X2 U2458 ( .A1(n4758), .A2(n3543), .B1(n3610), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2460 ( .A1(n4756), .A2(n3543), .B1(n3602), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U2462 ( .A1(n4754), .A2(n3543), .B1(n4486), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2464 ( .A1(n4752), .A2(n3543), .B1(n3983), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2466 ( .A1(n4750), .A2(n3543), .B1(n3975), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2468 ( .A1(n4748), .A2(n3543), .B1(n3967), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2470 ( .A1(n4746), .A2(n3543), .B1(n3959), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2472 ( .A1(n4744), .A2(n3543), .B1(n3951), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2474 ( .A1(n4742), .A2(n3543), .B1(n3943), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2476 ( .A1(n4740), .A2(n3543), .B1(n3935), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2478 ( .A1(n4738), .A2(n3543), .B1(n3927), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2480 ( .A1(n4736), .A2(n3543), .B1(n3919), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2482 ( .A1(n4734), .A2(n3543), .B1(n3911), .B2(n4609), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 )
         );
  OAI22_X2 U2484 ( .A1(n4732), .A2(n3543), .B1(n3903), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2486 ( .A1(n4730), .A2(n3543), .B1(n4480), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2488 ( .A1(n4728), .A2(n3543), .B1(n4474), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2490 ( .A1(n4726), .A2(n3543), .B1(n3891), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2492 ( .A1(n4724), .A2(n3543), .B1(n3886), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2494 ( .A1(n4722), .A2(n3543), .B1(n3881), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2496 ( .A1(n4720), .A2(n3543), .B1(n4467), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2498 ( .A1(n4718), .A2(n3543), .B1(n4461), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2500 ( .A1(n4716), .A2(n3543), .B1(n4455), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2502 ( .A1(n4714), .A2(n3543), .B1(n4449), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U2504 ( .A1(n4712), .A2(n3543), .B1(n4443), .B2(n4608), .ZN(
        \REGISTER_FILE_32[0].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 )
         );
  AND3_X2 U2508 ( .A1(n1025), .A2(n1026), .A3(n3447), .ZN(n3426) );
  INV_X4 U2511 ( .A(rd[0]), .ZN(n1025) );
  INV_X4 U2512 ( .A(rd[1]), .ZN(n1026) );
  INV_X4 U2513 ( .A(rd[4]), .ZN(n1027) );
  INV_X4 U2514 ( .A(ra[0]), .ZN(n1028) );
  INV_X4 U2515 ( .A(ra[1]), .ZN(n1029) );
  INV_X4 U2516 ( .A(ra[2]), .ZN(n1030) );
  INV_X4 U2517 ( .A(ra[3]), .ZN(n1031) );
  INV_X4 U2518 ( .A(rb[0]), .ZN(n1032) );
  INV_X4 U2519 ( .A(rb[1]), .ZN(n1033) );
  INV_X4 U2520 ( .A(rb[2]), .ZN(n1034) );
  INV_X4 U2521 ( .A(rb[3]), .ZN(n1035) );
  INV_X4 U2522 ( .A(writeEnable), .ZN(n1036) );
  OAI21_X2 U3547 ( .B1(n2217), .B2(n2218), .A(n4907), .ZN(n2216) );
  OAI21_X2 U3548 ( .B1(n2237), .B2(n2238), .A(n4907), .ZN(n2236) );
  OAI21_X2 U3549 ( .B1(n2277), .B2(n2278), .A(n4907), .ZN(n2276) );
  OAI21_X2 U3550 ( .B1(n2297), .B2(n2298), .A(n4907), .ZN(n2296) );
  OAI21_X2 U3551 ( .B1(n2317), .B2(n2318), .A(n4908), .ZN(n2316) );
  OAI21_X2 U3552 ( .B1(n2337), .B2(n2338), .A(n4908), .ZN(n2336) );
  OAI21_X2 U3553 ( .B1(n2357), .B2(n2358), .A(n4908), .ZN(n2356) );
  OAI21_X2 U3554 ( .B1(n2385), .B2(n2386), .A(n4849), .ZN(n2374) );
  OAI21_X2 U3555 ( .B1(n2397), .B2(n2398), .A(n4908), .ZN(n2396) );
  OAI21_X2 U3556 ( .B1(n2417), .B2(n2418), .A(n4908), .ZN(n2416) );
  OAI21_X2 U3557 ( .B1(n2437), .B2(n2438), .A(n4908), .ZN(n2436) );
  OAI21_X2 U3558 ( .B1(n2457), .B2(n2458), .A(n4908), .ZN(n2456) );
  OAI21_X2 U3559 ( .B1(n2497), .B2(n2498), .A(n4908), .ZN(n2496) );
  OAI21_X2 U3560 ( .B1(n2517), .B2(n2518), .A(n4908), .ZN(n2516) );
  OAI21_X2 U3561 ( .B1(n2537), .B2(n2538), .A(n4908), .ZN(n2536) );
  OAI21_X2 U3562 ( .B1(n2557), .B2(n2558), .A(n4908), .ZN(n2556) );
  OAI21_X2 U3563 ( .B1(n2577), .B2(n2578), .A(n4907), .ZN(n2576) );
  OAI21_X2 U3564 ( .B1(n2597), .B2(n2598), .A(n4908), .ZN(n2596) );
  OAI21_X2 U3565 ( .B1(n2617), .B2(n2618), .A(n4907), .ZN(n2616) );
  OAI21_X2 U3566 ( .B1(n2637), .B2(n2638), .A(n4908), .ZN(n2636) );
  OAI21_X2 U3567 ( .B1(n2657), .B2(n2658), .A(n4907), .ZN(n2656) );
  OAI21_X2 U3568 ( .B1(n2677), .B2(n2678), .A(n4908), .ZN(n2676) );
  OAI21_X2 U3569 ( .B1(n2065), .B2(n2066), .A(n4907), .ZN(n2064) );
  OAI21_X2 U3570 ( .B1(n2097), .B2(n2098), .A(n4907), .ZN(n2096) );
  OAI21_X2 U3571 ( .B1(n2117), .B2(n2118), .A(n4907), .ZN(n2116) );
  OAI21_X2 U3572 ( .B1(n2137), .B2(n2138), .A(n4907), .ZN(n2136) );
  OAI21_X2 U3573 ( .B1(n2157), .B2(n2158), .A(n4907), .ZN(n2156) );
  OAI21_X2 U3574 ( .B1(n2177), .B2(n2178), .A(n4907), .ZN(n2176) );
  OAI21_X2 U3575 ( .B1(n2197), .B2(n2198), .A(n4907), .ZN(n2196) );
  OAI21_X2 U3576 ( .B1(n2265), .B2(n2266), .A(n4848), .ZN(n2254) );
  OAI21_X2 U3577 ( .B1(n2477), .B2(n2478), .A(n4908), .ZN(n2476) );
  OAI21_X2 U3578 ( .B1(n2697), .B2(n2698), .A(n4907), .ZN(n2696) );
  OAI21_X2 U3579 ( .B1(n2873), .B2(n2874), .A(n4844), .ZN(n2872) );
  OAI21_X2 U3580 ( .B1(n2893), .B2(n2894), .A(n4844), .ZN(n2892) );
  OAI21_X2 U3581 ( .B1(n2933), .B2(n2934), .A(n4844), .ZN(n2932) );
  OAI21_X2 U3582 ( .B1(n2953), .B2(n2954), .A(n4844), .ZN(n2952) );
  OAI21_X2 U3583 ( .B1(n2985), .B2(n2986), .A(n4781), .ZN(n2969) );
  OAI21_X2 U3584 ( .B1(n2993), .B2(n2994), .A(n4845), .ZN(n2992) );
  OAI21_X2 U3585 ( .B1(n3013), .B2(n3014), .A(n4845), .ZN(n3012) );
  OAI21_X2 U3586 ( .B1(n3033), .B2(n3034), .A(n4845), .ZN(n3032) );
  OAI21_X2 U3587 ( .B1(n3053), .B2(n3054), .A(n4845), .ZN(n3052) );
  OAI21_X2 U3588 ( .B1(n3073), .B2(n3074), .A(n4845), .ZN(n3072) );
  OAI21_X2 U3589 ( .B1(n3093), .B2(n3094), .A(n4845), .ZN(n3092) );
  OAI21_X2 U3590 ( .B1(n3113), .B2(n3114), .A(n4845), .ZN(n3112) );
  OAI21_X2 U3591 ( .B1(n3153), .B2(n3154), .A(n4845), .ZN(n3152) );
  OAI21_X2 U3592 ( .B1(n3173), .B2(n3174), .A(n4845), .ZN(n3172) );
  OAI21_X2 U3593 ( .B1(n3205), .B2(n3206), .A(n4781), .ZN(n3189) );
  OAI21_X2 U3594 ( .B1(n3213), .B2(n3214), .A(n4845), .ZN(n3212) );
  OAI21_X2 U3595 ( .B1(n3233), .B2(n3234), .A(n4844), .ZN(n3232) );
  OAI21_X2 U3596 ( .B1(n3253), .B2(n3254), .A(n4845), .ZN(n3252) );
  OAI21_X2 U3597 ( .B1(n3273), .B2(n3274), .A(n4844), .ZN(n3272) );
  OAI21_X2 U3598 ( .B1(n3293), .B2(n3294), .A(n4845), .ZN(n3292) );
  OAI21_X2 U3599 ( .B1(n3313), .B2(n3314), .A(n4844), .ZN(n3312) );
  OAI21_X2 U3600 ( .B1(n3333), .B2(n3334), .A(n4845), .ZN(n3332) );
  OAI21_X2 U3601 ( .B1(n2744), .B2(n2745), .A(n4780), .ZN(n2717) );
  OAI21_X2 U3602 ( .B1(n2761), .B2(n2762), .A(n4782), .ZN(n2750) );
  OAI21_X2 U3603 ( .B1(n2773), .B2(n2774), .A(n4844), .ZN(n2772) );
  OAI21_X2 U3604 ( .B1(n2793), .B2(n2794), .A(n4844), .ZN(n2792) );
  OAI21_X2 U3605 ( .B1(n2813), .B2(n2814), .A(n4844), .ZN(n2812) );
  OAI21_X2 U3606 ( .B1(n2833), .B2(n2834), .A(n4844), .ZN(n2832) );
  OAI21_X2 U3607 ( .B1(n2853), .B2(n2854), .A(n4844), .ZN(n2852) );
  OAI21_X2 U3608 ( .B1(n2925), .B2(n2926), .A(n4780), .ZN(n2909) );
  OAI21_X2 U3609 ( .B1(n3133), .B2(n3134), .A(n4845), .ZN(n3132) );
  OAI21_X2 U3610 ( .B1(n3357), .B2(n3358), .A(n4784), .ZN(n3351) );
  NOR2_X2 U3611 ( .A1(rb[3]), .A2(rb[4]), .ZN(n2715) );
  NOR2_X2 U3612 ( .A1(n1035), .A2(rb[4]), .ZN(n2714) );
  NOR2_X2 U3613 ( .A1(n1031), .A2(ra[4]), .ZN(n3370) );
  NOR2_X2 U3614 ( .A1(ra[3]), .A2(ra[4]), .ZN(n3371) );
  NOR2_X2 U3615 ( .A1(n1036), .A2(rd[2]), .ZN(n3447) );
  NOR2_X2 U3616 ( .A1(n1027), .A2(rd[3]), .ZN(n3408) );
  NOR2_X2 U3617 ( .A1(rd[3]), .A2(rd[4]), .ZN(n3411) );
  OAI21_X2 U3618 ( .B1(n2229), .B2(n2230), .A(n4846), .ZN(n2213) );
  OAI21_X2 U3619 ( .B1(n2225), .B2(n2226), .A(n4848), .ZN(n2214) );
  OAI21_X2 U3620 ( .B1(n2221), .B2(n2222), .A(n4850), .ZN(n2215) );
  OAI21_X2 U3621 ( .B1(n2249), .B2(n2250), .A(n4846), .ZN(n2233) );
  OAI21_X2 U3622 ( .B1(n2245), .B2(n2246), .A(n4848), .ZN(n2234) );
  OAI21_X2 U3623 ( .B1(n2241), .B2(n2242), .A(n4850), .ZN(n2235) );
  OAI21_X2 U3624 ( .B1(n2289), .B2(n2290), .A(n4846), .ZN(n2273) );
  OAI21_X2 U3625 ( .B1(n2285), .B2(n2286), .A(n4848), .ZN(n2274) );
  OAI21_X2 U3626 ( .B1(n2281), .B2(n2282), .A(n4850), .ZN(n2275) );
  OAI21_X2 U3627 ( .B1(n2309), .B2(n2310), .A(n4846), .ZN(n2293) );
  OAI21_X2 U3628 ( .B1(n2305), .B2(n2306), .A(n4848), .ZN(n2294) );
  OAI21_X2 U3629 ( .B1(n2301), .B2(n2302), .A(n4850), .ZN(n2295) );
  OAI21_X2 U3630 ( .B1(n2329), .B2(n2330), .A(n4847), .ZN(n2313) );
  OAI21_X2 U3631 ( .B1(n2325), .B2(n2326), .A(n4849), .ZN(n2314) );
  OAI21_X2 U3632 ( .B1(n2321), .B2(n2322), .A(n4851), .ZN(n2315) );
  OAI21_X2 U3633 ( .B1(n2349), .B2(n2350), .A(n4847), .ZN(n2333) );
  OAI21_X2 U3634 ( .B1(n2345), .B2(n2346), .A(n4849), .ZN(n2334) );
  OAI21_X2 U3635 ( .B1(n2341), .B2(n2342), .A(n4851), .ZN(n2335) );
  OAI21_X2 U3636 ( .B1(n2369), .B2(n2370), .A(n4847), .ZN(n2353) );
  OAI21_X2 U3637 ( .B1(n2365), .B2(n2366), .A(n4849), .ZN(n2354) );
  OAI21_X2 U3638 ( .B1(n2361), .B2(n2362), .A(n4851), .ZN(n2355) );
  OAI21_X2 U3639 ( .B1(n2389), .B2(n2390), .A(n4847), .ZN(n2373) );
  OAI21_X2 U3640 ( .B1(n2381), .B2(n2382), .A(n4851), .ZN(n2375) );
  OAI21_X2 U3641 ( .B1(n2377), .B2(n2378), .A(n4908), .ZN(n2376) );
  OAI21_X2 U3642 ( .B1(n2409), .B2(n2410), .A(n4847), .ZN(n2393) );
  OAI21_X2 U3643 ( .B1(n2405), .B2(n2406), .A(n4849), .ZN(n2394) );
  OAI21_X2 U3644 ( .B1(n2401), .B2(n2402), .A(n4851), .ZN(n2395) );
  OAI21_X2 U3645 ( .B1(n2429), .B2(n2430), .A(n4847), .ZN(n2413) );
  OAI21_X2 U3646 ( .B1(n2425), .B2(n2426), .A(n4849), .ZN(n2414) );
  OAI21_X2 U3647 ( .B1(n2421), .B2(n2422), .A(n4851), .ZN(n2415) );
  OAI21_X2 U3648 ( .B1(n2449), .B2(n2450), .A(n4847), .ZN(n2433) );
  OAI21_X2 U3649 ( .B1(n2445), .B2(n2446), .A(n4849), .ZN(n2434) );
  OAI21_X2 U3650 ( .B1(n2441), .B2(n2442), .A(n4851), .ZN(n2435) );
  OAI21_X2 U3651 ( .B1(n2469), .B2(n2470), .A(n4847), .ZN(n2453) );
  OAI21_X2 U3652 ( .B1(n2465), .B2(n2466), .A(n4849), .ZN(n2454) );
  OAI21_X2 U3653 ( .B1(n2461), .B2(n2462), .A(n4851), .ZN(n2455) );
  OAI21_X2 U3654 ( .B1(n2509), .B2(n2510), .A(n4847), .ZN(n2493) );
  OAI21_X2 U3655 ( .B1(n2505), .B2(n2506), .A(n4849), .ZN(n2494) );
  OAI21_X2 U3656 ( .B1(n2501), .B2(n2502), .A(n4851), .ZN(n2495) );
  OAI21_X2 U3657 ( .B1(n2529), .B2(n2530), .A(n4847), .ZN(n2513) );
  OAI21_X2 U3658 ( .B1(n2525), .B2(n2526), .A(n4849), .ZN(n2514) );
  OAI21_X2 U3659 ( .B1(n2521), .B2(n2522), .A(n4851), .ZN(n2515) );
  OAI21_X2 U3660 ( .B1(n2549), .B2(n2550), .A(n4847), .ZN(n2533) );
  OAI21_X2 U3661 ( .B1(n2545), .B2(n2546), .A(n4849), .ZN(n2534) );
  OAI21_X2 U3662 ( .B1(n2541), .B2(n2542), .A(n4851), .ZN(n2535) );
  OAI21_X2 U3663 ( .B1(n2569), .B2(n2570), .A(n4847), .ZN(n2553) );
  OAI21_X2 U3664 ( .B1(n2565), .B2(n2566), .A(n4849), .ZN(n2554) );
  OAI21_X2 U3665 ( .B1(n2561), .B2(n2562), .A(n4851), .ZN(n2555) );
  OAI21_X2 U3666 ( .B1(n2589), .B2(n2590), .A(n4846), .ZN(n2573) );
  OAI21_X2 U3667 ( .B1(n2585), .B2(n2586), .A(n4848), .ZN(n2574) );
  OAI21_X2 U3668 ( .B1(n2581), .B2(n2582), .A(n4850), .ZN(n2575) );
  OAI21_X2 U3669 ( .B1(n2609), .B2(n2610), .A(n4847), .ZN(n2593) );
  OAI21_X2 U3670 ( .B1(n2605), .B2(n2606), .A(n4849), .ZN(n2594) );
  OAI21_X2 U3671 ( .B1(n2601), .B2(n2602), .A(n4851), .ZN(n2595) );
  OAI21_X2 U3672 ( .B1(n2629), .B2(n2630), .A(n4846), .ZN(n2613) );
  OAI21_X2 U3673 ( .B1(n2625), .B2(n2626), .A(n4848), .ZN(n2614) );
  OAI21_X2 U3674 ( .B1(n2621), .B2(n2622), .A(n4850), .ZN(n2615) );
  OAI21_X2 U3675 ( .B1(n2649), .B2(n2650), .A(n4847), .ZN(n2633) );
  OAI21_X2 U3676 ( .B1(n2641), .B2(n2642), .A(n4851), .ZN(n2635) );
  OAI21_X2 U3677 ( .B1(n2645), .B2(n2646), .A(n4849), .ZN(n2634) );
  OAI21_X2 U3678 ( .B1(n2669), .B2(n2670), .A(n4846), .ZN(n2653) );
  OAI21_X2 U3679 ( .B1(n2665), .B2(n2666), .A(n4848), .ZN(n2654) );
  OAI21_X2 U3680 ( .B1(n2661), .B2(n2662), .A(n4850), .ZN(n2655) );
  OAI21_X2 U3681 ( .B1(n2689), .B2(n2690), .A(n4847), .ZN(n2673) );
  OAI21_X2 U3682 ( .B1(n2685), .B2(n2686), .A(n4849), .ZN(n2674) );
  OAI21_X2 U3683 ( .B1(n2681), .B2(n2682), .A(n4851), .ZN(n2675) );
  OAI21_X2 U3684 ( .B1(n2088), .B2(n2089), .A(n4846), .ZN(n2061) );
  OAI21_X2 U3685 ( .B1(n2083), .B2(n2084), .A(n4848), .ZN(n2062) );
  OAI21_X2 U3686 ( .B1(n2078), .B2(n2079), .A(n4850), .ZN(n2063) );
  OAI21_X2 U3687 ( .B1(n2109), .B2(n2110), .A(n4846), .ZN(n2093) );
  OAI21_X2 U3688 ( .B1(n2105), .B2(n2106), .A(n4848), .ZN(n2094) );
  OAI21_X2 U3689 ( .B1(n2101), .B2(n2102), .A(n4850), .ZN(n2095) );
  OAI21_X2 U3690 ( .B1(n2129), .B2(n2130), .A(n4846), .ZN(n2113) );
  OAI21_X2 U3691 ( .B1(n2125), .B2(n2126), .A(n4848), .ZN(n2114) );
  OAI21_X2 U3692 ( .B1(n2121), .B2(n2122), .A(n4850), .ZN(n2115) );
  OAI21_X2 U3693 ( .B1(n2149), .B2(n2150), .A(n4846), .ZN(n2133) );
  OAI21_X2 U3694 ( .B1(n2145), .B2(n2146), .A(n4848), .ZN(n2134) );
  OAI21_X2 U3695 ( .B1(n2141), .B2(n2142), .A(n4850), .ZN(n2135) );
  OAI21_X2 U3696 ( .B1(n2169), .B2(n2170), .A(n4846), .ZN(n2153) );
  OAI21_X2 U3697 ( .B1(n2165), .B2(n2166), .A(n4848), .ZN(n2154) );
  OAI21_X2 U3698 ( .B1(n2161), .B2(n2162), .A(n4850), .ZN(n2155) );
  OAI21_X2 U3699 ( .B1(n2189), .B2(n2190), .A(n4846), .ZN(n2173) );
  OAI21_X2 U3700 ( .B1(n2185), .B2(n2186), .A(n4848), .ZN(n2174) );
  OAI21_X2 U3701 ( .B1(n2181), .B2(n2182), .A(n4850), .ZN(n2175) );
  OAI21_X2 U3702 ( .B1(n2209), .B2(n2210), .A(n4846), .ZN(n2193) );
  OAI21_X2 U3703 ( .B1(n2205), .B2(n2206), .A(n4848), .ZN(n2194) );
  OAI21_X2 U3704 ( .B1(n2201), .B2(n2202), .A(n4850), .ZN(n2195) );
  OAI21_X2 U3705 ( .B1(n2269), .B2(n2270), .A(n4846), .ZN(n2253) );
  OAI21_X2 U3706 ( .B1(n2261), .B2(n2262), .A(n4850), .ZN(n2255) );
  OAI21_X2 U3707 ( .B1(n2257), .B2(n2258), .A(n4907), .ZN(n2256) );
  OAI21_X2 U3708 ( .B1(n2489), .B2(n2490), .A(n4847), .ZN(n2473) );
  OAI21_X2 U3709 ( .B1(n2485), .B2(n2486), .A(n4849), .ZN(n2474) );
  OAI21_X2 U3710 ( .B1(n2481), .B2(n2482), .A(n4851), .ZN(n2475) );
  OAI21_X2 U3711 ( .B1(n2709), .B2(n2710), .A(n4846), .ZN(n2693) );
  OAI21_X2 U3712 ( .B1(n2705), .B2(n2706), .A(n4848), .ZN(n2694) );
  OAI21_X2 U3713 ( .B1(n2701), .B2(n2702), .A(n4850), .ZN(n2695) );
  OAI21_X2 U3714 ( .B1(n2885), .B2(n2886), .A(n4780), .ZN(n2869) );
  OAI21_X2 U3715 ( .B1(n2877), .B2(n2878), .A(n4784), .ZN(n2871) );
  OAI21_X2 U3716 ( .B1(n2881), .B2(n2882), .A(n4782), .ZN(n2870) );
  OAI21_X2 U3717 ( .B1(n2905), .B2(n2906), .A(n4780), .ZN(n2889) );
  OAI21_X2 U3718 ( .B1(n2901), .B2(n2902), .A(n4782), .ZN(n2890) );
  OAI21_X2 U3719 ( .B1(n2897), .B2(n2898), .A(n4784), .ZN(n2891) );
  OAI21_X2 U3720 ( .B1(n2945), .B2(n2946), .A(n4780), .ZN(n2929) );
  OAI21_X2 U3721 ( .B1(n2941), .B2(n2942), .A(n4782), .ZN(n2930) );
  OAI21_X2 U3722 ( .B1(n2937), .B2(n2938), .A(n4784), .ZN(n2931) );
  OAI21_X2 U3723 ( .B1(n2965), .B2(n2966), .A(n4780), .ZN(n2949) );
  OAI21_X2 U3724 ( .B1(n2961), .B2(n2962), .A(n4782), .ZN(n2950) );
  OAI21_X2 U3725 ( .B1(n2957), .B2(n2958), .A(n4784), .ZN(n2951) );
  OAI21_X2 U3726 ( .B1(n2981), .B2(n2982), .A(n4783), .ZN(n2970) );
  OAI21_X2 U3727 ( .B1(n2977), .B2(n2978), .A(n4785), .ZN(n2971) );
  OAI21_X2 U3728 ( .B1(n2973), .B2(n2974), .A(n4845), .ZN(n2972) );
  OAI21_X2 U3729 ( .B1(n3005), .B2(n3006), .A(n4781), .ZN(n2989) );
  OAI21_X2 U3730 ( .B1(n3001), .B2(n3002), .A(n4783), .ZN(n2990) );
  OAI21_X2 U3731 ( .B1(n2997), .B2(n2998), .A(n4785), .ZN(n2991) );
  OAI21_X2 U3732 ( .B1(n3025), .B2(n3026), .A(n4781), .ZN(n3009) );
  OAI21_X2 U3733 ( .B1(n3021), .B2(n3022), .A(n4783), .ZN(n3010) );
  OAI21_X2 U3734 ( .B1(n3017), .B2(n3018), .A(n4785), .ZN(n3011) );
  OAI21_X2 U3735 ( .B1(n3045), .B2(n3046), .A(n4781), .ZN(n3029) );
  OAI21_X2 U3736 ( .B1(n3041), .B2(n3042), .A(n4783), .ZN(n3030) );
  OAI21_X2 U3737 ( .B1(n3037), .B2(n3038), .A(n4785), .ZN(n3031) );
  OAI21_X2 U3738 ( .B1(n3065), .B2(n3066), .A(n4781), .ZN(n3049) );
  OAI21_X2 U3739 ( .B1(n3061), .B2(n3062), .A(n4783), .ZN(n3050) );
  OAI21_X2 U3740 ( .B1(n3057), .B2(n3058), .A(n4785), .ZN(n3051) );
  OAI21_X2 U3741 ( .B1(n3085), .B2(n3086), .A(n4781), .ZN(n3069) );
  OAI21_X2 U3742 ( .B1(n3081), .B2(n3082), .A(n4783), .ZN(n3070) );
  OAI21_X2 U3743 ( .B1(n3077), .B2(n3078), .A(n4785), .ZN(n3071) );
  OAI21_X2 U3744 ( .B1(n3105), .B2(n3106), .A(n4781), .ZN(n3089) );
  OAI21_X2 U3745 ( .B1(n3101), .B2(n3102), .A(n4783), .ZN(n3090) );
  OAI21_X2 U3746 ( .B1(n3097), .B2(n3098), .A(n4785), .ZN(n3091) );
  OAI21_X2 U3747 ( .B1(n3125), .B2(n3126), .A(n4781), .ZN(n3109) );
  OAI21_X2 U3748 ( .B1(n3121), .B2(n3122), .A(n4783), .ZN(n3110) );
  OAI21_X2 U3749 ( .B1(n3117), .B2(n3118), .A(n4785), .ZN(n3111) );
  OAI21_X2 U3750 ( .B1(n3165), .B2(n3166), .A(n4781), .ZN(n3149) );
  OAI21_X2 U3751 ( .B1(n3161), .B2(n3162), .A(n4783), .ZN(n3150) );
  OAI21_X2 U3752 ( .B1(n3157), .B2(n3158), .A(n4785), .ZN(n3151) );
  OAI21_X2 U3753 ( .B1(n3185), .B2(n3186), .A(n4781), .ZN(n3169) );
  OAI21_X2 U3754 ( .B1(n3181), .B2(n3182), .A(n4783), .ZN(n3170) );
  OAI21_X2 U3755 ( .B1(n3177), .B2(n3178), .A(n4785), .ZN(n3171) );
  OAI21_X2 U3756 ( .B1(n3201), .B2(n3202), .A(n4783), .ZN(n3190) );
  OAI21_X2 U3757 ( .B1(n3197), .B2(n3198), .A(n4785), .ZN(n3191) );
  OAI21_X2 U3758 ( .B1(n3193), .B2(n3194), .A(n4845), .ZN(n3192) );
  OAI21_X2 U3759 ( .B1(n3225), .B2(n3226), .A(n4781), .ZN(n3209) );
  OAI21_X2 U3760 ( .B1(n3221), .B2(n3222), .A(n4783), .ZN(n3210) );
  OAI21_X2 U3761 ( .B1(n3217), .B2(n3218), .A(n4785), .ZN(n3211) );
  OAI21_X2 U3762 ( .B1(n3245), .B2(n3246), .A(n4780), .ZN(n3229) );
  OAI21_X2 U3763 ( .B1(n3241), .B2(n3242), .A(n4782), .ZN(n3230) );
  OAI21_X2 U3764 ( .B1(n3237), .B2(n3238), .A(n4784), .ZN(n3231) );
  OAI21_X2 U3765 ( .B1(n3265), .B2(n3266), .A(n4781), .ZN(n3249) );
  OAI21_X2 U3766 ( .B1(n3261), .B2(n3262), .A(n4783), .ZN(n3250) );
  OAI21_X2 U3767 ( .B1(n3257), .B2(n3258), .A(n4785), .ZN(n3251) );
  OAI21_X2 U3768 ( .B1(n3285), .B2(n3286), .A(n4780), .ZN(n3269) );
  OAI21_X2 U3769 ( .B1(n3281), .B2(n3282), .A(n4782), .ZN(n3270) );
  OAI21_X2 U3770 ( .B1(n3277), .B2(n3278), .A(n4784), .ZN(n3271) );
  OAI21_X2 U3771 ( .B1(n3305), .B2(n3306), .A(n4781), .ZN(n3289) );
  OAI21_X2 U3772 ( .B1(n3301), .B2(n3302), .A(n4783), .ZN(n3290) );
  OAI21_X2 U3773 ( .B1(n3297), .B2(n3298), .A(n4785), .ZN(n3291) );
  OAI21_X2 U3774 ( .B1(n3325), .B2(n3326), .A(n4780), .ZN(n3309) );
  OAI21_X2 U3775 ( .B1(n3317), .B2(n3318), .A(n4784), .ZN(n3311) );
  OAI21_X2 U3776 ( .B1(n3321), .B2(n3322), .A(n4782), .ZN(n3310) );
  OAI21_X2 U3777 ( .B1(n3345), .B2(n3346), .A(n4781), .ZN(n3329) );
  OAI21_X2 U3778 ( .B1(n3341), .B2(n3342), .A(n4783), .ZN(n3330) );
  OAI21_X2 U3779 ( .B1(n3337), .B2(n3338), .A(n4785), .ZN(n3331) );
  OAI21_X2 U3780 ( .B1(n2739), .B2(n2740), .A(n4782), .ZN(n2718) );
  OAI21_X2 U3781 ( .B1(n2734), .B2(n2735), .A(n4784), .ZN(n2719) );
  OAI21_X2 U3782 ( .B1(n2721), .B2(n2722), .A(n4844), .ZN(n2720) );
  OAI21_X2 U3783 ( .B1(n2757), .B2(n2758), .A(n4784), .ZN(n2751) );
  OAI21_X2 U3784 ( .B1(n2753), .B2(n2754), .A(n4844), .ZN(n2752) );
  OAI21_X2 U3785 ( .B1(n2765), .B2(n2766), .A(n4780), .ZN(n2749) );
  OAI21_X2 U3786 ( .B1(n2785), .B2(n2786), .A(n4780), .ZN(n2769) );
  OAI21_X2 U3787 ( .B1(n2781), .B2(n2782), .A(n4782), .ZN(n2770) );
  OAI21_X2 U3788 ( .B1(n2777), .B2(n2778), .A(n4784), .ZN(n2771) );
  OAI21_X2 U3789 ( .B1(n2805), .B2(n2806), .A(n4780), .ZN(n2789) );
  OAI21_X2 U3790 ( .B1(n2801), .B2(n2802), .A(n4782), .ZN(n2790) );
  OAI21_X2 U3791 ( .B1(n2797), .B2(n2798), .A(n4784), .ZN(n2791) );
  OAI21_X2 U3792 ( .B1(n2825), .B2(n2826), .A(n4780), .ZN(n2809) );
  OAI21_X2 U3793 ( .B1(n2821), .B2(n2822), .A(n4782), .ZN(n2810) );
  OAI21_X2 U3794 ( .B1(n2817), .B2(n2818), .A(n4784), .ZN(n2811) );
  OAI21_X2 U3795 ( .B1(n2845), .B2(n2846), .A(n4780), .ZN(n2829) );
  OAI21_X2 U3796 ( .B1(n2841), .B2(n2842), .A(n4782), .ZN(n2830) );
  OAI21_X2 U3797 ( .B1(n2837), .B2(n2838), .A(n4784), .ZN(n2831) );
  OAI21_X2 U3798 ( .B1(n2865), .B2(n2866), .A(n4780), .ZN(n2849) );
  OAI21_X2 U3799 ( .B1(n2861), .B2(n2862), .A(n4782), .ZN(n2850) );
  OAI21_X2 U3800 ( .B1(n2857), .B2(n2858), .A(n4784), .ZN(n2851) );
  OAI21_X2 U3801 ( .B1(n2921), .B2(n2922), .A(n4782), .ZN(n2910) );
  OAI21_X2 U3802 ( .B1(n2917), .B2(n2918), .A(n4784), .ZN(n2911) );
  OAI21_X2 U3803 ( .B1(n2913), .B2(n2914), .A(n4844), .ZN(n2912) );
  OAI21_X2 U3804 ( .B1(n3145), .B2(n3146), .A(n4781), .ZN(n3129) );
  OAI21_X2 U3805 ( .B1(n3141), .B2(n3142), .A(n4783), .ZN(n3130) );
  OAI21_X2 U3806 ( .B1(n3137), .B2(n3138), .A(n4785), .ZN(n3131) );
  OAI21_X2 U3807 ( .B1(n3365), .B2(n3366), .A(n4780), .ZN(n3349) );
  OAI21_X2 U3808 ( .B1(n3361), .B2(n3362), .A(n4782), .ZN(n3350) );
  OAI21_X2 U3809 ( .B1(n3353), .B2(n3354), .A(n4844), .ZN(n3352) );
  NAND2_X2 U3810 ( .A1(n2713), .A2(n1034), .ZN(n3483) );
  NAND2_X2 U3811 ( .A1(rb[2]), .A2(n2713), .ZN(n3484) );
  AND2_X4 U3812 ( .A1(rb[2]), .A2(n2714), .ZN(n3485) );
  AND2_X4 U3813 ( .A1(ra[2]), .A2(n3370), .ZN(n3486) );
  AND2_X4 U3814 ( .A1(ra[2]), .A2(n3371), .ZN(n3487) );
  AND2_X4 U3815 ( .A1(rb[2]), .A2(n2715), .ZN(n3488) );
  AND2_X4 U3816 ( .A1(n3370), .A2(n1030), .ZN(n3489) );
  AND2_X4 U3817 ( .A1(n3371), .A2(n1030), .ZN(n3490) );
  NAND2_X2 U3818 ( .A1(n3368), .A2(n1030), .ZN(n3491) );
  NAND2_X2 U3819 ( .A1(ra[2]), .A2(n3368), .ZN(n3492) );
  AND2_X4 U3820 ( .A1(n2714), .A2(n1034), .ZN(n3493) );
  NAND2_X2 U3821 ( .A1(n2712), .A2(n1034), .ZN(n3494) );
  AND2_X4 U3822 ( .A1(n2715), .A2(n1034), .ZN(n3495) );
  NAND2_X2 U3823 ( .A1(rb[2]), .A2(n2712), .ZN(n3496) );
  INV_X4 U3824 ( .A(n3483), .ZN(n4860) );
  INV_X4 U3825 ( .A(n3485), .ZN(n4893) );
  INV_X4 U3826 ( .A(n3542), .ZN(n4794) );
  INV_X4 U3827 ( .A(n3541), .ZN(n4823) );
  INV_X4 U3828 ( .A(n3483), .ZN(n4865) );
  INV_X4 U3829 ( .A(n4425), .ZN(n4778) );
  INV_X4 U3830 ( .A(n4425), .ZN(n4779) );
  NAND2_X2 U3831 ( .A1(ra[2]), .A2(n3369), .ZN(n3541) );
  NAND2_X2 U3832 ( .A1(n3369), .A2(n1030), .ZN(n3542) );
  INV_X4 U3833 ( .A(n3490), .ZN(n4814) );
  INV_X4 U3834 ( .A(n3487), .ZN(n4843) );
  INV_X4 U3835 ( .A(n3493), .ZN(n4872) );
  INV_X4 U3836 ( .A(n3485), .ZN(n4899) );
  INV_X4 U3837 ( .A(n3491), .ZN(n4792) );
  INV_X4 U3838 ( .A(n3492), .ZN(n4821) );
  NAND2_X4 U3839 ( .A1(n3426), .A2(n3411), .ZN(n3543) );
  NAND2_X4 U3840 ( .A1(n3418), .A2(n3407), .ZN(n3544) );
  NAND2_X4 U3841 ( .A1(n3415), .A2(n3407), .ZN(n3545) );
  NAND2_X4 U3842 ( .A1(n3470), .A2(n3411), .ZN(n3546) );
  NAND2_X4 U3843 ( .A1(n3470), .A2(n3408), .ZN(n3547) );
  NAND2_X4 U3844 ( .A1(n3470), .A2(n3418), .ZN(n3548) );
  NAND2_X4 U3845 ( .A1(n3470), .A2(n3415), .ZN(n3549) );
  NAND2_X4 U3846 ( .A1(n3461), .A2(n3411), .ZN(n3550) );
  NAND2_X4 U3847 ( .A1(n3461), .A2(n3408), .ZN(n3551) );
  NAND2_X4 U3848 ( .A1(n3461), .A2(n3418), .ZN(n3552) );
  AND2_X4 U3849 ( .A1(n4910), .A2(n3543), .ZN(n3553) );
  AND2_X4 U3850 ( .A1(n4910), .A2(n3544), .ZN(n3554) );
  AND2_X4 U3851 ( .A1(n4910), .A2(n3545), .ZN(n3555) );
  AND2_X4 U3852 ( .A1(n4910), .A2(n3546), .ZN(n3556) );
  AND2_X4 U3853 ( .A1(n4910), .A2(n3547), .ZN(n3557) );
  AND2_X4 U3854 ( .A1(n4910), .A2(n3548), .ZN(n3558) );
  AND2_X4 U3855 ( .A1(n4910), .A2(n3549), .ZN(n3559) );
  AND2_X4 U3856 ( .A1(n4910), .A2(n3550), .ZN(n3560) );
  AND2_X4 U3857 ( .A1(n4910), .A2(n3551), .ZN(n3561) );
  AND2_X4 U3858 ( .A1(n4910), .A2(n3552), .ZN(n3562) );
  INV_X4 U3859 ( .A(n3542), .ZN(n4797) );
  INV_X4 U3860 ( .A(n3541), .ZN(n4826) );
  INV_X4 U3861 ( .A(n3489), .ZN(n4802) );
  INV_X4 U3862 ( .A(n3489), .ZN(n4803) );
  INV_X4 U3863 ( .A(n3486), .ZN(n4831) );
  INV_X4 U3864 ( .A(n3486), .ZN(n4832) );
  INV_X4 U3865 ( .A(n3495), .ZN(n4874) );
  INV_X4 U3866 ( .A(n3495), .ZN(n4875) );
  INV_X4 U3867 ( .A(n3488), .ZN(n4901) );
  INV_X4 U3868 ( .A(n3488), .ZN(n4902) );
  INV_X4 U3869 ( .A(n3496), .ZN(n4882) );
  INV_X4 U3870 ( .A(n3496), .ZN(n4881) );
  INV_X4 U3871 ( .A(n3494), .ZN(n4854) );
  INV_X4 U3872 ( .A(n4428), .ZN(n4776) );
  INV_X4 U3873 ( .A(n4428), .ZN(n4777) );
  INV_X4 U3874 ( .A(n4420), .ZN(n4686) );
  INV_X4 U3875 ( .A(n4420), .ZN(n4687) );
  INV_X4 U3876 ( .A(n4421), .ZN(n4690) );
  INV_X4 U3877 ( .A(n4421), .ZN(n4691) );
  INV_X4 U3878 ( .A(n4422), .ZN(n4706) );
  INV_X4 U3879 ( .A(n4422), .ZN(n4707) );
  INV_X4 U3880 ( .A(n4426), .ZN(n4694) );
  INV_X4 U3881 ( .A(n4426), .ZN(n4695) );
  INV_X4 U3882 ( .A(n4427), .ZN(n4698) );
  INV_X4 U3883 ( .A(n4427), .ZN(n4699) );
  INV_X4 U3884 ( .A(n4417), .ZN(n4710) );
  INV_X4 U3885 ( .A(n4417), .ZN(n4711) );
  INV_X4 U3886 ( .A(n4423), .ZN(n4756) );
  INV_X4 U3887 ( .A(n4423), .ZN(n4757) );
  INV_X4 U3888 ( .A(n4424), .ZN(n4758) );
  INV_X4 U3889 ( .A(n4424), .ZN(n4759) );
  AND2_X4 U3890 ( .A1(n4910), .A2(n3459), .ZN(n3779) );
  AND2_X4 U3891 ( .A1(n4910), .A2(n3457), .ZN(n3780) );
  AND2_X4 U3892 ( .A1(n4910), .A2(n3455), .ZN(n3781) );
  AND2_X4 U3893 ( .A1(n4910), .A2(n3453), .ZN(n3782) );
  AND2_X4 U3894 ( .A1(n4910), .A2(n3451), .ZN(n3783) );
  AND2_X4 U3895 ( .A1(n4910), .A2(n3448), .ZN(n3784) );
  AND2_X4 U3896 ( .A1(n4910), .A2(n3445), .ZN(n3785) );
  AND2_X4 U3897 ( .A1(n4910), .A2(n3443), .ZN(n3786) );
  AND2_X4 U3898 ( .A1(n4910), .A2(n3441), .ZN(n3787) );
  AND2_X4 U3899 ( .A1(n4910), .A2(n3438), .ZN(n3788) );
  AND2_X4 U3900 ( .A1(n4910), .A2(n3436), .ZN(n3789) );
  AND2_X4 U3901 ( .A1(n4909), .A2(n3434), .ZN(n3790) );
  INV_X4 U3902 ( .A(n3542), .ZN(n4798) );
  INV_X4 U3903 ( .A(n3542), .ZN(n4795) );
  INV_X4 U3904 ( .A(n3542), .ZN(n4796) );
  INV_X4 U3905 ( .A(n3541), .ZN(n4827) );
  INV_X4 U3906 ( .A(n3541), .ZN(n4824) );
  INV_X4 U3907 ( .A(n3541), .ZN(n4825) );
  INV_X4 U3908 ( .A(n3489), .ZN(n4805) );
  INV_X4 U3909 ( .A(n3489), .ZN(n4804) );
  INV_X4 U3910 ( .A(n3486), .ZN(n4833) );
  INV_X4 U3911 ( .A(n3486), .ZN(n4834) );
  INV_X4 U3912 ( .A(n3490), .ZN(n4809) );
  INV_X4 U3913 ( .A(n3490), .ZN(n4810) );
  INV_X4 U3914 ( .A(n3487), .ZN(n4838) );
  INV_X4 U3915 ( .A(n3487), .ZN(n4839) );
  INV_X4 U3916 ( .A(n3495), .ZN(n4877) );
  INV_X4 U3917 ( .A(n3495), .ZN(n4876) );
  INV_X4 U3918 ( .A(n3488), .ZN(n4903) );
  INV_X4 U3919 ( .A(n3488), .ZN(n4904) );
  INV_X4 U3920 ( .A(n3493), .ZN(n4867) );
  INV_X4 U3921 ( .A(n3493), .ZN(n4868) );
  INV_X4 U3922 ( .A(n3485), .ZN(n4894) );
  INV_X4 U3923 ( .A(n3485), .ZN(n4895) );
  INV_X4 U3924 ( .A(n3494), .ZN(n4853) );
  INV_X4 U3925 ( .A(n3494), .ZN(n4855) );
  INV_X4 U3926 ( .A(n3494), .ZN(n4856) );
  INV_X4 U3927 ( .A(n3496), .ZN(n4883) );
  INV_X4 U3928 ( .A(n3496), .ZN(n4884) );
  INV_X4 U3929 ( .A(n3491), .ZN(n4788) );
  INV_X4 U3930 ( .A(n3491), .ZN(n4787) );
  INV_X4 U3931 ( .A(n3492), .ZN(n4816) );
  INV_X4 U3932 ( .A(n3492), .ZN(n4817) );
  INV_X4 U3933 ( .A(n3483), .ZN(n4862) );
  INV_X4 U3934 ( .A(n3484), .ZN(n4889) );
  INV_X4 U3935 ( .A(n4418), .ZN(n4679) );
  INV_X4 U3936 ( .A(n4418), .ZN(n4678) );
  INV_X4 U3937 ( .A(n4419), .ZN(n4683) );
  INV_X4 U3938 ( .A(n4419), .ZN(n4682) );
  INV_X4 U3939 ( .A(n4416), .ZN(n4702) );
  INV_X4 U3940 ( .A(n4416), .ZN(n4703) );
  AND2_X4 U3941 ( .A1(busW[10]), .A2(n4909), .ZN(n4020) );
  AND2_X4 U3942 ( .A1(busW[11]), .A2(n4909), .ZN(n4021) );
  AND2_X4 U3943 ( .A1(busW[12]), .A2(n4911), .ZN(n4022) );
  AND2_X4 U3944 ( .A1(busW[13]), .A2(n4909), .ZN(n4023) );
  AND2_X4 U3945 ( .A1(busW[14]), .A2(reset), .ZN(n4024) );
  AND2_X4 U3946 ( .A1(busW[15]), .A2(reset), .ZN(n4025) );
  AND2_X4 U3947 ( .A1(busW[16]), .A2(reset), .ZN(n4026) );
  AND2_X4 U3948 ( .A1(busW[17]), .A2(reset), .ZN(n4027) );
  AND2_X4 U3949 ( .A1(busW[18]), .A2(reset), .ZN(n4028) );
  AND2_X4 U3950 ( .A1(busW[19]), .A2(n4909), .ZN(n4029) );
  AND2_X4 U3951 ( .A1(busW[1]), .A2(n4909), .ZN(n4030) );
  AND2_X4 U3952 ( .A1(busW[20]), .A2(n4909), .ZN(n4031) );
  AND2_X4 U3953 ( .A1(busW[0]), .A2(n4911), .ZN(n4032) );
  AND2_X4 U3954 ( .A1(busW[21]), .A2(n4911), .ZN(n4033) );
  AND2_X4 U3955 ( .A1(busW[22]), .A2(n4911), .ZN(n4034) );
  AND2_X4 U3956 ( .A1(busW[23]), .A2(n4911), .ZN(n4035) );
  AND2_X4 U3957 ( .A1(busW[24]), .A2(n4911), .ZN(n4036) );
  AND2_X4 U3958 ( .A1(busW[25]), .A2(n4911), .ZN(n4037) );
  AND2_X4 U3959 ( .A1(busW[26]), .A2(n4911), .ZN(n4038) );
  AND2_X4 U3960 ( .A1(busW[27]), .A2(n4911), .ZN(n4039) );
  AND2_X4 U3961 ( .A1(busW[28]), .A2(n4911), .ZN(n4040) );
  AND2_X4 U3962 ( .A1(busW[29]), .A2(n4911), .ZN(n4041) );
  AND2_X4 U3963 ( .A1(n4909), .A2(n4679), .ZN(n4398) );
  AND2_X4 U3964 ( .A1(n4909), .A2(n4683), .ZN(n4399) );
  AND2_X4 U3965 ( .A1(n4909), .A2(n4686), .ZN(n4400) );
  AND2_X4 U3966 ( .A1(n4909), .A2(n4690), .ZN(n4401) );
  AND2_X4 U3967 ( .A1(n4909), .A2(n4694), .ZN(n4402) );
  AND2_X4 U3968 ( .A1(n4909), .A2(n4698), .ZN(n4403) );
  AND2_X4 U3969 ( .A1(n4909), .A2(n4702), .ZN(n4404) );
  AND2_X4 U3970 ( .A1(n4909), .A2(n4706), .ZN(n4405) );
  AND2_X4 U3971 ( .A1(n4909), .A2(n4710), .ZN(n4406) );
  AND2_X4 U3972 ( .A1(n4909), .A2(n4776), .ZN(n4407) );
  OR2_X4 U3973 ( .A1(n1029), .A2(n1028), .ZN(n4408) );
  OR2_X4 U3974 ( .A1(n1033), .A2(n1032), .ZN(n4409) );
  OR2_X4 U3975 ( .A1(n1028), .A2(ra[1]), .ZN(n4410) );
  OR2_X4 U3976 ( .A1(n1032), .A2(rb[1]), .ZN(n4411) );
  OR2_X4 U3977 ( .A1(n1029), .A2(ra[0]), .ZN(n4412) );
  OR2_X4 U3978 ( .A1(n1033), .A2(rb[0]), .ZN(n4413) );
  OR2_X4 U3979 ( .A1(ra[0]), .A2(ra[1]), .ZN(n4414) );
  OR2_X4 U3980 ( .A1(rb[0]), .A2(rb[1]), .ZN(n4415) );
  INV_X4 U3981 ( .A(n3382), .ZN(n4761) );
  INV_X4 U3982 ( .A(n4761), .ZN(n4760) );
  INV_X4 U3983 ( .A(n3381), .ZN(n4763) );
  INV_X4 U3984 ( .A(n4763), .ZN(n4762) );
  INV_X4 U3985 ( .A(n3380), .ZN(n4765) );
  INV_X4 U3986 ( .A(n4765), .ZN(n4764) );
  INV_X4 U3987 ( .A(n3379), .ZN(n4767) );
  INV_X4 U3988 ( .A(n4767), .ZN(n4766) );
  INV_X4 U3989 ( .A(n3378), .ZN(n4769) );
  INV_X4 U3990 ( .A(n4769), .ZN(n4768) );
  INV_X4 U3991 ( .A(n3377), .ZN(n4771) );
  INV_X4 U3992 ( .A(n4771), .ZN(n4770) );
  INV_X4 U3993 ( .A(n3376), .ZN(n4773) );
  INV_X4 U3994 ( .A(n4773), .ZN(n4772) );
  INV_X4 U3995 ( .A(n3490), .ZN(n4811) );
  INV_X4 U3996 ( .A(n3490), .ZN(n4812) );
  INV_X4 U3997 ( .A(n3487), .ZN(n4840) );
  INV_X4 U3998 ( .A(n3487), .ZN(n4841) );
  INV_X4 U3999 ( .A(n3493), .ZN(n4870) );
  INV_X4 U4000 ( .A(n3493), .ZN(n4869) );
  INV_X4 U4001 ( .A(n3485), .ZN(n4896) );
  INV_X4 U4002 ( .A(n3485), .ZN(n4897) );
  INV_X4 U4003 ( .A(n3491), .ZN(n4789) );
  INV_X4 U4004 ( .A(n3491), .ZN(n4790) );
  INV_X4 U4005 ( .A(n3492), .ZN(n4818) );
  INV_X4 U4006 ( .A(n3492), .ZN(n4819) );
  INV_X4 U4007 ( .A(n3483), .ZN(n4863) );
  INV_X4 U4008 ( .A(n3483), .ZN(n4864) );
  INV_X4 U4009 ( .A(n3483), .ZN(n4861) );
  INV_X4 U4010 ( .A(n3484), .ZN(n4890) );
  INV_X4 U4011 ( .A(n3484), .ZN(n4891) );
  INV_X4 U4012 ( .A(n3484), .ZN(n4888) );
  INV_X4 U4013 ( .A(n4912), .ZN(n4909) );
  INV_X4 U4014 ( .A(n4912), .ZN(n4910) );
  INV_X4 U4015 ( .A(n3489), .ZN(n4806) );
  INV_X4 U4016 ( .A(n3489), .ZN(n4807) );
  INV_X4 U4017 ( .A(n3486), .ZN(n4835) );
  INV_X4 U4018 ( .A(n3486), .ZN(n4836) );
  INV_X4 U4019 ( .A(n3495), .ZN(n4878) );
  INV_X4 U4020 ( .A(n3495), .ZN(n4879) );
  INV_X4 U4021 ( .A(n3488), .ZN(n4905) );
  INV_X4 U4022 ( .A(n3488), .ZN(n4906) );
  INV_X4 U4023 ( .A(n3542), .ZN(n4800) );
  INV_X4 U4024 ( .A(n3542), .ZN(n4799) );
  INV_X4 U4025 ( .A(n3541), .ZN(n4829) );
  INV_X4 U4026 ( .A(n3541), .ZN(n4828) );
  INV_X4 U4027 ( .A(n3494), .ZN(n4857) );
  INV_X4 U4028 ( .A(n3494), .ZN(n4858) );
  INV_X4 U4029 ( .A(n3496), .ZN(n4885) );
  INV_X4 U4030 ( .A(n3496), .ZN(n4886) );
  AND2_X4 U4031 ( .A1(n3418), .A2(n3414), .ZN(n4416) );
  AND2_X4 U4032 ( .A1(n3411), .A2(n3407), .ZN(n4417) );
  AND2_X4 U4033 ( .A1(n3426), .A2(n3418), .ZN(n4418) );
  AND2_X4 U4034 ( .A1(n3429), .A2(n3418), .ZN(n4419) );
  AND2_X4 U4035 ( .A1(n3429), .A2(n3415), .ZN(n4420) );
  AND2_X4 U4036 ( .A1(n3426), .A2(n3415), .ZN(n4421) );
  AND2_X4 U4037 ( .A1(n3414), .A2(n3415), .ZN(n4422) );
  AND2_X4 U4038 ( .A1(busW[2]), .A2(n4911), .ZN(n4423) );
  AND2_X4 U4039 ( .A1(busW[30]), .A2(n4911), .ZN(n4424) );
  AND2_X4 U4040 ( .A1(busW[9]), .A2(n4909), .ZN(n4425) );
  AND2_X4 U4041 ( .A1(n3414), .A2(n3411), .ZN(n4426) );
  AND2_X4 U4042 ( .A1(n3414), .A2(n3408), .ZN(n4427) );
  AND2_X4 U4043 ( .A1(n3407), .A2(n3408), .ZN(n4428) );
  INV_X4 U4044 ( .A(n3459), .ZN(n4631) );
  INV_X4 U4045 ( .A(n4631), .ZN(n4630) );
  INV_X4 U4046 ( .A(n3451), .ZN(n4647) );
  INV_X4 U4047 ( .A(n4647), .ZN(n4646) );
  INV_X4 U4048 ( .A(n3448), .ZN(n4651) );
  INV_X4 U4049 ( .A(n4651), .ZN(n4650) );
  INV_X4 U4050 ( .A(n3441), .ZN(n4663) );
  INV_X4 U4051 ( .A(n4663), .ZN(n4662) );
  INV_X4 U4052 ( .A(n3438), .ZN(n4667) );
  INV_X4 U4053 ( .A(n4667), .ZN(n4666) );
  INV_X4 U4054 ( .A(n3457), .ZN(n4635) );
  INV_X4 U4055 ( .A(n4635), .ZN(n4634) );
  INV_X4 U4056 ( .A(n3455), .ZN(n4639) );
  INV_X4 U4057 ( .A(n4639), .ZN(n4638) );
  INV_X4 U4058 ( .A(n3453), .ZN(n4643) );
  INV_X4 U4059 ( .A(n4643), .ZN(n4642) );
  INV_X4 U4060 ( .A(n3445), .ZN(n4655) );
  INV_X4 U4061 ( .A(n4655), .ZN(n4654) );
  INV_X4 U4062 ( .A(n3443), .ZN(n4659) );
  INV_X4 U4063 ( .A(n4659), .ZN(n4658) );
  INV_X4 U4064 ( .A(n3436), .ZN(n4671) );
  INV_X4 U4065 ( .A(n4671), .ZN(n4670) );
  INV_X4 U4066 ( .A(n3434), .ZN(n4675) );
  INV_X4 U4067 ( .A(n4675), .ZN(n4674) );
  INV_X4 U4068 ( .A(n4032), .ZN(n4712) );
  INV_X4 U4069 ( .A(n4032), .ZN(n4713) );
  INV_X4 U4070 ( .A(n4020), .ZN(n4714) );
  INV_X4 U4071 ( .A(n4020), .ZN(n4715) );
  INV_X4 U4072 ( .A(n4021), .ZN(n4716) );
  INV_X4 U4073 ( .A(n4021), .ZN(n4717) );
  INV_X4 U4074 ( .A(n4022), .ZN(n4718) );
  INV_X4 U4075 ( .A(n4022), .ZN(n4719) );
  INV_X4 U4076 ( .A(n4023), .ZN(n4720) );
  INV_X4 U4077 ( .A(n4023), .ZN(n4721) );
  INV_X4 U4078 ( .A(n4024), .ZN(n4722) );
  INV_X4 U4079 ( .A(n4024), .ZN(n4723) );
  INV_X4 U4080 ( .A(n4025), .ZN(n4724) );
  INV_X4 U4081 ( .A(n4025), .ZN(n4725) );
  INV_X4 U4082 ( .A(n4026), .ZN(n4726) );
  INV_X4 U4083 ( .A(n4026), .ZN(n4727) );
  INV_X4 U4084 ( .A(n4027), .ZN(n4728) );
  INV_X4 U4085 ( .A(n4027), .ZN(n4729) );
  INV_X4 U4086 ( .A(n4028), .ZN(n4730) );
  INV_X4 U4087 ( .A(n4028), .ZN(n4731) );
  INV_X4 U4088 ( .A(n4029), .ZN(n4732) );
  INV_X4 U4089 ( .A(n4029), .ZN(n4733) );
  INV_X4 U4090 ( .A(n4030), .ZN(n4734) );
  INV_X4 U4091 ( .A(n4030), .ZN(n4735) );
  INV_X4 U4092 ( .A(n4031), .ZN(n4736) );
  INV_X4 U4093 ( .A(n4031), .ZN(n4737) );
  INV_X4 U4094 ( .A(n4033), .ZN(n4738) );
  INV_X4 U4095 ( .A(n4033), .ZN(n4739) );
  INV_X4 U4096 ( .A(n4034), .ZN(n4740) );
  INV_X4 U4097 ( .A(n4034), .ZN(n4741) );
  INV_X4 U4098 ( .A(n4035), .ZN(n4742) );
  INV_X4 U4099 ( .A(n4035), .ZN(n4743) );
  INV_X4 U4100 ( .A(n4036), .ZN(n4744) );
  INV_X4 U4101 ( .A(n4036), .ZN(n4745) );
  INV_X4 U4102 ( .A(n4037), .ZN(n4746) );
  INV_X4 U4103 ( .A(n4037), .ZN(n4747) );
  INV_X4 U4104 ( .A(n4038), .ZN(n4748) );
  INV_X4 U4105 ( .A(n4038), .ZN(n4749) );
  INV_X4 U4106 ( .A(n4039), .ZN(n4750) );
  INV_X4 U4107 ( .A(n4039), .ZN(n4751) );
  INV_X4 U4108 ( .A(n4040), .ZN(n4752) );
  INV_X4 U4109 ( .A(n4040), .ZN(n4753) );
  INV_X4 U4110 ( .A(n4041), .ZN(n4754) );
  INV_X4 U4111 ( .A(n4041), .ZN(n4755) );
  INV_X4 U4112 ( .A(n3553), .ZN(n4608) );
  INV_X4 U4113 ( .A(n3553), .ZN(n4609) );
  INV_X4 U4114 ( .A(n3554), .ZN(n4610) );
  INV_X4 U4115 ( .A(n3554), .ZN(n4611) );
  INV_X4 U4116 ( .A(n3555), .ZN(n4612) );
  INV_X4 U4117 ( .A(n3555), .ZN(n4613) );
  INV_X4 U4118 ( .A(n3556), .ZN(n4614) );
  INV_X4 U4119 ( .A(n3556), .ZN(n4615) );
  INV_X4 U4120 ( .A(n3557), .ZN(n4616) );
  INV_X4 U4121 ( .A(n3557), .ZN(n4617) );
  INV_X4 U4122 ( .A(n3558), .ZN(n4618) );
  INV_X4 U4123 ( .A(n3558), .ZN(n4619) );
  INV_X4 U4124 ( .A(n3559), .ZN(n4620) );
  INV_X4 U4125 ( .A(n3559), .ZN(n4621) );
  INV_X4 U4126 ( .A(n3560), .ZN(n4622) );
  INV_X4 U4127 ( .A(n3560), .ZN(n4623) );
  INV_X4 U4128 ( .A(n3561), .ZN(n4624) );
  INV_X4 U4129 ( .A(n3561), .ZN(n4625) );
  INV_X4 U4130 ( .A(n3562), .ZN(n4626) );
  INV_X4 U4131 ( .A(n3562), .ZN(n4627) );
  INV_X4 U4132 ( .A(n3779), .ZN(n4628) );
  INV_X4 U4133 ( .A(n3779), .ZN(n4629) );
  INV_X4 U4134 ( .A(n3780), .ZN(n4632) );
  INV_X4 U4135 ( .A(n3780), .ZN(n4633) );
  INV_X4 U4136 ( .A(n3781), .ZN(n4636) );
  INV_X4 U4137 ( .A(n3781), .ZN(n4637) );
  INV_X4 U4138 ( .A(n3782), .ZN(n4640) );
  INV_X4 U4139 ( .A(n3782), .ZN(n4641) );
  INV_X4 U4140 ( .A(n3783), .ZN(n4644) );
  INV_X4 U4141 ( .A(n3783), .ZN(n4645) );
  INV_X4 U4142 ( .A(n3784), .ZN(n4648) );
  INV_X4 U4143 ( .A(n3784), .ZN(n4649) );
  INV_X4 U4144 ( .A(n3785), .ZN(n4652) );
  INV_X4 U4145 ( .A(n3785), .ZN(n4653) );
  INV_X4 U4146 ( .A(n3786), .ZN(n4656) );
  INV_X4 U4147 ( .A(n3786), .ZN(n4657) );
  INV_X4 U4148 ( .A(n3787), .ZN(n4660) );
  INV_X4 U4149 ( .A(n3787), .ZN(n4661) );
  INV_X4 U4150 ( .A(n3788), .ZN(n4664) );
  INV_X4 U4151 ( .A(n3788), .ZN(n4665) );
  INV_X4 U4152 ( .A(n3789), .ZN(n4668) );
  INV_X4 U4153 ( .A(n3789), .ZN(n4669) );
  INV_X4 U4154 ( .A(n3790), .ZN(n4672) );
  INV_X4 U4155 ( .A(n3790), .ZN(n4673) );
  INV_X4 U4156 ( .A(n4398), .ZN(n4676) );
  INV_X4 U4157 ( .A(n4398), .ZN(n4677) );
  INV_X4 U4158 ( .A(n4399), .ZN(n4680) );
  INV_X4 U4159 ( .A(n4399), .ZN(n4681) );
  INV_X4 U4160 ( .A(n4400), .ZN(n4684) );
  INV_X4 U4161 ( .A(n4400), .ZN(n4685) );
  INV_X4 U4162 ( .A(n4401), .ZN(n4688) );
  INV_X4 U4163 ( .A(n4401), .ZN(n4689) );
  INV_X4 U4164 ( .A(n4402), .ZN(n4692) );
  INV_X4 U4165 ( .A(n4402), .ZN(n4693) );
  INV_X4 U4166 ( .A(n4403), .ZN(n4696) );
  INV_X4 U4167 ( .A(n4403), .ZN(n4697) );
  INV_X4 U4168 ( .A(n4404), .ZN(n4700) );
  INV_X4 U4169 ( .A(n4404), .ZN(n4701) );
  INV_X4 U4170 ( .A(n4405), .ZN(n4704) );
  INV_X4 U4171 ( .A(n4405), .ZN(n4705) );
  INV_X4 U4172 ( .A(n4406), .ZN(n4708) );
  INV_X4 U4173 ( .A(n4406), .ZN(n4709) );
  INV_X4 U4174 ( .A(n4407), .ZN(n4774) );
  INV_X4 U4175 ( .A(n4407), .ZN(n4775) );
  INV_X4 U4176 ( .A(n4408), .ZN(n4780) );
  INV_X4 U4177 ( .A(n4408), .ZN(n4781) );
  INV_X4 U4178 ( .A(n4412), .ZN(n4782) );
  INV_X4 U4179 ( .A(n4412), .ZN(n4783) );
  INV_X4 U4180 ( .A(n4410), .ZN(n4784) );
  INV_X4 U4181 ( .A(n4410), .ZN(n4785) );
  INV_X4 U4182 ( .A(n4414), .ZN(n4844) );
  INV_X4 U4183 ( .A(n4414), .ZN(n4845) );
  INV_X4 U4184 ( .A(n4409), .ZN(n4846) );
  INV_X4 U4185 ( .A(n4409), .ZN(n4847) );
  INV_X4 U4186 ( .A(n4413), .ZN(n4848) );
  INV_X4 U4187 ( .A(n4413), .ZN(n4849) );
  INV_X4 U4188 ( .A(n4411), .ZN(n4850) );
  INV_X4 U4189 ( .A(n4411), .ZN(n4851) );
  INV_X4 U4190 ( .A(n4415), .ZN(n4907) );
  INV_X4 U4191 ( .A(n4415), .ZN(n4908) );
  INV_X4 U4192 ( .A(n3489), .ZN(n4801) );
  INV_X4 U4193 ( .A(n3486), .ZN(n4830) );
  INV_X4 U4194 ( .A(n3495), .ZN(n4873) );
  INV_X4 U4195 ( .A(n3488), .ZN(n4900) );
  INV_X4 U4196 ( .A(n3542), .ZN(n4793) );
  INV_X4 U4197 ( .A(n3541), .ZN(n4822) );
  INV_X4 U4198 ( .A(n3494), .ZN(n4852) );
  INV_X4 U4199 ( .A(n3496), .ZN(n4880) );
  INV_X4 U4200 ( .A(n3490), .ZN(n4808) );
  INV_X4 U4201 ( .A(n3490), .ZN(n4813) );
  INV_X4 U4202 ( .A(n3487), .ZN(n4837) );
  INV_X4 U4203 ( .A(n3487), .ZN(n4842) );
  INV_X4 U4204 ( .A(n3493), .ZN(n4866) );
  INV_X4 U4205 ( .A(n3493), .ZN(n4871) );
  INV_X4 U4206 ( .A(n3485), .ZN(n4892) );
  INV_X4 U4207 ( .A(n3485), .ZN(n4898) );
  INV_X4 U4208 ( .A(n3491), .ZN(n4786) );
  INV_X4 U4209 ( .A(n3491), .ZN(n4791) );
  INV_X4 U4210 ( .A(n3492), .ZN(n4815) );
  INV_X4 U4211 ( .A(n3492), .ZN(n4820) );
  INV_X4 U4212 ( .A(n3483), .ZN(n4859) );
  INV_X4 U4213 ( .A(n3484), .ZN(n4887) );
  INV_X4 U4214 ( .A(reset), .ZN(n4912) );
  INV_X4 U4215 ( .A(n4912), .ZN(n4911) );
endmodule

