module testbench;
    reg [0:31] in0;
    reg [0:31] in1;
    reg [0:31] in2;
    reg [0:31] in3;
    reg [0:31] in4;
    reg [0:31] in5;
    reg [0:31] in6;
    reg [0:31] in7;

    reg [0:2] SEL;
    wire [0:31] Z;

    mux8to1_32bit MUX8TO1_32BIT (
        .in0(in0),
        .in1(in1),
        .in2(in2),
        .in3(in3),
        .in4(in4),
        .in5(in5),
        .in6(in6),
        .in7(in7),
        .sel(SEL),
        .Z(Z)
    );
    
    initial begin
        $monitor("in0=%h in1=%h in2=%h in3=%h in4=%h in5=%h in6=%h in7=%h sel=%h Z=%h",in0,in1,in2,in3,in4,in5,in6,in7,SEL,Z);

        #0 in0 = 32'h00000000; in1 = 32'h11111111; in2 = 32'h22222222; in3 = 32'h33333333; in4 = 32'h44444444; in5 = 32'h55555555; in6 = 32'h66666666; in7 = 32'h77777777; SEL=3'h0;
        #1 in0 = 32'h00000000; in1 = 32'h11111111; in2 = 32'h22222222; in3 = 32'h33333333; in4 = 32'h44444444; in5 = 32'h55555555; in6 = 32'h66666666; in7 = 32'h77777777; SEL=3'h1;
        #1 in0 = 32'h00000000; in1 = 32'h11111111; in2 = 32'h22222222; in3 = 32'h33333333; in4 = 32'h44444444; in5 = 32'h55555555; in6 = 32'h66666666; in7 = 32'h77777777; SEL=3'h2;
        #1 in0 = 32'h00000000; in1 = 32'h11111111; in2 = 32'h22222222; in3 = 32'h33333333; in4 = 32'h44444444; in5 = 32'h55555555; in6 = 32'h66666666; in7 = 32'h77777777; SEL=3'h3;

        #1 in0 = 32'h00000000; in1 = 32'h11111111; in2 = 32'h22222222; in3 = 32'h33333333; in4 = 32'h44444444; in5 = 32'h55555555; in6 = 32'h66666666; in7 = 32'h77777777; SEL=3'h4;
        #1 in0 = 32'h00000000; in1 = 32'h11111111; in2 = 32'h22222222; in3 = 32'h33333333; in4 = 32'h44444444; in5 = 32'h55555555; in6 = 32'h66666666; in7 = 32'h77777777; SEL=3'h5;
        #1 in0 = 32'h00000000; in1 = 32'h11111111; in2 = 32'h22222222; in3 = 32'h33333333; in4 = 32'h44444444; in5 = 32'h55555555; in6 = 32'h66666666; in7 = 32'h77777777; SEL=3'h6;
        #1 in0 = 32'h00000000; in1 = 32'h11111111; in2 = 32'h22222222; in3 = 32'h33333333; in4 = 32'h44444444; in5 = 32'h55555555; in6 = 32'h66666666; in7 = 32'h77777777; SEL=3'h7;

    end
endmodule // testbench