
module single_cycle_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   \ab[28][2] , \ab[27][3] , \ab[27][0] , \ab[26][4] , \ab[26][3] ,
         \ab[26][2] , \ab[26][1] , \ab[26][0] , \ab[25][4] , \ab[25][1] ,
         \ab[25][0] , \ab[24][6] , \ab[24][5] , \ab[24][2] , \ab[24][0] ,
         \ab[23][8] , \ab[23][6] , \ab[23][5] , \ab[23][2] , \ab[23][0] ,
         \ab[22][8] , \ab[22][6] , \ab[22][4] , \ab[22][2] , \ab[22][1] ,
         \ab[22][0] , \ab[21][10] , \ab[21][9] , \ab[21][7] , \ab[21][6] ,
         \ab[21][4] , \ab[21][3] , \ab[21][2] , \ab[21][1] , \ab[21][0] ,
         \ab[20][10] , \ab[20][8] , \ab[20][7] , \ab[20][6] , \ab[20][4] ,
         \ab[20][3] , \ab[20][2] , \ab[20][1] , \ab[20][0] , \ab[19][12] ,
         \ab[19][11] , \ab[19][9] , \ab[19][8] , \ab[19][7] , \ab[19][5] ,
         \ab[19][4] , \ab[19][3] , \ab[19][2] , \ab[19][0] , \ab[18][13] ,
         \ab[18][12] , \ab[18][10] , \ab[18][9] , \ab[18][7] , \ab[18][6] ,
         \ab[18][5] , \ab[18][4] , \ab[18][3] , \ab[18][2] , \ab[18][1] ,
         \ab[18][0] , \ab[17][13] , \ab[17][11] , \ab[17][10] , \ab[17][8] ,
         \ab[17][7] , \ab[17][5] , \ab[17][4] , \ab[17][3] , \ab[17][2] ,
         \ab[17][1] , \ab[17][0] , \ab[16][15] , \ab[16][14] , \ab[16][12] ,
         \ab[16][11] , \ab[16][8] , \ab[16][6] , \ab[16][5] , \ab[16][4] ,
         \ab[16][3] , \ab[16][2] , \ab[16][0] , \ab[15][16] , \ab[15][15] ,
         \ab[15][14] , \ab[15][12] , \ab[15][11] , \ab[15][9] , \ab[15][8] ,
         \ab[15][7] , \ab[15][6] , \ab[15][5] , \ab[15][4] , \ab[15][3] ,
         \ab[15][2] , \ab[15][0] , \ab[14][16] , \ab[14][15] , \ab[14][13] ,
         \ab[14][12] , \ab[14][11] , \ab[14][9] , \ab[14][7] , \ab[14][6] ,
         \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][1] , \ab[14][0] ,
         \ab[13][18] , \ab[13][17] , \ab[13][16] , \ab[13][15] , \ab[13][13] ,
         \ab[13][12] , \ab[13][10] , \ab[13][9] , \ab[13][7] , \ab[13][6] ,
         \ab[13][5] , \ab[13][4] , \ab[13][3] , \ab[13][2] , \ab[13][0] ,
         \ab[12][19] , \ab[12][18] , \ab[12][17] , \ab[12][16] , \ab[12][14] ,
         \ab[12][13] , \ab[12][12] , \ab[12][9] , \ab[12][7] , \ab[12][6] ,
         \ab[12][5] , \ab[12][4] , \ab[12][3] , \ab[12][2] , \ab[12][0] ,
         \ab[11][20] , \ab[11][19] , \ab[11][18] , \ab[11][17] , \ab[11][16] ,
         \ab[11][15] , \ab[11][14] , \ab[11][13] , \ab[11][11] , \ab[11][10] ,
         \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] , \ab[11][4] ,
         \ab[11][3] , \ab[11][1] , \ab[11][0] , \ab[10][21] , \ab[10][20] ,
         \ab[10][19] , \ab[10][18] , \ab[10][16] , \ab[10][15] , \ab[10][14] ,
         \ab[10][13] , \ab[10][11] , \ab[10][9] , \ab[10][8] , \ab[10][7] ,
         \ab[10][6] , \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][1] ,
         \ab[10][0] , \ab[9][22] , \ab[9][21] , \ab[9][20] , \ab[9][19] ,
         \ab[9][16] , \ab[9][15] , \ab[9][14] , \ab[9][11] , \ab[9][9] ,
         \ab[9][8] , \ab[9][7] , \ab[9][6] , \ab[9][5] , \ab[9][4] ,
         \ab[9][3] , \ab[9][2] , \ab[9][1] , \ab[9][0] , \ab[8][23] ,
         \ab[8][22] , \ab[8][21] , \ab[8][20] , \ab[8][18] , \ab[8][16] ,
         \ab[8][15] , \ab[8][14] , \ab[8][13] , \ab[8][11] , \ab[8][9] ,
         \ab[8][8] , \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][24] , \ab[7][23] ,
         \ab[7][22] , \ab[7][21] , \ab[7][20] , \ab[7][19] , \ab[7][18] ,
         \ab[7][17] , \ab[7][16] , \ab[7][15] , \ab[7][14] , \ab[7][13] ,
         \ab[7][12] , \ab[7][10] , \ab[7][9] , \ab[7][8] , \ab[7][7] ,
         \ab[7][6] , \ab[7][5] , \ab[7][3] , \ab[7][2] , \ab[7][1] ,
         \ab[7][0] , \ab[6][25] , \ab[6][24] , \ab[6][23] , \ab[6][22] ,
         \ab[6][20] , \ab[6][19] , \ab[6][18] , \ab[6][17] , \ab[6][16] ,
         \ab[6][15] , \ab[6][13] , \ab[6][12] , \ab[6][10] , \ab[6][9] ,
         \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] ,
         \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][26] ,
         \ab[5][25] , \ab[5][24] , \ab[5][23] , \ab[5][21] , \ab[5][20] ,
         \ab[5][19] , \ab[5][18] , \ab[5][17] , \ab[5][16] , \ab[5][13] ,
         \ab[5][12] , \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] ,
         \ab[5][6] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][27] , \ab[4][26] , \ab[4][25] , \ab[4][24] ,
         \ab[4][23] , \ab[4][21] , \ab[4][20] , \ab[4][19] , \ab[4][18] ,
         \ab[4][17] , \ab[4][14] , \ab[4][13] , \ab[4][12] , \ab[4][11] ,
         \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] , \ab[4][6] ,
         \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] , \ab[4][1] ,
         \ab[4][0] , \ab[3][28] , \ab[3][27] , \ab[3][26] , \ab[3][25] ,
         \ab[3][24] , \ab[3][22] , \ab[3][21] , \ab[3][20] , \ab[3][19] ,
         \ab[3][18] , \ab[3][17] , \ab[3][14] , \ab[3][12] , \ab[3][11] ,
         \ab[3][10] , \ab[3][9] , \ab[3][8] , \ab[3][7] , \ab[3][6] ,
         \ab[3][5] , \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] ,
         \ab[3][0] , \ab[2][29] , \ab[2][28] , \ab[2][27] , \ab[2][26] ,
         \ab[2][25] , \ab[2][22] , \ab[2][21] , \ab[2][20] , \ab[2][19] ,
         \ab[2][18] , \ab[2][17] , \ab[2][15] , \ab[2][14] , \ab[2][12] ,
         \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] , \ab[2][5] ,
         \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] ,
         \ab[1][30] , \ab[1][29] , \ab[1][28] , \ab[1][27] , \ab[1][26] ,
         \ab[1][25] , \ab[1][21] , \ab[1][20] , \ab[1][19] , \ab[1][18] ,
         \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] ,
         \ab[0][31] , \ab[0][30] , \ab[0][29] , \ab[0][28] , \ab[0][27] ,
         \ab[0][24] , \ab[0][23] , \ab[0][22] , \ab[0][21] , \ab[0][20] ,
         \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][9] , \ab[0][6] ,
         \ab[0][5] , \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[15][15] ,
         \CARRYB[15][14] , \CARRYB[15][12] , \CARRYB[15][11] , \CARRYB[15][8] ,
         \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][3] , \CARRYB[15][2] ,
         \CARRYB[15][0] , \CARRYB[14][16] , \CARRYB[14][15] , \CARRYB[14][14] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][9] , \CARRYB[14][7] ,
         \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] , \CARRYB[14][3] ,
         \CARRYB[14][2] , \CARRYB[14][0] , \CARRYB[13][17] , \CARRYB[13][16] ,
         \CARRYB[13][15] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][0] , \CARRYB[12][18] ,
         \CARRYB[12][17] , \CARRYB[12][16] , \CARRYB[12][15] ,
         \CARRYB[12][13] , \CARRYB[12][12] , \CARRYB[12][7] , \CARRYB[12][6] ,
         \CARRYB[12][5] , \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] ,
         \CARRYB[12][0] , \CARRYB[11][19] , \CARRYB[11][18] , \CARRYB[11][17] ,
         \CARRYB[11][16] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][9] , \CARRYB[11][7] , \CARRYB[11][6] ,
         \CARRYB[11][5] , \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] ,
         \CARRYB[11][0] , \CARRYB[10][20] , \CARRYB[10][19] , \CARRYB[10][18] ,
         \CARRYB[10][17] , \CARRYB[10][16] , \CARRYB[10][15] ,
         \CARRYB[10][14] , \CARRYB[10][13] , \CARRYB[10][10] , \CARRYB[10][8] ,
         \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] ,
         \CARRYB[10][3] , \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][21] ,
         \CARRYB[9][20] , \CARRYB[9][19] , \CARRYB[9][18] , \CARRYB[9][16] ,
         \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][11] ,
         \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] ,
         \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][1] ,
         \CARRYB[9][0] , \CARRYB[8][22] , \CARRYB[8][21] , \CARRYB[8][20] ,
         \CARRYB[8][19] , \CARRYB[8][16] , \CARRYB[8][15] , \CARRYB[8][14] ,
         \CARRYB[8][11] , \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] ,
         \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][23] , \CARRYB[7][22] , \CARRYB[7][21] ,
         \CARRYB[7][20] , \CARRYB[7][16] , \CARRYB[7][15] , \CARRYB[7][14] ,
         \CARRYB[7][13] , \CARRYB[7][11] , \CARRYB[7][9] , \CARRYB[7][8] ,
         \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][2] ,
         \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][24] , \CARRYB[6][23] ,
         \CARRYB[6][22] , \CARRYB[6][19] , \CARRYB[6][18] , \CARRYB[6][17] ,
         \CARRYB[6][16] , \CARRYB[6][15] , \CARRYB[6][13] , \CARRYB[6][12] ,
         \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][7] , \CARRYB[6][6] ,
         \CARRYB[6][5] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][25] , \CARRYB[5][24] , \CARRYB[5][23] ,
         \CARRYB[5][22] , \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] ,
         \CARRYB[5][17] , \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][13] ,
         \CARRYB[5][12] , \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] ,
         \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] ,
         \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] ,
         \CARRYB[4][26] , \CARRYB[4][25] , \CARRYB[4][24] , \CARRYB[4][23] ,
         \CARRYB[4][21] , \CARRYB[4][20] , \CARRYB[4][19] , \CARRYB[4][18] ,
         \CARRYB[4][17] , \CARRYB[4][16] , \CARRYB[4][13] , \CARRYB[4][12] ,
         \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] , \CARRYB[4][7] ,
         \CARRYB[4][6] , \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] ,
         \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][27] , \CARRYB[3][26] ,
         \CARRYB[3][25] , \CARRYB[3][24] , \CARRYB[3][23] , \CARRYB[3][21] ,
         \CARRYB[3][20] , \CARRYB[3][19] , \CARRYB[3][18] , \CARRYB[3][17] ,
         \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][11] , \CARRYB[3][10] ,
         \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][28] , \CARRYB[2][27] , \CARRYB[2][26] ,
         \CARRYB[2][25] , \CARRYB[2][24] , \CARRYB[2][22] , \CARRYB[2][21] ,
         \CARRYB[2][20] , \CARRYB[2][19] , \CARRYB[2][18] , \CARRYB[2][17] ,
         \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][11] , \CARRYB[2][10] ,
         \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \CARRYB[1][26] , \CARRYB[1][22] , \CARRYB[1][21] , \CARRYB[1][20] ,
         \CARRYB[1][19] , \CARRYB[1][18] , \CARRYB[1][15] , \CARRYB[1][12] ,
         \CARRYB[1][11] , \CARRYB[1][10] , \CARRYB[1][9] , \CARRYB[1][5] ,
         \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] , \CARRYB[1][0] ,
         \SUMB[15][15] , \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][9] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[14][17] , \SUMB[14][16] , \SUMB[14][15] , \SUMB[14][13] ,
         \SUMB[14][12] , \SUMB[14][7] , \SUMB[14][6] , \SUMB[14][5] ,
         \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][1] , \SUMB[13][18] ,
         \SUMB[13][17] , \SUMB[13][16] , \SUMB[13][14] , \SUMB[13][13] ,
         \SUMB[13][12] , \SUMB[13][10] , \SUMB[13][8] , \SUMB[13][7] ,
         \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][2] ,
         \SUMB[13][1] , \SUMB[12][19] , \SUMB[12][18] , \SUMB[12][17] ,
         \SUMB[12][16] , \SUMB[12][15] , \SUMB[12][14] , \SUMB[12][13] ,
         \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][8] , \SUMB[12][7] ,
         \SUMB[12][6] , \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] ,
         \SUMB[11][20] , \SUMB[11][19] , \SUMB[11][18] , \SUMB[11][17] ,
         \SUMB[11][15] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][10] ,
         \SUMB[11][8] , \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] ,
         \SUMB[11][4] , \SUMB[11][3] , \SUMB[11][1] , \SUMB[10][21] ,
         \SUMB[10][20] , \SUMB[10][19] , \SUMB[10][18] , \SUMB[10][16] ,
         \SUMB[10][15] , \SUMB[10][14] , \SUMB[10][12] , \SUMB[10][9] ,
         \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][2] , \SUMB[10][1] , \SUMB[9][22] ,
         \SUMB[9][21] , \SUMB[9][20] , \SUMB[9][19] , \SUMB[9][16] ,
         \SUMB[9][15] , \SUMB[9][14] , \SUMB[9][12] , \SUMB[9][10] ,
         \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] ,
         \SUMB[9][4] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][23] ,
         \SUMB[8][22] , \SUMB[8][21] , \SUMB[8][20] , \SUMB[8][16] ,
         \SUMB[8][15] , \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] ,
         \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][2] , \SUMB[8][1] ,
         \SUMB[7][24] , \SUMB[7][23] , \SUMB[7][22] , \SUMB[7][21] ,
         \SUMB[7][19] , \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] ,
         \SUMB[7][14] , \SUMB[7][12] , \SUMB[7][10] , \SUMB[7][9] ,
         \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][25] , \SUMB[6][24] , \SUMB[6][23] , \SUMB[6][22] ,
         \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][17] , \SUMB[6][16] ,
         \SUMB[6][15] , \SUMB[6][13] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][4] ,
         \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][26] ,
         \SUMB[5][25] , \SUMB[5][24] , \SUMB[5][23] , \SUMB[5][21] ,
         \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] , \SUMB[5][17] ,
         \SUMB[5][16] , \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][11] ,
         \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][27] ,
         \SUMB[4][26] , \SUMB[4][24] , \SUMB[4][22] , \SUMB[4][21] ,
         \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] , \SUMB[4][17] ,
         \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][5] , \SUMB[4][4] ,
         \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][28] ,
         \SUMB[3][27] , \SUMB[3][26] , \SUMB[3][25] , \SUMB[3][24] ,
         \SUMB[3][22] , \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] ,
         \SUMB[3][18] , \SUMB[3][15] , \SUMB[3][14] , \SUMB[3][12] ,
         \SUMB[3][11] , \SUMB[3][10] , \SUMB[3][9] , \SUMB[3][8] ,
         \SUMB[3][7] , \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] ,
         \SUMB[3][1] , \SUMB[2][29] , \SUMB[2][28] , \SUMB[2][27] ,
         \SUMB[2][26] , \SUMB[2][25] , \SUMB[2][23] , \SUMB[2][22] ,
         \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] ,
         \SUMB[2][15] , \SUMB[2][14] , \SUMB[2][13] , \SUMB[2][12] ,
         \SUMB[2][11] , \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] ,
         \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] ,
         \SUMB[2][1] , \SUMB[1][29] , \SUMB[1][28] , \SUMB[1][27] ,
         \SUMB[1][26] , \SUMB[1][23] , \SUMB[1][21] , \SUMB[1][20] ,
         \SUMB[1][19] , \SUMB[1][16] , \SUMB[1][13] , \SUMB[1][12] ,
         \SUMB[1][11] , \SUMB[1][10] , \SUMB[1][9] , \SUMB[1][6] ,
         \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] ,
         \CARRYB[27][2] , \CARRYB[27][1] , \CARRYB[26][3] , \CARRYB[26][0] ,
         \CARRYB[25][4] , \CARRYB[25][3] , \CARRYB[25][2] , \CARRYB[25][0] ,
         \CARRYB[24][5] , \CARRYB[24][4] , \CARRYB[24][1] , \CARRYB[24][0] ,
         \CARRYB[23][7] , \CARRYB[23][6] , \CARRYB[23][5] , \CARRYB[23][2] ,
         \CARRYB[23][0] , \CARRYB[22][8] , \CARRYB[22][6] , \CARRYB[22][4] ,
         \CARRYB[22][2] , \CARRYB[22][0] , \CARRYB[21][9] , \CARRYB[21][8] ,
         \CARRYB[21][6] , \CARRYB[21][4] , \CARRYB[21][2] , \CARRYB[21][1] ,
         \CARRYB[21][0] , \CARRYB[20][10] , \CARRYB[20][9] , \CARRYB[20][7] ,
         \CARRYB[20][6] , \CARRYB[20][4] , \CARRYB[20][2] , \CARRYB[20][1] ,
         \CARRYB[20][0] , \CARRYB[19][11] , \CARRYB[19][10] , \CARRYB[19][8] ,
         \CARRYB[19][7] , \CARRYB[19][6] , \CARRYB[19][4] , \CARRYB[19][3] ,
         \CARRYB[19][2] , \CARRYB[19][0] , \CARRYB[18][12] , \CARRYB[18][11] ,
         \CARRYB[18][9] , \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][0] ,
         \CARRYB[17][13] , \CARRYB[17][10] , \CARRYB[17][9] , \CARRYB[17][5] ,
         \CARRYB[17][4] , \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][0] ,
         \CARRYB[16][14] , \CARRYB[16][13] , \CARRYB[16][11] , \CARRYB[16][8] ,
         \CARRYB[16][7] , \CARRYB[16][5] , \CARRYB[16][3] , \CARRYB[16][2] ,
         \CARRYB[16][0] , \SUMB[26][4] , \SUMB[26][1] , \SUMB[25][5] ,
         \SUMB[25][4] , \SUMB[24][5] , \SUMB[23][8] , \SUMB[23][6] ,
         \SUMB[23][1] , \SUMB[22][9] , \SUMB[22][7] , \SUMB[22][3] ,
         \SUMB[22][1] , \SUMB[21][10] , \SUMB[21][9] , \SUMB[21][7] ,
         \SUMB[21][4] , \SUMB[21][3] , \SUMB[21][2] , \SUMB[21][1] ,
         \SUMB[20][11] , \SUMB[20][10] , \SUMB[20][8] , \SUMB[20][4] ,
         \SUMB[20][3] , \SUMB[20][2] , \SUMB[20][1] , \SUMB[19][11] ,
         \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] , \SUMB[19][2] ,
         \SUMB[19][1] , \SUMB[18][12] , \SUMB[18][8] , \SUMB[18][5] ,
         \SUMB[18][4] , \SUMB[18][3] , \SUMB[18][1] , \SUMB[17][14] ,
         \SUMB[17][13] , \SUMB[17][11] , \SUMB[17][10] , \SUMB[17][5] ,
         \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][1] , \SUMB[16][14] ,
         \SUMB[16][12] , \SUMB[16][11] , \SUMB[16][9] , \SUMB[16][8] ,
         \SUMB[16][6] , \SUMB[16][5] , \SUMB[16][4] , \SUMB[16][3] ,
         \SUMB[16][2] , net70435, net70441, net70443, net70445, net70447,
         net70449, net70451, net70452, net70453, net70454, net70455, net70456,
         net70457, net70459, net70460, net70461, net70463, net70465, net70467,
         net70469, net70470, net70471, net70472, net70473, net70474, net70475,
         net70476, net70477, net70478, net70482, net70486, net70491, net70492,
         net77860, net77858, net77868, net77866, net77878, net77886, net77882,
         net77892, net77900, net77898, net77908, net77906, net77914, net77912,
         net77920, net77926, net77924, net77932, net77930, net77940, net77938,
         net77948, net77946, net77956, net77966, net77964, net77970,
         \*UDW_*112679/net78533 , \*UDW_*112684/net78547 ,
         \*UDW_*112694/net78575 , \*UDW_*112704/net78605 ,
         \*UDW_*112739/net78703 , net79906, net79905, net79904, net79893,
         net79892, net79891, net79939, net79937, net79936, net79935, net79961,
         net79960, net79959, net79957, net79956, net79955, net79953, net79952,
         net79951, net79970, net79969, net79968, net79993, net79992, net80258,
         net80255, net80254, net80248, net80247, net80246, net80275, net80274,
         net80273, net80264, net80356, net80355, net80350, net80349, net80348,
         net80392, net80409, net80451, net80449, net80480, net80479, net80478,
         net80510, net80523, net80522, net80521, net80520, net80519, net80518,
         net80566, net80565, net80563, net80562, net80561, net80643, net80676,
         net80675, net80674, net80673, net80672, net80671, net80694, net80727,
         net80769, net80768, net80767, net80796, net80795, net80793, net80792,
         net80791, net80818, net80817, net80816, net80814, net80813, net80812,
         net80806, net80805, net80852, net80850, net80845, net80844, net80840,
         net80839, net80838, net80836, net80835, net80880, net80879, net80926,
         net80925, net80924, net80922, net80921, net80920, net80958, net80957,
         net80956, net80942, net80941, net80940, net80983, net80993, net80992,
         net80991, net80990, net81038, net81037, net81036, net81035, net81034,
         net81033, net81069, net81068, net81067, net81066, net81065, net81060,
         net81059, net81058, net81057, net81056, net81053, net81052, net81080,
         net81112, net81111, net81110, net81180, net81179, net81178, net81169,
         net81206, net81205, net81204, net81213, net81212, net81211, net81267,
         net81266, net81265, net81262, net81261, net81260, net81259, net81258,
         net81354, net81367, net81365, net81424, net81431, net81491, net81493,
         net81535, net81533, net81531, net81530, net81515, net81514, net81513,
         net81548, net81581, net81586, net81617, net81616, net81615, net81663,
         net81673, net81714, net81713, net81756, net81781, net81780, net81779,
         net81782, net81815, net81945, net81956, net81955, net81958, net81983,
         net81995, net82031, net82029, net82028, net82027, net82024, net82046,
         net82045, net82089, net82101, net82099, net82149, net82154, net82159,
         net82239, net82238, net82247, net82408, net82407, net82534, net82532,
         net82548, net82558, net82557, net82556, net82551, net82550, net82601,
         net82641, net82669, net82668, net82667, net82666, net82665, net82664,
         net82678, net82723, net82760, net82759, net82757, net82834, net82850,
         net82849, net82848, net82890, net83121, net83120, net83134, net83151,
         net83175, net83174, net83172, net83263, net83296, net83351, net83358,
         net83357, net83445, net83535, net83736, net83784, net83797, net83796,
         net83850, net83866, net83919, net84007, net84118, net84116, net84163,
         net84212, net84211, net84209, net84309, net84308, net84305, net84304,
         net84303, net84302, net84301, net84300, net84299, net84298, net84297,
         net84348, net84358, net84481, net84657, net84698, net84712, net84711,
         net84710, net84708, net84707, net84706, net84746, net84826, net84825,
         net84818, net84817, net84891, net84902, net84926, net84925, net84924,
         net84948, net84947, net85000, net84999, net84998, net85017, net85036,
         net85035, net85044, net85043, net85212, net85254, net85251, net85325,
         net85373, net85469, net85465, net85457, net85456, net85455, net85543,
         net85540, net85603, net85602, net85716, net85732, net85734, net85979,
         net86054, net86101, net86159, net86158, net86172, net86171, net86170,
         net86385, net86414, net86413, net86412, net86427, net86440, net86464,
         net86557, net86565, net86601, net86630, net86629, net86656, net86654,
         net86653, net86652, net86651, net86649, net86662, net86661, net86704,
         net86703, net86702, net86699, net86698, net86697, net86844, net86864,
         net86896, net86895, net86894, net86893, net87012, net87011, net87010,
         net87005, net87004, net87003, net87045, net87064, net87136, net87133,
         net87310, net87309, net87308, net87411, net87465, net87464, net87573,
         net87619, net87683, net87682, net87874, net88086, net88157, net88156,
         net88165, net88166, net88177, net88211, net88210, net88209, net88208,
         net88207, net88206, net88297, net88296, net88295, net88344, net88410,
         net88408, net88407, net88444, net88449, net88455, net88525, net88638,
         net88656, net88655, net88692, net88702, net88704, net88703, net88712,
         net88800, net88860, net88859, net88868, net88867, net88887, net88928,
         net88934, net89026, net89255, net89289, net89402, net89467, net89819,
         net89876, net89997, net90174, net90347, net90433, net90687, net90702,
         net90731, net91001, net91088, net91118, net91243, net91301, net91660,
         \SUMB[25][1] , net92341, net92322, net92314, net92311, net92378,
         net92405, net92542, net92724, net92718, net92717, net92716, net92863,
         net92862, net92884, net93203, net93243, net93309, net93308, net93713,
         net93747, net93840, net93878, net93880, \ab[6][21] , \SUMB[6][21] ,
         \CARRYB[6][21] , \CARRYB[6][20] , \CARRYB[5][21] , net84883,
         \ab[2][24] , \ab[0][26] , \SUMB[1][25] , \*UDW_*112644/net78437 ,
         \ab[19][10] , \CARRYB[18][10] , \ab[0][25] , net80303, net80302,
         \ab[9][18] , \CARRYB[8][18] , \CARRYB[7][18] , net93674,
         \SUMB[13][15] , \ab[23][7] , \ab[16][13] , net89353, net88647,
         \ab[18][11] , \SUMB[18][11] , \CARRYB[17][11] , net86231, net81340,
         \ab[8][19] , \SUMB[8][19] , \SUMB[7][20] , \CARRYB[7][19] ,
         \ab[2][23] , \ab[1][23] , net80803, net80802, net80801, net79950,
         \ab[10][17] , \SUMB[9][18] , \CARRYB[9][17] , \ab[21][8] ,
         \SUMB[19][9] , \CARRYB[20][8] , net88961, \SUMB[22][8] , \ab[13][14] ,
         net89461, net80267, \ab[22][7] , \CARRYB[22][7] , \ab[15][13] ,
         \CARRYB[15][13] , \ab[12][15] , \CARRYB[11][15] , net89094, net83116,
         net83115, net80110, net79863, \SUMB[23][7] , \SUMB[5][22] ,
         \SUMB[4][23] , \ab[1][24] , \ab[14][14] , \CARRYB[13][14] , net90525,
         net90103, net81290, \ab[17][12] , \SUMB[17][12] , \SUMB[16][13] ,
         \SUMB[15][14] , \CARRYB[17][12] , \CARRYB[16][12] , net84357,
         net70480, \ab[3][23] , \CARRYB[2][23] , net81946, net79865, net79864,
         \ab[24][7] , \CARRYB[24][6] , net84978, net92323, net92321, net92320,
         net92319, net86937, net84979, net82807, \ab[31][0] , \ab[27][4] ,
         \ab[26][5] , \SUMB[26][5] , \CARRYB[26][4] , net88004, net83576,
         net83575, net83044, net82124, net82044, net82043, net90801, net81113,
         net80268, \SUMB[21][8] , \CARRYB[21][7] , \SUMB[2][24] , net79867,
         \ab[25][5] , \SUMB[24][6] , \CARRYB[25][5] , \SUMB[11][16] , net90671,
         net87855, \ab[4][22] , \SUMB[3][23] , \CARRYB[3][22] , net80825,
         net80794, net88756, net82658, net82657, \CARRYB[12][14] , net88916,
         net86696, net79868, net93107, net85119, net80485, net80484,
         \SUMB[14][14] , \CARRYB[14][13] , net84313, net84312, net84311,
         net81285, net81284, \ab[5][22] , \CARRYB[4][22] , net88226, net88225,
         net86409, net86407, net81394, net80517, \SUMB[10][17] , net80257,
         \ab[25][2] , net83755, \SUMB[15][7] , net83202, \SUMB[20][5] ,
         net93792, net93791, net81070, \SUMB[26][2] , \CARRYB[26][1] ,
         net119817, net119855, net119949, net119921, net119920, net119982,
         net119979, net120174, net120359, net120468, net120467, net120466,
         net120464, net120463, net120501, net120519, net120518, net120517,
         net120515, net120514, net120513, net120586, net120585, net120628,
         net120627, net120653, net120652, net120651, net120922, net121150,
         net121285, net121380, net121455, net121454, net121453, net121523,
         net121607, net121606, net121785, net121814, net121859, net121926,
         net122087, net90802, net87134, net87009, net86404, net86403, net82396,
         net82255, net81954, net81953, \ab[20][9] , \SUMB[20][9] ,
         \SUMB[19][10] , \CARRYB[19][9] , net80660, net80658, net80657,
         net80366, \CARRYB[7][17] , net123000, net123072, net123062, net123055,
         net123028, net123019, net123143, net123142, net123303, net123430,
         net123429, net123428, net123427, net123509, net123592, net123591,
         net123843, net123842, net123899, net123898, net123897, net124104,
         net124367, net124434, net124563, net124618, net124723, net124757,
         net124874, net125062, net125375, net90817, net88668, net93672,
         net92325, net92318, net92317, net87655, net87654, net81157,
         \CARRYB[29][1] , net86884, net83030, \SUMB[26][3] , net84447,
         \SUMB[8][14] , net83438, net80346, \ab[9][13] , \SUMB[10][13] ,
         net93756, net87942, net82263, \SUMB[14][10] , \CARRYB[15][9] ,
         \SUMB[18][9] , \ab[15][10] , net87797, net124392, net87068, net87067,
         net87065, net81371, \CARRYB[8][13] , net88700, \ab[5][15] , net88079,
         net124908, net120511, net83630, net83629, net83628, net80251,
         net80250, \ab[11][12] , \ab[2][16] , net93813, net89008, net84434,
         net79909, \SUMB[23][5] , net82030, net86799, \ab[16][9] ,
         \SUMB[15][10] , \ab[23][4] , net87944, net87688, net86801, net82561,
         net82560, net82559, net125934, \ab[16][10] , \SUMB[15][11] ,
         \SUMB[14][11] , \CARRYB[15][10] , net93410, net87945, net85808,
         net85807, \ab[18][8] , \SUMB[17][9] , \CARRYB[17][8] , net87490,
         net83631, net81168, net81167, net81166, net81087, \ab[12][11] ,
         net84213, net80290, net79991, net79990, net79989, \CARRYB[21][5] ,
         net93918, net80686, \ab[27][2] , net89453, net80474, net80473,
         net80472, net80989, net80988, net80987, net80263, net80262, net80261,
         \CARRYB[26][2] , net90604, net90262, net89670, net84824, net82022,
         net82021, \ab[13][11] , \SUMB[11][12] , \CARRYB[12][11] ,
         \CARRYB[11][11] , net84680, net84679, net84678, \CARRYB[24][3] ,
         net89109, net90996, net89982, net89065, net85399, net84822, net84820,
         net84819, net80353, net80352, net80351, \ab[10][12] , \SUMB[9][13] ,
         \CARRYB[9][12] , \CARRYB[10][12] , net88123, net87941, net87940,
         net87939, net87938, net86024, net86023, net86022, net82544, net81007,
         net81006, \ab[25][3] , \SUMB[24][4] , net80021, net79908, net79907,
         net84208, net81992, net79981, net79980, net121214, net120657,
         net120656, net120655, \ab[17][9] , \CARRYB[16][9] , net85096,
         net80668, net80667, net86162, net84445, net80834, net80833, net119976,
         net119953, \ab[4][16] , \SUMB[3][17] , \CARRYB[3][16] , net93800,
         net89356, net88943, net88881, net88880, net87066, net81372, net83057,
         net83055, net83054, net80927, net123363, net121770, net121452,
         net121451, net121450, net121449, \SUMB[25][3] , net82162, net82161,
         net82160, \ab[14][10] , \CARRYB[14][10] , \CARRYB[13][10] ,
         \CARRYB[12][10] , net93277, net120649, \SUMB[13][11] , net88906,
         net84349, net81560, net81559, net87937, net87936, net87935, net87934,
         net84059, net82158, net120648, net120647, net84001, net84000,
         net124635, \ab[24][4] , \CARRYB[23][4] , net87681, net81555, net81553,
         net81552, net81042, net93683, net93279, net90818, net90022, net88699,
         net87950, net87949, net87391, net123293, net123291, net89110,
         net89104, net89103, net85094, net79882, net79881, net79880,
         \CARRYB[28][1] , net124610, \ab[1][7] , \ab[0][8] , net125691,
         \SUMB[5][5] , \SUMB[4][6] , net88199, net88198, \ab[7][4] ,
         \SUMB[8][3] , \CARRYB[8][3] , \CARRYB[7][3] , \ab[1][8] , net89958,
         \ab[5][5] , net88776, net85903, net85902, net122156, \ab[24][1] ,
         \SUMB[24][1] , \SUMB[23][2] , \ab[11][2] , \SUMB[10][3] , net88200,
         \ab[8][4] , \SUMB[8][4] , \SUMB[7][5] , \SUMB[7][4] , \SUMB[6][5] ,
         \CARRYB[8][4] , \CARRYB[7][4] , \CARRYB[6][4] , net86135, net86134,
         \ab[15][1] , \ab[14][2] , \SUMB[15][1] , \SUMB[14][2] , \SUMB[13][3] ,
         \CARRYB[15][1] , \CARRYB[14][1] , \CARRYB[13][2] , \ab[2][6] ,
         \ab[0][7] , \SUMB[1][7] , \CARRYB[2][6] , net93676, net81097,
         net81095, \ab[19][1] , \SUMB[18][2] , \CARRYB[19][1] , net82543,
         net82542, net82541, \ab[23][1] , \SUMB[22][2] , \CARRYB[23][1] ,
         \CARRYB[22][1] , \ab[16][1] , \SUMB[17][2] , \SUMB[16][1] ,
         \SUMB[15][2] , \CARRYB[18][1] , \CARRYB[17][1] , \CARRYB[16][1] ,
         net86131, net86129, net85032, net122130, \ab[13][1] , \ab[12][1] ,
         \SUMB[12][2] , \SUMB[12][1] , \SUMB[11][2] , \CARRYB[13][1] ,
         \CARRYB[12][1] , \CARRYB[11][1] , net87962, net87961, net84929,
         net84928, net77976, \ab[2][7] , \SUMB[3][6] , \SUMB[2][7] ,
         \SUMB[1][8] , \CARRYB[4][5] , \CARRYB[3][5] , \CARRYB[2][7] ,
         \CARRYB[1][7] , \*UDW_*112734/net78687 , net147451, net147444,
         net147421, net147940, net147939, net147938, net147936, net147930,
         net147929, net147928, net147922, net147920, net147999, net147998,
         net148015, net148053, net148051, net148179, net148235, net148233,
         net148230, net148302, net148582, net148754, net149004, net149526,
         net149530, net149580, net149605, net149611, net149917, net149916,
         net88856, net84374, net83776, \SUMB[18][7] , \SUMB[17][8] ,
         \SUMB[20][6] , net80511, net80509, \ab[22][3] , \CARRYB[20][3] ,
         net124949, \ab[24][3] , net84327, \SUMB[1][18] , net119952, net119901,
         net119899, \ab[0][17] , \CARRYB[1][16] , \*UDW_*112689/net78561 ,
         net92337, net86055, net81158, \ab[29][1] , \SUMB[28][2] , \ab[27][1] ,
         net84946, net84945, \CARRYB[4][14] , net83536, net36614, \ab[30][0] ,
         \ab[21][5] , net84856, net84446, net82297, \ab[6][14] , \SUMB[5][15] ,
         \SUMB[4][16] , net81630, net77988, \*UDW_*112684/net78549 , net90897,
         net90348, net88660, \SUMB[6][14] , \CARRYB[6][14] , \CARRYB[5][14] ,
         net83977, net83976, net83975, \SUMB[24][2] , \CARRYB[25][1] ,
         net81269, net80541, net80540, \SUMB[17][7] , \CARRYB[16][6] ,
         net92790, \SUMB[25][2] , \ab[17][6] , \ab[9][12] , net87050, net86959,
         net85688, net82286, \ab[1][17] , \SUMB[10][11] , net93914, net90810,
         net82009, net81947, net81270, net81268, net124627, \ab[19][6] ,
         net82405, net77904, net70444, net120626, \ab[20][5] , \SUMB[19][6] ,
         \CARRYB[20][5] , net89149, net88841, net85461, net85460, net85459,
         net84870, net84868, net84867, net84672, net84671, net84670, net84669,
         net82837, net81375, net81374, net81373, \SUMB[8][13] , net91003,
         net87367, net87366, net87365, net87364, net83876, net82838, net77864,
         net70436, \CARRYB[28][0] , net80564, net84873, net83882, net83881,
         net83880, net121898, \ab[12][10] , \CARRYB[11][10] , net80773,
         net80771, \SUMB[27][1] , \CARRYB[27][0] , net91377, net90576,
         net88878, net86806, net85611, net85610, net82748, net82404, net82403,
         net81264, net124589, net120625, \SUMB[18][6] , \SUMB[17][6] ,
         \CARRYB[17][6] , net92622, net86145, net86144, net86142, net83848,
         net82295, net82294, net82292, net81182, \SUMB[12][10] ,
         \CARRYB[12][9] , net92553, net92552, net92551, net92550, net89840,
         net89447, net89369, net89167, net88303, net88302, net87043, net85539,
         net85537, net84874, net81165, \SUMB[11][11] , \CARRYB[10][11] ,
         net92569, net92568, net88665, net86520, net86519, \ab[23][3] ,
         \SUMB[22][4] , \CARRYB[24][2] , \CARRYB[22][3] , \CARRYB[21][3] ,
         net80848, net80847, net70458, \ab[8][12] , \SUMB[7][13] ,
         \CARRYB[8][12] , \CARRYB[7][12] , net82152, net123752, net119951,
         net119928, net89652, net87363, net148829, net148828, \ab[14][8] ,
         \SUMB[13][9] , net86375, net86374, net80538, net80537, net80536,
         net77916, net70448, \ab[16][7] , \CARRYB[15][7] , net123269,
         net123268, net123267, net123266, net119974, net119960, net119955,
         net119910, net119909, net89455, net88648, net86109, net85109,
         net84668, net84667, net84666, net83101, net120366, net120364,
         \ab[22][5] , \SUMB[23][4] , \SUMB[22][5] , \SUMB[21][6] ,
         \CARRYB[22][5] , net85372, net82289, net82288, net80906,
         \SUMB[16][7] , net89460, net83625, net83624, net83623, net81867,
         net80986, net123365, net83705, net80862, net149133, net147926,
         net147925, net147924, \SUMB[21][5] , net88904, net86537, net86536,
         net83273, net81668, net81667, net81666, \SUMB[15][8] , \SUMB[14][9] ,
         \SUMB[14][8] , \CARRYB[14][8] , net83918, net148838, net148837,
         net148836, net119948, net119927, net119908, \ab[5][14] , net92331,
         net92330, net87798, net86792, net85287, net79885, net79884, net79883,
         \ab[28][1] , net87396, \ab[1][15] , \ab[8][10] , net89168, net122062,
         \SUMB[12][9] , \CARRYB[13][8] , \CARRYB[7][10] , \ab[3][13] ,
         \ab[1][13] , \ab[0][15] , net91419, net84656, net84654, \ab[11][9] ,
         net93307, net93306, net93305, net93304, net90735, net84268, net84267,
         \CARRYB[10][9] , net84072, net84069, net83042, \SUMB[9][11] ,
         \SUMB[10][10] , net91259, net84071, net84070, net77984, net70493,
         \ab[1][14] , net86151, \ab[6][11] , net89537, net121447, net121446,
         net121445, \ab[12][8] , \CARRYB[11][8] , net81216, net81215,
         \ab[9][10] , \SUMB[8][11] , \CARRYB[8][10] , net88104, net81116,
         net81115, net80507, net80506, net80505, net77922, net70450,
         \ab[13][8] , \SUMB[11][9] , \CARRYB[12][8] , net91298, net87459,
         net87458, net87457, net87456, net83062, net83061, net81643, net81256,
         net81001, \ab[10][10] , \CARRYB[9][10] , \SUMB[7][11] , net70462,
         net124833, net120392, net120391, \ab[2][13] , \ab[0][14] ,
         \SUMB[1][14] , \CARRYB[2][13] , \CARRYB[1][13] ,
         \*UDW_*112699/net78591 , net88085, net88084, net82763, net82762,
         net124527, \ab[5][11] , \SUMB[4][12] , \CARRYB[5][11] ,
         \CARRYB[4][11] , net84652, \ab[7][11] , \SUMB[5][12] ,
         \CARRYB[6][11] , net89227, net88010, net85493, net84270, net81694,
         net81416, net70466, \ab[0][16] , \SUMB[3][13] , \SUMB[1][15] ,
         \CARRYB[1][14] , \*UDW_*112699/net78589 , net89021, net88107,
         net88106, net88105, net87462, net87461, net87460, net83045, net81209,
         \SUMB[6][12] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378;

  FA_X1 S2_13_18 ( .A(\ab[13][18] ), .B(\CARRYB[12][18] ), .CI(\SUMB[12][19] ), 
        .S(\SUMB[13][18] ) );
  FA_X1 S2_12_18 ( .A(\ab[12][18] ), .B(\CARRYB[11][18] ), .CI(\SUMB[11][19] ), 
        .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FA_X1 S2_12_19 ( .A(\ab[12][19] ), .B(\CARRYB[11][19] ), .CI(\SUMB[11][20] ), 
        .S(\SUMB[12][19] ) );
  FA_X1 S2_11_6 ( .A(\CARRYB[10][6] ), .B(\ab[11][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA_X1 S2_11_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(\SUMB[10][20] ), 
        .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FA_X1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(PRODUCT[10]) );
  FA_X1 S2_10_5 ( .A(\CARRYB[9][5] ), .B(\ab[10][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA_X1 S2_10_7 ( .A(\CARRYB[9][7] ), .B(\ab[10][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(PRODUCT[9]) );
  FA_X1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA_X1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(PRODUCT[8]) );
  FA_X1 S2_8_2 ( .A(\CARRYB[7][2] ), .B(\ab[8][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA_X1 S2_8_5 ( .A(\CARRYB[7][5] ), .B(\ab[8][5] ), .CI(n2375), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_8_21 ( .A(\ab[8][21] ), .B(\CARRYB[7][21] ), .CI(\SUMB[7][22] ), 
        .CO(\CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FA_X1 S2_8_23 ( .A(\ab[8][23] ), .B(\CARRYB[7][23] ), .CI(\SUMB[7][24] ), 
        .S(\SUMB[8][23] ) );
  FA_X1 S1_7_0 ( .A(\ab[7][0] ), .B(\SUMB[6][1] ), .CI(\CARRYB[6][0] ), .CO(
        \CARRYB[7][0] ), .S(PRODUCT[7]) );
  FA_X1 S2_7_2 ( .A(\CARRYB[6][2] ), .B(\ab[7][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA_X1 S2_7_24 ( .A(\ab[7][24] ), .B(\CARRYB[6][24] ), .CI(\SUMB[6][25] ), 
        .S(\SUMB[7][24] ) );
  FA_X1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(PRODUCT[6]) );
  FA_X1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA_X1 S2_6_9 ( .A(\CARRYB[5][9] ), .B(\ab[6][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA_X1 S2_6_22 ( .A(\CARRYB[5][22] ), .B(\ab[6][22] ), .CI(\SUMB[5][23] ), 
        .CO(\CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FA_X1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(PRODUCT[5]) );
  FA_X1 S2_5_2 ( .A(\CARRYB[4][2] ), .B(\ab[5][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA_X1 S2_5_4 ( .A(\CARRYB[4][4] ), .B(\ab[5][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA_X1 S2_5_6 ( .A(\CARRYB[4][6] ), .B(\ab[5][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .CI(n1185), .CO(
        \CARRYB[5][24] ), .S(\SUMB[5][24] ) );
  FA_X1 S1_4_0 ( .A(\CARRYB[3][0] ), .B(\ab[4][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(PRODUCT[4]) );
  FA_X1 S2_4_2 ( .A(\CARRYB[3][2] ), .B(\ab[4][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA_X1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA_X1 S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .CI(\SUMB[3][27] ), 
        .CO(\CARRYB[4][26] ), .S(\SUMB[4][26] ) );
  FA_X1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(PRODUCT[3]) );
  FA_X1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA_X1 S2_3_2 ( .A(\CARRYB[2][2] ), .B(\ab[3][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA_X1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA_X1 S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .CI(\SUMB[2][29] ), 
        .S(\SUMB[3][28] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(n40), .CO(
        \CARRYB[2][0] ), .S(PRODUCT[2]) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(n41), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(n43), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA_X1 S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA_X1 S2_2_26 ( .A(\ab[2][26] ), .B(\CARRYB[1][26] ), .CI(\SUMB[1][27] ), 
        .CO(\CARRYB[2][26] ), .S(\SUMB[2][26] ) );
  FA_X1 S2_2_27 ( .A(\ab[2][27] ), .B(n44), .CI(\SUMB[1][28] ), .CO(
        \CARRYB[2][27] ), .S(\SUMB[2][27] ) );
  FA_X1 S2_2_29 ( .A(\ab[2][29] ), .B(n42), .CI(n355), .S(\SUMB[2][29] ) );
  FA_X1 S2_6_21 ( .A(\CARRYB[5][21] ), .B(\ab[6][21] ), .CI(\SUMB[5][22] ), 
        .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FA_X1 S2_12_15 ( .A(\CARRYB[11][15] ), .B(\ab[12][15] ), .CI(\SUMB[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA_X1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA_X1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA_X1 S2_20_3 ( .A(\SUMB[19][4] ), .B(\ab[20][3] ), .CI(\CARRYB[19][3] ), 
        .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FA_X1 S2_6_14 ( .A(\SUMB[5][15] ), .B(\ab[6][14] ), .CI(\CARRYB[5][14] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA_X1 S2_22_5 ( .A(\CARRYB[21][5] ), .B(\ab[22][5] ), .CI(\SUMB[21][6] ), 
        .CO(\CARRYB[22][5] ), .S(\SUMB[22][5] ) );
  FA_X1 S2_17_6 ( .A(\CARRYB[16][6] ), .B(\ab[17][6] ), .CI(\SUMB[16][7] ), 
        .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FA_X1 S2_14_8 ( .A(\SUMB[13][9] ), .B(\ab[14][8] ), .CI(\CARRYB[13][8] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  INV_X4 U2 ( .A(\CARRYB[10][12] ), .ZN(net83629) );
  INV_X2 U3 ( .A(net85094), .ZN(net148179) );
  NAND2_X2 U4 ( .A1(net89453), .A2(\ab[30][0] ), .ZN(net80473) );
  NAND2_X2 U5 ( .A1(\SUMB[13][11] ), .A2(\CARRYB[13][10] ), .ZN(net82162) );
  NAND2_X2 U6 ( .A1(net123427), .A2(\ab[26][3] ), .ZN(n2116) );
  NAND2_X2 U7 ( .A1(\CARRYB[29][1] ), .A2(net81548), .ZN(n836) );
  NAND2_X2 U8 ( .A1(net86024), .A2(net86023), .ZN(n3) );
  NAND2_X4 U9 ( .A1(n534), .A2(n535), .ZN(n4) );
  NAND2_X2 U10 ( .A1(\ab[5][17] ), .A2(\SUMB[4][18] ), .ZN(n2202) );
  NAND2_X1 U11 ( .A1(\ab[23][7] ), .A2(n949), .ZN(net86413) );
  NAND2_X2 U12 ( .A1(n399), .A2(net86629), .ZN(n1412) );
  INV_X2 U13 ( .A(\CARRYB[16][7] ), .ZN(n5) );
  INV_X2 U14 ( .A(n5), .ZN(n6) );
  INV_X8 U16 ( .A(\CARRYB[8][9] ), .ZN(n1172) );
  INV_X2 U18 ( .A(\CARRYB[24][3] ), .ZN(net121450) );
  NAND2_X2 U19 ( .A1(\CARRYB[24][3] ), .A2(\ab[25][3] ), .ZN(net81007) );
  NAND2_X4 U20 ( .A1(net123303), .A2(\ab[4][16] ), .ZN(net80835) );
  NAND2_X2 U21 ( .A1(n1323), .A2(\SUMB[12][14] ), .ZN(n87) );
  INV_X2 U22 ( .A(\SUMB[18][6] ), .ZN(n7) );
  INV_X4 U23 ( .A(n7), .ZN(n8) );
  INV_X8 U24 ( .A(\CARRYB[3][16] ), .ZN(n654) );
  NAND2_X2 U25 ( .A1(\ab[3][22] ), .A2(\CARRYB[2][22] ), .ZN(n1068) );
  CLKBUF_X3 U26 ( .A(net87411), .Z(net86385) );
  XNOR2_X2 U27 ( .A(\CARRYB[24][2] ), .B(n10), .ZN(n9) );
  INV_X32 U28 ( .A(\ab[25][2] ), .ZN(n10) );
  NAND2_X4 U31 ( .A1(net148302), .A2(net149605), .ZN(n626) );
  NAND2_X2 U32 ( .A1(n476), .A2(net85287), .ZN(n14) );
  NAND2_X4 U33 ( .A1(n12), .A2(n13), .ZN(n15) );
  NAND2_X4 U34 ( .A1(n14), .A2(n15), .ZN(net86792) );
  INV_X4 U36 ( .A(net85287), .ZN(n13) );
  INV_X16 U37 ( .A(B[16]), .ZN(net70466) );
  NAND2_X2 U38 ( .A1(net82255), .A2(\SUMB[19][10] ), .ZN(net81035) );
  INV_X2 U39 ( .A(net89110), .ZN(net148015) );
  XNOR2_X2 U41 ( .A(n360), .B(\SUMB[20][1] ), .ZN(PRODUCT[21]) );
  CLKBUF_X3 U42 ( .A(\SUMB[17][1] ), .Z(n16) );
  NAND3_X2 U43 ( .A1(n1969), .A2(n1968), .A3(n1967), .ZN(n17) );
  NAND2_X2 U44 ( .A1(\CARRYB[13][2] ), .A2(\SUMB[13][3] ), .ZN(net81781) );
  XOR2_X2 U45 ( .A(n1808), .B(n16), .Z(PRODUCT[18]) );
  XNOR2_X2 U46 ( .A(n18), .B(n1280), .ZN(PRODUCT[22]) );
  XNOR2_X2 U47 ( .A(\ab[22][0] ), .B(\CARRYB[21][0] ), .ZN(n18) );
  NAND3_X2 U48 ( .A1(n1995), .A2(n1996), .A3(n1997), .ZN(n19) );
  CLKBUF_X2 U49 ( .A(\CARRYB[19][2] ), .Z(n20) );
  NAND2_X2 U50 ( .A1(\CARRYB[13][4] ), .A2(\SUMB[13][5] ), .ZN(n2150) );
  NAND2_X2 U51 ( .A1(\CARRYB[19][2] ), .A2(\SUMB[19][3] ), .ZN(n1916) );
  NAND2_X2 U52 ( .A1(\ab[6][3] ), .A2(\CARRYB[5][3] ), .ZN(n1566) );
  XNOR2_X2 U53 ( .A(n425), .B(n21), .ZN(\SUMB[20][1] ) );
  INV_X4 U54 ( .A(\SUMB[19][2] ), .ZN(n21) );
  XNOR2_X2 U55 ( .A(\SUMB[17][2] ), .B(\ab[18][1] ), .ZN(n396) );
  INV_X2 U56 ( .A(n36), .ZN(n962) );
  NAND3_X4 U57 ( .A1(n732), .A2(n733), .A3(n734), .ZN(\CARRYB[3][5] ) );
  NAND2_X2 U58 ( .A1(\CARRYB[21][0] ), .A2(\SUMB[21][1] ), .ZN(n1798) );
  INV_X4 U59 ( .A(n962), .ZN(n963) );
  XNOR2_X2 U60 ( .A(n22), .B(n963), .ZN(PRODUCT[23]) );
  XNOR2_X2 U61 ( .A(\SUMB[22][1] ), .B(\ab[23][0] ), .ZN(n22) );
  XNOR2_X2 U62 ( .A(net93713), .B(net83358), .ZN(n23) );
  CLKBUF_X2 U63 ( .A(\SUMB[18][3] ), .Z(n24) );
  XNOR2_X2 U64 ( .A(n2171), .B(net122087), .ZN(n25) );
  XNOR2_X2 U66 ( .A(n2026), .B(n1134), .ZN(PRODUCT[26]) );
  XNOR2_X2 U68 ( .A(n27), .B(n597), .ZN(PRODUCT[25]) );
  XNOR2_X2 U69 ( .A(\CARRYB[24][0] ), .B(\ab[25][0] ), .ZN(n27) );
  INV_X8 U70 ( .A(net70491), .ZN(net77976) );
  NAND2_X2 U71 ( .A1(n1973), .A2(n1308), .ZN(n226) );
  XNOR2_X2 U72 ( .A(n28), .B(\ab[26][0] ), .ZN(n2026) );
  INV_X4 U73 ( .A(n940), .ZN(n28) );
  XNOR2_X2 U74 ( .A(\CARRYB[26][0] ), .B(\ab[27][0] ), .ZN(n192) );
  INV_X2 U75 ( .A(\CARRYB[11][6] ), .ZN(n1192) );
  INV_X4 U76 ( .A(n47), .ZN(n29) );
  INV_X4 U77 ( .A(net120359), .ZN(n30) );
  INV_X4 U78 ( .A(\CARRYB[25][2] ), .ZN(net120359) );
  INV_X4 U79 ( .A(\SUMB[20][4] ), .ZN(net148233) );
  NOR2_X4 U80 ( .A1(net70450), .A2(net86101), .ZN(\ab[1][8] ) );
  NOR2_X4 U81 ( .A1(net70460), .A2(n331), .ZN(net124833) );
  INV_X8 U82 ( .A(net77976), .ZN(n331) );
  NAND2_X2 U83 ( .A1(\SUMB[2][12] ), .A2(\CARRYB[2][11] ), .ZN(n2028) );
  NAND2_X2 U84 ( .A1(n248), .A2(n249), .ZN(n251) );
  NAND2_X2 U85 ( .A1(net124949), .A2(\SUMB[21][4] ), .ZN(n503) );
  NAND2_X4 U86 ( .A1(n1024), .A2(n1025), .ZN(n2335) );
  NAND2_X2 U87 ( .A1(n1764), .A2(n371), .ZN(n254) );
  NAND2_X2 U88 ( .A1(net123897), .A2(net123898), .ZN(n872) );
  CLKBUF_X3 U89 ( .A(\SUMB[6][15] ), .Z(net93800) );
  NAND2_X1 U90 ( .A1(net88881), .A2(\SUMB[6][15] ), .ZN(net81367) );
  INV_X4 U91 ( .A(\ab[4][12] ), .ZN(n316) );
  XNOR2_X2 U92 ( .A(\CARRYB[13][17] ), .B(n31), .ZN(n1532) );
  OR2_X4 U93 ( .A1(net70467), .A2(net123000), .ZN(n31) );
  INV_X8 U94 ( .A(n1196), .ZN(n1197) );
  XNOR2_X2 U95 ( .A(\SUMB[7][20] ), .B(net86231), .ZN(n32) );
  INV_X2 U96 ( .A(\SUMB[2][23] ), .ZN(n33) );
  INV_X4 U97 ( .A(n33), .ZN(n34) );
  NAND2_X1 U98 ( .A1(\ab[9][19] ), .A2(\SUMB[8][20] ), .ZN(n2290) );
  CLKBUF_X2 U99 ( .A(\CARRYB[13][1] ), .Z(n35) );
  NAND3_X2 U100 ( .A1(n1796), .A2(n1797), .A3(n1798), .ZN(n36) );
  XNOR2_X2 U101 ( .A(n2112), .B(\SUMB[5][18] ), .ZN(n37) );
  XNOR2_X2 U102 ( .A(\SUMB[11][14] ), .B(n1753), .ZN(n38) );
  NOR2_X4 U103 ( .A1(net88344), .A2(net77964), .ZN(n817) );
  AND2_X2 U104 ( .A1(\ab[1][24] ), .A2(\ab[0][25] ), .ZN(n39) );
  NOR2_X2 U106 ( .A1(net81673), .A2(net77892), .ZN(n870) );
  INV_X4 U107 ( .A(net92311), .ZN(\ab[28][2] ) );
  NAND2_X4 U108 ( .A1(\ab[5][22] ), .A2(\CARRYB[4][22] ), .ZN(net80794) );
  XOR2_X2 U109 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(n40) );
  AND2_X2 U110 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .ZN(n41) );
  NOR2_X1 U111 ( .A1(net77914), .A2(net70451), .ZN(\ab[22][7] ) );
  INV_X8 U112 ( .A(n406), .ZN(n420) );
  INV_X2 U113 ( .A(\ab[24][5] ), .ZN(n2195) );
  NOR2_X1 U114 ( .A1(net77898), .A2(net70447), .ZN(\ab[24][5] ) );
  AND2_X2 U115 ( .A1(\ab[0][30] ), .A2(\ab[1][29] ), .ZN(n42) );
  NAND2_X2 U116 ( .A1(\ab[5][7] ), .A2(\CARRYB[4][7] ), .ZN(n143) );
  NAND2_X4 U117 ( .A1(\ab[4][8] ), .A2(\CARRYB[3][8] ), .ZN(n1944) );
  AND2_X2 U118 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .ZN(n43) );
  AND2_X2 U119 ( .A1(\ab[0][28] ), .A2(\ab[1][27] ), .ZN(n44) );
  INV_X4 U120 ( .A(net70458), .ZN(n491) );
  INV_X8 U121 ( .A(n452), .ZN(\CARRYB[1][13] ) );
  AND3_X4 U122 ( .A1(n2007), .A2(n2008), .A3(n2009), .ZN(n45) );
  NAND2_X4 U123 ( .A1(\CARRYB[11][4] ), .A2(\ab[12][4] ), .ZN(n667) );
  INV_X8 U124 ( .A(n194), .ZN(\SUMB[10][6] ) );
  NAND2_X4 U125 ( .A1(\ab[2][15] ), .A2(\CARRYB[1][15] ), .ZN(n1984) );
  NAND2_X4 U126 ( .A1(\CARRYB[9][9] ), .A2(\ab[10][9] ), .ZN(n325) );
  NAND2_X4 U127 ( .A1(net85602), .A2(net85603), .ZN(\SUMB[2][18] ) );
  NAND2_X4 U128 ( .A1(n1127), .A2(n1128), .ZN(n1256) );
  INV_X4 U129 ( .A(net89168), .ZN(net123142) );
  NAND2_X4 U130 ( .A1(\CARRYB[15][5] ), .A2(\ab[16][5] ), .ZN(n2071) );
  XOR2_X2 U131 ( .A(net88881), .B(\ab[7][14] ), .Z(n46) );
  INV_X8 U132 ( .A(net88878), .ZN(\SUMB[18][6] ) );
  NAND3_X4 U133 ( .A1(net81267), .A2(net81266), .A3(net81265), .ZN(net87619)
         );
  NAND2_X4 U134 ( .A1(\ab[16][9] ), .A2(\CARRYB[15][9] ), .ZN(n805) );
  INV_X8 U135 ( .A(\SUMB[12][12] ), .ZN(net120648) );
  NAND2_X4 U136 ( .A1(n391), .A2(n384), .ZN(n390) );
  NAND2_X2 U137 ( .A1(\ab[20][9] ), .A2(\CARRYB[19][9] ), .ZN(net81033) );
  NAND2_X4 U138 ( .A1(n1511), .A2(n1510), .ZN(n1190) );
  NAND2_X4 U139 ( .A1(n2156), .A2(n2157), .ZN(n896) );
  NAND2_X4 U141 ( .A1(\ab[12][13] ), .A2(\CARRYB[11][13] ), .ZN(n1795) );
  NAND2_X2 U142 ( .A1(net93813), .A2(\ab[24][4] ), .ZN(net79908) );
  NAND2_X2 U143 ( .A1(n312), .A2(\ab[9][5] ), .ZN(n1786) );
  INV_X4 U144 ( .A(\CARRYB[1][18] ), .ZN(n709) );
  NAND2_X4 U145 ( .A1(net87949), .A2(net87950), .ZN(n311) );
  NAND2_X4 U146 ( .A1(\SUMB[16][9] ), .A2(net93410), .ZN(n812) );
  NAND2_X2 U147 ( .A1(n1765), .A2(\SUMB[2][21] ), .ZN(n1433) );
  XNOR2_X2 U149 ( .A(net93203), .B(n1901), .ZN(\SUMB[5][14] ) );
  INV_X8 U150 ( .A(B[19]), .ZN(net70472) );
  NAND2_X2 U151 ( .A1(\ab[25][4] ), .A2(net90433), .ZN(n2113) );
  NAND2_X2 U152 ( .A1(\CARRYB[1][14] ), .A2(\ab[2][14] ), .ZN(net86172) );
  INV_X2 U153 ( .A(\CARRYB[4][8] ), .ZN(n1514) );
  INV_X1 U154 ( .A(net84000), .ZN(net84434) );
  NAND3_X2 U155 ( .A1(n738), .A2(n739), .A3(n740), .ZN(\CARRYB[11][1] ) );
  NAND2_X1 U156 ( .A1(\ab[15][1] ), .A2(\SUMB[14][2] ), .ZN(n652) );
  BUF_X4 U157 ( .A(\SUMB[4][10] ), .Z(n1258) );
  BUF_X8 U158 ( .A(\SUMB[3][10] ), .Z(n1259) );
  NAND2_X2 U159 ( .A1(\ab[14][3] ), .A2(\SUMB[13][4] ), .ZN(n1968) );
  NAND2_X2 U161 ( .A1(\SUMB[23][5] ), .A2(net84434), .ZN(net79909) );
  NAND2_X1 U162 ( .A1(\CARRYB[5][7] ), .A2(n1313), .ZN(n49) );
  NAND2_X4 U163 ( .A1(n47), .A2(n48), .ZN(n50) );
  NAND2_X2 U164 ( .A1(n49), .A2(n50), .ZN(n1329) );
  INV_X4 U165 ( .A(\CARRYB[5][7] ), .ZN(n47) );
  INV_X4 U166 ( .A(n1313), .ZN(n48) );
  NAND3_X2 U167 ( .A1(n1673), .A2(n1674), .A3(n1675), .ZN(n51) );
  NAND2_X2 U168 ( .A1(\SUMB[3][10] ), .A2(\CARRYB[3][9] ), .ZN(n1963) );
  NAND2_X1 U169 ( .A1(\CARRYB[22][7] ), .A2(\ab[23][7] ), .ZN(n54) );
  NAND2_X2 U170 ( .A1(n52), .A2(n53), .ZN(n55) );
  NAND2_X2 U171 ( .A1(n54), .A2(n55), .ZN(net88961) );
  INV_X1 U172 ( .A(\CARRYB[22][7] ), .ZN(n52) );
  INV_X1 U173 ( .A(\ab[23][7] ), .ZN(n53) );
  NAND3_X2 U174 ( .A1(n2241), .A2(n2240), .A3(n2242), .ZN(n56) );
  XNOR2_X2 U175 ( .A(\ab[2][21] ), .B(\CARRYB[1][21] ), .ZN(n57) );
  NAND2_X2 U176 ( .A1(net87009), .A2(\SUMB[17][11] ), .ZN(n60) );
  INV_X4 U179 ( .A(net87009), .ZN(n58) );
  INV_X4 U180 ( .A(\SUMB[17][11] ), .ZN(n59) );
  NOR2_X2 U181 ( .A1(net77912), .A2(net70449), .ZN(\ab[23][7] ) );
  NAND2_X2 U182 ( .A1(\SUMB[4][20] ), .A2(\ab[5][19] ), .ZN(n2241) );
  NAND2_X4 U183 ( .A1(\SUMB[2][14] ), .A2(n99), .ZN(net81513) );
  NAND3_X2 U184 ( .A1(net82667), .A2(net82668), .A3(net82669), .ZN(
        \CARRYB[19][10] ) );
  NAND2_X4 U185 ( .A1(net80657), .A2(net80658), .ZN(net80660) );
  NAND2_X4 U186 ( .A1(net123055), .A2(n927), .ZN(n928) );
  NAND2_X2 U187 ( .A1(\ab[8][18] ), .A2(n1109), .ZN(n1105) );
  NAND2_X2 U188 ( .A1(\ab[14][15] ), .A2(\SUMB[13][16] ), .ZN(n1871) );
  NAND2_X4 U189 ( .A1(\SUMB[1][15] ), .A2(\CARRYB[1][14] ), .ZN(net86171) );
  INV_X4 U190 ( .A(\CARRYB[8][16] ), .ZN(n1599) );
  NAND2_X1 U191 ( .A1(net90702), .A2(\CARRYB[6][17] ), .ZN(n932) );
  INV_X2 U192 ( .A(\CARRYB[4][18] ), .ZN(n1767) );
  INV_X4 U193 ( .A(n1927), .ZN(n1524) );
  NAND2_X4 U194 ( .A1(n216), .A2(n217), .ZN(n219) );
  NAND2_X4 U195 ( .A1(\SUMB[14][6] ), .A2(\ab[15][5] ), .ZN(n1978) );
  NAND2_X2 U196 ( .A1(\ab[1][17] ), .A2(net85688), .ZN(net82286) );
  INV_X8 U197 ( .A(net83736), .ZN(net121606) );
  BUF_X8 U198 ( .A(\SUMB[7][11] ), .Z(net120922) );
  NAND2_X4 U199 ( .A1(n1562), .A2(n94), .ZN(n911) );
  NAND2_X2 U200 ( .A1(net83705), .A2(n71), .ZN(n64) );
  NAND2_X4 U201 ( .A1(n62), .A2(n63), .ZN(n65) );
  NAND2_X4 U202 ( .A1(n64), .A2(n65), .ZN(n366) );
  INV_X4 U203 ( .A(net83705), .ZN(n62) );
  INV_X4 U204 ( .A(n71), .ZN(n63) );
  BUF_X4 U205 ( .A(\SUMB[20][6] ), .Z(n71) );
  NAND2_X2 U206 ( .A1(n366), .A2(net86464), .ZN(n2302) );
  NAND2_X4 U207 ( .A1(n148), .A2(n149), .ZN(net82154) );
  NOR2_X4 U208 ( .A1(n392), .A2(n2355), .ZN(\ab[0][27] ) );
  NAND2_X2 U209 ( .A1(n1598), .A2(n1597), .ZN(n91) );
  CLKBUF_X2 U210 ( .A(\SUMB[25][4] ), .Z(net83030) );
  NAND2_X2 U211 ( .A1(\SUMB[25][4] ), .A2(\ab[26][3] ), .ZN(net81052) );
  NAND2_X4 U212 ( .A1(n1271), .A2(\SUMB[10][6] ), .ZN(n2061) );
  NAND2_X2 U213 ( .A1(\SUMB[13][5] ), .A2(\ab[14][4] ), .ZN(n2151) );
  XNOR2_X2 U214 ( .A(\CARRYB[20][4] ), .B(n945), .ZN(n66) );
  CLKBUF_X2 U215 ( .A(\SUMB[6][11] ), .Z(net149004) );
  NAND3_X4 U216 ( .A1(n1874), .A2(n1875), .A3(n1876), .ZN(\CARRYB[10][18] ) );
  NAND2_X2 U218 ( .A1(\SUMB[6][11] ), .A2(\CARRYB[6][10] ), .ZN(n473) );
  INV_X2 U219 ( .A(n1699), .ZN(n67) );
  INV_X4 U220 ( .A(n491), .ZN(n68) );
  NOR2_X4 U221 ( .A1(net70478), .A2(net86101), .ZN(n2196) );
  NAND2_X4 U222 ( .A1(n1385), .A2(net87005), .ZN(net82641) );
  INV_X4 U223 ( .A(net82551), .ZN(net90433) );
  INV_X2 U224 ( .A(net86893), .ZN(n229) );
  OR2_X4 U225 ( .A1(net85251), .A2(n497), .ZN(n494) );
  INV_X1 U226 ( .A(net81553), .ZN(n69) );
  INV_X8 U227 ( .A(\CARRYB[20][6] ), .ZN(net81553) );
  NOR2_X4 U228 ( .A1(net120391), .A2(net80409), .ZN(\ab[1][13] ) );
  INV_X8 U229 ( .A(B[13]), .ZN(net120391) );
  CLKBUF_X3 U230 ( .A(\SUMB[9][11] ), .Z(n70) );
  NAND2_X2 U231 ( .A1(n1742), .A2(n852), .ZN(n240) );
  XNOR2_X2 U232 ( .A(\ab[2][18] ), .B(\CARRYB[1][18] ), .ZN(n397) );
  INV_X8 U233 ( .A(\CARRYB[10][10] ), .ZN(n201) );
  NAND2_X2 U234 ( .A1(\SUMB[26][3] ), .A2(\ab[27][2] ), .ZN(n809) );
  NAND2_X2 U235 ( .A1(\SUMB[23][4] ), .A2(n417), .ZN(net84678) );
  NAND2_X2 U237 ( .A1(\CARRYB[24][0] ), .A2(\SUMB[24][1] ), .ZN(net81530) );
  NAND2_X2 U238 ( .A1(\CARRYB[12][5] ), .A2(\ab[13][5] ), .ZN(n1920) );
  NAND3_X4 U239 ( .A1(net80484), .A2(net80485), .A3(n1058), .ZN(
        \CARRYB[15][13] ) );
  NAND2_X4 U240 ( .A1(\SUMB[14][14] ), .A2(\CARRYB[14][13] ), .ZN(net80485) );
  NAND2_X2 U241 ( .A1(\CARRYB[14][6] ), .A2(\ab[15][6] ), .ZN(n1438) );
  NAND2_X2 U242 ( .A1(\ab[15][13] ), .A2(\SUMB[14][14] ), .ZN(net80484) );
  XNOR2_X2 U243 ( .A(\CARRYB[22][7] ), .B(\ab[23][7] ), .ZN(n867) );
  NAND2_X4 U244 ( .A1(n777), .A2(net87391), .ZN(n72) );
  NAND2_X2 U245 ( .A1(n777), .A2(net87391), .ZN(net87949) );
  INV_X8 U246 ( .A(net90022), .ZN(n777) );
  INV_X8 U247 ( .A(net120625), .ZN(net86806) );
  BUF_X8 U248 ( .A(\SUMB[12][18] ), .Z(n1240) );
  INV_X4 U249 ( .A(\CARRYB[6][22] ), .ZN(n876) );
  NAND2_X2 U250 ( .A1(\CARRYB[21][4] ), .A2(\ab[22][4] ), .ZN(n75) );
  NAND2_X4 U251 ( .A1(n73), .A2(n74), .ZN(n76) );
  NAND2_X4 U252 ( .A1(n76), .A2(n75), .ZN(net80862) );
  INV_X4 U254 ( .A(\ab[22][4] ), .ZN(n74) );
  NAND2_X2 U255 ( .A1(\CARRYB[3][11] ), .A2(\ab[4][11] ), .ZN(net88086) );
  NAND2_X4 U256 ( .A1(n1543), .A2(n1542), .ZN(n362) );
  NAND2_X2 U257 ( .A1(n1845), .A2(n1255), .ZN(n1542) );
  XNOR2_X2 U258 ( .A(\ab[2][18] ), .B(\*UDW_*112679/net78533 ), .ZN(n287) );
  AND2_X4 U259 ( .A1(B[15]), .A2(A[2]), .ZN(\ab[2][15] ) );
  NAND2_X4 U260 ( .A1(n323), .A2(n324), .ZN(n326) );
  INV_X4 U261 ( .A(\CARRYB[9][9] ), .ZN(n323) );
  CLKBUF_X3 U263 ( .A(n1207), .Z(n1324) );
  INV_X2 U264 ( .A(\SUMB[11][13] ), .ZN(n785) );
  NAND2_X2 U265 ( .A1(net85325), .A2(n682), .ZN(n79) );
  NAND2_X4 U266 ( .A1(n77), .A2(n78), .ZN(n80) );
  NAND2_X4 U267 ( .A1(n79), .A2(n80), .ZN(\SUMB[17][10] ) );
  INV_X4 U268 ( .A(net85325), .ZN(n77) );
  INV_X4 U269 ( .A(n682), .ZN(n78) );
  NAND2_X2 U270 ( .A1(n1226), .A2(n556), .ZN(n83) );
  NAND2_X4 U271 ( .A1(n81), .A2(n82), .ZN(n84) );
  NAND2_X4 U272 ( .A1(n83), .A2(n84), .ZN(\SUMB[11][14] ) );
  INV_X4 U273 ( .A(n1226), .ZN(n81) );
  INV_X4 U274 ( .A(n556), .ZN(n82) );
  NAND2_X2 U275 ( .A1(n85), .A2(n86), .ZN(n88) );
  NAND2_X4 U276 ( .A1(n87), .A2(n88), .ZN(\SUMB[13][13] ) );
  INV_X4 U277 ( .A(n1323), .ZN(n85) );
  INV_X2 U278 ( .A(\SUMB[12][14] ), .ZN(n86) );
  INV_X8 U279 ( .A(\SUMB[17][10] ), .ZN(n825) );
  NAND2_X4 U280 ( .A1(n562), .A2(\SUMB[11][14] ), .ZN(n1793) );
  NAND2_X4 U281 ( .A1(\SUMB[13][13] ), .A2(n1345), .ZN(n2120) );
  NAND2_X2 U282 ( .A1(\SUMB[13][13] ), .A2(n134), .ZN(n135) );
  INV_X2 U283 ( .A(\SUMB[13][13] ), .ZN(n133) );
  INV_X8 U284 ( .A(\CARRYB[1][11] ), .ZN(n586) );
  NAND2_X4 U285 ( .A1(\ab[11][4] ), .A2(n563), .ZN(n1833) );
  NAND3_X4 U286 ( .A1(n2104), .A2(n2103), .A3(n2105), .ZN(n176) );
  NAND2_X4 U288 ( .A1(net82029), .A2(n490), .ZN(net82152) );
  NAND3_X2 U289 ( .A1(n2007), .A2(n2008), .A3(n2009), .ZN(n89) );
  NAND2_X4 U291 ( .A1(n641), .A2(n622), .ZN(n624) );
  NAND2_X4 U292 ( .A1(\ab[21][2] ), .A2(n596), .ZN(n2187) );
  NAND3_X4 U293 ( .A1(n1590), .A2(n1747), .A3(n1748), .ZN(\CARRYB[6][10] ) );
  CLKBUF_X3 U294 ( .A(n1425), .Z(n1157) );
  NAND2_X4 U295 ( .A1(\CARRYB[18][3] ), .A2(\ab[19][3] ), .ZN(n2275) );
  NOR2_X4 U296 ( .A1(net92314), .A2(n1181), .ZN(n1182) );
  NAND2_X4 U297 ( .A1(\ab[5][18] ), .A2(\SUMB[4][19] ), .ZN(n2140) );
  INV_X4 U298 ( .A(n1742), .ZN(n238) );
  NAND2_X4 U299 ( .A1(\CARRYB[4][14] ), .A2(net84946), .ZN(net84947) );
  INV_X4 U300 ( .A(n1901), .ZN(n1126) );
  INV_X4 U301 ( .A(net119948), .ZN(n477) );
  INV_X8 U302 ( .A(net119974), .ZN(net119910) );
  NAND2_X4 U303 ( .A1(net84817), .A2(net84818), .ZN(n1743) );
  NOR2_X2 U304 ( .A1(net70486), .A2(net80409), .ZN(\ab[1][26] ) );
  NAND2_X4 U305 ( .A1(\ab[17][10] ), .A2(\SUMB[16][11] ), .ZN(n1580) );
  NAND2_X2 U306 ( .A1(\SUMB[9][16] ), .A2(\CARRYB[9][15] ), .ZN(n1841) );
  NAND2_X2 U307 ( .A1(\ab[10][15] ), .A2(\SUMB[9][16] ), .ZN(n1840) );
  NOR2_X2 U308 ( .A1(net84698), .A2(net77932), .ZN(\ab[7][14] ) );
  INV_X2 U310 ( .A(\SUMB[18][7] ), .ZN(net90576) );
  NOR2_X4 U311 ( .A1(n68), .A2(net70491), .ZN(\ab[2][12] ) );
  NAND2_X4 U312 ( .A1(\ab[17][2] ), .A2(\CARRYB[16][2] ), .ZN(n1668) );
  INV_X2 U313 ( .A(net87396), .ZN(n90) );
  INV_X4 U314 ( .A(net87050), .ZN(\ab[1][17] ) );
  NOR2_X2 U315 ( .A1(net123000), .A2(net82247), .ZN(net149526) );
  NAND2_X1 U316 ( .A1(\CARRYB[3][21] ), .A2(\SUMB[3][22] ), .ZN(n2276) );
  NAND2_X4 U317 ( .A1(n1516), .A2(net90174), .ZN(n1518) );
  NOR2_X4 U318 ( .A1(net70458), .A2(net80409), .ZN(n237) );
  INV_X2 U319 ( .A(\SUMB[7][8] ), .ZN(n1864) );
  NAND2_X4 U320 ( .A1(\SUMB[16][9] ), .A2(\ab[17][8] ), .ZN(n811) );
  NAND2_X1 U321 ( .A1(\ab[13][16] ), .A2(\SUMB[12][17] ), .ZN(n2317) );
  NAND2_X2 U322 ( .A1(\CARRYB[28][0] ), .A2(n344), .ZN(n250) );
  NAND2_X2 U323 ( .A1(\ab[5][10] ), .A2(n181), .ZN(n1746) );
  NAND2_X2 U324 ( .A1(n181), .A2(n228), .ZN(n1745) );
  NAND2_X2 U325 ( .A1(\CARRYB[4][10] ), .A2(\ab[5][10] ), .ZN(n1031) );
  INV_X1 U326 ( .A(net88079), .ZN(n92) );
  INV_X2 U327 ( .A(n92), .ZN(n93) );
  NAND2_X4 U328 ( .A1(n1126), .A2(n174), .ZN(n1127) );
  INV_X2 U329 ( .A(n910), .ZN(n94) );
  INV_X8 U331 ( .A(n917), .ZN(n927) );
  NAND2_X4 U332 ( .A1(net147920), .A2(\ab[5][11] ), .ZN(n677) );
  INV_X2 U333 ( .A(\SUMB[2][15] ), .ZN(n1557) );
  INV_X1 U334 ( .A(n799), .ZN(n95) );
  INV_X4 U335 ( .A(net87936), .ZN(n96) );
  INV_X8 U336 ( .A(n96), .ZN(n97) );
  INV_X8 U337 ( .A(\SUMB[22][7] ), .ZN(n697) );
  NAND2_X4 U338 ( .A1(\ab[9][15] ), .A2(n151), .ZN(n2049) );
  XNOR2_X2 U339 ( .A(\SUMB[15][2] ), .B(n98), .ZN(n646) );
  INV_X32 U340 ( .A(\ab[16][1] ), .ZN(n98) );
  NAND2_X2 U341 ( .A1(\CARRYB[25][2] ), .A2(\ab[26][2] ), .ZN(n1033) );
  NAND2_X2 U342 ( .A1(\ab[17][0] ), .A2(\SUMB[16][1] ), .ZN(net86654) );
  NOR2_X4 U343 ( .A1(net124610), .A2(net77906), .ZN(\ab[0][6] ) );
  INV_X8 U344 ( .A(B[6]), .ZN(net77906) );
  XNOR2_X1 U345 ( .A(\CARRYB[24][1] ), .B(\ab[25][1] ), .ZN(net93880) );
  NAND2_X4 U346 ( .A1(\CARRYB[20][6] ), .A2(net81042), .ZN(n781) );
  NAND3_X2 U347 ( .A1(n454), .A2(n453), .A3(n455), .ZN(n99) );
  INV_X8 U348 ( .A(A[1]), .ZN(net70493) );
  NAND2_X4 U349 ( .A1(n818), .A2(\ab[22][6] ), .ZN(n820) );
  NAND2_X2 U351 ( .A1(\ab[2][17] ), .A2(\*UDW_*112684/net78547 ), .ZN(n1343)
         );
  NAND2_X2 U352 ( .A1(n1882), .A2(net82408), .ZN(n100) );
  NAND2_X2 U353 ( .A1(n101), .A2(net82407), .ZN(net86464) );
  INV_X4 U354 ( .A(n100), .ZN(n101) );
  NAND2_X4 U355 ( .A1(\ab[8][10] ), .A2(\SUMB[7][11] ), .ZN(net81215) );
  NAND2_X4 U356 ( .A1(n280), .A2(n281), .ZN(n283) );
  INV_X4 U357 ( .A(net88648), .ZN(n102) );
  INV_X4 U358 ( .A(\SUMB[22][5] ), .ZN(net88648) );
  NAND2_X4 U359 ( .A1(net86702), .A2(net86703), .ZN(n1401) );
  INV_X4 U360 ( .A(n869), .ZN(net86703) );
  XNOR2_X1 U361 ( .A(net125934), .B(net86801), .ZN(\SUMB[14][11] ) );
  NAND2_X1 U362 ( .A1(\SUMB[13][12] ), .A2(\ab[14][11] ), .ZN(net82557) );
  NAND2_X2 U363 ( .A1(n56), .A2(\ab[6][19] ), .ZN(n979) );
  NAND2_X2 U364 ( .A1(n1272), .A2(\SUMB[26][4] ), .ZN(net80816) );
  NAND2_X4 U365 ( .A1(n1031), .A2(n1032), .ZN(n1658) );
  NAND2_X1 U366 ( .A1(\CARRYB[3][6] ), .A2(\SUMB[3][7] ), .ZN(net88208) );
  NAND2_X4 U367 ( .A1(\ab[16][3] ), .A2(\CARRYB[15][3] ), .ZN(n1131) );
  NAND2_X4 U368 ( .A1(net88177), .A2(\ab[1][9] ), .ZN(n1517) );
  NAND2_X2 U369 ( .A1(\ab[21][0] ), .A2(\SUMB[20][1] ), .ZN(n1806) );
  NOR2_X2 U370 ( .A1(n247), .A2(n103), .ZN(n409) );
  NAND2_X2 U371 ( .A1(n405), .A2(n420), .ZN(n103) );
  INV_X4 U372 ( .A(\SUMB[22][4] ), .ZN(n405) );
  NAND2_X2 U373 ( .A1(\SUMB[22][4] ), .A2(n420), .ZN(n419) );
  OR2_X2 U374 ( .A1(\SUMB[22][4] ), .A2(\ab[23][3] ), .ZN(n422) );
  NAND2_X2 U375 ( .A1(\SUMB[3][9] ), .A2(\ab[4][8] ), .ZN(n1945) );
  NAND2_X4 U376 ( .A1(n1944), .A2(n1328), .ZN(n1551) );
  NAND2_X4 U377 ( .A1(\SUMB[16][3] ), .A2(\CARRYB[16][2] ), .ZN(n1669) );
  INV_X4 U378 ( .A(\CARRYB[2][11] ), .ZN(n913) );
  NAND2_X2 U379 ( .A1(\CARRYB[6][19] ), .A2(\SUMB[6][20] ), .ZN(n1103) );
  BUF_X8 U380 ( .A(net88079), .Z(n137) );
  NAND2_X4 U381 ( .A1(n279), .A2(net123267), .ZN(net120511) );
  NAND3_X4 U382 ( .A1(n1070), .A2(n1069), .A3(n1068), .ZN(\CARRYB[3][22] ) );
  NAND2_X4 U383 ( .A1(net85543), .A2(n484), .ZN(n104) );
  NAND3_X2 U384 ( .A1(net82561), .A2(net82560), .A3(net82559), .ZN(n105) );
  NAND2_X2 U385 ( .A1(\CARRYB[3][17] ), .A2(\ab[4][17] ), .ZN(n108) );
  NAND2_X4 U386 ( .A1(n106), .A2(n107), .ZN(n109) );
  NAND2_X4 U387 ( .A1(n108), .A2(n109), .ZN(n1742) );
  INV_X4 U388 ( .A(\CARRYB[3][17] ), .ZN(n106) );
  INV_X2 U389 ( .A(\ab[4][17] ), .ZN(n107) );
  CLKBUF_X3 U390 ( .A(net91088), .Z(net122062) );
  XNOR2_X2 U391 ( .A(\SUMB[6][21] ), .B(n110), .ZN(\SUMB[7][20] ) );
  XOR2_X2 U392 ( .A(\CARRYB[6][20] ), .B(net81340), .Z(n110) );
  NAND2_X2 U393 ( .A1(net119955), .A2(net119927), .ZN(net148838) );
  NAND2_X2 U394 ( .A1(\ab[16][11] ), .A2(\CARRYB[15][11] ), .ZN(n2097) );
  INV_X2 U395 ( .A(\CARRYB[15][11] ), .ZN(n1733) );
  NAND2_X2 U396 ( .A1(n814), .A2(\SUMB[14][12] ), .ZN(n815) );
  NAND2_X4 U397 ( .A1(n1599), .A2(\ab[9][16] ), .ZN(n1602) );
  NAND2_X2 U398 ( .A1(\CARRYB[7][11] ), .A2(\ab[8][11] ), .ZN(n2128) );
  NAND3_X2 U399 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n111) );
  NOR2_X4 U400 ( .A1(net87396), .A2(net80409), .ZN(n112) );
  INV_X32 U401 ( .A(net77984), .ZN(net80409) );
  NAND2_X4 U403 ( .A1(n700), .A2(n701), .ZN(n703) );
  NAND2_X1 U404 ( .A1(\ab[24][3] ), .A2(n417), .ZN(net84680) );
  INV_X4 U405 ( .A(\CARRYB[13][4] ), .ZN(n1631) );
  INV_X2 U406 ( .A(\SUMB[24][5] ), .ZN(n1596) );
  NAND2_X4 U407 ( .A1(n113), .A2(n114), .ZN(n116) );
  NAND2_X4 U408 ( .A1(n115), .A2(n116), .ZN(net84902) );
  INV_X4 U409 ( .A(\CARRYB[27][2] ), .ZN(n113) );
  INV_X4 U410 ( .A(\ab[28][2] ), .ZN(n114) );
  NAND2_X2 U411 ( .A1(n1658), .A2(\SUMB[4][11] ), .ZN(n119) );
  NAND2_X4 U412 ( .A1(n117), .A2(n118), .ZN(n120) );
  NAND2_X4 U413 ( .A1(n119), .A2(n120), .ZN(\SUMB[5][10] ) );
  INV_X4 U414 ( .A(n1658), .ZN(n117) );
  INV_X4 U415 ( .A(\SUMB[4][11] ), .ZN(n118) );
  NAND2_X2 U416 ( .A1(net84902), .A2(n402), .ZN(n534) );
  INV_X4 U417 ( .A(net84902), .ZN(n533) );
  NAND2_X4 U418 ( .A1(n46), .A2(n230), .ZN(n232) );
  INV_X8 U419 ( .A(n437), .ZN(\SUMB[1][15] ) );
  INV_X2 U420 ( .A(\SUMB[21][8] ), .ZN(n684) );
  NAND2_X1 U421 ( .A1(\SUMB[6][19] ), .A2(\ab[7][18] ), .ZN(net80303) );
  INV_X8 U422 ( .A(\CARRYB[13][12] ), .ZN(n1486) );
  NAND3_X4 U423 ( .A1(n2123), .A2(n2124), .A3(n2125), .ZN(\CARRYB[13][12] ) );
  NAND2_X4 U424 ( .A1(n1242), .A2(\ab[5][16] ), .ZN(n1897) );
  NAND2_X2 U425 ( .A1(\SUMB[12][13] ), .A2(\CARRYB[12][12] ), .ZN(n2123) );
  INV_X4 U426 ( .A(\CARRYB[16][9] ), .ZN(net120655) );
  NAND2_X2 U427 ( .A1(net82152), .A2(net84327), .ZN(n122) );
  NAND2_X4 U429 ( .A1(n123), .A2(n122), .ZN(net119951) );
  NAND2_X2 U431 ( .A1(\ab[1][18] ), .A2(n365), .ZN(n126) );
  NAND2_X4 U432 ( .A1(n124), .A2(n125), .ZN(n127) );
  NAND2_X4 U433 ( .A1(n127), .A2(n126), .ZN(n536) );
  INV_X8 U434 ( .A(\ab[1][18] ), .ZN(n124) );
  INV_X8 U435 ( .A(net81354), .ZN(n125) );
  NAND2_X2 U436 ( .A1(net119928), .A2(net119951), .ZN(net123268) );
  INV_X8 U437 ( .A(net119951), .ZN(net123266) );
  INV_X4 U438 ( .A(net87681), .ZN(net83101) );
  NAND2_X2 U439 ( .A1(\SUMB[13][12] ), .A2(\CARRYB[13][11] ), .ZN(net82558) );
  NAND2_X2 U440 ( .A1(\CARRYB[12][12] ), .A2(\ab[13][12] ), .ZN(n1373) );
  NAND2_X2 U441 ( .A1(n131), .A2(n132), .ZN(net88665) );
  NAND2_X2 U442 ( .A1(net92569), .A2(net88665), .ZN(n498) );
  NAND2_X4 U445 ( .A1(\CARRYB[17][1] ), .A2(\ab[18][1] ), .ZN(n746) );
  XNOR2_X1 U447 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .ZN(n736) );
  XNOR2_X1 U449 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .ZN(n2324) );
  INV_X4 U450 ( .A(\CARRYB[15][5] ), .ZN(n1454) );
  NAND2_X4 U451 ( .A1(n25), .A2(\ab[22][1] ), .ZN(net82543) );
  INV_X8 U452 ( .A(net77976), .ZN(n175) );
  INV_X4 U453 ( .A(\CARRYB[13][10] ), .ZN(net88408) );
  NAND2_X4 U454 ( .A1(n1533), .A2(n1534), .ZN(n1536) );
  CLKBUF_X3 U456 ( .A(\CARRYB[4][10] ), .Z(n228) );
  NAND2_X4 U457 ( .A1(net123428), .A2(net123429), .ZN(n895) );
  NAND2_X2 U458 ( .A1(\SUMB[2][23] ), .A2(\CARRYB[2][22] ), .ZN(n1070) );
  INV_X8 U459 ( .A(\CARRYB[28][1] ), .ZN(net85094) );
  NOR2_X4 U460 ( .A1(n955), .A2(net70491), .ZN(\ab[2][21] ) );
  NAND2_X2 U461 ( .A1(\CARRYB[2][10] ), .A2(\ab[3][10] ), .ZN(n186) );
  NAND2_X4 U462 ( .A1(\SUMB[5][11] ), .A2(\CARRYB[5][10] ), .ZN(n1748) );
  INV_X8 U463 ( .A(\CARRYB[9][8] ), .ZN(n1289) );
  CLKBUF_X3 U464 ( .A(\SUMB[2][11] ), .Z(n128) );
  NAND2_X2 U466 ( .A1(n129), .A2(n130), .ZN(n132) );
  INV_X1 U468 ( .A(\ab[25][2] ), .ZN(n130) );
  NOR2_X4 U469 ( .A1(net77878), .A2(net70445), .ZN(\ab[25][2] ) );
  INV_X8 U470 ( .A(\CARRYB[5][11] ), .ZN(n146) );
  CLKBUF_X3 U471 ( .A(\CARRYB[9][11] ), .Z(net82678) );
  XNOR2_X2 U472 ( .A(n2031), .B(n151), .ZN(n367) );
  NAND2_X4 U473 ( .A1(\ab[26][0] ), .A2(n152), .ZN(n2027) );
  INV_X2 U474 ( .A(n170), .ZN(net84978) );
  NAND2_X2 U475 ( .A1(\CARRYB[16][11] ), .A2(\SUMB[16][12] ), .ZN(net87011) );
  INV_X2 U476 ( .A(\SUMB[1][16] ), .ZN(n1352) );
  NAND2_X1 U477 ( .A1(n133), .A2(net83535), .ZN(n136) );
  NAND2_X2 U478 ( .A1(n135), .A2(n136), .ZN(n816) );
  INV_X1 U479 ( .A(net83535), .ZN(n134) );
  NAND2_X4 U480 ( .A1(n72), .A2(net87950), .ZN(net149530) );
  NAND2_X4 U481 ( .A1(net80264), .A2(n684), .ZN(n685) );
  INV_X4 U482 ( .A(\SUMB[4][16] ), .ZN(net86162) );
  INV_X8 U483 ( .A(n1937), .ZN(n1506) );
  INV_X8 U484 ( .A(\CARRYB[2][17] ), .ZN(n799) );
  INV_X8 U486 ( .A(net83866), .ZN(net85455) );
  NAND2_X1 U487 ( .A1(\CARRYB[7][5] ), .A2(n2375), .ZN(n138) );
  NAND2_X1 U488 ( .A1(\ab[8][5] ), .A2(n2375), .ZN(n139) );
  NAND2_X1 U489 ( .A1(\ab[8][5] ), .A2(\CARRYB[7][5] ), .ZN(n140) );
  NAND3_X2 U490 ( .A1(n138), .A2(n139), .A3(n140), .ZN(n312) );
  NOR2_X1 U491 ( .A1(net77898), .A2(net77924), .ZN(\ab[8][5] ) );
  BUF_X4 U492 ( .A(n312), .Z(n1206) );
  NAND2_X2 U493 ( .A1(n141), .A2(n142), .ZN(n144) );
  NAND2_X2 U494 ( .A1(n143), .A2(n144), .ZN(n1122) );
  INV_X2 U495 ( .A(\ab[5][7] ), .ZN(n141) );
  INV_X4 U496 ( .A(\CARRYB[4][7] ), .ZN(n142) );
  NOR2_X4 U497 ( .A1(net77912), .A2(net77946), .ZN(\ab[5][7] ) );
  NAND2_X4 U498 ( .A1(\SUMB[25][1] ), .A2(\CARRYB[25][0] ), .ZN(net81535) );
  NAND2_X2 U499 ( .A1(n1855), .A2(n1854), .ZN(n145) );
  NAND2_X1 U500 ( .A1(\CARRYB[5][11] ), .A2(\ab[6][11] ), .ZN(n148) );
  NAND2_X4 U501 ( .A1(n146), .A2(n147), .ZN(n149) );
  INV_X1 U502 ( .A(\ab[6][11] ), .ZN(n147) );
  NAND2_X2 U503 ( .A1(\CARRYB[7][12] ), .A2(\ab[8][12] ), .ZN(net87310) );
  NAND2_X4 U504 ( .A1(net87457), .A2(net87456), .ZN(net87459) );
  INV_X8 U506 ( .A(\CARRYB[4][14] ), .ZN(net84945) );
  NOR2_X2 U507 ( .A1(net77988), .A2(net70466), .ZN(net81416) );
  INV_X4 U508 ( .A(\SUMB[6][16] ), .ZN(n1375) );
  NAND2_X4 U509 ( .A1(n1387), .A2(n1388), .ZN(n151) );
  NAND2_X2 U510 ( .A1(n1387), .A2(n1388), .ZN(\SUMB[8][16] ) );
  INV_X8 U511 ( .A(\CARRYB[22][3] ), .ZN(n404) );
  INV_X8 U512 ( .A(net77904), .ZN(net77898) );
  NAND3_X4 U513 ( .A1(n1564), .A2(n1565), .A3(n1566), .ZN(\CARRYB[6][3] ) );
  NAND3_X2 U514 ( .A1(n2025), .A2(net81530), .A3(net81531), .ZN(n152) );
  XOR2_X2 U515 ( .A(\CARRYB[7][4] ), .B(\ab[8][4] ), .Z(n153) );
  XOR2_X2 U516 ( .A(\SUMB[7][5] ), .B(n153), .Z(\SUMB[8][4] ) );
  NAND2_X2 U517 ( .A1(\CARRYB[7][4] ), .A2(\SUMB[7][5] ), .ZN(n154) );
  NAND2_X2 U518 ( .A1(\ab[8][4] ), .A2(\SUMB[7][5] ), .ZN(n155) );
  NAND2_X2 U519 ( .A1(\ab[8][4] ), .A2(\CARRYB[7][4] ), .ZN(n156) );
  NAND3_X4 U520 ( .A1(n154), .A2(n155), .A3(n156), .ZN(\CARRYB[8][4] ) );
  NAND2_X2 U521 ( .A1(n1552), .A2(\SUMB[5][7] ), .ZN(n159) );
  NAND2_X4 U522 ( .A1(n157), .A2(n158), .ZN(n160) );
  NAND2_X4 U523 ( .A1(n159), .A2(n160), .ZN(\SUMB[6][6] ) );
  INV_X4 U524 ( .A(n1552), .ZN(n157) );
  INV_X1 U525 ( .A(\SUMB[5][7] ), .ZN(n158) );
  NOR2_X1 U526 ( .A1(net77892), .A2(net77924), .ZN(\ab[8][4] ) );
  NAND2_X2 U527 ( .A1(\ab[9][4] ), .A2(\CARRYB[8][4] ), .ZN(net82099) );
  NAND2_X2 U528 ( .A1(\SUMB[6][6] ), .A2(\ab[7][5] ), .ZN(n1521) );
  NAND2_X4 U529 ( .A1(n243), .A2(n244), .ZN(n246) );
  INV_X8 U530 ( .A(net119955), .ZN(net148836) );
  INV_X4 U531 ( .A(n549), .ZN(n307) );
  NAND2_X4 U532 ( .A1(\ab[2][10] ), .A2(\SUMB[1][11] ), .ZN(n1653) );
  NAND2_X4 U533 ( .A1(n256), .A2(n257), .ZN(n259) );
  NAND2_X1 U534 ( .A1(n2377), .A2(\ab[6][8] ), .ZN(n163) );
  NAND2_X4 U535 ( .A1(n161), .A2(n162), .ZN(n164) );
  NAND2_X4 U536 ( .A1(n163), .A2(n164), .ZN(n1994) );
  INV_X2 U537 ( .A(\CARRYB[5][8] ), .ZN(n161) );
  INV_X4 U538 ( .A(\ab[6][8] ), .ZN(n162) );
  NAND3_X2 U539 ( .A1(n1822), .A2(n1823), .A3(n1824), .ZN(n165) );
  NAND2_X1 U540 ( .A1(n398), .A2(\ab[24][1] ), .ZN(n168) );
  NAND2_X4 U541 ( .A1(n166), .A2(n167), .ZN(n169) );
  NAND2_X4 U542 ( .A1(n168), .A2(n169), .ZN(net88776) );
  INV_X4 U543 ( .A(n398), .ZN(n166) );
  INV_X1 U544 ( .A(\ab[24][1] ), .ZN(n167) );
  NOR2_X4 U545 ( .A1(net77920), .A2(net77938), .ZN(\ab[6][8] ) );
  INV_X8 U546 ( .A(n1994), .ZN(n1001) );
  NOR2_X2 U547 ( .A1(net77866), .A2(net70447), .ZN(\ab[24][1] ) );
  NAND3_X2 U548 ( .A1(net80925), .A2(net80924), .A3(net80926), .ZN(
        \CARRYB[22][2] ) );
  INV_X4 U549 ( .A(net89109), .ZN(net85287) );
  NAND2_X2 U550 ( .A1(\SUMB[25][5] ), .A2(\ab[26][4] ), .ZN(n1080) );
  NAND3_X4 U551 ( .A1(net84312), .A2(net84313), .A3(n1057), .ZN(
        \CARRYB[4][22] ) );
  NAND2_X2 U552 ( .A1(net121445), .A2(net121446), .ZN(n466) );
  XNOR2_X2 U553 ( .A(n171), .B(n1083), .ZN(n170) );
  XNOR2_X2 U554 ( .A(\SUMB[23][8] ), .B(n1084), .ZN(n171) );
  INV_X4 U555 ( .A(net81158), .ZN(n200) );
  NOR2_X2 U556 ( .A1(net70456), .A2(net77966), .ZN(\ab[3][11] ) );
  NAND2_X4 U557 ( .A1(\CARRYB[14][9] ), .A2(\ab[15][9] ), .ZN(net84817) );
  INV_X2 U558 ( .A(\CARRYB[2][9] ), .ZN(n1245) );
  NAND2_X4 U559 ( .A1(\SUMB[23][2] ), .A2(\ab[24][1] ), .ZN(net80921) );
  INV_X2 U560 ( .A(\SUMB[16][4] ), .ZN(n560) );
  NOR2_X1 U561 ( .A1(net70454), .A2(net77938), .ZN(\ab[6][10] ) );
  BUF_X16 U562 ( .A(net70454), .Z(net91660) );
  NAND3_X2 U563 ( .A1(n651), .A2(n652), .A3(n653), .ZN(\CARRYB[15][1] ) );
  INV_X2 U564 ( .A(\CARRYB[10][7] ), .ZN(n172) );
  INV_X4 U565 ( .A(n172), .ZN(n173) );
  INV_X8 U566 ( .A(net85035), .ZN(net85036) );
  INV_X4 U567 ( .A(net87363), .ZN(net148828) );
  NOR2_X4 U568 ( .A1(net70470), .A2(net86101), .ZN(\ab[1][18] ) );
  INV_X4 U570 ( .A(n91), .ZN(n578) );
  NAND2_X4 U571 ( .A1(n1362), .A2(net86440), .ZN(n1418) );
  XNOR2_X2 U572 ( .A(\CARRYB[3][13] ), .B(\ab[4][13] ), .ZN(n1562) );
  INV_X1 U573 ( .A(n1611), .ZN(n1368) );
  NOR2_X2 U574 ( .A1(net123000), .A2(net82247), .ZN(net88449) );
  NAND2_X4 U575 ( .A1(\ab[9][13] ), .A2(\SUMB[8][14] ), .ZN(net80349) );
  NAND2_X2 U576 ( .A1(\ab[30][0] ), .A2(net87797), .ZN(net80474) );
  NAND2_X4 U577 ( .A1(n198), .A2(n197), .ZN(\SUMB[9][8] ) );
  NAND2_X4 U578 ( .A1(n195), .A2(n196), .ZN(n198) );
  NAND2_X2 U580 ( .A1(n569), .A2(n1189), .ZN(n218) );
  NAND2_X4 U581 ( .A1(\CARRYB[7][6] ), .A2(\SUMB[7][7] ), .ZN(n1827) );
  AND2_X2 U582 ( .A1(B[10]), .A2(A[3]), .ZN(\ab[3][10] ) );
  INV_X2 U583 ( .A(\ab[0][12] ), .ZN(net120501) );
  BUF_X4 U584 ( .A(\CARRYB[27][0] ), .Z(n284) );
  NAND2_X4 U585 ( .A1(net84868), .A2(net84867), .ZN(net84870) );
  INV_X4 U586 ( .A(net93203), .ZN(n174) );
  INV_X4 U587 ( .A(net83919), .ZN(net93203) );
  INV_X8 U588 ( .A(\ab[0][24] ), .ZN(net82044) );
  NAND2_X2 U589 ( .A1(net82124), .A2(net83044), .ZN(net83576) );
  NAND2_X2 U590 ( .A1(\ab[2][23] ), .A2(n2357), .ZN(net83575) );
  NAND2_X2 U591 ( .A1(n319), .A2(n320), .ZN(n322) );
  NOR2_X4 U592 ( .A1(n2355), .A2(n242), .ZN(\ab[1][27] ) );
  NOR2_X4 U593 ( .A1(n392), .A2(n2354), .ZN(\ab[0][28] ) );
  NAND2_X4 U594 ( .A1(\ab[9][9] ), .A2(\CARRYB[8][9] ), .ZN(n1621) );
  XNOR2_X2 U595 ( .A(\CARRYB[13][11] ), .B(\ab[14][11] ), .ZN(net125934) );
  NAND2_X4 U596 ( .A1(net123291), .A2(n775), .ZN(n776) );
  NAND2_X2 U597 ( .A1(\CARRYB[16][9] ), .A2(\ab[17][9] ), .ZN(net120657) );
  NAND2_X2 U598 ( .A1(n1199), .A2(n558), .ZN(n179) );
  NAND2_X4 U599 ( .A1(n177), .A2(n178), .ZN(n180) );
  NAND2_X4 U600 ( .A1(n179), .A2(n180), .ZN(\SUMB[3][11] ) );
  INV_X4 U601 ( .A(n1199), .ZN(n177) );
  INV_X2 U602 ( .A(n558), .ZN(n178) );
  XNOR2_X2 U603 ( .A(net121785), .B(n1311), .ZN(n181) );
  BUF_X8 U604 ( .A(\SUMB[11][7] ), .Z(n371) );
  BUF_X4 U605 ( .A(\SUMB[3][12] ), .Z(net121785) );
  BUF_X8 U606 ( .A(net70470), .Z(n182) );
  INV_X2 U607 ( .A(net121445), .ZN(n183) );
  INV_X8 U608 ( .A(net90735), .ZN(net121445) );
  NAND2_X1 U609 ( .A1(\CARRYB[17][11] ), .A2(net88647), .ZN(net82666) );
  INV_X1 U610 ( .A(\SUMB[3][20] ), .ZN(n1420) );
  NAND2_X4 U611 ( .A1(n1768), .A2(\SUMB[4][19] ), .ZN(n2141) );
  NAND2_X2 U612 ( .A1(n1486), .A2(n1487), .ZN(n1489) );
  NAND2_X4 U613 ( .A1(net85808), .A2(net84208), .ZN(net87945) );
  NAND2_X4 U614 ( .A1(\ab[14][4] ), .A2(\CARRYB[13][4] ), .ZN(n2152) );
  NAND2_X4 U615 ( .A1(net123293), .A2(n776), .ZN(net93683) );
  NAND2_X4 U616 ( .A1(net147939), .A2(net147940), .ZN(\SUMB[24][2] ) );
  NAND2_X2 U618 ( .A1(n184), .A2(n185), .ZN(n187) );
  NAND2_X4 U619 ( .A1(n186), .A2(n187), .ZN(n1399) );
  INV_X4 U620 ( .A(\CARRYB[2][10] ), .ZN(n184) );
  INV_X1 U621 ( .A(\ab[3][10] ), .ZN(n185) );
  NAND2_X4 U622 ( .A1(net90022), .A2(net90818), .ZN(net87950) );
  NAND2_X1 U623 ( .A1(net81992), .A2(\SUMB[15][10] ), .ZN(n190) );
  NAND2_X2 U624 ( .A1(n188), .A2(n189), .ZN(n191) );
  NAND2_X4 U625 ( .A1(n190), .A2(n191), .ZN(\SUMB[16][9] ) );
  INV_X4 U626 ( .A(net81992), .ZN(n188) );
  INV_X2 U627 ( .A(\SUMB[15][10] ), .ZN(n189) );
  INV_X4 U629 ( .A(n290), .ZN(n1134) );
  INV_X2 U630 ( .A(\SUMB[11][11] ), .ZN(net89840) );
  NAND2_X2 U631 ( .A1(\SUMB[9][9] ), .A2(\CARRYB[9][8] ), .ZN(n1776) );
  NAND2_X4 U632 ( .A1(net87938), .A2(net87939), .ZN(net87941) );
  XNOR2_X2 U634 ( .A(n417), .B(net85109), .ZN(n364) );
  XNOR2_X2 U635 ( .A(n192), .B(\SUMB[26][1] ), .ZN(PRODUCT[27]) );
  INV_X4 U636 ( .A(n1429), .ZN(n288) );
  INV_X4 U638 ( .A(n193), .ZN(net121814) );
  INV_X4 U640 ( .A(net121450), .ZN(net121770) );
  XNOR2_X2 U641 ( .A(\SUMB[9][7] ), .B(n996), .ZN(n194) );
  BUF_X8 U642 ( .A(\SUMB[10][8] ), .Z(n1249) );
  XNOR2_X2 U643 ( .A(net88776), .B(net85903), .ZN(\SUMB[24][1] ) );
  NAND2_X4 U644 ( .A1(n594), .A2(n595), .ZN(\SUMB[11][4] ) );
  NAND2_X2 U645 ( .A1(n2015), .A2(n950), .ZN(n197) );
  INV_X4 U646 ( .A(n2015), .ZN(n195) );
  INV_X4 U647 ( .A(n950), .ZN(n196) );
  NAND2_X2 U648 ( .A1(net123142), .A2(n299), .ZN(n301) );
  NAND2_X1 U649 ( .A1(\ab[12][17] ), .A2(\SUMB[11][18] ), .ZN(n1468) );
  NAND3_X4 U650 ( .A1(net81038), .A2(net81037), .A3(net81036), .ZN(
        \CARRYB[21][8] ) );
  NAND2_X2 U651 ( .A1(\CARRYB[20][8] ), .A2(n859), .ZN(net81038) );
  NAND2_X4 U652 ( .A1(n643), .A2(n644), .ZN(net88699) );
  NAND2_X2 U653 ( .A1(n549), .A2(\SUMB[17][8] ), .ZN(n309) );
  NAND2_X4 U654 ( .A1(net121449), .A2(net121450), .ZN(n199) );
  NAND2_X2 U655 ( .A1(net121450), .A2(net121449), .ZN(net121452) );
  INV_X8 U656 ( .A(net82544), .ZN(net121449) );
  NAND2_X4 U657 ( .A1(n532), .A2(net85096), .ZN(net81158) );
  INV_X8 U659 ( .A(\CARRYB[8][8] ), .ZN(n1177) );
  INV_X2 U660 ( .A(\CARRYB[4][11] ), .ZN(net147920) );
  XNOR2_X1 U661 ( .A(\CARRYB[1][13] ), .B(\ab[2][13] ), .ZN(net124618) );
  NAND2_X4 U662 ( .A1(n1193), .A2(\ab[12][6] ), .ZN(n1917) );
  NAND2_X4 U663 ( .A1(n537), .A2(n538), .ZN(n540) );
  INV_X2 U664 ( .A(\SUMB[1][18] ), .ZN(n538) );
  NAND2_X2 U665 ( .A1(\CARRYB[10][10] ), .A2(net87045), .ZN(n203) );
  NAND2_X2 U666 ( .A1(n201), .A2(n202), .ZN(n204) );
  NAND2_X2 U667 ( .A1(n203), .A2(n204), .ZN(net85732) );
  INV_X1 U668 ( .A(net87045), .ZN(n202) );
  NAND2_X2 U669 ( .A1(net81694), .A2(net84270), .ZN(n207) );
  NAND2_X4 U670 ( .A1(n2366), .A2(n206), .ZN(n208) );
  NAND2_X4 U671 ( .A1(n208), .A2(n207), .ZN(\SUMB[3][13] ) );
  INV_X4 U673 ( .A(net84270), .ZN(n206) );
  INV_X8 U674 ( .A(net122062), .ZN(n299) );
  INV_X2 U675 ( .A(\ab[11][10] ), .ZN(net87045) );
  NAND2_X4 U676 ( .A1(\SUMB[3][13] ), .A2(\ab[4][12] ), .ZN(net82759) );
  BUF_X4 U677 ( .A(\SUMB[3][13] ), .Z(net85493) );
  NAND3_X2 U678 ( .A1(n2115), .A2(n2114), .A3(n2113), .ZN(\CARRYB[25][4] ) );
  OR2_X2 U679 ( .A1(n2361), .A2(n2359), .ZN(n209) );
  NAND2_X4 U680 ( .A1(n45), .A2(n316), .ZN(n318) );
  NAND2_X4 U681 ( .A1(n1507), .A2(n1508), .ZN(n210) );
  NAND2_X2 U683 ( .A1(n211), .A2(\ab[4][13] ), .ZN(n214) );
  INV_X2 U685 ( .A(\CARRYB[3][13] ), .ZN(n211) );
  INV_X1 U686 ( .A(\ab[4][13] ), .ZN(n212) );
  NAND2_X2 U687 ( .A1(n1507), .A2(n1508), .ZN(\SUMB[13][10] ) );
  NOR2_X4 U688 ( .A1(net70460), .A2(net119855), .ZN(\ab[4][13] ) );
  NAND2_X2 U689 ( .A1(n857), .A2(n910), .ZN(n912) );
  NAND2_X4 U690 ( .A1(n1604), .A2(n1605), .ZN(n215) );
  NAND2_X2 U691 ( .A1(n1604), .A2(n1605), .ZN(\SUMB[7][17] ) );
  NAND2_X2 U692 ( .A1(net92724), .A2(\*UDW_*112694/net78575 ), .ZN(n1163) );
  NAND2_X4 U694 ( .A1(n218), .A2(n219), .ZN(n1209) );
  INV_X4 U695 ( .A(n569), .ZN(n216) );
  INV_X1 U696 ( .A(n1189), .ZN(n217) );
  NAND2_X4 U697 ( .A1(\SUMB[12][6] ), .A2(\ab[13][5] ), .ZN(n1921) );
  XNOR2_X2 U698 ( .A(n11), .B(n1270), .ZN(n1189) );
  NAND2_X1 U699 ( .A1(n221), .A2(n2001), .ZN(n222) );
  NAND2_X2 U700 ( .A1(n220), .A2(n939), .ZN(n223) );
  NAND2_X2 U701 ( .A1(n222), .A2(n223), .ZN(\SUMB[8][8] ) );
  INV_X1 U702 ( .A(n2001), .ZN(n220) );
  NAND2_X4 U705 ( .A1(n226), .A2(n227), .ZN(n864) );
  INV_X2 U706 ( .A(n1973), .ZN(n224) );
  INV_X1 U707 ( .A(n1308), .ZN(n225) );
  INV_X4 U708 ( .A(\SUMB[13][7] ), .ZN(n1308) );
  NOR2_X2 U709 ( .A1(net70470), .A2(net86101), .ZN(n401) );
  INV_X4 U710 ( .A(n2095), .ZN(n1725) );
  NAND2_X4 U711 ( .A1(net87682), .A2(net87683), .ZN(n1344) );
  NAND2_X4 U712 ( .A1(n1343), .A2(n1344), .ZN(net82024) );
  NOR2_X2 U713 ( .A1(net82239), .A2(n175), .ZN(\ab[2][25] ) );
  NAND2_X4 U714 ( .A1(net83061), .A2(\ab[10][10] ), .ZN(n458) );
  NAND2_X4 U715 ( .A1(n1684), .A2(n1685), .ZN(\SUMB[2][20] ) );
  INV_X8 U717 ( .A(\CARRYB[8][11] ), .ZN(net86893) );
  NAND2_X1 U718 ( .A1(n797), .A2(net93800), .ZN(n231) );
  NAND2_X2 U719 ( .A1(n231), .A2(n232), .ZN(\SUMB[7][14] ) );
  INV_X2 U720 ( .A(net93800), .ZN(n230) );
  NAND2_X2 U721 ( .A1(n941), .A2(n1618), .ZN(n235) );
  NAND2_X4 U722 ( .A1(n233), .A2(n234), .ZN(n236) );
  NAND2_X4 U723 ( .A1(n235), .A2(n236), .ZN(n1230) );
  INV_X4 U724 ( .A(n941), .ZN(n233) );
  INV_X4 U725 ( .A(n1618), .ZN(n234) );
  XNOR2_X1 U726 ( .A(net81581), .B(net120922), .ZN(n941) );
  INV_X8 U727 ( .A(n1230), .ZN(\SUMB[9][9] ) );
  NAND2_X4 U728 ( .A1(net91301), .A2(\ab[13][8] ), .ZN(net80506) );
  NAND2_X4 U729 ( .A1(\SUMB[11][10] ), .A2(\ab[12][9] ), .ZN(net88296) );
  NAND2_X2 U730 ( .A1(n869), .A2(net83134), .ZN(net86704) );
  INV_X2 U731 ( .A(net88123), .ZN(net123429) );
  NAND2_X2 U732 ( .A1(\ab[10][9] ), .A2(\SUMB[9][10] ), .ZN(n471) );
  INV_X2 U733 ( .A(B[16]), .ZN(net89652) );
  NAND2_X4 U734 ( .A1(\ab[22][4] ), .A2(net86464), .ZN(net79992) );
  NAND2_X4 U735 ( .A1(n940), .A2(\ab[26][0] ), .ZN(net81533) );
  NAND2_X4 U736 ( .A1(\CARRYB[23][0] ), .A2(\ab[24][0] ), .ZN(n1569) );
  NAND2_X2 U737 ( .A1(\ab[4][7] ), .A2(\SUMB[3][8] ), .ZN(n1909) );
  NAND2_X4 U738 ( .A1(n1211), .A2(\SUMB[14][5] ), .ZN(n1707) );
  INV_X16 U739 ( .A(net80392), .ZN(net81673) );
  INV_X16 U740 ( .A(B[15]), .ZN(net87396) );
  CLKBUF_X3 U741 ( .A(\SUMB[1][15] ), .Z(net93243) );
  NAND2_X1 U742 ( .A1(\SUMB[5][18] ), .A2(n1490), .ZN(n2245) );
  NAND2_X2 U743 ( .A1(n238), .A2(n239), .ZN(n241) );
  NAND2_X2 U744 ( .A1(n240), .A2(n241), .ZN(\SUMB[4][17] ) );
  INV_X1 U745 ( .A(n852), .ZN(n239) );
  INV_X4 U746 ( .A(n341), .ZN(n242) );
  INV_X2 U747 ( .A(net80409), .ZN(n341) );
  NAND2_X4 U748 ( .A1(\SUMB[2][15] ), .A2(n1186), .ZN(n1989) );
  INV_X4 U749 ( .A(net81581), .ZN(net123842) );
  NAND2_X1 U750 ( .A1(net149611), .A2(net121859), .ZN(n245) );
  NAND2_X4 U751 ( .A1(n245), .A2(n246), .ZN(\SUMB[3][15] ) );
  INV_X1 U752 ( .A(net149611), .ZN(n243) );
  INV_X2 U753 ( .A(net121859), .ZN(n244) );
  NAND2_X4 U754 ( .A1(net124367), .A2(net123303), .ZN(n2158) );
  NAND2_X4 U755 ( .A1(\CARRYB[11][7] ), .A2(\ab[12][7] ), .ZN(n2019) );
  XNOR2_X2 U756 ( .A(\CARRYB[19][8] ), .B(\ab[20][8] ), .ZN(n368) );
  NAND3_X2 U757 ( .A1(n503), .A2(n501), .A3(n502), .ZN(n247) );
  NAND2_X4 U758 ( .A1(n250), .A2(n251), .ZN(net81431) );
  INV_X2 U759 ( .A(\CARRYB[28][0] ), .ZN(n248) );
  INV_X4 U760 ( .A(n344), .ZN(n249) );
  NAND2_X4 U761 ( .A1(n252), .A2(n253), .ZN(n255) );
  NAND2_X4 U762 ( .A1(n255), .A2(n254), .ZN(\SUMB[12][6] ) );
  INV_X4 U763 ( .A(n1764), .ZN(n252) );
  INV_X4 U764 ( .A(n371), .ZN(n253) );
  BUF_X4 U765 ( .A(\SUMB[12][6] ), .Z(n1260) );
  NAND2_X2 U766 ( .A1(\SUMB[12][7] ), .A2(\ab[13][6] ), .ZN(n258) );
  NAND2_X2 U767 ( .A1(n258), .A2(n259), .ZN(n1899) );
  INV_X4 U768 ( .A(\SUMB[12][7] ), .ZN(n256) );
  INV_X1 U769 ( .A(\ab[13][6] ), .ZN(n257) );
  NOR2_X2 U770 ( .A1(net77908), .A2(net70469), .ZN(\ab[13][6] ) );
  NOR2_X1 U771 ( .A1(net77878), .A2(net86101), .ZN(\ab[1][2] ) );
  NAND2_X4 U772 ( .A1(net88692), .A2(net121150), .ZN(n1390) );
  NOR2_X4 U773 ( .A1(\ab[28][2] ), .A2(n260), .ZN(n261) );
  NOR2_X2 U774 ( .A1(n530), .A2(n261), .ZN(net92314) );
  INV_X4 U775 ( .A(n348), .ZN(n260) );
  INV_X1 U776 ( .A(net83116), .ZN(n262) );
  NAND2_X2 U777 ( .A1(n1609), .A2(n866), .ZN(n265) );
  NAND2_X4 U778 ( .A1(n263), .A2(n264), .ZN(n266) );
  NAND2_X4 U779 ( .A1(n265), .A2(n266), .ZN(n1233) );
  INV_X4 U780 ( .A(n1609), .ZN(n263) );
  INV_X2 U781 ( .A(n866), .ZN(n264) );
  NAND2_X2 U782 ( .A1(n859), .A2(net90801), .ZN(n269) );
  NAND2_X4 U783 ( .A1(n267), .A2(n268), .ZN(n270) );
  NAND2_X4 U784 ( .A1(n269), .A2(n270), .ZN(net89461) );
  INV_X4 U785 ( .A(n859), .ZN(n267) );
  INV_X4 U786 ( .A(net90801), .ZN(n268) );
  NAND2_X2 U787 ( .A1(net85119), .A2(\SUMB[13][15] ), .ZN(n273) );
  NAND2_X4 U788 ( .A1(n271), .A2(n272), .ZN(n274) );
  NAND2_X4 U789 ( .A1(n273), .A2(n274), .ZN(\SUMB[14][14] ) );
  INV_X4 U790 ( .A(net85119), .ZN(n271) );
  INV_X2 U791 ( .A(\SUMB[13][15] ), .ZN(n272) );
  NAND2_X2 U792 ( .A1(\SUMB[14][14] ), .A2(net93107), .ZN(n277) );
  NAND2_X4 U793 ( .A1(n275), .A2(n276), .ZN(n278) );
  NAND2_X4 U794 ( .A1(n277), .A2(n278), .ZN(\SUMB[15][13] ) );
  INV_X2 U795 ( .A(\SUMB[14][14] ), .ZN(n275) );
  INV_X4 U796 ( .A(net93107), .ZN(n276) );
  NAND2_X1 U797 ( .A1(B[2]), .A2(A[28]), .ZN(net92311) );
  NAND2_X2 U798 ( .A1(n56), .A2(\SUMB[5][20] ), .ZN(n2281) );
  NAND2_X2 U799 ( .A1(\ab[6][19] ), .A2(\SUMB[5][20] ), .ZN(n2280) );
  NAND2_X2 U800 ( .A1(n1233), .A2(\ab[4][20] ), .ZN(n2238) );
  NAND2_X2 U801 ( .A1(net120625), .A2(net120626), .ZN(net120628) );
  NAND2_X4 U802 ( .A1(\ab[10][8] ), .A2(\SUMB[9][9] ), .ZN(n1775) );
  INV_X4 U803 ( .A(n38), .ZN(n1628) );
  OAI21_X4 U805 ( .B1(net119909), .B2(net119910), .A(n477), .ZN(n279) );
  NAND2_X2 U806 ( .A1(\ab[2][16] ), .A2(\CARRYB[1][16] ), .ZN(n282) );
  NAND2_X4 U807 ( .A1(n283), .A2(n282), .ZN(net119952) );
  INV_X4 U809 ( .A(\CARRYB[1][16] ), .ZN(n281) );
  XNOR2_X2 U810 ( .A(net119952), .B(\*UDW_*112684/net78549 ), .ZN(net149611)
         );
  NAND2_X2 U811 ( .A1(n728), .A2(\SUMB[8][4] ), .ZN(net82850) );
  NAND2_X4 U812 ( .A1(\CARRYB[28][0] ), .A2(n344), .ZN(net79883) );
  NAND2_X4 U813 ( .A1(\SUMB[25][2] ), .A2(\ab[26][1] ), .ZN(net83977) );
  NAND2_X2 U814 ( .A1(n944), .A2(net87874), .ZN(n1337) );
  XNOR2_X2 U815 ( .A(n417), .B(n286), .ZN(n285) );
  INV_X32 U816 ( .A(net85109), .ZN(n286) );
  INV_X4 U817 ( .A(\SUMB[24][4] ), .ZN(net87938) );
  NAND2_X2 U818 ( .A1(n300), .A2(n301), .ZN(\SUMB[12][9] ) );
  BUF_X4 U819 ( .A(\SUMB[8][11] ), .Z(net125375) );
  NAND2_X1 U820 ( .A1(\ab[3][12] ), .A2(n1207), .ZN(n2009) );
  NAND2_X1 U821 ( .A1(\ab[15][12] ), .A2(\SUMB[14][13] ), .ZN(n2199) );
  CLKBUF_X3 U822 ( .A(\CARRYB[13][13] ), .Z(n695) );
  INV_X8 U823 ( .A(n933), .ZN(n936) );
  NAND2_X4 U824 ( .A1(\SUMB[10][15] ), .A2(\CARRYB[10][14] ), .ZN(n1844) );
  NAND3_X4 U825 ( .A1(n1106), .A2(n1105), .A3(n1107), .ZN(\CARRYB[8][18] ) );
  INV_X2 U826 ( .A(n1118), .ZN(net80643) );
  INV_X8 U827 ( .A(\CARRYB[18][7] ), .ZN(n1615) );
  NAND2_X2 U829 ( .A1(\CARRYB[1][15] ), .A2(\SUMB[1][16] ), .ZN(n1986) );
  NAND2_X2 U830 ( .A1(\SUMB[9][10] ), .A2(\CARRYB[9][9] ), .ZN(n472) );
  INV_X2 U831 ( .A(net83755), .ZN(net120518) );
  NAND2_X2 U833 ( .A1(\SUMB[7][11] ), .A2(\CARRYB[7][10] ), .ZN(net81216) );
  INV_X2 U834 ( .A(\SUMB[1][13] ), .ZN(net123509) );
  XNOR2_X2 U835 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .ZN(n849) );
  XNOR2_X2 U836 ( .A(n1216), .B(n1220), .ZN(n556) );
  INV_X4 U838 ( .A(\SUMB[6][9] ), .ZN(n1429) );
  INV_X8 U839 ( .A(\ab[2][11] ), .ZN(n585) );
  NOR2_X4 U840 ( .A1(n405), .A2(n421), .ZN(n410) );
  XOR2_X2 U841 ( .A(\ab[13][0] ), .B(\SUMB[12][1] ), .Z(n291) );
  XOR2_X2 U842 ( .A(n291), .B(\CARRYB[12][0] ), .Z(PRODUCT[13]) );
  NAND2_X2 U843 ( .A1(\ab[13][0] ), .A2(\SUMB[12][1] ), .ZN(n292) );
  NAND2_X2 U844 ( .A1(\ab[13][0] ), .A2(\CARRYB[12][0] ), .ZN(n293) );
  NAND2_X2 U845 ( .A1(\SUMB[12][1] ), .A2(\CARRYB[12][0] ), .ZN(n294) );
  NAND3_X4 U846 ( .A1(n292), .A2(n293), .A3(n294), .ZN(\CARRYB[13][0] ) );
  XOR2_X1 U847 ( .A(\ab[14][0] ), .B(\SUMB[13][1] ), .Z(n295) );
  XOR2_X1 U848 ( .A(n295), .B(\CARRYB[13][0] ), .Z(PRODUCT[14]) );
  NAND2_X2 U849 ( .A1(\ab[14][0] ), .A2(\SUMB[13][1] ), .ZN(n296) );
  NAND2_X1 U850 ( .A1(\ab[14][0] ), .A2(\CARRYB[13][0] ), .ZN(n297) );
  NAND2_X2 U851 ( .A1(\SUMB[13][1] ), .A2(\CARRYB[13][0] ), .ZN(n298) );
  NAND3_X4 U852 ( .A1(n296), .A2(n297), .A3(n298), .ZN(\CARRYB[14][0] ) );
  NAND2_X1 U853 ( .A1(net89168), .A2(net122062), .ZN(n300) );
  INV_X8 U854 ( .A(net84327), .ZN(net119921) );
  NAND2_X4 U855 ( .A1(net84672), .A2(net84671), .ZN(\SUMB[9][12] ) );
  NAND2_X4 U856 ( .A1(net82759), .A2(n1829), .ZN(n1734) );
  INV_X1 U857 ( .A(n393), .ZN(net84979) );
  NAND2_X2 U858 ( .A1(\SUMB[10][16] ), .A2(\CARRYB[10][15] ), .ZN(n1091) );
  NAND2_X2 U859 ( .A1(n112), .A2(\ab[0][16] ), .ZN(n304) );
  NAND2_X4 U860 ( .A1(n302), .A2(n303), .ZN(n305) );
  NAND2_X4 U861 ( .A1(n304), .A2(n305), .ZN(n437) );
  INV_X4 U862 ( .A(\ab[1][15] ), .ZN(n302) );
  INV_X8 U863 ( .A(\ab[0][16] ), .ZN(n303) );
  XNOR2_X2 U864 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .ZN(n774) );
  NOR2_X4 U865 ( .A1(net82043), .A2(net82044), .ZN(net82124) );
  XNOR2_X2 U866 ( .A(\SUMB[14][15] ), .B(net86054), .ZN(net90525) );
  NAND2_X4 U867 ( .A1(net123269), .A2(net123268), .ZN(net119955) );
  NAND3_X4 U868 ( .A1(n1954), .A2(n1953), .A3(n1952), .ZN(\CARRYB[16][14] ) );
  NAND2_X2 U869 ( .A1(\SUMB[22][2] ), .A2(\ab[23][1] ), .ZN(n751) );
  NAND2_X2 U870 ( .A1(\SUMB[6][6] ), .A2(\CARRYB[6][5] ), .ZN(n1519) );
  NAND2_X4 U871 ( .A1(n1615), .A2(n1614), .ZN(n1616) );
  NAND2_X2 U872 ( .A1(\ab[4][12] ), .A2(n89), .ZN(n1829) );
  NAND2_X1 U873 ( .A1(net88916), .A2(net86696), .ZN(net79868) );
  NAND2_X4 U874 ( .A1(n819), .A2(n820), .ZN(n822) );
  NAND2_X2 U875 ( .A1(\SUMB[18][9] ), .A2(net93683), .ZN(n643) );
  NAND2_X4 U876 ( .A1(n575), .A2(n679), .ZN(n681) );
  NAND2_X4 U877 ( .A1(net85808), .A2(\ab[17][9] ), .ZN(net80813) );
  INV_X4 U878 ( .A(net86374), .ZN(n306) );
  INV_X4 U879 ( .A(net86374), .ZN(net86375) );
  NAND2_X2 U880 ( .A1(\ab[8][10] ), .A2(\CARRYB[7][10] ), .ZN(n461) );
  NAND2_X4 U881 ( .A1(n307), .A2(n308), .ZN(n310) );
  NAND2_X4 U882 ( .A1(n309), .A2(n310), .ZN(\SUMB[18][7] ) );
  INV_X2 U883 ( .A(\SUMB[17][8] ), .ZN(n308) );
  NAND2_X2 U885 ( .A1(\ab[22][0] ), .A2(\SUMB[21][1] ), .ZN(n1797) );
  NOR2_X1 U887 ( .A1(n2354), .A2(n175), .ZN(\ab[2][28] ) );
  NOR2_X1 U888 ( .A1(n2355), .A2(n175), .ZN(\ab[2][27] ) );
  NAND2_X2 U889 ( .A1(net81416), .A2(n112), .ZN(\*UDW_*112694/net78575 ) );
  NOR2_X2 U890 ( .A1(net88344), .A2(net77948), .ZN(\ab[5][16] ) );
  BUF_X8 U891 ( .A(net88344), .Z(net124723) );
  INV_X8 U892 ( .A(net93914), .ZN(net82009) );
  INV_X16 U893 ( .A(B[18]), .ZN(net70470) );
  NAND2_X2 U894 ( .A1(B[18]), .A2(net81630), .ZN(net86959) );
  NAND2_X4 U895 ( .A1(\SUMB[1][13] ), .A2(\ab[2][12] ), .ZN(n2080) );
  NOR2_X1 U896 ( .A1(net70486), .A2(net77966), .ZN(\ab[3][26] ) );
  NAND2_X4 U897 ( .A1(n313), .A2(n314), .ZN(n315) );
  NAND2_X4 U898 ( .A1(n2022), .A2(n315), .ZN(n1732) );
  INV_X1 U900 ( .A(\ab[13][7] ), .ZN(n314) );
  NAND2_X1 U901 ( .A1(n89), .A2(\ab[4][12] ), .ZN(n317) );
  NAND2_X4 U902 ( .A1(n317), .A2(n318), .ZN(net89227) );
  NAND2_X1 U903 ( .A1(\CARRYB[7][10] ), .A2(\ab[8][10] ), .ZN(n321) );
  NAND2_X4 U904 ( .A1(n321), .A2(n322), .ZN(net81581) );
  INV_X2 U905 ( .A(\CARRYB[7][10] ), .ZN(n319) );
  INV_X1 U906 ( .A(\ab[8][10] ), .ZN(n320) );
  NAND2_X4 U907 ( .A1(n325), .A2(n326), .ZN(net82723) );
  INV_X1 U908 ( .A(\ab[10][9] ), .ZN(n324) );
  NOR2_X1 U909 ( .A1(net77914), .A2(net70469), .ZN(\ab[13][7] ) );
  NAND2_X2 U910 ( .A1(net81581), .A2(net120922), .ZN(n873) );
  NOR2_X2 U911 ( .A1(net70452), .A2(net70475), .ZN(\ab[10][9] ) );
  INV_X4 U912 ( .A(net82723), .ZN(net120513) );
  CLKBUF_X3 U913 ( .A(\SUMB[4][13] ), .Z(n448) );
  NOR2_X4 U914 ( .A1(net70476), .A2(net86101), .ZN(\ab[1][21] ) );
  NAND2_X4 U915 ( .A1(net80302), .A2(net80660), .ZN(net80366) );
  NAND2_X2 U916 ( .A1(n351), .A2(net89402), .ZN(n2285) );
  NAND2_X2 U917 ( .A1(\ab[23][6] ), .A2(net89402), .ZN(n2284) );
  NOR2_X4 U918 ( .A1(net70474), .A2(net82149), .ZN(\ab[0][20] ) );
  NAND2_X4 U919 ( .A1(net93840), .A2(\ab[25][2] ), .ZN(net80263) );
  INV_X8 U920 ( .A(n2329), .ZN(\CARRYB[1][5] ) );
  NAND2_X4 U921 ( .A1(\SUMB[16][8] ), .A2(\ab[17][7] ), .ZN(net81266) );
  NAND2_X2 U922 ( .A1(n1376), .A2(\SUMB[6][16] ), .ZN(n1377) );
  NOR2_X4 U923 ( .A1(net70454), .A2(net86101), .ZN(\ab[1][10] ) );
  NAND2_X2 U924 ( .A1(\CARRYB[3][7] ), .A2(\SUMB[3][8] ), .ZN(n1910) );
  NAND2_X4 U925 ( .A1(n639), .A2(n640), .ZN(n1741) );
  NAND2_X1 U926 ( .A1(\CARRYB[7][15] ), .A2(\ab[8][15] ), .ZN(n329) );
  NAND2_X2 U927 ( .A1(n327), .A2(n328), .ZN(n330) );
  NAND2_X2 U928 ( .A1(n329), .A2(n330), .ZN(n1736) );
  INV_X4 U929 ( .A(\CARRYB[7][15] ), .ZN(n327) );
  INV_X1 U930 ( .A(\ab[8][15] ), .ZN(n328) );
  NOR2_X2 U931 ( .A1(net81424), .A2(net77926), .ZN(\ab[8][15] ) );
  NAND2_X4 U932 ( .A1(net83175), .A2(net83174), .ZN(n2244) );
  NAND2_X4 U933 ( .A1(n542), .A2(net82834), .ZN(net83174) );
  INV_X1 U934 ( .A(n375), .ZN(n332) );
  INV_X4 U935 ( .A(n332), .ZN(n333) );
  INV_X2 U936 ( .A(net147938), .ZN(n334) );
  NAND2_X4 U937 ( .A1(n404), .A2(n406), .ZN(n421) );
  NAND2_X4 U939 ( .A1(n915), .A2(n916), .ZN(n1199) );
  NAND2_X4 U940 ( .A1(\CARRYB[17][4] ), .A2(\ab[18][4] ), .ZN(n2040) );
  NAND2_X2 U941 ( .A1(net81087), .A2(net90262), .ZN(n337) );
  NAND2_X4 U942 ( .A1(n335), .A2(n336), .ZN(n338) );
  NAND2_X4 U943 ( .A1(n337), .A2(n338), .ZN(net89670) );
  INV_X2 U944 ( .A(net81087), .ZN(n335) );
  INV_X2 U945 ( .A(net90262), .ZN(n336) );
  BUF_X4 U946 ( .A(\SUMB[10][13] ), .Z(net90262) );
  OR2_X2 U947 ( .A1(\SUMB[15][11] ), .A2(\CARRYB[15][10] ), .ZN(n339) );
  INV_X8 U948 ( .A(n2248), .ZN(n1592) );
  NAND2_X2 U949 ( .A1(\ab[8][14] ), .A2(\SUMB[7][15] ), .ZN(n2272) );
  INV_X2 U950 ( .A(n929), .ZN(n918) );
  INV_X4 U951 ( .A(n675), .ZN(n340) );
  NAND2_X4 U952 ( .A1(n1855), .A2(n1854), .ZN(n675) );
  NAND2_X4 U953 ( .A1(net84945), .A2(\ab[5][14] ), .ZN(net84948) );
  INV_X2 U954 ( .A(\SUMB[6][12] ), .ZN(net88106) );
  NOR2_X4 U955 ( .A1(net124610), .A2(net77912), .ZN(\ab[0][7] ) );
  XNOR2_X2 U956 ( .A(n343), .B(\ab[6][4] ), .ZN(net92884) );
  NAND2_X4 U957 ( .A1(\SUMB[20][6] ), .A2(\ab[21][5] ), .ZN(net79990) );
  NAND2_X4 U958 ( .A1(\SUMB[4][14] ), .A2(\ab[5][13] ), .ZN(n1981) );
  BUF_X4 U959 ( .A(net80564), .Z(net83296) );
  INV_X8 U960 ( .A(\*UDW_*112644/net78437 ), .ZN(\SUMB[1][25] ) );
  NOR2_X4 U962 ( .A1(n392), .A2(net70456), .ZN(\ab[0][11] ) );
  NAND2_X4 U963 ( .A1(\ab[3][14] ), .A2(\SUMB[2][15] ), .ZN(n1988) );
  NAND2_X1 U964 ( .A1(\SUMB[16][13] ), .A2(\ab[17][12] ), .ZN(n893) );
  NAND2_X4 U965 ( .A1(net92790), .A2(\ab[25][2] ), .ZN(net80262) );
  INV_X2 U966 ( .A(net81663), .ZN(n577) );
  BUF_X4 U967 ( .A(\CARRYB[19][8] ), .Z(net89467) );
  INV_X4 U968 ( .A(n825), .ZN(n826) );
  NOR2_X4 U969 ( .A1(net70482), .A2(net80409), .ZN(\ab[1][24] ) );
  NAND3_X4 U970 ( .A1(n1579), .A2(n1580), .A3(net84746), .ZN(\CARRYB[17][10] )
         );
  INV_X8 U971 ( .A(\CARRYB[14][9] ), .ZN(n831) );
  NOR2_X4 U972 ( .A1(n392), .A2(net70482), .ZN(\ab[0][24] ) );
  INV_X16 U973 ( .A(net80392), .ZN(n392) );
  NAND3_X4 U974 ( .A1(n1390), .A2(n1391), .A3(n1392), .ZN(\CARRYB[19][8] ) );
  NAND2_X4 U975 ( .A1(net88692), .A2(\ab[19][8] ), .ZN(n1391) );
  NAND2_X2 U976 ( .A1(\CARRYB[5][20] ), .A2(\SUMB[5][21] ), .ZN(net79935) );
  NAND2_X4 U977 ( .A1(\ab[5][8] ), .A2(\CARRYB[4][8] ), .ZN(n1964) );
  NAND2_X4 U978 ( .A1(n542), .A2(\ab[21][3] ), .ZN(net80509) );
  INV_X2 U979 ( .A(\CARRYB[5][4] ), .ZN(n342) );
  INV_X4 U980 ( .A(n342), .ZN(n343) );
  NAND3_X4 U981 ( .A1(n1295), .A2(n1296), .A3(n667), .ZN(\CARRYB[12][4] ) );
  NAND2_X2 U982 ( .A1(\CARRYB[11][4] ), .A2(\SUMB[11][5] ), .ZN(n1295) );
  INV_X2 U983 ( .A(net123365), .ZN(net83623) );
  BUF_X16 U984 ( .A(\SUMB[10][2] ), .Z(n730) );
  NAND2_X2 U985 ( .A1(\CARRYB[5][3] ), .A2(\SUMB[5][4] ), .ZN(n1564) );
  NAND2_X4 U986 ( .A1(n1155), .A2(n1156), .ZN(n1651) );
  NAND2_X4 U987 ( .A1(net82544), .A2(net121770), .ZN(net121451) );
  NOR2_X4 U988 ( .A1(net70474), .A2(net80409), .ZN(\ab[1][20] ) );
  NOR2_X4 U989 ( .A1(net70462), .A2(net82149), .ZN(\ab[0][14] ) );
  NOR2_X2 U990 ( .A1(n404), .A2(n419), .ZN(n412) );
  INV_X1 U991 ( .A(\SUMB[18][5] ), .ZN(n1347) );
  NOR2_X4 U992 ( .A1(n407), .A2(n408), .ZN(n413) );
  NOR2_X4 U993 ( .A1(net89652), .A2(net70491), .ZN(\ab[2][16] ) );
  INV_X1 U994 ( .A(\SUMB[28][2] ), .ZN(n531) );
  NAND2_X1 U996 ( .A1(\SUMB[4][22] ), .A2(\ab[5][21] ), .ZN(n1116) );
  NOR2_X4 U998 ( .A1(net123000), .A2(net82247), .ZN(\ab[0][17] ) );
  NOR2_X4 U999 ( .A1(net82247), .A2(net70480), .ZN(\ab[0][23] ) );
  INV_X16 U1000 ( .A(net81630), .ZN(net82247) );
  NOR2_X2 U1001 ( .A1(net77866), .A2(net77970), .ZN(\ab[2][1] ) );
  NOR2_X2 U1002 ( .A1(net77878), .A2(net77930), .ZN(\ab[7][2] ) );
  NOR2_X1 U1003 ( .A1(net77860), .A2(net77970), .ZN(\ab[2][0] ) );
  NOR2_X2 U1004 ( .A1(net77860), .A2(net77930), .ZN(\ab[7][0] ) );
  NAND2_X2 U1005 ( .A1(\ab[12][4] ), .A2(\SUMB[11][5] ), .ZN(n1296) );
  NOR2_X2 U1006 ( .A1(net77892), .A2(net77930), .ZN(\ab[7][4] ) );
  NOR2_X1 U1007 ( .A1(net77882), .A2(net77966), .ZN(\ab[3][3] ) );
  NOR2_X2 U1008 ( .A1(net77878), .A2(net77924), .ZN(\ab[8][2] ) );
  INV_X8 U1009 ( .A(A[11]), .ZN(net70473) );
  NOR2_X1 U1010 ( .A1(net77878), .A2(net77966), .ZN(\ab[3][2] ) );
  NOR2_X1 U1011 ( .A1(net77860), .A2(net70467), .ZN(\ab[14][0] ) );
  NOR2_X1 U1012 ( .A1(net77858), .A2(net119855), .ZN(\ab[4][0] ) );
  NOR2_X1 U1013 ( .A1(net77860), .A2(net70477), .ZN(\ab[9][0] ) );
  NOR2_X2 U1014 ( .A1(net81424), .A2(net70477), .ZN(\ab[9][15] ) );
  INV_X4 U1015 ( .A(B[30]), .ZN(n2353) );
  NOR2_X2 U1016 ( .A1(net81673), .A2(n2353), .ZN(\ab[0][30] ) );
  NOR2_X2 U1017 ( .A1(net77920), .A2(net70467), .ZN(\ab[14][8] ) );
  NOR2_X1 U1018 ( .A1(net77908), .A2(net70461), .ZN(\ab[17][6] ) );
  NAND2_X2 U1019 ( .A1(n673), .A2(n674), .ZN(n1198) );
  NAND2_X2 U1020 ( .A1(n671), .A2(n672), .ZN(n674) );
  NOR2_X1 U1021 ( .A1(net77906), .A2(net77946), .ZN(\ab[5][6] ) );
  NOR2_X1 U1022 ( .A1(net77892), .A2(net77956), .ZN(\ab[4][4] ) );
  INV_X4 U1023 ( .A(\ab[11][2] ), .ZN(net85032) );
  NOR2_X1 U1024 ( .A1(net77878), .A2(net77946), .ZN(\ab[5][2] ) );
  INV_X4 U1025 ( .A(A[8]), .ZN(net77924) );
  NOR2_X1 U1026 ( .A1(net81673), .A2(net77866), .ZN(\ab[0][1] ) );
  NOR2_X1 U1027 ( .A1(net77858), .A2(net77946), .ZN(\ab[5][0] ) );
  NOR2_X1 U1028 ( .A1(net77860), .A2(net70475), .ZN(\ab[10][0] ) );
  INV_X4 U1029 ( .A(n2344), .ZN(\SUMB[1][21] ) );
  INV_X4 U1030 ( .A(\*UDW_*112694/net78575 ), .ZN(\CARRYB[1][15] ) );
  NAND3_X2 U1031 ( .A1(n1931), .A2(n1930), .A3(n1932), .ZN(\CARRYB[2][22] ) );
  NOR2_X2 U1032 ( .A1(net80727), .A2(net77956), .ZN(\ab[4][20] ) );
  NAND3_X2 U1033 ( .A1(n2165), .A2(n2166), .A3(n2167), .ZN(\CARRYB[2][25] ) );
  INV_X4 U1034 ( .A(\ab[10][15] ), .ZN(n1624) );
  NAND3_X2 U1035 ( .A1(n2260), .A2(n2261), .A3(n2262), .ZN(\CARRYB[2][28] ) );
  INV_X4 U1036 ( .A(\ab[9][20] ), .ZN(n1889) );
  NOR2_X2 U1037 ( .A1(net81424), .A2(net70469), .ZN(\ab[13][15] ) );
  INV_X4 U1038 ( .A(n1830), .ZN(n1760) );
  INV_X4 U1039 ( .A(n1553), .ZN(n628) );
  INV_X2 U1040 ( .A(\ab[18][10] ), .ZN(n897) );
  INV_X4 U1041 ( .A(n1588), .ZN(n1445) );
  NOR2_X2 U1042 ( .A1(net77908), .A2(net70459), .ZN(\ab[18][6] ) );
  NAND3_X2 U1043 ( .A1(n1948), .A2(n1947), .A3(n143), .ZN(\CARRYB[5][7] ) );
  NOR2_X2 U1044 ( .A1(net77892), .A2(net70469), .ZN(\ab[13][4] ) );
  NOR2_X1 U1045 ( .A1(net77898), .A2(net70475), .ZN(\ab[10][5] ) );
  INV_X4 U1046 ( .A(n592), .ZN(n563) );
  INV_X4 U1047 ( .A(net87961), .ZN(net87962) );
  NAND2_X2 U1048 ( .A1(\ab[2][6] ), .A2(\SUMB[1][7] ), .ZN(n760) );
  NOR2_X2 U1049 ( .A1(net77886), .A2(net77924), .ZN(\ab[8][3] ) );
  NOR2_X2 U1050 ( .A1(net77898), .A2(net77956), .ZN(\ab[4][5] ) );
  NOR2_X1 U1051 ( .A1(net77858), .A2(net70445), .ZN(\ab[25][0] ) );
  NOR2_X1 U1052 ( .A1(net77866), .A2(net77966), .ZN(\ab[3][1] ) );
  NOR2_X1 U1053 ( .A1(net77866), .A2(net70477), .ZN(\ab[9][1] ) );
  INV_X4 U1054 ( .A(\ab[17][1] ), .ZN(net88712) );
  NOR2_X1 U1055 ( .A1(net77858), .A2(net77966), .ZN(\ab[3][0] ) );
  NOR2_X2 U1056 ( .A1(net77860), .A2(net77924), .ZN(\ab[8][0] ) );
  NOR2_X1 U1057 ( .A1(net77860), .A2(net70469), .ZN(\ab[13][0] ) );
  NAND2_X2 U1058 ( .A1(net82024), .A2(\SUMB[1][18] ), .ZN(n539) );
  NAND2_X2 U1059 ( .A1(n95), .A2(\SUMB[2][18] ), .ZN(n1716) );
  NOR2_X2 U1060 ( .A1(net86565), .A2(net77964), .ZN(\ab[3][19] ) );
  NAND3_X2 U1061 ( .A1(n2146), .A2(n2147), .A3(n1548), .ZN(\CARRYB[3][18] ) );
  NAND2_X2 U1062 ( .A1(\ab[4][13] ), .A2(\CARRYB[3][13] ), .ZN(n2089) );
  NOR2_X2 U1063 ( .A1(net84358), .A2(n331), .ZN(\ab[2][23] ) );
  INV_X4 U1064 ( .A(n2043), .ZN(n1749) );
  NOR2_X2 U1065 ( .A1(net81424), .A2(net77932), .ZN(\ab[7][15] ) );
  NAND2_X2 U1066 ( .A1(n2360), .A2(\ab[9][12] ), .ZN(net81374) );
  CLKBUF_X3 U1067 ( .A(\SUMB[3][24] ), .Z(n1089) );
  NAND2_X2 U1068 ( .A1(n957), .A2(n958), .ZN(n960) );
  INV_X16 U1069 ( .A(n444), .ZN(net77932) );
  INV_X4 U1070 ( .A(\CARRYB[4][12] ), .ZN(net87465) );
  NOR2_X2 U1071 ( .A1(net91660), .A2(net70477), .ZN(\ab[9][10] ) );
  NAND2_X2 U1072 ( .A1(\SUMB[9][14] ), .A2(\CARRYB[9][13] ), .ZN(net80248) );
  NAND2_X2 U1073 ( .A1(n1040), .A2(n1039), .ZN(n1227) );
  NOR2_X2 U1074 ( .A1(net124723), .A2(net70475), .ZN(\ab[10][16] ) );
  NAND3_X2 U1075 ( .A1(n1843), .A2(n1842), .A3(n1844), .ZN(\CARRYB[11][14] )
         );
  NAND2_X2 U1076 ( .A1(net121447), .A2(n466), .ZN(net89537) );
  INV_X4 U1077 ( .A(\ab[10][19] ), .ZN(n1886) );
  NOR2_X2 U1078 ( .A1(net77920), .A2(net70475), .ZN(\ab[10][8] ) );
  INV_X4 U1079 ( .A(net84007), .ZN(net84209) );
  INV_X2 U1080 ( .A(\ab[14][13] ), .ZN(n400) );
  NAND3_X2 U1081 ( .A1(net79891), .A2(net79892), .A3(net79893), .ZN(
        \CARRYB[13][15] ) );
  NAND2_X2 U1082 ( .A1(\ab[14][13] ), .A2(\SUMB[13][14] ), .ZN(n1060) );
  NAND2_X2 U1083 ( .A1(n615), .A2(n616), .ZN(n618) );
  INV_X8 U1084 ( .A(net77988), .ZN(net81630) );
  NOR2_X2 U1085 ( .A1(net77908), .A2(net70453), .ZN(\ab[21][6] ) );
  BUF_X8 U1086 ( .A(net70456), .Z(net85716) );
  INV_X4 U1087 ( .A(n1429), .ZN(n1430) );
  NOR2_X1 U1088 ( .A1(net77906), .A2(net70473), .ZN(\ab[11][6] ) );
  CLKBUF_X3 U1089 ( .A(\SUMB[14][7] ), .Z(n1123) );
  NAND2_X2 U1090 ( .A1(\CARRYB[14][5] ), .A2(\ab[15][5] ), .ZN(n1977) );
  INV_X4 U1091 ( .A(\ab[23][6] ), .ZN(n1234) );
  NAND2_X2 U1092 ( .A1(n683), .A2(\SUMB[21][8] ), .ZN(n686) );
  INV_X4 U1093 ( .A(\ab[18][6] ), .ZN(net82748) );
  NAND2_X2 U1094 ( .A1(\ab[22][2] ), .A2(\SUMB[21][3] ), .ZN(net80925) );
  INV_X4 U1095 ( .A(\ab[24][3] ), .ZN(net85109) );
  NOR2_X2 U1096 ( .A1(net77914), .A2(net86101), .ZN(\ab[1][7] ) );
  INV_X4 U1097 ( .A(n1650), .ZN(n363) );
  INV_X4 U1098 ( .A(\ab[13][4] ), .ZN(n1530) );
  NOR2_X1 U1099 ( .A1(net77878), .A2(net70441), .ZN(\ab[27][2] ) );
  NOR2_X2 U1100 ( .A1(net77886), .A2(net70455), .ZN(\ab[20][3] ) );
  NOR2_X1 U1101 ( .A1(net77866), .A2(net70441), .ZN(\ab[27][1] ) );
  NOR2_X1 U1102 ( .A1(n1078), .A2(net77858), .ZN(\ab[31][0] ) );
  NOR2_X2 U1103 ( .A1(net81673), .A2(net77882), .ZN(\ab[0][3] ) );
  INV_X8 U1104 ( .A(A[23]), .ZN(net70449) );
  INV_X4 U1105 ( .A(n2325), .ZN(\CARRYB[1][3] ) );
  NOR2_X2 U1106 ( .A1(net77886), .A2(net77946), .ZN(\ab[5][3] ) );
  NOR2_X1 U1107 ( .A1(net77892), .A2(net77946), .ZN(\ab[5][4] ) );
  NAND3_X2 U1108 ( .A1(n744), .A2(net82534), .A3(n743), .ZN(\CARRYB[17][1] )
         );
  NAND2_X2 U1109 ( .A1(\CARRYB[16][1] ), .A2(\SUMB[16][2] ), .ZN(n744) );
  INV_X4 U1110 ( .A(\ab[20][1] ), .ZN(net89997) );
  NOR2_X1 U1111 ( .A1(net77858), .A2(net70441), .ZN(\ab[27][0] ) );
  NOR2_X2 U1112 ( .A1(net77866), .A2(net77956), .ZN(\ab[4][1] ) );
  NOR2_X1 U1113 ( .A1(net77858), .A2(net70443), .ZN(\ab[26][0] ) );
  AND2_X2 U1114 ( .A1(A[29]), .A2(net77864), .ZN(n344) );
  AND2_X2 U1115 ( .A1(A[28]), .A2(net77864), .ZN(n345) );
  INV_X16 U1116 ( .A(B[1]), .ZN(net77866) );
  INV_X4 U1117 ( .A(n215), .ZN(n428) );
  NAND3_X1 U1118 ( .A1(net84998), .A2(net84999), .A3(net85000), .ZN(n346) );
  AND2_X2 U1119 ( .A1(\ab[0][29] ), .A2(\ab[1][28] ), .ZN(n347) );
  AND3_X4 U1120 ( .A1(n809), .A2(net80686), .A3(net93918), .ZN(n348) );
  INV_X4 U1121 ( .A(\CARRYB[4][10] ), .ZN(n1029) );
  AND2_X2 U1122 ( .A1(\ab[0][26] ), .A2(\ab[1][25] ), .ZN(n349) );
  AND2_X2 U1123 ( .A1(\ab[0][7] ), .A2(\ab[1][6] ), .ZN(n350) );
  NAND3_X1 U1124 ( .A1(net80942), .A2(net80941), .A3(net80940), .ZN(n351) );
  OR2_X2 U1125 ( .A1(\ab[16][10] ), .A2(\CARRYB[15][10] ), .ZN(n352) );
  INV_X4 U1127 ( .A(net90174), .ZN(net88177) );
  INV_X4 U1128 ( .A(n2332), .ZN(\CARRYB[1][10] ) );
  OR2_X4 U1129 ( .A1(net82850), .A2(n714), .ZN(n354) );
  INV_X4 U1130 ( .A(n2346), .ZN(n1692) );
  XOR2_X2 U1131 ( .A(\ab[1][30] ), .B(\ab[0][31] ), .Z(n355) );
  OR2_X2 U1132 ( .A1(\ab[9][3] ), .A2(n728), .ZN(n356) );
  INV_X1 U1133 ( .A(n1111), .ZN(net82238) );
  INV_X4 U1134 ( .A(net82238), .ZN(net82239) );
  INV_X2 U1135 ( .A(\ab[5][11] ), .ZN(net83351) );
  INV_X8 U1136 ( .A(n449), .ZN(n450) );
  INV_X8 U1137 ( .A(n450), .ZN(net77948) );
  INV_X8 U1138 ( .A(n450), .ZN(net77946) );
  NOR2_X2 U1139 ( .A1(net91660), .A2(net70473), .ZN(\ab[11][10] ) );
  AND2_X2 U1140 ( .A1(B[2]), .A2(A[10]), .ZN(n357) );
  INV_X16 U1141 ( .A(A[6]), .ZN(net77940) );
  INV_X16 U1142 ( .A(n443), .ZN(n444) );
  INV_X16 U1143 ( .A(n444), .ZN(net77930) );
  INV_X4 U1144 ( .A(\ab[26][2] ), .ZN(net93792) );
  INV_X2 U1145 ( .A(\ab[19][6] ), .ZN(net81947) );
  INV_X2 U1146 ( .A(\ab[17][8] ), .ZN(net83776) );
  INV_X16 U1147 ( .A(net77864), .ZN(net77858) );
  INV_X8 U1148 ( .A(net70436), .ZN(net77864) );
  INV_X2 U1149 ( .A(\ab[22][6] ), .ZN(n824) );
  NAND2_X1 U1150 ( .A1(A[29]), .A2(net92331), .ZN(net92337) );
  NAND2_X1 U1151 ( .A1(A[28]), .A2(net92331), .ZN(net92330) );
  XOR2_X1 U1152 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  NAND2_X2 U1154 ( .A1(\SUMB[5][9] ), .A2(\CARRYB[5][8] ), .ZN(n2077) );
  NAND2_X2 U1155 ( .A1(n2377), .A2(\ab[6][8] ), .ZN(n2079) );
  XNOR2_X1 U1157 ( .A(\CARRYB[20][0] ), .B(\ab[21][0] ), .ZN(n360) );
  XNOR2_X2 U1158 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .ZN(n423) );
  XNOR2_X2 U1159 ( .A(\ab[17][2] ), .B(\SUMB[16][3] ), .ZN(n742) );
  INV_X4 U1160 ( .A(\CARRYB[2][7] ), .ZN(n566) );
  NAND2_X2 U1161 ( .A1(n1271), .A2(n1835), .ZN(n1783) );
  NAND2_X4 U1162 ( .A1(n1458), .A2(\SUMB[10][6] ), .ZN(n1460) );
  OR2_X2 U1163 ( .A1(n405), .A2(n406), .ZN(n418) );
  INV_X8 U1164 ( .A(\CARRYB[11][7] ), .ZN(n1286) );
  XNOR2_X2 U1166 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .ZN(n2328) );
  NAND3_X2 U1167 ( .A1(n1972), .A2(n1971), .A3(n1970), .ZN(\CARRYB[15][2] ) );
  NAND2_X1 U1168 ( .A1(\ab[1][11] ), .A2(\ab[0][12] ), .ZN(n1024) );
  NAND2_X4 U1169 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .ZN(n2329) );
  NAND2_X2 U1170 ( .A1(\ab[4][6] ), .A2(\CARRYB[3][6] ), .ZN(net88206) );
  NAND2_X4 U1171 ( .A1(n1633), .A2(n1634), .ZN(n1993) );
  NAND2_X4 U1172 ( .A1(n1631), .A2(n1632), .ZN(n1634) );
  XNOR2_X1 U1173 ( .A(\SUMB[2][6] ), .B(n361), .ZN(\SUMB[3][5] ) );
  XNOR2_X2 U1174 ( .A(\CARRYB[2][5] ), .B(\ab[3][5] ), .ZN(n361) );
  XNOR2_X2 U1175 ( .A(n765), .B(\CARRYB[13][2] ), .ZN(\SUMB[14][2] ) );
  INV_X2 U1176 ( .A(n395), .ZN(n1224) );
  NAND2_X2 U1177 ( .A1(\ab[8][15] ), .A2(n858), .ZN(n2252) );
  INV_X2 U1179 ( .A(\CARRYB[17][6] ), .ZN(net85610) );
  NAND2_X4 U1180 ( .A1(net92550), .A2(net92551), .ZN(net92553) );
  INV_X2 U1182 ( .A(n566), .ZN(n567) );
  BUF_X8 U1183 ( .A(net86101), .Z(net83263) );
  INV_X8 U1184 ( .A(\CARRYB[15][9] ), .ZN(n658) );
  NAND2_X2 U1185 ( .A1(\ab[15][2] ), .A2(\CARRYB[14][2] ), .ZN(n1970) );
  NAND3_X4 U1186 ( .A1(net81779), .A2(net81780), .A3(net81781), .ZN(
        \CARRYB[14][2] ) );
  INV_X8 U1187 ( .A(n389), .ZN(net85807) );
  NAND2_X4 U1188 ( .A1(\SUMB[13][11] ), .A2(\ab[14][10] ), .ZN(net82161) );
  INV_X4 U1189 ( .A(n1224), .ZN(n1225) );
  XNOR2_X2 U1190 ( .A(n1266), .B(\CARRYB[20][1] ), .ZN(\SUMB[21][1] ) );
  NAND2_X4 U1191 ( .A1(n401), .A2(n365), .ZN(\*UDW_*112679/net78533 ) );
  INV_X8 U1192 ( .A(\*UDW_*112679/net78533 ), .ZN(\CARRYB[1][18] ) );
  XNOR2_X2 U1193 ( .A(\CARRYB[7][6] ), .B(n363), .ZN(n561) );
  NAND2_X4 U1194 ( .A1(\CARRYB[21][7] ), .A2(\SUMB[21][8] ), .ZN(net80268) );
  NAND3_X1 U1195 ( .A1(n2209), .A2(n2208), .A3(n2210), .ZN(n858) );
  INV_X8 U1196 ( .A(\*UDW_*112684/net78547 ), .ZN(net87683) );
  NAND2_X4 U1197 ( .A1(\CARRYB[19][2] ), .A2(\ab[20][2] ), .ZN(n1915) );
  NAND2_X2 U1198 ( .A1(\ab[7][7] ), .A2(\CARRYB[6][7] ), .ZN(n1822) );
  INV_X4 U1199 ( .A(net87067), .ZN(n554) );
  NOR2_X4 U1200 ( .A1(net70472), .A2(net82149), .ZN(n365) );
  CLKBUF_X3 U1201 ( .A(\CARRYB[7][14] ), .Z(n833) );
  CLKBUF_X3 U1202 ( .A(n1185), .Z(n844) );
  NAND2_X1 U1203 ( .A1(\ab[13][14] ), .A2(net88756), .ZN(net82657) );
  NAND2_X1 U1204 ( .A1(\CARRYB[12][14] ), .A2(net88756), .ZN(net82658) );
  CLKBUF_X3 U1205 ( .A(\SUMB[20][3] ), .Z(net122087) );
  XNOR2_X2 U1206 ( .A(net88881), .B(\ab[7][14] ), .ZN(n797) );
  NAND2_X4 U1207 ( .A1(n602), .A2(n603), .ZN(n605) );
  BUF_X4 U1208 ( .A(n1195), .Z(n863) );
  NAND2_X4 U1209 ( .A1(\SUMB[25][3] ), .A2(\ab[26][2] ), .ZN(net80988) );
  INV_X1 U1210 ( .A(\CARRYB[20][9] ), .ZN(n369) );
  INV_X2 U1211 ( .A(n369), .ZN(n370) );
  NAND2_X4 U1212 ( .A1(\SUMB[3][11] ), .A2(\CARRYB[3][10] ), .ZN(n1394) );
  NAND2_X4 U1213 ( .A1(n604), .A2(n605), .ZN(net81995) );
  INV_X2 U1216 ( .A(\SUMB[7][14] ), .ZN(net85460) );
  INV_X2 U1217 ( .A(net122156), .ZN(net85902) );
  NAND2_X4 U1218 ( .A1(net122156), .A2(\CARRYB[23][1] ), .ZN(net80920) );
  INV_X8 U1219 ( .A(\*UDW_*112699/net78589 ), .ZN(\CARRYB[1][14] ) );
  NAND2_X4 U1220 ( .A1(\ab[1][14] ), .A2(\ab[0][15] ), .ZN(
        \*UDW_*112699/net78589 ) );
  NAND3_X2 U1221 ( .A1(n2186), .A2(n2185), .A3(n2187), .ZN(n372) );
  INV_X16 U1222 ( .A(net82149), .ZN(net80392) );
  INV_X2 U1223 ( .A(\ab[9][16] ), .ZN(n1600) );
  NOR2_X4 U1224 ( .A1(net124723), .A2(net70477), .ZN(\ab[9][16] ) );
  XNOR2_X2 U1225 ( .A(n373), .B(\SUMB[9][19] ), .ZN(\SUMB[10][18] ) );
  XNOR2_X2 U1226 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .ZN(n373) );
  INV_X2 U1227 ( .A(\ab[10][10] ), .ZN(net81643) );
  NOR2_X4 U1228 ( .A1(net91660), .A2(net70475), .ZN(\ab[10][10] ) );
  INV_X1 U1229 ( .A(\ab[7][20] ), .ZN(net81340) );
  NAND2_X4 U1230 ( .A1(n1590), .A2(n1591), .ZN(n1694) );
  NAND2_X2 U1231 ( .A1(n1035), .A2(n1036), .ZN(\SUMB[26][5] ) );
  XNOR2_X2 U1232 ( .A(net88776), .B(net85903), .ZN(n597) );
  INV_X4 U1233 ( .A(n105), .ZN(n374) );
  INV_X8 U1234 ( .A(\SUMB[15][11] ), .ZN(n375) );
  INV_X1 U1235 ( .A(\ab[16][10] ), .ZN(n376) );
  NOR2_X2 U1236 ( .A1(n374), .A2(n375), .ZN(n377) );
  NOR2_X2 U1237 ( .A1(n374), .A2(n376), .ZN(n378) );
  NOR2_X4 U1238 ( .A1(n376), .A2(n339), .ZN(n379) );
  NOR2_X4 U1239 ( .A1(n333), .A2(n352), .ZN(n380) );
  NOR2_X4 U1240 ( .A1(n383), .A2(n376), .ZN(n382) );
  NOR2_X2 U1241 ( .A1(n377), .A2(n378), .ZN(n384) );
  NOR2_X2 U1242 ( .A1(\SUMB[15][11] ), .A2(\ab[16][10] ), .ZN(n385) );
  NOR2_X4 U1243 ( .A1(n374), .A2(n375), .ZN(n386) );
  INV_X4 U1244 ( .A(n386), .ZN(n383) );
  NOR2_X4 U1245 ( .A1(n379), .A2(n380), .ZN(n387) );
  NOR2_X4 U1246 ( .A1(n381), .A2(n382), .ZN(n388) );
  NAND2_X4 U1247 ( .A1(n387), .A2(n388), .ZN(n389) );
  OR2_X4 U1248 ( .A1(n375), .A2(n376), .ZN(n391) );
  AND2_X2 U1249 ( .A1(n105), .A2(n385), .ZN(n381) );
  NAND2_X4 U1250 ( .A1(\ab[22][7] ), .A2(net89461), .ZN(net80267) );
  XNOR2_X2 U1251 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .ZN(n754) );
  INV_X2 U1252 ( .A(n279), .ZN(net119927) );
  AND2_X2 U1253 ( .A1(n247), .A2(\SUMB[22][4] ), .ZN(n407) );
  INV_X8 U1254 ( .A(n416), .ZN(net86519) );
  NAND2_X4 U1255 ( .A1(\CARRYB[23][1] ), .A2(\ab[24][1] ), .ZN(net80922) );
  NAND2_X4 U1256 ( .A1(\SUMB[20][4] ), .A2(\ab[21][3] ), .ZN(net80510) );
  INV_X4 U1257 ( .A(\ab[21][3] ), .ZN(net82834) );
  NAND2_X2 U1258 ( .A1(\ab[19][2] ), .A2(n2373), .ZN(n1911) );
  OAI21_X2 U1259 ( .B1(n1499), .B2(\CARRYB[6][7] ), .A(n1443), .ZN(n1821) );
  NAND3_X4 U1260 ( .A1(n1330), .A2(n1331), .A3(n1332), .ZN(\CARRYB[6][7] ) );
  NAND2_X1 U1261 ( .A1(\ab[6][6] ), .A2(\SUMB[5][7] ), .ZN(n1950) );
  XNOR2_X2 U1262 ( .A(\CARRYB[25][5] ), .B(\ab[26][5] ), .ZN(n393) );
  INV_X4 U1263 ( .A(net85902), .ZN(net85903) );
  INV_X2 U1264 ( .A(\SUMB[1][20] ), .ZN(n1012) );
  NAND3_X2 U1265 ( .A1(net80925), .A2(net80924), .A3(net80926), .ZN(n394) );
  NAND2_X4 U1266 ( .A1(n972), .A2(n1256), .ZN(n2070) );
  INV_X1 U1267 ( .A(n1160), .ZN(n972) );
  INV_X4 U1268 ( .A(\SUMB[7][15] ), .ZN(n602) );
  NAND2_X2 U1269 ( .A1(\SUMB[7][15] ), .A2(\ab[8][14] ), .ZN(n604) );
  XNOR2_X2 U1270 ( .A(\SUMB[13][17] ), .B(n2188), .ZN(\SUMB[14][16] ) );
  INV_X4 U1271 ( .A(\ab[13][8] ), .ZN(net80694) );
  NOR2_X4 U1272 ( .A1(net77920), .A2(net70469), .ZN(\ab[13][8] ) );
  NOR2_X4 U1273 ( .A1(net70452), .A2(net70471), .ZN(\ab[12][9] ) );
  NAND2_X4 U1274 ( .A1(n1159), .A2(n1160), .ZN(n1162) );
  INV_X8 U1276 ( .A(net89103), .ZN(net89104) );
  NAND2_X4 U1277 ( .A1(n506), .A2(n507), .ZN(net89447) );
  NAND2_X4 U1278 ( .A1(n504), .A2(n505), .ZN(n507) );
  NAND2_X4 U1279 ( .A1(n2248), .A2(n1593), .ZN(n1594) );
  XNOR2_X2 U1280 ( .A(n1584), .B(n1202), .ZN(n395) );
  NAND2_X4 U1281 ( .A1(n395), .A2(\ab[15][4] ), .ZN(n1706) );
  NOR2_X2 U1282 ( .A1(n411), .A2(n412), .ZN(n415) );
  NAND2_X2 U1283 ( .A1(\SUMB[1][21] ), .A2(\CARRYB[1][20] ), .ZN(n2053) );
  INV_X1 U1284 ( .A(\SUMB[1][21] ), .ZN(n1683) );
  NAND3_X4 U1285 ( .A1(net82030), .A2(net82029), .A3(net82031), .ZN(
        \CARRYB[3][16] ) );
  NAND2_X4 U1286 ( .A1(net148828), .A2(net148829), .ZN(n490) );
  NAND2_X4 U1287 ( .A1(n1536), .A2(n1535), .ZN(n1758) );
  INV_X4 U1288 ( .A(net92318), .ZN(n607) );
  NAND2_X4 U1289 ( .A1(n366), .A2(\ab[22][4] ), .ZN(net79993) );
  NAND3_X2 U1290 ( .A1(n1406), .A2(net86651), .A3(net86652), .ZN(
        \CARRYB[16][0] ) );
  NOR2_X4 U1291 ( .A1(net77866), .A2(net70445), .ZN(\ab[25][1] ) );
  INV_X4 U1292 ( .A(\ab[6][17] ), .ZN(n2045) );
  NAND2_X4 U1293 ( .A1(n1490), .A2(\ab[6][17] ), .ZN(n2046) );
  NAND2_X2 U1294 ( .A1(\ab[6][17] ), .A2(n1490), .ZN(n2247) );
  NOR2_X4 U1295 ( .A1(net123000), .A2(net77940), .ZN(\ab[6][17] ) );
  INV_X2 U1296 ( .A(net120585), .ZN(net124434) );
  NAND2_X4 U1297 ( .A1(net120585), .A2(net120586), .ZN(n1020) );
  INV_X4 U1298 ( .A(\ab[10][14] ), .ZN(n1037) );
  NOR2_X2 U1299 ( .A1(net84698), .A2(net70475), .ZN(\ab[10][14] ) );
  NAND2_X4 U1300 ( .A1(n710), .A2(\SUMB[1][19] ), .ZN(n1713) );
  NAND2_X4 U1301 ( .A1(\SUMB[1][19] ), .A2(\ab[2][18] ), .ZN(n1712) );
  INV_X2 U1302 ( .A(\SUMB[1][19] ), .ZN(n1498) );
  INV_X8 U1303 ( .A(n2340), .ZN(\SUMB[1][19] ) );
  NAND2_X4 U1304 ( .A1(\SUMB[1][14] ), .A2(net124833), .ZN(n454) );
  INV_X2 U1305 ( .A(net87935), .ZN(net121285) );
  NAND2_X4 U1306 ( .A1(\ab[15][9] ), .A2(\SUMB[14][10] ), .ZN(n828) );
  INV_X4 U1307 ( .A(\ab[15][9] ), .ZN(n830) );
  NOR2_X4 U1308 ( .A1(net70452), .A2(net70465), .ZN(\ab[15][9] ) );
  NAND2_X4 U1309 ( .A1(n1592), .A2(n570), .ZN(n1595) );
  NAND2_X4 U1310 ( .A1(net86162), .A2(net80834), .ZN(net84445) );
  NOR2_X4 U1311 ( .A1(net70470), .A2(net70491), .ZN(\ab[2][18] ) );
  NAND2_X4 U1312 ( .A1(n414), .A2(n415), .ZN(n416) );
  NOR2_X4 U1313 ( .A1(n409), .A2(n410), .ZN(n414) );
  INV_X2 U1314 ( .A(net124949), .ZN(net88867) );
  NOR2_X1 U1315 ( .A1(net77878), .A2(net77970), .ZN(\ab[2][2] ) );
  NAND2_X4 U1316 ( .A1(net147928), .A2(net147929), .ZN(n678) );
  INV_X1 U1317 ( .A(n795), .ZN(n796) );
  NAND2_X2 U1318 ( .A1(net84209), .A2(n795), .ZN(net84212) );
  NOR2_X1 U1319 ( .A1(net77868), .A2(net70473), .ZN(\ab[11][1] ) );
  NOR2_X1 U1320 ( .A1(net77868), .A2(net70471), .ZN(\ab[12][1] ) );
  NAND2_X1 U1321 ( .A1(\CARRYB[4][20] ), .A2(\SUMB[4][21] ), .ZN(n1883) );
  NAND3_X2 U1322 ( .A1(n750), .A2(n751), .A3(n752), .ZN(n398) );
  XNOR2_X2 U1323 ( .A(\CARRYB[13][13] ), .B(n400), .ZN(n399) );
  INV_X4 U1324 ( .A(n399), .ZN(net83445) );
  XNOR2_X2 U1325 ( .A(n736), .B(\SUMB[12][2] ), .ZN(\SUMB[13][1] ) );
  NAND3_X2 U1326 ( .A1(net81110), .A2(net81111), .A3(net81112), .ZN(
        \CARRYB[18][2] ) );
  XNOR2_X2 U1327 ( .A(\SUMB[26][4] ), .B(n1758), .ZN(n402) );
  XNOR2_X2 U1328 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .ZN(n574) );
  NAND2_X4 U1329 ( .A1(n1529), .A2(n2064), .ZN(n1496) );
  INV_X8 U1330 ( .A(n1486), .ZN(n1345) );
  XNOR2_X2 U1331 ( .A(n683), .B(net89461), .ZN(net89402) );
  INV_X8 U1332 ( .A(net80264), .ZN(n683) );
  NAND2_X2 U1333 ( .A1(\ab[15][3] ), .A2(\SUMB[14][4] ), .ZN(n1992) );
  NAND2_X2 U1334 ( .A1(\ab[13][2] ), .A2(n19), .ZN(n762) );
  NOR2_X1 U1335 ( .A1(net77878), .A2(net70469), .ZN(\ab[13][2] ) );
  NOR2_X4 U1336 ( .A1(net85716), .A2(net70467), .ZN(\ab[14][11] ) );
  NAND2_X2 U1337 ( .A1(\CARRYB[20][5] ), .A2(\ab[21][5] ), .ZN(net79989) );
  INV_X4 U1338 ( .A(\ab[12][11] ), .ZN(net84824) );
  NAND2_X2 U1339 ( .A1(net90604), .A2(\ab[12][11] ), .ZN(net84825) );
  NAND2_X1 U1340 ( .A1(\ab[12][11] ), .A2(net90604), .ZN(n806) );
  NOR2_X4 U1341 ( .A1(net85716), .A2(net70471), .ZN(\ab[12][11] ) );
  NAND2_X2 U1342 ( .A1(\ab[3][19] ), .A2(\SUMB[2][20] ), .ZN(n2055) );
  NAND2_X2 U1343 ( .A1(\ab[2][21] ), .A2(\CARRYB[1][21] ), .ZN(n2189) );
  NAND2_X2 U1344 ( .A1(net80862), .A2(\SUMB[21][5] ), .ZN(net147926) );
  INV_X4 U1345 ( .A(\ab[14][6] ), .ZN(n1607) );
  NOR2_X2 U1346 ( .A1(net77908), .A2(net70467), .ZN(\ab[14][6] ) );
  NAND3_X4 U1347 ( .A1(n1414), .A2(n1415), .A3(n1416), .ZN(\CARRYB[18][3] ) );
  XNOR2_X2 U1348 ( .A(\SUMB[13][3] ), .B(\ab[14][2] ), .ZN(n765) );
  NAND2_X4 U1349 ( .A1(\CARRYB[25][1] ), .A2(\ab[26][1] ), .ZN(net83976) );
  NAND2_X4 U1350 ( .A1(n1363), .A2(net148754), .ZN(n1365) );
  NAND2_X2 U1351 ( .A1(net92317), .A2(net92318), .ZN(n608) );
  NAND2_X4 U1352 ( .A1(\CARRYB[20][4] ), .A2(\ab[21][4] ), .ZN(n1882) );
  INV_X4 U1353 ( .A(\ab[21][4] ), .ZN(n945) );
  NAND2_X4 U1354 ( .A1(\CARRYB[17][3] ), .A2(n424), .ZN(n1414) );
  NAND2_X4 U1355 ( .A1(\SUMB[16][4] ), .A2(\CARRYB[16][3] ), .ZN(n2108) );
  XNOR2_X2 U1356 ( .A(\CARRYB[16][3] ), .B(n2013), .ZN(n559) );
  NAND3_X4 U1357 ( .A1(n1130), .A2(n1129), .A3(n1131), .ZN(\CARRYB[16][3] ) );
  NAND2_X2 U1358 ( .A1(net93747), .A2(n826), .ZN(net80879) );
  XNOR2_X2 U1359 ( .A(\SUMB[2][5] ), .B(n403), .ZN(\SUMB[3][4] ) );
  XNOR2_X2 U1360 ( .A(\CARRYB[2][4] ), .B(\ab[3][4] ), .ZN(n403) );
  NAND2_X4 U1361 ( .A1(\SUMB[25][3] ), .A2(n30), .ZN(net80989) );
  INV_X4 U1362 ( .A(\ab[23][3] ), .ZN(n406) );
  NOR2_X4 U1363 ( .A1(n404), .A2(n406), .ZN(n408) );
  NOR2_X2 U1364 ( .A1(n422), .A2(n404), .ZN(n411) );
  NAND2_X4 U1365 ( .A1(n418), .A2(n413), .ZN(n417) );
  NOR2_X1 U1366 ( .A1(net77886), .A2(net70449), .ZN(\ab[23][3] ) );
  NAND2_X2 U1367 ( .A1(\CARRYB[15][3] ), .A2(\SUMB[15][4] ), .ZN(n1129) );
  INV_X4 U1368 ( .A(net91003), .ZN(net87364) );
  NAND2_X4 U1369 ( .A1(\SUMB[9][12] ), .A2(\ab[10][11] ), .ZN(net80957) );
  NAND2_X4 U1370 ( .A1(net123143), .A2(n909), .ZN(net91301) );
  NAND2_X4 U1371 ( .A1(\SUMB[1][18] ), .A2(net87683), .ZN(net82028) );
  NAND2_X4 U1372 ( .A1(n641), .A2(n642), .ZN(n644) );
  AND3_X4 U1373 ( .A1(net88295), .A2(net88296), .A3(net88297), .ZN(n510) );
  INV_X4 U1374 ( .A(\ab[10][11] ), .ZN(net83876) );
  NOR2_X4 U1375 ( .A1(net85716), .A2(net70475), .ZN(\ab[10][11] ) );
  NAND2_X1 U1376 ( .A1(\SUMB[2][20] ), .A2(\CARRYB[2][19] ), .ZN(n2056) );
  NAND3_X4 U1377 ( .A1(n747), .A2(n746), .A3(n745), .ZN(\CARRYB[18][1] ) );
  NAND2_X2 U1378 ( .A1(\SUMB[17][2] ), .A2(\ab[18][1] ), .ZN(n745) );
  INV_X4 U1379 ( .A(\ab[12][9] ), .ZN(n1054) );
  XNOR2_X1 U1380 ( .A(n1902), .B(n1248), .ZN(n553) );
  XNOR2_X2 U1381 ( .A(n423), .B(n571), .ZN(\SUMB[16][2] ) );
  NAND2_X4 U1382 ( .A1(\ab[8][6] ), .A2(\SUMB[7][7] ), .ZN(n1826) );
  INV_X2 U1383 ( .A(\ab[8][6] ), .ZN(n1650) );
  NOR2_X1 U1384 ( .A1(net77906), .A2(net77924), .ZN(\ab[8][6] ) );
  NAND2_X4 U1385 ( .A1(\SUMB[17][4] ), .A2(\ab[18][3] ), .ZN(n1415) );
  NAND2_X4 U1386 ( .A1(n1721), .A2(n1228), .ZN(n1152) );
  INV_X4 U1387 ( .A(n1228), .ZN(n1151) );
  BUF_X4 U1388 ( .A(n864), .Z(n1228) );
  XNOR2_X2 U1389 ( .A(n1936), .B(n863), .ZN(n424) );
  INV_X2 U1390 ( .A(\ab[9][11] ), .ZN(net86894) );
  NOR2_X2 U1391 ( .A1(net70456), .A2(net70477), .ZN(\ab[9][11] ) );
  INV_X4 U1392 ( .A(net87874), .ZN(net88638) );
  INV_X2 U1393 ( .A(\SUMB[20][5] ), .ZN(net87874) );
  NAND2_X2 U1394 ( .A1(\ab[2][10] ), .A2(\CARRYB[1][10] ), .ZN(n1652) );
  NAND2_X4 U1395 ( .A1(net92321), .A2(net92325), .ZN(n834) );
  XNOR2_X2 U1396 ( .A(\CARRYB[19][1] ), .B(net89997), .ZN(n425) );
  NAND2_X2 U1397 ( .A1(\ab[21][8] ), .A2(\SUMB[20][9] ), .ZN(net81037) );
  NAND2_X4 U1398 ( .A1(n1642), .A2(n587), .ZN(n1485) );
  NAND2_X2 U1399 ( .A1(\CARRYB[20][0] ), .A2(\SUMB[20][1] ), .ZN(n1805) );
  INV_X4 U1400 ( .A(\ab[27][1] ), .ZN(net81867) );
  NAND2_X2 U1401 ( .A1(n1023), .A2(net120501), .ZN(n1025) );
  NAND2_X4 U1402 ( .A1(\ab[4][13] ), .A2(\SUMB[3][14] ), .ZN(n2090) );
  NAND2_X4 U1403 ( .A1(\SUMB[18][5] ), .A2(\ab[19][4] ), .ZN(n2235) );
  INV_X4 U1404 ( .A(net86884), .ZN(net89103) );
  NOR2_X4 U1405 ( .A1(net82247), .A2(net120391), .ZN(\ab[0][13] ) );
  INV_X2 U1406 ( .A(n1190), .ZN(n544) );
  NAND2_X4 U1407 ( .A1(\SUMB[20][5] ), .A2(\CARRYB[20][4] ), .ZN(net82408) );
  INV_X4 U1408 ( .A(net82009), .ZN(net88856) );
  NAND2_X2 U1409 ( .A1(\CARRYB[3][13] ), .A2(\SUMB[3][14] ), .ZN(n2091) );
  XNOR2_X2 U1410 ( .A(n35), .B(n426), .ZN(\SUMB[14][1] ) );
  XNOR2_X2 U1411 ( .A(\SUMB[13][2] ), .B(\ab[14][1] ), .ZN(n426) );
  XNOR2_X2 U1412 ( .A(\ab[20][2] ), .B(\SUMB[19][3] ), .ZN(n1232) );
  NAND2_X4 U1413 ( .A1(\SUMB[1][14] ), .A2(\CARRYB[1][13] ), .ZN(n453) );
  NOR2_X1 U1414 ( .A1(net83784), .A2(net77932), .ZN(\ab[7][12] ) );
  INV_X2 U1415 ( .A(\ab[7][12] ), .ZN(net85251) );
  NAND2_X4 U1416 ( .A1(n895), .A2(net123430), .ZN(n2338) );
  NAND2_X4 U1417 ( .A1(\SUMB[10][12] ), .A2(\ab[11][11] ), .ZN(net81167) );
  INV_X4 U1418 ( .A(\SUMB[9][13] ), .ZN(net120652) );
  NAND2_X4 U1419 ( .A1(net119976), .A2(\SUMB[4][16] ), .ZN(net84446) );
  INV_X4 U1420 ( .A(\ab[24][2] ), .ZN(net121380) );
  NAND2_X2 U1421 ( .A1(net124627), .A2(net81947), .ZN(n518) );
  NAND2_X2 U1422 ( .A1(\SUMB[4][10] ), .A2(n943), .ZN(n1398) );
  INV_X4 U1423 ( .A(\ab[11][9] ), .ZN(net93305) );
  NOR2_X2 U1424 ( .A1(net70452), .A2(net70473), .ZN(\ab[11][9] ) );
  BUF_X8 U1425 ( .A(n424), .Z(n1241) );
  NAND2_X4 U1426 ( .A1(\SUMB[16][4] ), .A2(\ab[17][3] ), .ZN(n2107) );
  INV_X4 U1427 ( .A(\ab[17][3] ), .ZN(n2013) );
  XNOR2_X2 U1428 ( .A(\CARRYB[18][2] ), .B(\ab[19][2] ), .ZN(n1254) );
  NAND2_X2 U1429 ( .A1(\ab[14][2] ), .A2(\SUMB[13][3] ), .ZN(net81779) );
  INV_X4 U1430 ( .A(net92317), .ZN(n606) );
  NAND2_X4 U1431 ( .A1(net82009), .A2(\ab[19][6] ), .ZN(n519) );
  NAND2_X4 U1432 ( .A1(n4), .A2(net148179), .ZN(net80668) );
  NAND3_X4 U1433 ( .A1(net80472), .A2(net80473), .A3(net80474), .ZN(n427) );
  INV_X8 U1434 ( .A(n427), .ZN(net92318) );
  NAND3_X2 U1435 ( .A1(net86022), .A2(net79907), .A3(n784), .ZN(net86024) );
  NAND3_X2 U1436 ( .A1(n250), .A2(net79885), .A3(net79884), .ZN(net87797) );
  NAND3_X2 U1437 ( .A1(net81157), .A2(n690), .A3(n689), .ZN(n835) );
  NAND2_X2 U1438 ( .A1(n584), .A2(n583), .ZN(net89110) );
  OAI211_X4 U1439 ( .C1(n428), .C2(n429), .A(n2298), .B(n2297), .ZN(
        \CARRYB[8][16] ) );
  INV_X1 U1440 ( .A(\ab[8][16] ), .ZN(n429) );
  XNOR2_X2 U1441 ( .A(n1094), .B(\SUMB[10][16] ), .ZN(\SUMB[11][15] ) );
  XNOR2_X2 U1442 ( .A(n926), .B(\CARRYB[7][17] ), .ZN(net88703) );
  NAND3_X2 U1443 ( .A1(n1528), .A2(n1892), .A3(n2205), .ZN(n1497) );
  NAND2_X2 U1444 ( .A1(\CARRYB[24][3] ), .A2(\SUMB[24][4] ), .ZN(net81006) );
  NAND2_X4 U1445 ( .A1(net88105), .A2(net89021), .ZN(n436) );
  NAND2_X4 U1446 ( .A1(net88107), .A2(n436), .ZN(\SUMB[7][11] ) );
  INV_X4 U1447 ( .A(net88106), .ZN(net89021) );
  NAND2_X2 U1448 ( .A1(net88106), .A2(net81209), .ZN(net88107) );
  INV_X4 U1449 ( .A(net81209), .ZN(net88105) );
  NAND2_X4 U1450 ( .A1(n432), .A2(n433), .ZN(\SUMB[6][12] ) );
  NAND2_X2 U1451 ( .A1(\ab[7][11] ), .A2(\SUMB[6][12] ), .ZN(net81212) );
  NAND2_X2 U1452 ( .A1(\SUMB[6][12] ), .A2(\CARRYB[6][11] ), .ZN(net81213) );
  NAND2_X4 U1453 ( .A1(n430), .A2(n431), .ZN(n433) );
  INV_X2 U1454 ( .A(\SUMB[5][13] ), .ZN(n431) );
  INV_X2 U1455 ( .A(n431), .ZN(n434) );
  INV_X4 U1456 ( .A(net82089), .ZN(n430) );
  NAND2_X2 U1457 ( .A1(net82089), .A2(n434), .ZN(n432) );
  NAND2_X4 U1458 ( .A1(net87462), .A2(n435), .ZN(net81209) );
  NAND2_X4 U1459 ( .A1(net87460), .A2(net87461), .ZN(n435) );
  INV_X4 U1460 ( .A(net83045), .ZN(net87461) );
  INV_X1 U1461 ( .A(\ab[7][11] ), .ZN(net83045) );
  NAND2_X2 U1462 ( .A1(net83045), .A2(\CARRYB[6][11] ), .ZN(net87462) );
  INV_X4 U1463 ( .A(\CARRYB[6][11] ), .ZN(net87460) );
  NAND2_X2 U1464 ( .A1(\SUMB[5][13] ), .A2(n1439), .ZN(net81714) );
  NAND2_X2 U1465 ( .A1(\SUMB[5][13] ), .A2(\ab[6][12] ), .ZN(net81713) );
  NAND2_X2 U1466 ( .A1(\ab[7][11] ), .A2(\CARRYB[6][11] ), .ZN(net81211) );
  NAND2_X4 U1467 ( .A1(n439), .A2(net88010), .ZN(n442) );
  NAND2_X4 U1468 ( .A1(n441), .A2(n442), .ZN(\SUMB[4][12] ) );
  INV_X4 U1469 ( .A(net85493), .ZN(net88010) );
  NAND2_X2 U1470 ( .A1(net89227), .A2(net85493), .ZN(n441) );
  INV_X4 U1471 ( .A(net89227), .ZN(n439) );
  NAND2_X1 U1472 ( .A1(\SUMB[3][13] ), .A2(n89), .ZN(net82760) );
  XNOR2_X2 U1473 ( .A(n438), .B(n440), .ZN(net84270) );
  CLKBUF_X3 U1474 ( .A(\SUMB[1][15] ), .Z(n440) );
  NAND2_X2 U1475 ( .A1(\SUMB[1][15] ), .A2(\ab[2][14] ), .ZN(net86170) );
  NOR2_X4 U1476 ( .A1(net70466), .A2(net82149), .ZN(\ab[0][16] ) );
  INV_X16 U1477 ( .A(A[0]), .ZN(net82149) );
  NOR2_X4 U1478 ( .A1(net70466), .A2(net80409), .ZN(net88123) );
  XNOR2_X1 U1479 ( .A(\CARRYB[1][14] ), .B(\ab[2][14] ), .ZN(n438) );
  XNOR2_X2 U1480 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .ZN(net86864) );
  XNOR2_X2 U1481 ( .A(\CARRYB[2][13] ), .B(\ab[3][13] ), .ZN(net81694) );
  INV_X8 U1482 ( .A(A[0]), .ZN(net77988) );
  NOR2_X1 U1483 ( .A1(net70456), .A2(net77930), .ZN(\ab[7][11] ) );
  INV_X4 U1484 ( .A(A[7]), .ZN(n443) );
  INV_X16 U1485 ( .A(B[11]), .ZN(net70456) );
  NAND3_X4 U1486 ( .A1(n445), .A2(n447), .A3(n446), .ZN(\CARRYB[6][11] ) );
  NAND2_X4 U1487 ( .A1(net84652), .A2(\ab[6][11] ), .ZN(n447) );
  INV_X4 U1488 ( .A(n146), .ZN(net84652) );
  NAND2_X4 U1489 ( .A1(net90731), .A2(net84652), .ZN(n445) );
  NAND2_X4 U1490 ( .A1(\SUMB[5][12] ), .A2(\ab[6][11] ), .ZN(n446) );
  XNOR2_X2 U1491 ( .A(net86151), .B(n448), .ZN(\SUMB[5][12] ) );
  NAND2_X2 U1492 ( .A1(net86151), .A2(n448), .ZN(net121455) );
  INV_X2 U1493 ( .A(n448), .ZN(net121454) );
  INV_X2 U1494 ( .A(net86151), .ZN(net121453) );
  NAND2_X2 U1495 ( .A1(\SUMB[4][13] ), .A2(\CARRYB[4][12] ), .ZN(net81206) );
  NAND2_X2 U1496 ( .A1(\ab[5][12] ), .A2(\SUMB[4][13] ), .ZN(net81205) );
  NAND3_X4 U1497 ( .A1(net82762), .A2(net82763), .A3(n451), .ZN(
        \CARRYB[5][11] ) );
  NAND2_X1 U1498 ( .A1(\ab[5][11] ), .A2(\CARRYB[4][11] ), .ZN(n451) );
  NAND2_X4 U1499 ( .A1(\SUMB[4][12] ), .A2(\ab[5][11] ), .ZN(net82763) );
  NAND2_X4 U1500 ( .A1(\SUMB[4][12] ), .A2(net124527), .ZN(net82762) );
  NAND3_X1 U1501 ( .A1(net88084), .A2(net88085), .A3(net88086), .ZN(net124527)
         );
  NAND3_X2 U1502 ( .A1(net88084), .A2(net88085), .A3(net88086), .ZN(
        \CARRYB[4][11] ) );
  NAND2_X1 U1503 ( .A1(\CARRYB[4][11] ), .A2(net83351), .ZN(net147922) );
  NOR2_X4 U1504 ( .A1(net70456), .A2(net77946), .ZN(\ab[5][11] ) );
  INV_X8 U1505 ( .A(A[5]), .ZN(n449) );
  NAND2_X1 U1506 ( .A1(net82757), .A2(\SUMB[4][12] ), .ZN(net123899) );
  INV_X2 U1507 ( .A(\SUMB[4][12] ), .ZN(net123898) );
  NAND2_X2 U1508 ( .A1(\SUMB[3][12] ), .A2(\CARRYB[3][11] ), .ZN(net88084) );
  NAND2_X4 U1509 ( .A1(\SUMB[3][12] ), .A2(\ab[4][11] ), .ZN(net88085) );
  NAND3_X4 U1510 ( .A1(n454), .A2(n453), .A3(n455), .ZN(\CARRYB[2][13] ) );
  NAND2_X2 U1511 ( .A1(n99), .A2(\ab[3][13] ), .ZN(net81515) );
  NAND2_X2 U1512 ( .A1(net124833), .A2(\CARRYB[1][13] ), .ZN(n455) );
  XNOR2_X2 U1513 ( .A(\CARRYB[1][13] ), .B(\ab[2][13] ), .ZN(n456) );
  NAND2_X2 U1514 ( .A1(\ab[0][14] ), .A2(\ab[1][13] ), .ZN(n452) );
  INV_X8 U1515 ( .A(\*UDW_*112699/net78591 ), .ZN(\SUMB[1][14] ) );
  XNOR2_X2 U1516 ( .A(n456), .B(\SUMB[1][14] ), .ZN(\SUMB[2][13] ) );
  XNOR2_X2 U1517 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .ZN(
        \*UDW_*112699/net78591 ) );
  NOR2_X4 U1518 ( .A1(net80727), .A2(n175), .ZN(\ab[2][20] ) );
  NOR2_X4 U1519 ( .A1(net70460), .A2(net70491), .ZN(\ab[2][13] ) );
  INV_X16 U1520 ( .A(A[2]), .ZN(net70491) );
  INV_X16 U1521 ( .A(net120392), .ZN(net70460) );
  INV_X4 U1522 ( .A(net120391), .ZN(net120392) );
  XNOR2_X2 U1523 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .ZN(
        \*UDW_*112704/net78605 ) );
  INV_X8 U1524 ( .A(B[14]), .ZN(net70462) );
  NOR2_X4 U1525 ( .A1(net70462), .A2(net86101), .ZN(\ab[1][14] ) );
  NAND2_X4 U1526 ( .A1(n458), .A2(net83062), .ZN(net81256) );
  INV_X4 U1528 ( .A(net81256), .ZN(net84069) );
  NAND2_X2 U1529 ( .A1(\CARRYB[9][10] ), .A2(net81643), .ZN(net83062) );
  INV_X4 U1530 ( .A(\CARRYB[9][10] ), .ZN(net83061) );
  NAND3_X4 U1531 ( .A1(net81001), .A2(n457), .A3(net87458), .ZN(
        \CARRYB[9][10] ) );
  NAND2_X2 U1532 ( .A1(\CARRYB[9][10] ), .A2(\ab[10][10] ), .ZN(net81260) );
  NAND2_X2 U1533 ( .A1(\SUMB[9][11] ), .A2(\CARRYB[9][10] ), .ZN(net81262) );
  NAND2_X4 U1534 ( .A1(\SUMB[8][11] ), .A2(\ab[9][10] ), .ZN(n457) );
  NAND2_X4 U1535 ( .A1(net91298), .A2(\SUMB[8][11] ), .ZN(net81001) );
  INV_X4 U1536 ( .A(net87457), .ZN(net91298) );
  INV_X4 U1537 ( .A(n2378), .ZN(net87457) );
  NAND2_X4 U1538 ( .A1(net91259), .A2(\ab[10][10] ), .ZN(net81261) );
  INV_X4 U1539 ( .A(A[10]), .ZN(net70475) );
  INV_X8 U1540 ( .A(B[10]), .ZN(net70454) );
  NAND2_X4 U1541 ( .A1(net87458), .A2(net87459), .ZN(net83736) );
  NAND2_X2 U1542 ( .A1(\CARRYB[8][10] ), .A2(\ab[9][10] ), .ZN(net87458) );
  INV_X1 U1543 ( .A(\ab[9][10] ), .ZN(net87456) );
  NAND3_X4 U1544 ( .A1(A[10]), .A2(B[2]), .A3(net147421), .ZN(net147451) );
  NAND2_X2 U1545 ( .A1(net81630), .A2(B[10]), .ZN(net90174) );
  NAND2_X2 U1546 ( .A1(\CARRYB[12][8] ), .A2(\ab[13][8] ), .ZN(net80507) );
  NAND3_X2 U1547 ( .A1(net80506), .A2(net80505), .A3(net80507), .ZN(
        \CARRYB[13][8] ) );
  NAND3_X4 U1548 ( .A1(net81115), .A2(n459), .A3(net81116), .ZN(
        \CARRYB[12][8] ) );
  NAND2_X2 U1549 ( .A1(net80694), .A2(\CARRYB[12][8] ), .ZN(net84712) );
  INV_X4 U1550 ( .A(\CARRYB[12][8] ), .ZN(net84710) );
  NAND2_X2 U1551 ( .A1(\SUMB[12][9] ), .A2(\CARRYB[12][8] ), .ZN(net80505) );
  NAND2_X4 U1552 ( .A1(net89537), .A2(\ab[12][8] ), .ZN(net81116) );
  NAND2_X2 U1553 ( .A1(\ab[12][8] ), .A2(\CARRYB[11][8] ), .ZN(n459) );
  NAND2_X2 U1554 ( .A1(\SUMB[11][9] ), .A2(\CARRYB[11][8] ), .ZN(net81115) );
  XNOR2_X2 U1555 ( .A(net90735), .B(net88104), .ZN(\SUMB[11][9] ) );
  BUF_X4 U1556 ( .A(\CARRYB[10][9] ), .Z(net88104) );
  INV_X2 U1557 ( .A(net88104), .ZN(net121446) );
  NAND2_X1 U1558 ( .A1(net90735), .A2(net88104), .ZN(net121447) );
  XNOR2_X1 U1559 ( .A(n183), .B(net88104), .ZN(net149580) );
  INV_X16 U1560 ( .A(A[13]), .ZN(net70469) );
  INV_X32 U1561 ( .A(net77922), .ZN(net77920) );
  INV_X4 U1562 ( .A(net70450), .ZN(net77922) );
  INV_X8 U1563 ( .A(B[8]), .ZN(net70450) );
  NOR2_X2 U1564 ( .A1(net124610), .A2(net70450), .ZN(\ab[0][8] ) );
  INV_X1 U1565 ( .A(net89537), .ZN(net93309) );
  XNOR2_X2 U1566 ( .A(\CARRYB[11][8] ), .B(\ab[12][8] ), .ZN(net82548) );
  NAND2_X2 U1567 ( .A1(\CARRYB[10][9] ), .A2(\ab[11][9] ), .ZN(net84268) );
  NAND2_X2 U1568 ( .A1(\SUMB[10][10] ), .A2(\CARRYB[10][9] ), .ZN(net84267) );
  INV_X4 U1569 ( .A(A[9]), .ZN(net70477) );
  NAND2_X4 U1570 ( .A1(n464), .A2(n465), .ZN(\SUMB[8][11] ) );
  NAND2_X4 U1571 ( .A1(n462), .A2(n460), .ZN(n465) );
  INV_X2 U1572 ( .A(n463), .ZN(n460) );
  INV_X2 U1573 ( .A(\SUMB[7][12] ), .ZN(n463) );
  NAND2_X2 U1574 ( .A1(n463), .A2(net80993), .ZN(n464) );
  INV_X4 U1575 ( .A(net80993), .ZN(n462) );
  NAND3_X2 U1576 ( .A1(net81216), .A2(n461), .A3(net81215), .ZN(
        \CARRYB[8][10] ) );
  NAND2_X2 U1577 ( .A1(net123072), .A2(A[9]), .ZN(net123055) );
  NOR2_X2 U1578 ( .A1(net77920), .A2(net70471), .ZN(\ab[12][8] ) );
  INV_X16 U1579 ( .A(A[12]), .ZN(net70471) );
  NAND3_X4 U1580 ( .A1(net84654), .A2(n467), .A3(net84656), .ZN(
        \CARRYB[11][8] ) );
  NAND2_X4 U1581 ( .A1(n468), .A2(\ab[11][8] ), .ZN(n467) );
  XNOR2_X2 U1582 ( .A(net82723), .B(net91419), .ZN(n468) );
  NAND2_X2 U1583 ( .A1(net91419), .A2(net82723), .ZN(net120515) );
  NOR2_X1 U1584 ( .A1(net70456), .A2(net77938), .ZN(\ab[6][11] ) );
  INV_X32 U1585 ( .A(A[6]), .ZN(net77938) );
  NAND2_X4 U1586 ( .A1(n469), .A2(net81204), .ZN(net86151) );
  NAND2_X4 U1587 ( .A1(net87465), .A2(net87464), .ZN(n469) );
  INV_X16 U1588 ( .A(net77984), .ZN(net86101) );
  INV_X16 U1589 ( .A(net70493), .ZN(net77984) );
  NAND2_X4 U1590 ( .A1(B[17]), .A2(net77984), .ZN(net87050) );
  INV_X8 U1591 ( .A(B[14]), .ZN(net84698) );
  NAND2_X4 U1592 ( .A1(net84072), .A2(net84071), .ZN(\SUMB[10][10] ) );
  INV_X1 U1593 ( .A(net91259), .ZN(net84070) );
  XNOR2_X2 U1594 ( .A(n470), .B(net90687), .ZN(net91259) );
  NAND2_X2 U1595 ( .A1(net86896), .A2(net86895), .ZN(n470) );
  NAND2_X2 U1596 ( .A1(net90687), .A2(n229), .ZN(net81259) );
  NAND2_X4 U1597 ( .A1(net86895), .A2(net86896), .ZN(net83042) );
  INV_X4 U1598 ( .A(\SUMB[10][10] ), .ZN(net93304) );
  NAND2_X4 U1599 ( .A1(\SUMB[10][10] ), .A2(\ab[11][9] ), .ZN(net93306) );
  NAND2_X4 U1600 ( .A1(net84069), .A2(n70), .ZN(net84072) );
  XNOR2_X2 U1601 ( .A(net91118), .B(net83042), .ZN(\SUMB[9][11] ) );
  NAND2_X2 U1602 ( .A1(net91118), .A2(\ab[9][11] ), .ZN(net81258) );
  NAND2_X4 U1603 ( .A1(net93306), .A2(net93307), .ZN(net90735) );
  NAND2_X4 U1604 ( .A1(net93304), .A2(net93305), .ZN(net93307) );
  NAND3_X2 U1605 ( .A1(n471), .A2(n325), .A3(n472), .ZN(\CARRYB[10][9] ) );
  NAND3_X4 U1606 ( .A1(net84267), .A2(net84268), .A3(net93306), .ZN(
        \CARRYB[11][9] ) );
  INV_X16 U1607 ( .A(B[9]), .ZN(net70452) );
  INV_X4 U1608 ( .A(net91419), .ZN(net120514) );
  NAND2_X4 U1609 ( .A1(\CARRYB[10][8] ), .A2(\SUMB[10][9] ), .ZN(net84654) );
  NAND2_X4 U1610 ( .A1(net120466), .A2(net84656), .ZN(net86844) );
  NAND2_X4 U1611 ( .A1(net147936), .A2(\ab[11][8] ), .ZN(net84656) );
  INV_X1 U1612 ( .A(\ab[11][8] ), .ZN(net120464) );
  AND2_X2 U1613 ( .A1(B[6]), .A2(n341), .ZN(\ab[1][6] ) );
  NOR2_X4 U1614 ( .A1(net87396), .A2(net82149), .ZN(\ab[0][15] ) );
  NOR2_X2 U1615 ( .A1(net70460), .A2(net77964), .ZN(\ab[3][13] ) );
  NAND2_X4 U1616 ( .A1(\ab[3][13] ), .A2(\SUMB[2][14] ), .ZN(net81514) );
  INV_X16 U1617 ( .A(A[3]), .ZN(net77964) );
  INV_X32 U1618 ( .A(A[3]), .ZN(net77966) );
  NAND3_X2 U1619 ( .A1(n473), .A2(n474), .A3(n475), .ZN(\CARRYB[7][10] ) );
  NAND2_X1 U1620 ( .A1(\ab[7][10] ), .A2(\CARRYB[6][10] ), .ZN(n475) );
  NAND2_X2 U1621 ( .A1(\SUMB[6][11] ), .A2(\ab[7][10] ), .ZN(n474) );
  XNOR2_X2 U1622 ( .A(\CARRYB[6][10] ), .B(\ab[7][10] ), .ZN(net81586) );
  NAND2_X1 U1623 ( .A1(net122062), .A2(net89168), .ZN(net123143) );
  NAND2_X4 U1624 ( .A1(net119982), .A2(net88297), .ZN(net89168) );
  NOR2_X2 U1625 ( .A1(net91660), .A2(net77924), .ZN(\ab[8][10] ) );
  NAND2_X2 U1626 ( .A1(net123072), .A2(A[8]), .ZN(net123019) );
  INV_X4 U1627 ( .A(A[8]), .ZN(net77926) );
  NOR2_X4 U1628 ( .A1(net87396), .A2(net80409), .ZN(\ab[1][15] ) );
  NAND3_X4 U1630 ( .A1(net79885), .A2(net79884), .A3(net79883), .ZN(net87798)
         );
  XNOR2_X2 U1631 ( .A(net87798), .B(\ab[30][0] ), .ZN(net83536) );
  NAND2_X4 U1632 ( .A1(\CARRYB[28][0] ), .A2(net86792), .ZN(net79885) );
  XNOR2_X2 U1633 ( .A(\CARRYB[27][1] ), .B(net92330), .ZN(n476) );
  INV_X4 U1634 ( .A(net92330), .ZN(\ab[28][1] ) );
  XNOR2_X2 U1635 ( .A(\CARRYB[27][1] ), .B(\ab[28][1] ), .ZN(net149605) );
  NAND2_X4 U1636 ( .A1(net89110), .A2(\ab[28][1] ), .ZN(net79881) );
  INV_X4 U1637 ( .A(net77866), .ZN(net92331) );
  INV_X32 U1638 ( .A(B[1]), .ZN(net77868) );
  NAND2_X4 U1639 ( .A1(net87411), .A2(n344), .ZN(net79884) );
  NAND3_X2 U1640 ( .A1(net82297), .A2(n479), .A3(n480), .ZN(\CARRYB[5][14] )
         );
  INV_X8 U1641 ( .A(net83918), .ZN(net83919) );
  NAND2_X4 U1642 ( .A1(n478), .A2(net148838), .ZN(net83918) );
  NAND2_X4 U1643 ( .A1(net148836), .A2(net148837), .ZN(n478) );
  INV_X4 U1644 ( .A(net119927), .ZN(net148837) );
  NOR2_X4 U1645 ( .A1(net84698), .A2(net77948), .ZN(\ab[5][14] ) );
  INV_X1 U1646 ( .A(\ab[5][14] ), .ZN(net84946) );
  OAI21_X4 U1647 ( .B1(net119909), .B2(net119910), .A(n477), .ZN(net119908) );
  OAI21_X4 U1648 ( .B1(net119908), .B2(net123267), .A(net123266), .ZN(
        net124908) );
  NOR2_X2 U1649 ( .A1(net119949), .A2(n353), .ZN(net119948) );
  XNOR2_X2 U1650 ( .A(\CARRYB[2][15] ), .B(n353), .ZN(net121859) );
  NAND2_X2 U1651 ( .A1(n353), .A2(net119949), .ZN(net119960) );
  NAND2_X4 U1652 ( .A1(net81666), .A2(net81667), .ZN(n481) );
  NAND2_X4 U1653 ( .A1(n481), .A2(net81668), .ZN(\SUMB[16][7] ) );
  INV_X4 U1654 ( .A(n104), .ZN(net81667) );
  INV_X4 U1655 ( .A(net80906), .ZN(net81666) );
  NAND2_X4 U1656 ( .A1(net85543), .A2(n484), .ZN(\SUMB[15][8] ) );
  NAND2_X2 U1657 ( .A1(\SUMB[15][8] ), .A2(net85372), .ZN(net80566) );
  NAND2_X2 U1658 ( .A1(net80906), .A2(n104), .ZN(net81668) );
  NAND2_X2 U1659 ( .A1(\ab[16][7] ), .A2(\SUMB[15][8] ), .ZN(net80565) );
  NAND2_X4 U1660 ( .A1(net83273), .A2(\SUMB[14][9] ), .ZN(n484) );
  INV_X8 U1661 ( .A(net88904), .ZN(\SUMB[14][9] ) );
  NAND2_X4 U1662 ( .A1(\SUMB[14][9] ), .A2(\ab[15][8] ), .ZN(net80562) );
  NAND2_X4 U1663 ( .A1(net86537), .A2(\SUMB[14][9] ), .ZN(net80563) );
  XNOR2_X2 U1664 ( .A(n482), .B(n210), .ZN(net88904) );
  XNOR2_X2 U1665 ( .A(n483), .B(net85043), .ZN(n482) );
  INV_X4 U1666 ( .A(\ab[14][9] ), .ZN(n483) );
  XNOR2_X2 U1667 ( .A(\ab[15][8] ), .B(net86537), .ZN(net83273) );
  INV_X4 U1668 ( .A(net86536), .ZN(net86537) );
  NAND2_X2 U1669 ( .A1(\ab[15][8] ), .A2(net86537), .ZN(net80561) );
  XNOR2_X2 U1670 ( .A(\ab[15][8] ), .B(net86537), .ZN(net93878) );
  INV_X2 U1671 ( .A(\CARRYB[14][8] ), .ZN(net86536) );
  INV_X4 U1672 ( .A(\SUMB[14][8] ), .ZN(net86374) );
  NAND2_X4 U1673 ( .A1(net147924), .A2(net147925), .ZN(n485) );
  NAND2_X4 U1674 ( .A1(n485), .A2(net147926), .ZN(\SUMB[22][4] ) );
  INV_X4 U1675 ( .A(\SUMB[21][5] ), .ZN(net147925) );
  INV_X4 U1676 ( .A(net80862), .ZN(net147924) );
  XNOR2_X2 U1677 ( .A(net149133), .B(n71), .ZN(\SUMB[21][5] ) );
  XNOR2_X2 U1678 ( .A(\CARRYB[20][5] ), .B(\ab[21][5] ), .ZN(net149133) );
  NAND2_X2 U1679 ( .A1(\SUMB[20][6] ), .A2(\CARRYB[20][5] ), .ZN(net79991) );
  XNOR2_X2 U1680 ( .A(\CARRYB[20][5] ), .B(\ab[21][5] ), .ZN(net83705) );
  OR2_X2 U1681 ( .A1(net80986), .A2(net83623), .ZN(net83625) );
  NAND2_X4 U1682 ( .A1(net83625), .A2(net83624), .ZN(\SUMB[27][1] ) );
  NAND2_X1 U1683 ( .A1(net80986), .A2(net83623), .ZN(net83624) );
  XNOR2_X2 U1684 ( .A(net89460), .B(net81867), .ZN(net80986) );
  NAND3_X2 U1685 ( .A1(net83975), .A2(net83977), .A3(net83976), .ZN(net89460)
         );
  NAND2_X4 U1686 ( .A1(n486), .A2(n487), .ZN(net123365) );
  NAND2_X4 U1687 ( .A1(net123365), .A2(\ab[27][1] ), .ZN(net80991) );
  NAND2_X4 U1688 ( .A1(\CARRYB[26][1] ), .A2(\ab[27][1] ), .ZN(net80990) );
  NAND3_X2 U1689 ( .A1(net83975), .A2(net83977), .A3(net83976), .ZN(
        \CARRYB[26][1] ) );
  NAND2_X2 U1690 ( .A1(n486), .A2(n487), .ZN(\SUMB[26][2] ) );
  NAND2_X4 U1691 ( .A1(net93791), .A2(net121814), .ZN(n487) );
  NAND2_X4 U1692 ( .A1(net80564), .A2(n488), .ZN(net80906) );
  NAND2_X4 U1693 ( .A1(net82289), .A2(net82288), .ZN(n488) );
  INV_X2 U1694 ( .A(\ab[16][7] ), .ZN(net82288) );
  INV_X8 U1695 ( .A(\CARRYB[15][7] ), .ZN(net82289) );
  INV_X1 U1696 ( .A(net82289), .ZN(net85372) );
  NAND2_X4 U1697 ( .A1(net120364), .A2(n285), .ZN(n489) );
  NAND2_X4 U1698 ( .A1(net120366), .A2(n489), .ZN(net92790) );
  INV_X4 U1699 ( .A(net89455), .ZN(net120364) );
  INV_X2 U1700 ( .A(\SUMB[23][4] ), .ZN(net89455) );
  NAND2_X2 U1701 ( .A1(n364), .A2(net89455), .ZN(net120366) );
  XNOR2_X2 U1702 ( .A(n102), .B(net86109), .ZN(\SUMB[23][4] ) );
  NAND2_X2 U1703 ( .A1(\SUMB[23][4] ), .A2(\ab[24][3] ), .ZN(net84679) );
  XNOR2_X2 U1704 ( .A(\CARRYB[22][4] ), .B(\ab[23][4] ), .ZN(net86109) );
  NAND2_X4 U1705 ( .A1(n102), .A2(net84213), .ZN(net80290) );
  INV_X4 U1706 ( .A(net88648), .ZN(net124635) );
  INV_X1 U1707 ( .A(\CARRYB[22][5] ), .ZN(net88859) );
  XNOR2_X2 U1708 ( .A(\CARRYB[22][5] ), .B(\ab[23][5] ), .ZN(net81983) );
  NAND2_X1 U1709 ( .A1(\ab[23][5] ), .A2(\CARRYB[22][5] ), .ZN(net79904) );
  NAND2_X4 U1710 ( .A1(net84668), .A2(net84667), .ZN(\SUMB[21][6] ) );
  NAND2_X4 U1711 ( .A1(net83101), .A2(n311), .ZN(net84667) );
  NAND2_X4 U1712 ( .A1(net84666), .A2(net87681), .ZN(net84668) );
  INV_X4 U1713 ( .A(net149530), .ZN(net84666) );
  NOR2_X4 U1714 ( .A1(net77900), .A2(net70451), .ZN(\ab[22][5] ) );
  INV_X16 U1715 ( .A(A[22]), .ZN(net70451) );
  INV_X32 U1716 ( .A(net77904), .ZN(net77900) );
  INV_X16 U1717 ( .A(net70444), .ZN(net77904) );
  BUF_X8 U1718 ( .A(\CARRYB[2][15] ), .Z(net119974) );
  INV_X4 U1719 ( .A(net119960), .ZN(net119909) );
  NAND2_X2 U1720 ( .A1(net123266), .A2(net123267), .ZN(net123269) );
  INV_X2 U1721 ( .A(net119928), .ZN(net123267) );
  NOR2_X2 U1722 ( .A1(net77914), .A2(net70463), .ZN(\ab[16][7] ) );
  NAND2_X2 U1723 ( .A1(\CARRYB[15][7] ), .A2(\ab[16][7] ), .ZN(net80564) );
  INV_X16 U1724 ( .A(A[16]), .ZN(net70463) );
  INV_X32 U1725 ( .A(net77916), .ZN(net77914) );
  INV_X16 U1726 ( .A(net70448), .ZN(net77916) );
  INV_X16 U1727 ( .A(net77916), .ZN(net77912) );
  INV_X8 U1728 ( .A(B[7]), .ZN(net70448) );
  NAND3_X4 U1729 ( .A1(net80537), .A2(net80538), .A3(net80536), .ZN(
        \CARRYB[15][7] ) );
  NAND2_X2 U1730 ( .A1(\ab[15][7] ), .A2(\CARRYB[14][7] ), .ZN(net80536) );
  NAND2_X4 U1731 ( .A1(n306), .A2(n346), .ZN(net80538) );
  NAND2_X4 U1732 ( .A1(net86375), .A2(\ab[15][7] ), .ZN(net80537) );
  NAND2_X1 U1733 ( .A1(net83755), .A2(net86375), .ZN(net120519) );
  INV_X1 U1734 ( .A(net86375), .ZN(net120517) );
  INV_X16 U1735 ( .A(A[14]), .ZN(net70467) );
  NAND2_X4 U1736 ( .A1(net82295), .A2(net82294), .ZN(\SUMB[13][9] ) );
  INV_X2 U1737 ( .A(n817), .ZN(net148829) );
  BUF_X8 U1739 ( .A(net89652), .Z(net88344) );
  AOI21_X4 U1740 ( .B1(net119899), .B2(\*UDW_*112684/net78549 ), .A(net119901), 
        .ZN(net87363) );
  NAND2_X1 U1741 ( .A1(\*UDW_*112684/net78549 ), .A2(net119899), .ZN(net119920) );
  XNOR2_X2 U1742 ( .A(net119952), .B(\*UDW_*112684/net78549 ), .ZN(net119949)
         );
  NAND2_X1 U1743 ( .A1(A[4]), .A2(net123752), .ZN(net119928) );
  INV_X1 U1744 ( .A(net81424), .ZN(net123752) );
  INV_X8 U1745 ( .A(A[4]), .ZN(net77956) );
  INV_X16 U1746 ( .A(A[4]), .ZN(net119855) );
  NAND3_X4 U1747 ( .A1(net80847), .A2(net80848), .A3(n493), .ZN(
        \CARRYB[8][12] ) );
  NAND2_X1 U1748 ( .A1(\ab[8][12] ), .A2(\CARRYB[7][12] ), .ZN(n493) );
  NAND2_X2 U1749 ( .A1(\SUMB[7][13] ), .A2(\CARRYB[7][12] ), .ZN(net80848) );
  NAND2_X2 U1750 ( .A1(\ab[8][12] ), .A2(net90348), .ZN(net80847) );
  NOR2_X2 U1751 ( .A1(net83784), .A2(net77926), .ZN(\ab[8][12] ) );
  INV_X1 U1752 ( .A(\ab[8][12] ), .ZN(net87308) );
  INV_X4 U1753 ( .A(n491), .ZN(net83784) );
  INV_X8 U1754 ( .A(B[12]), .ZN(net70458) );
  NOR2_X4 U1755 ( .A1(net82247), .A2(net70458), .ZN(\ab[0][12] ) );
  NAND3_X4 U1756 ( .A1(n494), .A2(n496), .A3(n495), .ZN(\CARRYB[7][12] ) );
  INV_X4 U1757 ( .A(\CARRYB[7][12] ), .ZN(net87309) );
  NAND2_X4 U1758 ( .A1(\SUMB[6][13] ), .A2(\ab[7][12] ), .ZN(n495) );
  NAND2_X4 U1759 ( .A1(net124104), .A2(n492), .ZN(n496) );
  INV_X2 U1760 ( .A(n497), .ZN(n492) );
  INV_X8 U1761 ( .A(\CARRYB[6][12] ), .ZN(n497) );
  NAND2_X4 U1762 ( .A1(n497), .A2(net85251), .ZN(net85254) );
  XNOR2_X2 U1763 ( .A(net90897), .B(net81756), .ZN(\SUMB[7][13] ) );
  XNOR2_X2 U1764 ( .A(\SUMB[7][13] ), .B(net85212), .ZN(net91118) );
  NAND2_X4 U1765 ( .A1(n499), .A2(n498), .ZN(\SUMB[25][2] ) );
  INV_X4 U1766 ( .A(net92568), .ZN(net92569) );
  NAND3_X4 U1768 ( .A1(net80257), .A2(n500), .A3(net80258), .ZN(
        \CARRYB[24][2] ) );
  NAND2_X4 U1769 ( .A1(net86520), .A2(\CARRYB[23][2] ), .ZN(n500) );
  INV_X8 U1770 ( .A(net86519), .ZN(net86520) );
  NAND2_X4 U1771 ( .A1(net86520), .A2(\ab[24][2] ), .ZN(net80257) );
  NAND3_X2 U1773 ( .A1(n503), .A2(n501), .A3(n502), .ZN(\CARRYB[22][3] ) );
  NAND3_X2 U1775 ( .A1(net80511), .A2(net80510), .A3(net80509), .ZN(
        \CARRYB[21][3] ) );
  NAND2_X2 U1776 ( .A1(\ab[22][3] ), .A2(\SUMB[21][4] ), .ZN(n501) );
  BUF_X32 U1777 ( .A(net77882), .Z(net77886) );
  INV_X8 U1778 ( .A(B[3]), .ZN(net77882) );
  NAND2_X4 U1779 ( .A1(net89840), .A2(net87043), .ZN(net84874) );
  NAND2_X4 U1780 ( .A1(net84874), .A2(net84873), .ZN(net83848) );
  AND2_X2 U1781 ( .A1(net84874), .A2(\CARRYB[12][9] ), .ZN(net85044) );
  INV_X4 U1782 ( .A(net88302), .ZN(net87043) );
  INV_X8 U1783 ( .A(net89447), .ZN(\SUMB[11][11] ) );
  NAND2_X4 U1784 ( .A1(\ab[12][10] ), .A2(\SUMB[11][11] ), .ZN(net81057) );
  NAND2_X2 U1785 ( .A1(\CARRYB[11][10] ), .A2(\SUMB[11][11] ), .ZN(net81058)
         );
  NAND2_X2 U1786 ( .A1(net88302), .A2(\SUMB[11][11] ), .ZN(net84873) );
  INV_X4 U1787 ( .A(net81165), .ZN(n505) );
  INV_X4 U1788 ( .A(net89167), .ZN(n504) );
  NAND2_X2 U1789 ( .A1(net81165), .A2(net89167), .ZN(n506) );
  NAND2_X4 U1790 ( .A1(net92552), .A2(net92553), .ZN(net88302) );
  INV_X4 U1791 ( .A(net88303), .ZN(net92551) );
  INV_X1 U1792 ( .A(\ab[12][10] ), .ZN(net88303) );
  INV_X4 U1793 ( .A(net89369), .ZN(net92550) );
  NAND3_X2 U1794 ( .A1(net83880), .A2(net83882), .A3(net83881), .ZN(net89369)
         );
  NAND2_X4 U1795 ( .A1(net85539), .A2(n509), .ZN(net81165) );
  NAND2_X2 U1796 ( .A1(net88525), .A2(net85537), .ZN(n509) );
  INV_X1 U1797 ( .A(\ab[11][11] ), .ZN(net85537) );
  NAND2_X4 U1798 ( .A1(n508), .A2(\ab[11][11] ), .ZN(net85539) );
  INV_X4 U1799 ( .A(\CARRYB[10][11] ), .ZN(n508) );
  INV_X1 U1800 ( .A(n508), .ZN(net87490) );
  NAND3_X2 U1801 ( .A1(net80957), .A2(net80956), .A3(net80958), .ZN(
        \CARRYB[10][11] ) );
  XNOR2_X2 U1802 ( .A(net89065), .B(net80983), .ZN(net89167) );
  NAND2_X1 U1803 ( .A1(\ab[12][10] ), .A2(\CARRYB[11][10] ), .ZN(net81056) );
  NAND2_X2 U1804 ( .A1(net92622), .A2(net83848), .ZN(net82294) );
  NAND2_X4 U1805 ( .A1(\SUMB[12][10] ), .A2(net82292), .ZN(net82295) );
  INV_X4 U1806 ( .A(net92622), .ZN(net82292) );
  INV_X4 U1807 ( .A(net83848), .ZN(\SUMB[12][10] ) );
  NAND2_X2 U1808 ( .A1(\SUMB[12][10] ), .A2(\ab[13][9] ), .ZN(net81060) );
  NAND2_X4 U1809 ( .A1(net86145), .A2(net86144), .ZN(net92622) );
  NAND2_X4 U1810 ( .A1(\CARRYB[12][9] ), .A2(net81182), .ZN(net86144) );
  INV_X1 U1811 ( .A(\ab[13][9] ), .ZN(net81182) );
  INV_X4 U1812 ( .A(net81182), .ZN(net86142) );
  NAND2_X4 U1813 ( .A1(n510), .A2(net86142), .ZN(net86145) );
  NAND2_X1 U1814 ( .A1(\ab[13][9] ), .A2(\CARRYB[12][9] ), .ZN(net81059) );
  NAND3_X2 U1815 ( .A1(net88295), .A2(net88296), .A3(net88297), .ZN(
        \CARRYB[12][9] ) );
  CLKBUF_X3 U1816 ( .A(net84873), .Z(net88455) );
  NAND2_X4 U1817 ( .A1(net124589), .A2(net86806), .ZN(net82404) );
  NAND3_X4 U1818 ( .A1(net82404), .A2(net82403), .A3(net82405), .ZN(
        \CARRYB[20][5] ) );
  NAND2_X4 U1819 ( .A1(net86806), .A2(\ab[20][5] ), .ZN(net82403) );
  INV_X8 U1820 ( .A(net91377), .ZN(net120625) );
  XNOR2_X2 U1821 ( .A(net90810), .B(net90576), .ZN(net124589) );
  NAND2_X2 U1822 ( .A1(net83202), .A2(net124589), .ZN(net147930) );
  INV_X2 U1823 ( .A(net124589), .ZN(net147929) );
  XNOR2_X2 U1824 ( .A(net90810), .B(net90576), .ZN(\SUMB[19][6] ) );
  NAND3_X4 U1825 ( .A1(n512), .A2(n511), .A3(net84708), .ZN(net91377) );
  NAND2_X2 U1826 ( .A1(net91377), .A2(\ab[20][5] ), .ZN(net120627) );
  NAND2_X4 U1827 ( .A1(\SUMB[18][6] ), .A2(\ab[19][5] ), .ZN(n511) );
  XNOR2_X2 U1828 ( .A(n8), .B(net92542), .ZN(\SUMB[19][5] ) );
  XNOR2_X2 U1829 ( .A(\SUMB[18][6] ), .B(net92542), .ZN(net88887) );
  NAND2_X4 U1830 ( .A1(\SUMB[18][6] ), .A2(net148582), .ZN(n512) );
  XNOR2_X2 U1831 ( .A(net81264), .B(\SUMB[17][7] ), .ZN(net88878) );
  XNOR2_X2 U1832 ( .A(net85611), .B(net82748), .ZN(net81264) );
  INV_X4 U1833 ( .A(net85610), .ZN(net85611) );
  INV_X4 U1834 ( .A(\SUMB[17][6] ), .ZN(net86661) );
  NAND2_X4 U1835 ( .A1(\SUMB[27][1] ), .A2(\CARRYB[27][0] ), .ZN(net80773) );
  NAND3_X4 U1836 ( .A1(net80773), .A2(n513), .A3(net80771), .ZN(
        \CARRYB[28][0] ) );
  NAND3_X4 U1837 ( .A1(net80768), .A2(net80769), .A3(net80767), .ZN(
        \CARRYB[27][0] ) );
  NAND2_X4 U1838 ( .A1(\CARRYB[27][0] ), .A2(n345), .ZN(n513) );
  NAND2_X4 U1839 ( .A1(\SUMB[27][1] ), .A2(n345), .ZN(net80771) );
  XNOR2_X2 U1840 ( .A(\SUMB[27][1] ), .B(n345), .ZN(net92378) );
  NOR2_X2 U1841 ( .A1(net91660), .A2(net70471), .ZN(\ab[12][10] ) );
  NAND2_X2 U1842 ( .A1(net121898), .A2(\SUMB[10][11] ), .ZN(net83880) );
  NAND3_X2 U1843 ( .A1(net83880), .A2(net83881), .A3(net83882), .ZN(
        \CARRYB[11][10] ) );
  INV_X1 U1844 ( .A(n201), .ZN(net121898) );
  NAND2_X2 U1845 ( .A1(n201), .A2(net87045), .ZN(net92863) );
  NAND2_X2 U1846 ( .A1(\SUMB[10][11] ), .A2(\ab[11][10] ), .ZN(net83881) );
  NAND2_X1 U1847 ( .A1(\ab[11][10] ), .A2(\CARRYB[10][10] ), .ZN(net83882) );
  INV_X2 U1848 ( .A(\SUMB[10][11] ), .ZN(net85373) );
  NAND2_X1 U1849 ( .A1(\CARRYB[10][10] ), .A2(\ab[11][10] ), .ZN(net92862) );
  INV_X32 U1850 ( .A(net77864), .ZN(net77860) );
  INV_X4 U1851 ( .A(B[0]), .ZN(net70436) );
  NAND2_X1 U1852 ( .A1(A[28]), .A2(B[3]), .ZN(net92320) );
  NAND2_X1 U1853 ( .A1(B[0]), .A2(net80392), .ZN(net70435) );
  NAND2_X4 U1854 ( .A1(net87365), .A2(net87364), .ZN(net87367) );
  NAND2_X4 U1855 ( .A1(net87367), .A2(net87366), .ZN(\SUMB[10][11] ) );
  NAND2_X2 U1856 ( .A1(net87366), .A2(net87367), .ZN(net91243) );
  INV_X4 U1857 ( .A(net82838), .ZN(net87365) );
  NAND2_X4 U1858 ( .A1(net84672), .A2(net84671), .ZN(net91003) );
  NAND2_X4 U1859 ( .A1(net82838), .A2(net91003), .ZN(net87366) );
  NAND2_X4 U1860 ( .A1(n516), .A2(n515), .ZN(net82838) );
  NAND2_X4 U1861 ( .A1(n514), .A2(net83876), .ZN(n516) );
  INV_X4 U1862 ( .A(\CARRYB[9][11] ), .ZN(n514) );
  NAND2_X2 U1863 ( .A1(\CARRYB[9][11] ), .A2(\ab[10][11] ), .ZN(n515) );
  NAND2_X1 U1864 ( .A1(\ab[10][11] ), .A2(\CARRYB[9][11] ), .ZN(net80958) );
  NAND2_X4 U1865 ( .A1(net84669), .A2(net84670), .ZN(net84672) );
  INV_X4 U1866 ( .A(n2360), .ZN(net84670) );
  INV_X4 U1867 ( .A(net84670), .ZN(net88841) );
  INV_X4 U1868 ( .A(net82837), .ZN(net84669) );
  NAND2_X4 U1870 ( .A1(net85459), .A2(net85460), .ZN(n517) );
  INV_X4 U1871 ( .A(net81958), .ZN(net85459) );
  NAND2_X2 U1872 ( .A1(net89356), .A2(net81958), .ZN(net85461) );
  NAND2_X4 U1873 ( .A1(net84870), .A2(net81373), .ZN(net82837) );
  NAND2_X4 U1874 ( .A1(net88841), .A2(net82837), .ZN(net84671) );
  INV_X1 U1875 ( .A(\ab[9][12] ), .ZN(net84867) );
  INV_X2 U1876 ( .A(net84868), .ZN(net89149) );
  NAND2_X4 U1877 ( .A1(\SUMB[7][14] ), .A2(\ab[8][13] ), .ZN(net81371) );
  NAND2_X4 U1878 ( .A1(net89356), .A2(net88943), .ZN(net81372) );
  NAND3_X2 U1879 ( .A1(net81374), .A2(net81375), .A3(net81373), .ZN(
        \CARRYB[9][12] ) );
  NAND2_X2 U1880 ( .A1(\SUMB[19][6] ), .A2(\ab[20][5] ), .ZN(net82405) );
  NOR2_X4 U1881 ( .A1(net77900), .A2(net70455), .ZN(\ab[20][5] ) );
  INV_X1 U1882 ( .A(\ab[20][5] ), .ZN(net120626) );
  INV_X16 U1883 ( .A(A[20]), .ZN(net70455) );
  INV_X8 U1884 ( .A(B[5]), .ZN(net70444) );
  NAND2_X4 U1885 ( .A1(n518), .A2(n519), .ZN(net90810) );
  NAND3_X2 U1886 ( .A1(net81270), .A2(net81269), .A3(net81268), .ZN(net93914)
         );
  NOR2_X4 U1887 ( .A1(net77908), .A2(net70457), .ZN(\ab[19][6] ) );
  NAND2_X2 U1888 ( .A1(\ab[19][6] ), .A2(net124627), .ZN(net81067) );
  NAND2_X4 U1889 ( .A1(\SUMB[18][7] ), .A2(\ab[19][6] ), .ZN(net81068) );
  INV_X16 U1890 ( .A(A[19]), .ZN(net70457) );
  INV_X4 U1891 ( .A(B[6]), .ZN(net77908) );
  NAND2_X2 U1892 ( .A1(\SUMB[17][7] ), .A2(net85611), .ZN(net81270) );
  NAND3_X2 U1893 ( .A1(net81270), .A2(net81269), .A3(net81268), .ZN(net124627)
         );
  NAND2_X2 U1894 ( .A1(\ab[18][6] ), .A2(net85611), .ZN(net81268) );
  NAND2_X4 U1895 ( .A1(net82286), .A2(n520), .ZN(\*UDW_*112684/net78549 ) );
  NAND2_X4 U1896 ( .A1(net85688), .A2(\ab[1][17] ), .ZN(
        \*UDW_*112684/net78547 ) );
  NOR2_X4 U1897 ( .A1(net70470), .A2(net82149), .ZN(net85688) );
  NAND2_X2 U1898 ( .A1(net86959), .A2(net87050), .ZN(n520) );
  INV_X16 U1899 ( .A(B[17]), .ZN(net123000) );
  NOR2_X2 U1900 ( .A1(net83784), .A2(net70477), .ZN(\ab[9][12] ) );
  XNOR2_X2 U1901 ( .A(net90348), .B(net85212), .ZN(net90687) );
  NAND2_X2 U1902 ( .A1(A[29]), .A2(B[2]), .ZN(net92341) );
  NAND2_X2 U1903 ( .A1(\CARRYB[25][1] ), .A2(\SUMB[25][2] ), .ZN(net83975) );
  XNOR2_X2 U1904 ( .A(\SUMB[25][2] ), .B(\ab[26][1] ), .ZN(net86427) );
  NAND2_X4 U1905 ( .A1(net92790), .A2(net93840), .ZN(net80261) );
  INV_X16 U1906 ( .A(A[17]), .ZN(net70461) );
  NAND3_X2 U1907 ( .A1(net80541), .A2(net80540), .A3(n521), .ZN(
        \CARRYB[16][6] ) );
  NAND2_X2 U1908 ( .A1(net90347), .A2(\ab[16][6] ), .ZN(n521) );
  NAND2_X2 U1909 ( .A1(\SUMB[15][7] ), .A2(\ab[16][6] ), .ZN(net80540) );
  NAND2_X2 U1910 ( .A1(\SUMB[15][7] ), .A2(net90347), .ZN(net80541) );
  XNOR2_X2 U1911 ( .A(n522), .B(\SUMB[16][8] ), .ZN(\SUMB[17][7] ) );
  NAND2_X2 U1912 ( .A1(\SUMB[17][7] ), .A2(\ab[18][6] ), .ZN(net81269) );
  XNOR2_X2 U1913 ( .A(\CARRYB[16][7] ), .B(\ab[17][7] ), .ZN(n522) );
  NAND3_X4 U1914 ( .A1(n523), .A2(n524), .A3(n525), .ZN(\CARRYB[25][1] ) );
  INV_X1 U1915 ( .A(\CARRYB[25][1] ), .ZN(net88655) );
  NAND2_X4 U1916 ( .A1(\CARRYB[24][1] ), .A2(\ab[25][1] ), .ZN(n525) );
  NAND2_X4 U1917 ( .A1(\CARRYB[24][1] ), .A2(\SUMB[24][2] ), .ZN(n523) );
  NAND2_X4 U1918 ( .A1(\SUMB[24][2] ), .A2(\ab[25][1] ), .ZN(n524) );
  XNOR2_X2 U1919 ( .A(\CARRYB[24][1] ), .B(\ab[25][1] ), .ZN(net124874) );
  XNOR2_X2 U1920 ( .A(net90897), .B(net81756), .ZN(net90348) );
  INV_X8 U1921 ( .A(net88660), .ZN(net90897) );
  NAND2_X4 U1922 ( .A1(net90897), .A2(net88444), .ZN(net80845) );
  NAND2_X4 U1923 ( .A1(net90897), .A2(\ab[7][13] ), .ZN(net80844) );
  INV_X4 U1924 ( .A(\SUMB[6][14] ), .ZN(net88660) );
  INV_X2 U1925 ( .A(\CARRYB[6][14] ), .ZN(net88880) );
  NAND2_X2 U1926 ( .A1(net83919), .A2(\CARRYB[4][14] ), .ZN(net82297) );
  NOR2_X1 U1927 ( .A1(net84698), .A2(net77940), .ZN(\ab[6][14] ) );
  NAND2_X4 U1928 ( .A1(net84445), .A2(net84446), .ZN(\SUMB[5][15] ) );
  INV_X8 U1929 ( .A(net84856), .ZN(\SUMB[4][16] ) );
  NAND2_X2 U1930 ( .A1(\SUMB[4][16] ), .A2(\ab[5][15] ), .ZN(net80839) );
  NAND2_X2 U1931 ( .A1(\SUMB[4][16] ), .A2(n137), .ZN(net80840) );
  NAND2_X4 U1932 ( .A1(n527), .A2(net148053), .ZN(net84856) );
  NAND2_X4 U1933 ( .A1(net148051), .A2(n526), .ZN(n527) );
  INV_X4 U1934 ( .A(net124367), .ZN(n526) );
  NOR2_X4 U1935 ( .A1(net77900), .A2(net70453), .ZN(\ab[21][5] ) );
  INV_X16 U1936 ( .A(A[21]), .ZN(net70453) );
  NAND2_X4 U1937 ( .A1(net88856), .A2(\SUMB[18][7] ), .ZN(net81069) );
  XNOR2_X2 U1938 ( .A(net83536), .B(net86055), .ZN(PRODUCT[30]) );
  NOR2_X1 U1939 ( .A1(net36614), .A2(net77858), .ZN(\ab[30][0] ) );
  INV_X4 U1940 ( .A(A[30]), .ZN(net36614) );
  NOR2_X1 U1941 ( .A1(net36614), .A2(net77866), .ZN(net81548) );
  NAND3_X4 U1942 ( .A1(n529), .A2(n528), .A3(net92718), .ZN(\CARRYB[4][14] )
         );
  NAND2_X4 U1943 ( .A1(net119817), .A2(\ab[4][14] ), .ZN(n528) );
  INV_X4 U1944 ( .A(A[27]), .ZN(net70441) );
  XNOR2_X2 U1945 ( .A(n531), .B(n200), .ZN(net86055) );
  NAND2_X4 U1946 ( .A1(n535), .A2(n534), .ZN(\SUMB[28][2] ) );
  XNOR2_X2 U1947 ( .A(net81158), .B(n4), .ZN(net89453) );
  NAND2_X2 U1948 ( .A1(\SUMB[28][2] ), .A2(\ab[29][1] ), .ZN(net80667) );
  NAND2_X4 U1949 ( .A1(n533), .A2(n530), .ZN(n535) );
  INV_X4 U1950 ( .A(n402), .ZN(n530) );
  NAND2_X4 U1951 ( .A1(net85094), .A2(net92337), .ZN(n532) );
  INV_X4 U1952 ( .A(net92337), .ZN(\ab[29][1] ) );
  NAND2_X4 U1953 ( .A1(\CARRYB[28][1] ), .A2(\ab[29][1] ), .ZN(net85096) );
  NAND2_X2 U1954 ( .A1(\CARRYB[1][16] ), .A2(\ab[2][16] ), .ZN(net119899) );
  INV_X8 U1955 ( .A(\*UDW_*112689/net78561 ), .ZN(\CARRYB[1][16] ) );
  NOR2_X4 U1956 ( .A1(\ab[2][16] ), .A2(\CARRYB[1][16] ), .ZN(net119901) );
  NAND2_X4 U1957 ( .A1(\ab[0][17] ), .A2(net88123), .ZN(
        \*UDW_*112689/net78561 ) );
  NAND2_X2 U1958 ( .A1(net149526), .A2(net88123), .ZN(net123430) );
  NAND2_X4 U1959 ( .A1(n540), .A2(n539), .ZN(net84327) );
  INV_X8 U1960 ( .A(n536), .ZN(\SUMB[1][18] ) );
  NAND2_X4 U1961 ( .A1(\SUMB[1][18] ), .A2(\ab[2][17] ), .ZN(net82027) );
  INV_X4 U1962 ( .A(net82024), .ZN(n537) );
  NOR2_X1 U1963 ( .A1(net77886), .A2(net70447), .ZN(\ab[24][3] ) );
  INV_X4 U1964 ( .A(A[24]), .ZN(net70447) );
  XNOR2_X2 U1965 ( .A(\SUMB[21][4] ), .B(\ab[22][3] ), .ZN(net81493) );
  NAND3_X2 U1966 ( .A1(net80509), .A2(net80511), .A3(net80510), .ZN(net124949)
         );
  NOR2_X4 U1967 ( .A1(net77886), .A2(net70451), .ZN(\ab[22][3] ) );
  NAND2_X4 U1968 ( .A1(n542), .A2(\SUMB[20][4] ), .ZN(net80511) );
  INV_X4 U1969 ( .A(\CARRYB[20][3] ), .ZN(n541) );
  NAND2_X1 U1970 ( .A1(net83172), .A2(n541), .ZN(net83175) );
  NAND2_X4 U1971 ( .A1(n546), .A2(n545), .ZN(\SUMB[20][6] ) );
  NAND2_X2 U1972 ( .A1(net84348), .A2(n547), .ZN(n545) );
  NAND2_X4 U1974 ( .A1(n543), .A2(n544), .ZN(n546) );
  INV_X4 U1975 ( .A(net84348), .ZN(n543) );
  INV_X4 U1976 ( .A(n552), .ZN(\SUMB[17][8] ) );
  NAND2_X4 U1977 ( .A1(\SUMB[17][8] ), .A2(net87619), .ZN(net81066) );
  NAND2_X4 U1978 ( .A1(\SUMB[17][8] ), .A2(\ab[18][7] ), .ZN(net81065) );
  XNOR2_X2 U1979 ( .A(n548), .B(\SUMB[16][9] ), .ZN(n552) );
  NAND2_X4 U1980 ( .A1(n551), .A2(net84374), .ZN(n548) );
  NAND2_X4 U1981 ( .A1(n550), .A2(\ab[17][8] ), .ZN(net84374) );
  INV_X8 U1982 ( .A(\CARRYB[16][8] ), .ZN(n550) );
  INV_X1 U1983 ( .A(n550), .ZN(net93410) );
  NAND2_X2 U1984 ( .A1(net83776), .A2(\CARRYB[16][8] ), .ZN(n551) );
  XNOR2_X2 U1985 ( .A(net87619), .B(\ab[18][7] ), .ZN(n549) );
  INV_X4 U1986 ( .A(net148015), .ZN(net148302) );
  INV_X4 U1987 ( .A(net85096), .ZN(net149916) );
  INV_X4 U1988 ( .A(net149916), .ZN(net149917) );
  NAND2_X2 U1989 ( .A1(n1699), .A2(n1698), .ZN(n1701) );
  NAND2_X2 U1990 ( .A1(\ab[20][2] ), .A2(\SUMB[19][3] ), .ZN(n1914) );
  INV_X4 U1991 ( .A(n554), .ZN(n555) );
  INV_X4 U1992 ( .A(\SUMB[9][16] ), .ZN(n1220) );
  XNOR2_X2 U1993 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .ZN(n557) );
  INV_X8 U1994 ( .A(\*UDW_*112704/net78605 ), .ZN(\SUMB[1][13] ) );
  NAND2_X2 U1996 ( .A1(net88407), .A2(net88408), .ZN(net88410) );
  NOR2_X2 U1997 ( .A1(net84698), .A2(net77926), .ZN(\ab[8][14] ) );
  NAND3_X4 U1998 ( .A1(n2048), .A2(n2049), .A3(n2050), .ZN(\CARRYB[9][15] ) );
  NAND2_X2 U1999 ( .A1(\CARRYB[8][15] ), .A2(n151), .ZN(n2048) );
  NAND2_X4 U2000 ( .A1(n1709), .A2(n1710), .ZN(n2031) );
  NAND2_X2 U2001 ( .A1(n886), .A2(n887), .ZN(n558) );
  INV_X4 U2003 ( .A(net149605), .ZN(net92405) );
  XNOR2_X2 U2004 ( .A(n559), .B(n560), .ZN(\SUMB[17][3] ) );
  XNOR2_X2 U2005 ( .A(\SUMB[7][7] ), .B(n561), .ZN(\SUMB[8][6] ) );
  INV_X1 U2006 ( .A(n1041), .ZN(n562) );
  NAND2_X2 U2007 ( .A1(\CARRYB[3][16] ), .A2(n803), .ZN(n656) );
  INV_X4 U2008 ( .A(\SUMB[10][5] ), .ZN(n592) );
  NAND2_X2 U2009 ( .A1(\ab[12][0] ), .A2(\SUMB[11][1] ), .ZN(n1144) );
  NAND2_X2 U2010 ( .A1(\SUMB[11][1] ), .A2(\CARRYB[11][0] ), .ZN(n1146) );
  XOR2_X2 U2011 ( .A(n1315), .B(n730), .Z(\SUMB[11][1] ) );
  CLKBUF_X3 U2012 ( .A(\SUMB[22][3] ), .Z(n564) );
  XNOR2_X2 U2013 ( .A(net81995), .B(n833), .ZN(n565) );
  NOR2_X2 U2014 ( .A1(net70456), .A2(net119855), .ZN(\ab[4][11] ) );
  NAND2_X2 U2015 ( .A1(n979), .A2(n980), .ZN(net86557) );
  OR2_X2 U2016 ( .A1(n1037), .A2(n1038), .ZN(n1302) );
  NAND3_X4 U2017 ( .A1(n1861), .A2(n1862), .A3(n1863), .ZN(\CARRYB[8][7] ) );
  NAND2_X2 U2018 ( .A1(\ab[8][7] ), .A2(\CARRYB[7][7] ), .ZN(n1863) );
  XNOR2_X2 U2019 ( .A(n1204), .B(\SUMB[19][11] ), .ZN(n568) );
  XNOR2_X2 U2020 ( .A(\CARRYB[17][4] ), .B(\ab[18][4] ), .ZN(n569) );
  INV_X4 U2021 ( .A(n1593), .ZN(n570) );
  INV_X4 U2022 ( .A(n37), .ZN(n1593) );
  NAND2_X4 U2023 ( .A1(\SUMB[19][5] ), .A2(\CARRYB[19][4] ), .ZN(n2230) );
  NAND2_X2 U2024 ( .A1(n1004), .A2(n1683), .ZN(n1685) );
  BUF_X8 U2025 ( .A(\SUMB[15][3] ), .Z(n571) );
  XNOR2_X2 U2026 ( .A(n1339), .B(n1229), .ZN(n572) );
  XOR2_X2 U2027 ( .A(\SUMB[8][19] ), .B(net79950), .Z(n573) );
  XNOR2_X2 U2028 ( .A(n574), .B(\SUMB[14][3] ), .ZN(\SUMB[15][2] ) );
  NAND2_X2 U2029 ( .A1(net92863), .A2(net92862), .ZN(n1617) );
  NAND2_X2 U2030 ( .A1(n1154), .A2(\CARRYB[1][10] ), .ZN(n1156) );
  NAND2_X1 U2031 ( .A1(\ab[9][8] ), .A2(\CARRYB[8][8] ), .ZN(n2086) );
  XOR2_X2 U2032 ( .A(n1207), .B(\ab[3][12] ), .Z(n575) );
  NOR2_X4 U2033 ( .A1(net83784), .A2(net77964), .ZN(\ab[3][12] ) );
  INV_X8 U2034 ( .A(net80392), .ZN(net124610) );
  INV_X2 U2035 ( .A(\SUMB[11][15] ), .ZN(n700) );
  NAND2_X4 U2036 ( .A1(n1366), .A2(n1708), .ZN(n1710) );
  NAND2_X4 U2037 ( .A1(\ab[2][11] ), .A2(\CARRYB[1][11] ), .ZN(n1642) );
  XNOR2_X2 U2038 ( .A(net81782), .B(n825), .ZN(n576) );
  INV_X4 U2039 ( .A(n576), .ZN(\SUMB[18][9] ) );
  INV_X8 U2040 ( .A(\SUMB[18][9] ), .ZN(n641) );
  NAND2_X4 U2041 ( .A1(\SUMB[5][14] ), .A2(\ab[6][13] ), .ZN(n2069) );
  NAND2_X2 U2042 ( .A1(\CARRYB[5][12] ), .A2(\ab[6][12] ), .ZN(n1417) );
  NAND2_X4 U2043 ( .A1(\SUMB[7][8] ), .A2(\ab[8][7] ), .ZN(n1862) );
  NAND2_X2 U2044 ( .A1(net83030), .A2(net81663), .ZN(n579) );
  NAND2_X4 U2045 ( .A1(n577), .A2(n578), .ZN(n580) );
  NAND2_X4 U2046 ( .A1(n579), .A2(n580), .ZN(net86884) );
  NAND2_X1 U2047 ( .A1(net80927), .A2(net89104), .ZN(n583) );
  INV_X2 U2048 ( .A(net80927), .ZN(n581) );
  NAND2_X4 U2049 ( .A1(n585), .A2(n586), .ZN(n587) );
  INV_X8 U2050 ( .A(n2334), .ZN(\CARRYB[1][11] ) );
  NAND2_X4 U2051 ( .A1(net80021), .A2(\SUMB[23][5] ), .ZN(net86023) );
  INV_X4 U2052 ( .A(n1118), .ZN(n955) );
  OR2_X4 U2053 ( .A1(n830), .A2(n831), .ZN(n827) );
  INV_X2 U2054 ( .A(net148233), .ZN(net148754) );
  NAND2_X1 U2055 ( .A1(\ab[15][12] ), .A2(\CARRYB[14][12] ), .ZN(n2200) );
  INV_X4 U2056 ( .A(n1044), .ZN(n588) );
  INV_X4 U2057 ( .A(n2337), .ZN(\SUMB[1][12] ) );
  CLKBUF_X3 U2058 ( .A(\SUMB[11][8] ), .Z(n1248) );
  NAND2_X2 U2059 ( .A1(n1551), .A2(n948), .ZN(n590) );
  NAND2_X4 U2060 ( .A1(n589), .A2(n947), .ZN(n591) );
  NAND2_X4 U2061 ( .A1(n590), .A2(n591), .ZN(\SUMB[4][8] ) );
  INV_X4 U2062 ( .A(n1551), .ZN(n589) );
  NAND2_X1 U2063 ( .A1(n563), .A2(n1276), .ZN(n594) );
  NAND2_X2 U2064 ( .A1(n592), .A2(n593), .ZN(n595) );
  INV_X4 U2065 ( .A(n1276), .ZN(n593) );
  INV_X4 U2066 ( .A(n947), .ZN(n948) );
  BUF_X4 U2067 ( .A(\SUMB[4][8] ), .Z(n1389) );
  XNOR2_X2 U2068 ( .A(\SUMB[11][4] ), .B(\ab[12][3] ), .ZN(n985) );
  NAND3_X2 U2069 ( .A1(n1914), .A2(n1916), .A3(n1915), .ZN(n596) );
  NAND2_X2 U2070 ( .A1(n1731), .A2(n1265), .ZN(n600) );
  NAND2_X4 U2071 ( .A1(n598), .A2(n599), .ZN(n601) );
  NAND2_X4 U2072 ( .A1(n600), .A2(n601), .ZN(\SUMB[16][4] ) );
  INV_X4 U2073 ( .A(n1731), .ZN(n598) );
  INV_X4 U2074 ( .A(n1265), .ZN(n599) );
  BUF_X8 U2075 ( .A(\SUMB[15][5] ), .Z(n1265) );
  NAND2_X4 U2076 ( .A1(\CARRYB[19][0] ), .A2(\ab[20][0] ), .ZN(n2100) );
  NAND2_X2 U2077 ( .A1(\CARRYB[10][0] ), .A2(\SUMB[10][1] ), .ZN(n1142) );
  NAND3_X4 U2078 ( .A1(n1471), .A2(n1472), .A3(n1473), .ZN(\CARRYB[10][1] ) );
  XNOR2_X2 U2079 ( .A(n350), .B(\ab[2][6] ), .ZN(n758) );
  INV_X1 U2080 ( .A(\ab[8][14] ), .ZN(n603) );
  NAND2_X4 U2081 ( .A1(n606), .A2(n607), .ZN(n609) );
  NAND2_X4 U2082 ( .A1(n609), .A2(n608), .ZN(PRODUCT[31]) );
  NAND2_X2 U2083 ( .A1(\CARRYB[18][8] ), .A2(\ab[19][8] ), .ZN(net123293) );
  BUF_X8 U2084 ( .A(\CARRYB[16][9] ), .Z(net89819) );
  BUF_X8 U2085 ( .A(\SUMB[13][6] ), .Z(n1202) );
  INV_X2 U2087 ( .A(net84707), .ZN(net148582) );
  NAND2_X1 U2088 ( .A1(\ab[25][5] ), .A2(\SUMB[24][6] ), .ZN(net79867) );
  INV_X4 U2089 ( .A(\SUMB[13][14] ), .ZN(net86629) );
  XNOR2_X2 U2090 ( .A(n610), .B(net87962), .ZN(\SUMB[3][6] ) );
  XNOR2_X2 U2091 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .ZN(n610) );
  XOR2_X2 U2092 ( .A(n1470), .B(net124757), .Z(\SUMB[10][1] ) );
  NAND2_X2 U2094 ( .A1(n1589), .A2(n1456), .ZN(n1591) );
  NAND3_X1 U2095 ( .A1(net86170), .A2(net86171), .A3(net86172), .ZN(n1186) );
  XNOR2_X1 U2096 ( .A(n1268), .B(n1241), .ZN(n868) );
  NAND2_X4 U2097 ( .A1(\CARRYB[17][3] ), .A2(\ab[18][3] ), .ZN(n1416) );
  NAND3_X2 U2098 ( .A1(n2236), .A2(n2235), .A3(n2234), .ZN(\CARRYB[19][4] ) );
  NAND2_X2 U2099 ( .A1(\SUMB[18][9] ), .A2(net88700), .ZN(n623) );
  NAND2_X2 U2100 ( .A1(net93203), .A2(n1901), .ZN(n1128) );
  NAND2_X4 U2101 ( .A1(net120655), .A2(net120656), .ZN(n804) );
  INV_X4 U2102 ( .A(n2197), .ZN(n1788) );
  NAND2_X2 U2103 ( .A1(\ab[16][12] ), .A2(\SUMB[15][13] ), .ZN(n1086) );
  NAND3_X2 U2104 ( .A1(n2206), .A2(n2207), .A3(n2205), .ZN(\CARRYB[6][16] ) );
  XOR2_X2 U2105 ( .A(\CARRYB[14][15] ), .B(\ab[15][15] ), .Z(n611) );
  XOR2_X2 U2106 ( .A(n1252), .B(n611), .Z(\SUMB[15][15] ) );
  NAND2_X1 U2107 ( .A1(\CARRYB[14][15] ), .A2(n1252), .ZN(n612) );
  NAND2_X1 U2108 ( .A1(\ab[15][15] ), .A2(n1252), .ZN(n613) );
  NAND2_X1 U2109 ( .A1(\ab[15][15] ), .A2(\CARRYB[14][15] ), .ZN(n614) );
  NAND3_X2 U2110 ( .A1(n612), .A2(n613), .A3(n614), .ZN(\CARRYB[15][15] ) );
  NAND2_X2 U2111 ( .A1(\SUMB[13][17] ), .A2(n2188), .ZN(n617) );
  NAND2_X4 U2112 ( .A1(n617), .A2(n618), .ZN(n1252) );
  INV_X2 U2113 ( .A(\SUMB[13][17] ), .ZN(n615) );
  INV_X2 U2114 ( .A(n2188), .ZN(n616) );
  NAND3_X4 U2115 ( .A1(n1870), .A2(n1871), .A3(n1872), .ZN(\CARRYB[14][15] )
         );
  NAND3_X4 U2116 ( .A1(n1071), .A2(net80267), .A3(net80268), .ZN(
        \CARRYB[22][7] ) );
  INV_X8 U2117 ( .A(\CARRYB[4][16] ), .ZN(n638) );
  NAND2_X4 U2118 ( .A1(\SUMB[7][9] ), .A2(\ab[8][8] ), .ZN(n2005) );
  NAND2_X2 U2119 ( .A1(\CARRYB[8][15] ), .A2(\ab[9][15] ), .ZN(n1709) );
  INV_X4 U2120 ( .A(\CARRYB[8][15] ), .ZN(n1366) );
  NAND2_X4 U2121 ( .A1(n1393), .A2(n890), .ZN(n1339) );
  XNOR2_X2 U2122 ( .A(n619), .B(n620), .ZN(n1413) );
  XNOR2_X2 U2123 ( .A(\SUMB[17][14] ), .B(n951), .ZN(n619) );
  XNOR2_X2 U2124 ( .A(\CARRYB[18][12] ), .B(\ab[19][12] ), .ZN(n620) );
  NAND2_X2 U2125 ( .A1(\ab[5][22] ), .A2(\SUMB[4][23] ), .ZN(net80795) );
  NAND3_X4 U2126 ( .A1(n2057), .A2(n2058), .A3(n2059), .ZN(n621) );
  NAND3_X2 U2127 ( .A1(n2057), .A2(n2058), .A3(n2059), .ZN(\CARRYB[7][8] ) );
  NAND2_X2 U2128 ( .A1(\ab[7][8] ), .A2(n1425), .ZN(n2059) );
  NAND2_X2 U2129 ( .A1(n1766), .A2(net90702), .ZN(n1604) );
  NAND2_X1 U2130 ( .A1(\ab[7][21] ), .A2(\SUMB[6][22] ), .ZN(n987) );
  NOR2_X1 U2131 ( .A1(net70478), .A2(net77964), .ZN(\ab[3][22] ) );
  NAND2_X2 U2132 ( .A1(\ab[4][22] ), .A2(n843), .ZN(net84313) );
  NAND2_X4 U2133 ( .A1(n1349), .A2(n1348), .ZN(\SUMB[19][4] ) );
  NAND2_X4 U2134 ( .A1(n623), .A2(n624), .ZN(net90818) );
  INV_X4 U2135 ( .A(net88700), .ZN(n622) );
  NAND2_X2 U2136 ( .A1(net92405), .A2(net148015), .ZN(n625) );
  NAND2_X4 U2137 ( .A1(n625), .A2(n626), .ZN(net87411) );
  XOR2_X1 U2138 ( .A(\CARRYB[10][0] ), .B(\ab[11][0] ), .Z(n1139) );
  NAND2_X2 U2139 ( .A1(\CARRYB[10][0] ), .A2(\ab[11][0] ), .ZN(n1140) );
  NAND2_X2 U2140 ( .A1(n704), .A2(\SUMB[9][9] ), .ZN(n707) );
  NAND2_X2 U2141 ( .A1(\CARRYB[15][12] ), .A2(\SUMB[15][13] ), .ZN(n1087) );
  NAND2_X4 U2142 ( .A1(\SUMB[20][5] ), .A2(\ab[21][4] ), .ZN(net82407) );
  INV_X2 U2143 ( .A(net90702), .ZN(net86601) );
  INV_X4 U2144 ( .A(n1218), .ZN(n1219) );
  NAND2_X2 U2145 ( .A1(n888), .A2(n889), .ZN(n890) );
  XNOR2_X2 U2146 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .ZN(n942) );
  NAND2_X2 U2147 ( .A1(n1284), .A2(n1553), .ZN(n629) );
  NAND2_X4 U2148 ( .A1(n627), .A2(n628), .ZN(n630) );
  NAND2_X4 U2149 ( .A1(n630), .A2(n629), .ZN(\SUMB[14][7] ) );
  INV_X8 U2150 ( .A(n1284), .ZN(n627) );
  NAND2_X2 U2151 ( .A1(n1856), .A2(net84657), .ZN(n632) );
  NAND2_X4 U2152 ( .A1(n631), .A2(net148230), .ZN(n633) );
  NAND2_X4 U2153 ( .A1(n632), .A2(n633), .ZN(\SUMB[16][6] ) );
  INV_X4 U2154 ( .A(n1856), .ZN(n631) );
  INV_X4 U2155 ( .A(net84657), .ZN(net148230) );
  NAND2_X1 U2156 ( .A1(n1718), .A2(net86662), .ZN(n635) );
  NAND2_X2 U2157 ( .A1(n634), .A2(net148235), .ZN(n636) );
  NAND2_X4 U2158 ( .A1(n635), .A2(n636), .ZN(\SUMB[18][5] ) );
  BUF_X4 U2161 ( .A(\SUMB[13][8] ), .Z(n1284) );
  BUF_X4 U2162 ( .A(\SUMB[15][7] ), .Z(net84657) );
  NAND2_X2 U2163 ( .A1(\SUMB[18][5] ), .A2(n2109), .ZN(n1348) );
  NAND2_X2 U2164 ( .A1(\ab[9][7] ), .A2(\CARRYB[8][7] ), .ZN(n2018) );
  XNOR2_X2 U2165 ( .A(n2111), .B(\SUMB[2][19] ), .ZN(n852) );
  NAND2_X4 U2166 ( .A1(\CARRYB[3][10] ), .A2(\ab[4][10] ), .ZN(n1393) );
  INV_X8 U2167 ( .A(\CARRYB[18][4] ), .ZN(n1858) );
  NAND2_X4 U2168 ( .A1(\SUMB[18][3] ), .A2(\ab[19][2] ), .ZN(n1912) );
  NAND2_X4 U2169 ( .A1(n1341), .A2(net88638), .ZN(n1336) );
  NAND2_X2 U2170 ( .A1(\CARRYB[13][4] ), .A2(\ab[14][4] ), .ZN(n1633) );
  INV_X4 U2171 ( .A(\SUMB[2][8] ), .ZN(net85035) );
  INV_X4 U2172 ( .A(n1504), .ZN(n885) );
  NAND2_X4 U2173 ( .A1(n638), .A2(n637), .ZN(n640) );
  INV_X4 U2174 ( .A(n1628), .ZN(n1191) );
  NAND2_X4 U2175 ( .A1(n830), .A2(n831), .ZN(net84818) );
  NAND2_X2 U2176 ( .A1(\ab[14][9] ), .A2(net85043), .ZN(n1938) );
  NAND2_X4 U2177 ( .A1(net120653), .A2(n1011), .ZN(\SUMB[10][12] ) );
  NAND2_X4 U2178 ( .A1(n678), .A2(net147930), .ZN(\SUMB[20][5] ) );
  NAND2_X2 U2179 ( .A1(\ab[5][16] ), .A2(\CARRYB[4][16] ), .ZN(n639) );
  INV_X1 U2180 ( .A(\ab[5][16] ), .ZN(n637) );
  INV_X4 U2181 ( .A(net93683), .ZN(n642) );
  AND3_X2 U2182 ( .A1(net86158), .A2(net86159), .A3(n1019), .ZN(n645) );
  NAND2_X2 U2183 ( .A1(\SUMB[11][13] ), .A2(\ab[12][12] ), .ZN(net86159) );
  NAND2_X2 U2184 ( .A1(net124434), .A2(\SUMB[11][13] ), .ZN(net86158) );
  INV_X8 U2185 ( .A(\CARRYB[18][5] ), .ZN(net84707) );
  NAND2_X4 U2186 ( .A1(n1205), .A2(n1576), .ZN(n1578) );
  NAND2_X2 U2187 ( .A1(net83445), .A2(\SUMB[13][14] ), .ZN(net86630) );
  NAND2_X4 U2188 ( .A1(\SUMB[3][11] ), .A2(\ab[4][10] ), .ZN(n1395) );
  XOR2_X2 U2189 ( .A(\CARRYB[15][1] ), .B(n646), .Z(\SUMB[16][1] ) );
  NAND2_X2 U2190 ( .A1(\SUMB[15][2] ), .A2(\CARRYB[15][1] ), .ZN(n647) );
  NAND2_X2 U2191 ( .A1(\ab[16][1] ), .A2(\SUMB[15][2] ), .ZN(n649) );
  NAND3_X4 U2192 ( .A1(n647), .A2(n648), .A3(n649), .ZN(\CARRYB[16][1] ) );
  NAND2_X2 U2195 ( .A1(\CARRYB[14][1] ), .A2(\SUMB[14][2] ), .ZN(n651) );
  NOR2_X2 U2196 ( .A1(net77868), .A2(net70465), .ZN(\ab[15][1] ) );
  NAND3_X4 U2197 ( .A1(n766), .A2(net86134), .A3(net86135), .ZN(
        \CARRYB[14][1] ) );
  INV_X8 U2198 ( .A(net89876), .ZN(\SUMB[20][4] ) );
  NAND2_X1 U2199 ( .A1(\ab[4][18] ), .A2(\SUMB[3][19] ), .ZN(n1724) );
  NAND2_X4 U2200 ( .A1(n654), .A2(n655), .ZN(n657) );
  NAND2_X4 U2201 ( .A1(n656), .A2(n657), .ZN(net80833) );
  INV_X4 U2202 ( .A(n803), .ZN(n655) );
  NAND2_X4 U2203 ( .A1(n658), .A2(n659), .ZN(n660) );
  INV_X1 U2204 ( .A(\ab[16][9] ), .ZN(n659) );
  NAND2_X2 U2205 ( .A1(net80833), .A2(\SUMB[3][17] ), .ZN(net148053) );
  INV_X4 U2206 ( .A(net80833), .ZN(net148051) );
  NAND2_X2 U2207 ( .A1(\CARRYB[8][13] ), .A2(net83438), .ZN(n663) );
  NAND2_X4 U2208 ( .A1(n661), .A2(n662), .ZN(n664) );
  NAND2_X4 U2209 ( .A1(n663), .A2(n664), .ZN(net80346) );
  INV_X4 U2210 ( .A(net84447), .ZN(n661) );
  INV_X4 U2211 ( .A(net83438), .ZN(n662) );
  INV_X2 U2212 ( .A(\ab[4][16] ), .ZN(n803) );
  INV_X1 U2213 ( .A(\ab[9][13] ), .ZN(net83438) );
  INV_X8 U2214 ( .A(\CARRYB[11][13] ), .ZN(n1041) );
  INV_X8 U2215 ( .A(\CARRYB[9][14] ), .ZN(n1038) );
  INV_X4 U2216 ( .A(net83202), .ZN(net147928) );
  NAND2_X4 U2217 ( .A1(net88887), .A2(\ab[20][4] ), .ZN(n2229) );
  NAND2_X2 U2218 ( .A1(\CARRYB[7][7] ), .A2(\SUMB[7][8] ), .ZN(n1861) );
  CLKBUF_X2 U2219 ( .A(\CARRYB[22][4] ), .Z(net84213) );
  NAND2_X4 U2220 ( .A1(n665), .A2(n666), .ZN(n668) );
  NAND2_X4 U2221 ( .A1(n667), .A2(n668), .ZN(n1243) );
  INV_X4 U2222 ( .A(\CARRYB[11][4] ), .ZN(n665) );
  INV_X1 U2223 ( .A(\ab[12][4] ), .ZN(n666) );
  NAND2_X2 U2224 ( .A1(net81431), .A2(net86385), .ZN(n669) );
  NAND2_X4 U2225 ( .A1(net147998), .A2(net147999), .ZN(n670) );
  NAND2_X4 U2226 ( .A1(n669), .A2(n670), .ZN(PRODUCT[29]) );
  INV_X4 U2227 ( .A(net81431), .ZN(net147998) );
  INV_X4 U2228 ( .A(net86385), .ZN(net147999) );
  NAND2_X1 U2229 ( .A1(\CARRYB[8][6] ), .A2(\ab[9][6] ), .ZN(n673) );
  INV_X4 U2230 ( .A(\CARRYB[8][6] ), .ZN(n671) );
  INV_X4 U2231 ( .A(\ab[9][6] ), .ZN(n672) );
  NOR2_X4 U2232 ( .A1(net77892), .A2(net70471), .ZN(\ab[12][4] ) );
  NOR2_X4 U2233 ( .A1(net77906), .A2(net70477), .ZN(\ab[9][6] ) );
  NAND2_X2 U2234 ( .A1(\CARRYB[14][0] ), .A2(\SUMB[14][1] ), .ZN(n1409) );
  NAND2_X4 U2235 ( .A1(\ab[17][1] ), .A2(\CARRYB[16][1] ), .ZN(n743) );
  NAND2_X4 U2236 ( .A1(\CARRYB[19][0] ), .A2(\SUMB[19][1] ), .ZN(n2102) );
  NAND2_X2 U2237 ( .A1(\SUMB[2][6] ), .A2(\CARRYB[2][5] ), .ZN(n732) );
  XNOR2_X2 U2238 ( .A(\CARRYB[15][3] ), .B(\ab[16][3] ), .ZN(n862) );
  NAND2_X2 U2239 ( .A1(\SUMB[11][4] ), .A2(\CARRYB[11][3] ), .ZN(n1675) );
  INV_X1 U2240 ( .A(n1750), .ZN(n676) );
  CLKBUF_X3 U2241 ( .A(n1261), .Z(n946) );
  XNOR2_X2 U2242 ( .A(\CARRYB[8][7] ), .B(\ab[9][7] ), .ZN(n1176) );
  XNOR2_X2 U2243 ( .A(n1222), .B(\ab[15][3] ), .ZN(n1010) );
  INV_X1 U2244 ( .A(\SUMB[6][13] ), .ZN(net88166) );
  INV_X1 U2245 ( .A(net83796), .ZN(net84891) );
  NAND2_X2 U2246 ( .A1(\CARRYB[11][5] ), .A2(\ab[12][5] ), .ZN(n1636) );
  NAND2_X2 U2247 ( .A1(n677), .A2(net147922), .ZN(net82757) );
  NAND2_X2 U2248 ( .A1(n1928), .A2(n1120), .ZN(n680) );
  NAND2_X4 U2249 ( .A1(n681), .A2(n680), .ZN(\SUMB[3][12] ) );
  INV_X4 U2250 ( .A(n1120), .ZN(n679) );
  NAND3_X2 U2251 ( .A1(n1776), .A2(n1775), .A3(n1774), .ZN(net147936) );
  NAND2_X4 U2253 ( .A1(n2364), .A2(net147938), .ZN(net147940) );
  INV_X8 U2255 ( .A(net86844), .ZN(net120468) );
  NAND2_X2 U2256 ( .A1(\ab[10][8] ), .A2(\CARRYB[9][8] ), .ZN(n1774) );
  NAND2_X4 U2257 ( .A1(n1728), .A2(n1727), .ZN(n682) );
  NAND2_X4 U2258 ( .A1(n685), .A2(n686), .ZN(\SUMB[22][7] ) );
  NAND2_X2 U2259 ( .A1(net92322), .A2(net92323), .ZN(n689) );
  NAND2_X4 U2260 ( .A1(n687), .A2(n688), .ZN(n690) );
  NAND2_X4 U2261 ( .A1(n689), .A2(n690), .ZN(net92321) );
  INV_X4 U2262 ( .A(net92322), .ZN(n687) );
  INV_X4 U2263 ( .A(net92323), .ZN(n688) );
  NAND2_X2 U2264 ( .A1(net81113), .A2(\SUMB[20][9] ), .ZN(n693) );
  NAND2_X4 U2265 ( .A1(n691), .A2(n692), .ZN(n694) );
  NAND2_X4 U2266 ( .A1(n693), .A2(n694), .ZN(\SUMB[21][8] ) );
  INV_X4 U2267 ( .A(\SUMB[20][9] ), .ZN(n691) );
  INV_X4 U2268 ( .A(net81113), .ZN(n692) );
  NAND2_X2 U2269 ( .A1(n2282), .A2(\SUMB[22][7] ), .ZN(n698) );
  NAND2_X4 U2270 ( .A1(n696), .A2(n697), .ZN(n699) );
  NAND2_X4 U2271 ( .A1(n698), .A2(n699), .ZN(n1780) );
  INV_X4 U2272 ( .A(n2282), .ZN(n696) );
  NAND2_X1 U2273 ( .A1(n1067), .A2(\SUMB[11][15] ), .ZN(n702) );
  NAND2_X4 U2274 ( .A1(n702), .A2(n703), .ZN(\SUMB[12][14] ) );
  INV_X2 U2275 ( .A(n1067), .ZN(n701) );
  NAND2_X2 U2276 ( .A1(n1727), .A2(n1728), .ZN(\SUMB[16][11] ) );
  NAND2_X1 U2277 ( .A1(\SUMB[12][14] ), .A2(\ab[13][13] ), .ZN(n1574) );
  NAND3_X4 U2278 ( .A1(n1639), .A2(n1641), .A3(n1640), .ZN(\CARRYB[13][4] ) );
  NAND2_X1 U2279 ( .A1(n1773), .A2(n705), .ZN(n706) );
  NAND2_X2 U2280 ( .A1(n706), .A2(n707), .ZN(\SUMB[10][8] ) );
  INV_X4 U2281 ( .A(n1773), .ZN(n704) );
  INV_X1 U2282 ( .A(\SUMB[9][9] ), .ZN(n705) );
  NAND2_X4 U2283 ( .A1(n1174), .A2(n1175), .ZN(n1618) );
  NAND2_X1 U2284 ( .A1(\CARRYB[16][12] ), .A2(\SUMB[16][13] ), .ZN(n892) );
  XNOR2_X2 U2285 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .ZN(n708) );
  INV_X4 U2286 ( .A(n708), .ZN(n1205) );
  NAND2_X2 U2287 ( .A1(n1419), .A2(\SUMB[3][20] ), .ZN(n1422) );
  NAND3_X1 U2288 ( .A1(n1714), .A2(n1715), .A3(n1716), .ZN(n861) );
  NAND2_X4 U2289 ( .A1(n1601), .A2(n1602), .ZN(n2303) );
  NAND2_X4 U2290 ( .A1(\ab[6][18] ), .A2(\SUMB[5][19] ), .ZN(n1681) );
  INV_X4 U2291 ( .A(\SUMB[5][17] ), .ZN(n1528) );
  BUF_X4 U2292 ( .A(\SUMB[7][10] ), .Z(n1325) );
  NAND3_X4 U2293 ( .A1(net81615), .A2(net81616), .A3(net81617), .ZN(
        \CARRYB[11][2] ) );
  NAND2_X2 U2294 ( .A1(\CARRYB[8][4] ), .A2(\SUMB[8][5] ), .ZN(net82101) );
  INV_X2 U2295 ( .A(n709), .ZN(n710) );
  INV_X4 U2296 ( .A(n1356), .ZN(n1262) );
  INV_X4 U2297 ( .A(\CARRYB[15][12] ), .ZN(net87004) );
  NAND2_X4 U2298 ( .A1(n210), .A2(\ab[14][9] ), .ZN(n1939) );
  NAND2_X2 U2299 ( .A1(n713), .A2(\ab[11][2] ), .ZN(net81617) );
  NAND2_X2 U2300 ( .A1(n713), .A2(\SUMB[10][3] ), .ZN(net81615) );
  INV_X4 U2301 ( .A(\ab[9][3] ), .ZN(n714) );
  NOR2_X4 U2302 ( .A1(n719), .A2(net147444), .ZN(n720) );
  XNOR2_X2 U2303 ( .A(n716), .B(net85032), .ZN(net122130) );
  XNOR2_X2 U2304 ( .A(n721), .B(n718), .ZN(\SUMB[10][2] ) );
  OAI21_X4 U2305 ( .B1(\ab[9][2] ), .B2(n726), .A(\CARRYB[8][2] ), .ZN(n712)
         );
  NAND2_X2 U2306 ( .A1(n726), .A2(\ab[9][2] ), .ZN(n711) );
  INV_X4 U2307 ( .A(n720), .ZN(n721) );
  XNOR2_X2 U2308 ( .A(n725), .B(n715), .ZN(n724) );
  INV_X4 U2309 ( .A(n724), .ZN(\SUMB[9][2] ) );
  MUX2_X2 U2310 ( .A(n723), .B(n356), .S(\SUMB[8][4] ), .Z(n722) );
  XNOR2_X2 U2311 ( .A(n726), .B(\ab[9][2] ), .ZN(n725) );
  INV_X32 U2312 ( .A(B[2]), .ZN(net77878) );
  OAI211_X1 U2313 ( .C1(net77878), .C2(net70475), .A(n711), .B(n712), .ZN(n717) );
  XNOR2_X1 U2314 ( .A(\ab[9][3] ), .B(n728), .ZN(n723) );
  NAND2_X1 U2315 ( .A1(\ab[9][3] ), .A2(n728), .ZN(net82848) );
  INV_X4 U2316 ( .A(n727), .ZN(n726) );
  INV_X2 U2317 ( .A(\SUMB[8][3] ), .ZN(n727) );
  INV_X4 U2318 ( .A(n729), .ZN(n728) );
  INV_X2 U2319 ( .A(\CARRYB[8][3] ), .ZN(n729) );
  NAND2_X1 U2320 ( .A1(\ab[9][3] ), .A2(\SUMB[8][4] ), .ZN(net82849) );
  NAND2_X4 U2321 ( .A1(n722), .A2(n354), .ZN(n718) );
  INV_X8 U2322 ( .A(net147451), .ZN(net147444) );
  INV_X1 U2323 ( .A(\CARRYB[8][2] ), .ZN(n715) );
  AOI21_X4 U2324 ( .B1(n717), .B2(n718), .A(net147444), .ZN(n716) );
  INV_X2 U2325 ( .A(n716), .ZN(n713) );
  NAND2_X4 U2326 ( .A1(n711), .A2(n712), .ZN(net147421) );
  NOR2_X2 U2327 ( .A1(net147421), .A2(n357), .ZN(n719) );
  NAND3_X2 U2328 ( .A1(n735), .A2(net84928), .A3(net84929), .ZN(\CARRYB[4][5] ) );
  NAND2_X1 U2329 ( .A1(\ab[5][5] ), .A2(\CARRYB[4][5] ), .ZN(net88209) );
  XNOR2_X1 U2330 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .ZN(net89958) );
  NAND2_X2 U2331 ( .A1(\CARRYB[4][5] ), .A2(\SUMB[4][6] ), .ZN(net88211) );
  NAND2_X1 U2332 ( .A1(\CARRYB[3][5] ), .A2(\SUMB[3][6] ), .ZN(net84929) );
  NAND2_X1 U2333 ( .A1(\ab[4][5] ), .A2(\SUMB[3][6] ), .ZN(net84928) );
  NAND2_X1 U2334 ( .A1(\ab[4][5] ), .A2(\CARRYB[3][5] ), .ZN(n735) );
  NAND2_X1 U2336 ( .A1(\ab[3][5] ), .A2(\CARRYB[2][5] ), .ZN(n734) );
  NAND2_X2 U2337 ( .A1(\ab[3][5] ), .A2(\SUMB[2][6] ), .ZN(n733) );
  NAND2_X2 U2339 ( .A1(\ab[3][6] ), .A2(net87962), .ZN(net84925) );
  NAND2_X2 U2340 ( .A1(\CARRYB[2][6] ), .A2(net87962), .ZN(net84926) );
  INV_X2 U2341 ( .A(\SUMB[2][7] ), .ZN(net87961) );
  NAND2_X2 U2342 ( .A1(net85036), .A2(n567), .ZN(net84116) );
  NAND2_X2 U2343 ( .A1(\ab[3][7] ), .A2(n567), .ZN(net84118) );
  INV_X4 U2344 ( .A(n731), .ZN(\SUMB[1][8] ) );
  XNOR2_X2 U2345 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .ZN(n731) );
  INV_X4 U2346 ( .A(\*UDW_*112734/net78687 ), .ZN(\CARRYB[1][7] ) );
  NAND2_X2 U2347 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .ZN(
        \*UDW_*112734/net78687 ) );
  NOR2_X2 U2348 ( .A1(net77912), .A2(net77970), .ZN(\ab[2][7] ) );
  INV_X16 U2349 ( .A(n26), .ZN(net77970) );
  NAND3_X2 U2350 ( .A1(net86129), .A2(n737), .A3(net86131), .ZN(
        \CARRYB[13][1] ) );
  NAND2_X2 U2351 ( .A1(\ab[14][1] ), .A2(\CARRYB[13][1] ), .ZN(net86134) );
  NAND2_X2 U2352 ( .A1(\CARRYB[13][1] ), .A2(\SUMB[13][2] ), .ZN(net86135) );
  NAND2_X2 U2353 ( .A1(\CARRYB[12][1] ), .A2(\SUMB[12][2] ), .ZN(net86131) );
  NAND2_X2 U2354 ( .A1(\ab[13][1] ), .A2(\SUMB[12][2] ), .ZN(n737) );
  NAND2_X2 U2355 ( .A1(\CARRYB[12][1] ), .A2(\ab[13][1] ), .ZN(net86129) );
  XNOR2_X2 U2356 ( .A(\SUMB[10][3] ), .B(net122130), .ZN(\SUMB[11][2] ) );
  NAND2_X2 U2357 ( .A1(\CARRYB[10][1] ), .A2(\SUMB[10][2] ), .ZN(n740) );
  NAND2_X2 U2358 ( .A1(\ab[11][1] ), .A2(\SUMB[10][2] ), .ZN(n739) );
  NAND2_X2 U2359 ( .A1(\CARRYB[10][1] ), .A2(\ab[11][1] ), .ZN(n738) );
  XNOR2_X2 U2360 ( .A(n741), .B(\SUMB[11][3] ), .ZN(\SUMB[12][2] ) );
  XNOR2_X2 U2361 ( .A(\CARRYB[11][2] ), .B(\ab[12][2] ), .ZN(n741) );
  NOR2_X4 U2362 ( .A1(net77868), .A2(net70469), .ZN(\ab[13][1] ) );
  NAND2_X2 U2363 ( .A1(\ab[19][1] ), .A2(\CARRYB[18][1] ), .ZN(net81095) );
  XNOR2_X1 U2364 ( .A(\CARRYB[18][1] ), .B(\ab[19][1] ), .ZN(net93676) );
  NAND2_X2 U2365 ( .A1(\CARRYB[17][1] ), .A2(\SUMB[17][2] ), .ZN(n747) );
  XNOR2_X2 U2366 ( .A(n742), .B(\CARRYB[16][2] ), .ZN(\SUMB[17][2] ) );
  XNOR2_X2 U2367 ( .A(\CARRYB[16][1] ), .B(net88712), .ZN(net82532) );
  NAND2_X2 U2368 ( .A1(\SUMB[16][1] ), .A2(\CARRYB[16][0] ), .ZN(net86656) );
  XOR2_X1 U2369 ( .A(\ab[17][0] ), .B(\SUMB[16][1] ), .Z(net86653) );
  NOR2_X4 U2370 ( .A1(net77868), .A2(net70463), .ZN(\ab[16][1] ) );
  NAND3_X2 U2371 ( .A1(n750), .A2(n751), .A3(n752), .ZN(\CARRYB[23][1] ) );
  NAND2_X2 U2372 ( .A1(\ab[23][1] ), .A2(\CARRYB[22][1] ), .ZN(n752) );
  NAND3_X2 U2373 ( .A1(net82541), .A2(net82542), .A3(net82543), .ZN(
        \CARRYB[22][1] ) );
  NAND2_X2 U2374 ( .A1(n748), .A2(\SUMB[22][2] ), .ZN(n750) );
  NOR2_X2 U2375 ( .A1(net77866), .A2(net70449), .ZN(\ab[23][1] ) );
  XNOR2_X2 U2376 ( .A(n748), .B(\ab[23][1] ), .ZN(net93713) );
  NAND2_X2 U2377 ( .A1(\CARRYB[21][1] ), .A2(\SUMB[21][2] ), .ZN(net82541) );
  NAND3_X2 U2378 ( .A1(net82541), .A2(net82542), .A3(net82543), .ZN(n748) );
  XNOR2_X2 U2380 ( .A(\SUMB[21][3] ), .B(n749), .ZN(\SUMB[22][2] ) );
  INV_X1 U2381 ( .A(\SUMB[22][2] ), .ZN(net83357) );
  XNOR2_X2 U2382 ( .A(\CARRYB[21][2] ), .B(\ab[22][2] ), .ZN(n749) );
  XNOR2_X2 U2383 ( .A(n753), .B(\CARRYB[21][1] ), .ZN(\SUMB[22][1] ) );
  XNOR2_X2 U2384 ( .A(\SUMB[21][2] ), .B(\ab[22][1] ), .ZN(n753) );
  NAND2_X2 U2385 ( .A1(\SUMB[21][3] ), .A2(n372), .ZN(net80924) );
  NAND3_X2 U2386 ( .A1(net81095), .A2(n756), .A3(net81097), .ZN(
        \CARRYB[19][1] ) );
  NAND2_X2 U2387 ( .A1(\ab[20][1] ), .A2(\CARRYB[19][1] ), .ZN(net80850) );
  NAND2_X2 U2388 ( .A1(\CARRYB[19][1] ), .A2(\SUMB[19][2] ), .ZN(net80852) );
  NAND2_X2 U2389 ( .A1(\ab[19][1] ), .A2(\SUMB[18][2] ), .ZN(n756) );
  XNOR2_X2 U2390 ( .A(n754), .B(n755), .ZN(\SUMB[18][2] ) );
  XNOR2_X2 U2391 ( .A(net93676), .B(n359), .ZN(\SUMB[19][1] ) );
  BUF_X8 U2392 ( .A(\SUMB[17][3] ), .Z(n755) );
  NOR2_X4 U2393 ( .A1(net77868), .A2(net70457), .ZN(\ab[19][1] ) );
  NAND2_X2 U2394 ( .A1(\CARRYB[17][2] ), .A2(\SUMB[17][3] ), .ZN(net81112) );
  NAND2_X2 U2395 ( .A1(\ab[18][2] ), .A2(\SUMB[17][3] ), .ZN(net81111) );
  NAND2_X2 U2396 ( .A1(\ab[18][2] ), .A2(\CARRYB[17][2] ), .ZN(net81110) );
  NAND3_X2 U2397 ( .A1(n759), .A2(n760), .A3(n761), .ZN(\CARRYB[2][6] ) );
  NAND2_X2 U2398 ( .A1(\ab[3][6] ), .A2(\CARRYB[2][6] ), .ZN(net84924) );
  NAND2_X1 U2399 ( .A1(\ab[2][6] ), .A2(n350), .ZN(n761) );
  NAND2_X2 U2400 ( .A1(n350), .A2(\SUMB[1][7] ), .ZN(n759) );
  INV_X4 U2401 ( .A(n757), .ZN(\SUMB[1][7] ) );
  XNOR2_X2 U2402 ( .A(\SUMB[1][7] ), .B(n758), .ZN(\SUMB[2][6] ) );
  XNOR2_X1 U2403 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .ZN(n757) );
  NOR2_X2 U2404 ( .A1(net77906), .A2(net77970), .ZN(\ab[2][6] ) );
  XNOR2_X2 U2405 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .ZN(\*UDW_*112739/net78703 ) );
  NOR2_X2 U2406 ( .A1(net124610), .A2(net70492), .ZN(\ab[0][29] ) );
  NAND2_X2 U2407 ( .A1(\CARRYB[15][0] ), .A2(\SUMB[15][1] ), .ZN(net86652) );
  NAND2_X2 U2408 ( .A1(\ab[16][0] ), .A2(\SUMB[15][1] ), .ZN(net86651) );
  XOR2_X1 U2409 ( .A(net86649), .B(\SUMB[15][1] ), .Z(PRODUCT[16]) );
  NAND2_X2 U2410 ( .A1(\SUMB[13][2] ), .A2(\ab[14][1] ), .ZN(n766) );
  INV_X16 U2411 ( .A(A[15]), .ZN(net70465) );
  NAND3_X4 U2412 ( .A1(n764), .A2(n763), .A3(n762), .ZN(\CARRYB[13][2] ) );
  NAND2_X4 U2413 ( .A1(\ab[14][2] ), .A2(\CARRYB[13][2] ), .ZN(net81780) );
  NAND2_X2 U2414 ( .A1(n19), .A2(\SUMB[12][3] ), .ZN(n764) );
  NAND2_X2 U2415 ( .A1(\ab[13][2] ), .A2(\SUMB[12][3] ), .ZN(n763) );
  XNOR2_X2 U2416 ( .A(\SUMB[12][4] ), .B(n767), .ZN(\SUMB[13][3] ) );
  XNOR2_X2 U2417 ( .A(n51), .B(\ab[13][3] ), .ZN(n767) );
  NOR2_X4 U2418 ( .A1(net77878), .A2(net70467), .ZN(\ab[14][2] ) );
  XNOR2_X2 U2419 ( .A(\CARRYB[8][4] ), .B(\ab[9][4] ), .ZN(net82601) );
  XNOR2_X2 U2420 ( .A(n769), .B(\CARRYB[6][5] ), .ZN(\SUMB[7][5] ) );
  XNOR2_X2 U2421 ( .A(\SUMB[6][6] ), .B(\ab[7][5] ), .ZN(n769) );
  INV_X32 U2422 ( .A(B[4]), .ZN(net77892) );
  XNOR2_X2 U2423 ( .A(\SUMB[5][6] ), .B(n768), .ZN(\SUMB[6][5] ) );
  XNOR2_X2 U2424 ( .A(\CARRYB[5][5] ), .B(\ab[6][5] ), .ZN(n768) );
  NAND3_X4 U2425 ( .A1(net88198), .A2(net88199), .A3(net88200), .ZN(
        \CARRYB[6][4] ) );
  NAND2_X2 U2426 ( .A1(n343), .A2(\SUMB[5][5] ), .ZN(net88200) );
  XNOR2_X2 U2427 ( .A(n770), .B(\CARRYB[9][3] ), .ZN(\SUMB[10][3] ) );
  NAND2_X2 U2428 ( .A1(\ab[11][2] ), .A2(\SUMB[10][3] ), .ZN(net81616) );
  XNOR2_X2 U2429 ( .A(\SUMB[9][4] ), .B(\ab[10][3] ), .ZN(n770) );
  NOR2_X1 U2430 ( .A1(net77878), .A2(net70473), .ZN(\ab[11][2] ) );
  XNOR2_X2 U2431 ( .A(net121523), .B(n564), .ZN(net122156) );
  XNOR2_X2 U2432 ( .A(net121523), .B(n564), .ZN(\SUMB[23][2] ) );
  NAND2_X2 U2433 ( .A1(n394), .A2(\SUMB[22][3] ), .ZN(net80255) );
  NAND2_X2 U2434 ( .A1(\SUMB[22][3] ), .A2(\ab[23][2] ), .ZN(net80254) );
  XNOR2_X2 U2435 ( .A(net89958), .B(net125691), .ZN(\SUMB[5][5] ) );
  NOR2_X4 U2436 ( .A1(net77898), .A2(net77946), .ZN(\ab[5][5] ) );
  NAND2_X2 U2437 ( .A1(\ab[5][5] ), .A2(\SUMB[4][6] ), .ZN(net88210) );
  NAND2_X2 U2438 ( .A1(\ab[6][4] ), .A2(\SUMB[5][5] ), .ZN(net88199) );
  NAND2_X2 U2439 ( .A1(\ab[6][4] ), .A2(n343), .ZN(net88198) );
  NAND3_X2 U2440 ( .A1(n771), .A2(n772), .A3(n773), .ZN(\CARRYB[7][3] ) );
  NAND2_X2 U2441 ( .A1(\CARRYB[6][3] ), .A2(\SUMB[6][4] ), .ZN(n773) );
  NAND2_X2 U2442 ( .A1(\ab[7][3] ), .A2(\SUMB[6][4] ), .ZN(n772) );
  NAND2_X1 U2443 ( .A1(\ab[7][3] ), .A2(\CARRYB[6][3] ), .ZN(n771) );
  XNOR2_X2 U2444 ( .A(net92884), .B(\SUMB[5][5] ), .ZN(\SUMB[6][4] ) );
  CLKBUF_X3 U2445 ( .A(\SUMB[4][6] ), .Z(net125691) );
  XNOR2_X2 U2446 ( .A(n774), .B(\SUMB[3][7] ), .ZN(\SUMB[4][6] ) );
  NAND2_X1 U2447 ( .A1(\ab[4][6] ), .A2(\SUMB[3][7] ), .ZN(net88207) );
  NAND3_X4 U2448 ( .A1(net79882), .A2(net79881), .A3(net79880), .ZN(
        \CARRYB[28][1] ) );
  XNOR2_X2 U2449 ( .A(net80927), .B(net89104), .ZN(net89109) );
  NAND2_X4 U2450 ( .A1(net89109), .A2(net123363), .ZN(net79882) );
  INV_X4 U2451 ( .A(net88699), .ZN(net87391) );
  INV_X1 U2453 ( .A(\ab[19][8] ), .ZN(n775) );
  INV_X4 U2454 ( .A(\CARRYB[18][8] ), .ZN(net123291) );
  NAND2_X4 U2455 ( .A1(n779), .A2(n780), .ZN(net90022) );
  NAND2_X4 U2456 ( .A1(n778), .A2(net93279), .ZN(n780) );
  INV_X4 U2457 ( .A(\ab[20][7] ), .ZN(net93279) );
  NAND2_X2 U2458 ( .A1(\ab[20][7] ), .A2(\CARRYB[19][7] ), .ZN(n779) );
  INV_X4 U2459 ( .A(\CARRYB[19][7] ), .ZN(n778) );
  NAND2_X1 U2460 ( .A1(\ab[20][7] ), .A2(net91001), .ZN(net80671) );
  NAND2_X2 U2461 ( .A1(net90818), .A2(\ab[20][7] ), .ZN(net80672) );
  NAND2_X4 U2462 ( .A1(net81555), .A2(n781), .ZN(net87681) );
  INV_X1 U2463 ( .A(\ab[21][6] ), .ZN(net81042) );
  INV_X4 U2464 ( .A(net81042), .ZN(net81552) );
  NAND2_X4 U2465 ( .A1(net81553), .A2(net81552), .ZN(net81555) );
  NAND2_X1 U2466 ( .A1(net149530), .A2(n69), .ZN(net80676) );
  NAND2_X1 U2467 ( .A1(\ab[21][6] ), .A2(net149530), .ZN(net80675) );
  NAND2_X1 U2468 ( .A1(\ab[21][6] ), .A2(\CARRYB[20][6] ), .ZN(net80674) );
  NAND2_X4 U2469 ( .A1(net84000), .A2(net84001), .ZN(n784) );
  NAND2_X4 U2470 ( .A1(net79907), .A2(n784), .ZN(net80021) );
  INV_X2 U2471 ( .A(\ab[24][4] ), .ZN(net84001) );
  INV_X8 U2472 ( .A(\CARRYB[23][4] ), .ZN(net84000) );
  NOR2_X4 U2473 ( .A1(net77892), .A2(net70447), .ZN(\ab[24][4] ) );
  NAND2_X4 U2474 ( .A1(\CARRYB[23][4] ), .A2(\ab[24][4] ), .ZN(net79907) );
  NOR2_X4 U2475 ( .A1(net77892), .A2(net70445), .ZN(\ab[25][4] ) );
  NAND3_X4 U2476 ( .A1(net80290), .A2(n782), .A3(n783), .ZN(\CARRYB[23][4] )
         );
  NAND2_X2 U2477 ( .A1(\ab[23][4] ), .A2(\CARRYB[22][4] ), .ZN(n783) );
  NAND2_X4 U2478 ( .A1(net124635), .A2(\ab[23][4] ), .ZN(n782) );
  NAND2_X4 U2479 ( .A1(net120647), .A2(net120648), .ZN(n789) );
  NAND2_X4 U2480 ( .A1(net120649), .A2(n789), .ZN(\SUMB[13][11] ) );
  INV_X4 U2481 ( .A(net84059), .ZN(net120647) );
  NAND2_X2 U2482 ( .A1(net87937), .A2(net87936), .ZN(net84059) );
  NAND2_X4 U2483 ( .A1(n787), .A2(n788), .ZN(\SUMB[12][12] ) );
  NAND2_X2 U2484 ( .A1(n786), .A2(n785), .ZN(n788) );
  INV_X2 U2485 ( .A(net89026), .ZN(n786) );
  INV_X2 U2486 ( .A(n785), .ZN(n790) );
  NAND2_X2 U2487 ( .A1(n790), .A2(net89026), .ZN(n787) );
  NAND2_X4 U2488 ( .A1(net87935), .A2(net87934), .ZN(net87937) );
  NAND2_X4 U2489 ( .A1(net87936), .A2(net87937), .ZN(net93277) );
  INV_X8 U2490 ( .A(\CARRYB[12][11] ), .ZN(net87935) );
  INV_X2 U2491 ( .A(\ab[13][11] ), .ZN(net87934) );
  NAND2_X4 U2492 ( .A1(\CARRYB[12][11] ), .A2(\ab[13][11] ), .ZN(net87936) );
  NAND3_X4 U2493 ( .A1(net82158), .A2(net82159), .A3(n97), .ZN(
        \CARRYB[13][11] ) );
  NAND2_X4 U2494 ( .A1(\SUMB[12][12] ), .A2(\ab[13][11] ), .ZN(net82158) );
  NOR2_X4 U2495 ( .A1(net77920), .A2(net70457), .ZN(\ab[19][8] ) );
  NAND3_X4 U2496 ( .A1(net81559), .A2(net81560), .A3(n791), .ZN(
        \CARRYB[18][8] ) );
  NAND2_X1 U2497 ( .A1(\ab[18][8] ), .A2(\CARRYB[17][8] ), .ZN(n791) );
  NAND2_X2 U2498 ( .A1(\SUMB[17][9] ), .A2(\CARRYB[17][8] ), .ZN(net81560) );
  NAND2_X2 U2499 ( .A1(\SUMB[17][9] ), .A2(\ab[18][8] ), .ZN(net81559) );
  XNOR2_X2 U2500 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .ZN(net88906) );
  XNOR2_X2 U2501 ( .A(\CARRYB[17][8] ), .B(\ab[18][8] ), .ZN(net84349) );
  XNOR2_X2 U2502 ( .A(net84349), .B(\SUMB[17][9] ), .ZN(\SUMB[18][8] ) );
  XNOR2_X2 U2503 ( .A(net88906), .B(\SUMB[17][9] ), .ZN(net88702) );
  NAND2_X2 U2504 ( .A1(net93277), .A2(\SUMB[12][12] ), .ZN(net120649) );
  XNOR2_X2 U2505 ( .A(net93277), .B(net82263), .ZN(net87942) );
  XNOR2_X2 U2506 ( .A(net93277), .B(net82263), .ZN(net93756) );
  NAND3_X4 U2507 ( .A1(net82162), .A2(net82161), .A3(net82160), .ZN(
        \CARRYB[14][10] ) );
  XNOR2_X2 U2508 ( .A(\CARRYB[14][10] ), .B(\ab[15][10] ), .ZN(net86799) );
  NAND2_X1 U2509 ( .A1(\CARRYB[14][10] ), .A2(\ab[15][10] ), .ZN(net82559) );
  NAND2_X2 U2510 ( .A1(net88668), .A2(\CARRYB[14][10] ), .ZN(net82561) );
  NAND2_X4 U2511 ( .A1(\CARRYB[13][10] ), .A2(\ab[14][10] ), .ZN(net82160) );
  NAND2_X4 U2512 ( .A1(net82160), .A2(net88410), .ZN(net84163) );
  NOR2_X2 U2513 ( .A1(net91660), .A2(net70467), .ZN(\ab[14][10] ) );
  INV_X1 U2514 ( .A(\ab[14][10] ), .ZN(net88407) );
  NAND3_X4 U2515 ( .A1(n794), .A2(n793), .A3(n792), .ZN(\CARRYB[13][10] ) );
  NAND2_X2 U2516 ( .A1(\ab[13][10] ), .A2(net124392), .ZN(n792) );
  NAND2_X4 U2517 ( .A1(\SUMB[12][11] ), .A2(\ab[13][10] ), .ZN(n793) );
  NAND2_X4 U2518 ( .A1(n796), .A2(\SUMB[12][11] ), .ZN(n794) );
  INV_X4 U2519 ( .A(\CARRYB[12][10] ), .ZN(n795) );
  NAND3_X2 U2520 ( .A1(net81058), .A2(net81057), .A3(net81056), .ZN(
        \CARRYB[12][10] ) );
  NAND2_X4 U2521 ( .A1(n199), .A2(net121451), .ZN(\SUMB[25][3] ) );
  NAND3_X2 U2522 ( .A1(net80992), .A2(net80991), .A3(net80990), .ZN(net123363)
         );
  NAND2_X4 U2523 ( .A1(net83057), .A2(net93918), .ZN(net80927) );
  NAND2_X4 U2524 ( .A1(net83054), .A2(net83055), .ZN(net83057) );
  INV_X1 U2525 ( .A(\ab[27][2] ), .ZN(net83055) );
  NAND3_X2 U2527 ( .A1(net81372), .A2(net81371), .A3(n555), .ZN(
        \CARRYB[8][13] ) );
  NAND3_X2 U2528 ( .A1(net81372), .A2(net81371), .A3(n555), .ZN(net84447) );
  INV_X2 U2529 ( .A(net87066), .ZN(net88943) );
  INV_X8 U2530 ( .A(\CARRYB[7][13] ), .ZN(net87066) );
  NAND2_X4 U2531 ( .A1(net87066), .A2(net87065), .ZN(net87068) );
  XNOR2_X2 U2532 ( .A(n797), .B(net93800), .ZN(net89356) );
  INV_X4 U2533 ( .A(net88880), .ZN(net88881) );
  NAND2_X1 U2534 ( .A1(net88881), .A2(\ab[7][14] ), .ZN(net81365) );
  XNOR2_X2 U2535 ( .A(net88079), .B(\ab[5][15] ), .ZN(net119976) );
  XNOR2_X2 U2536 ( .A(net88079), .B(net119953), .ZN(net80834) );
  INV_X4 U2537 ( .A(\ab[5][15] ), .ZN(net119953) );
  NAND2_X4 U2538 ( .A1(n800), .A2(n801), .ZN(n802) );
  XNOR2_X2 U2539 ( .A(n802), .B(\SUMB[2][18] ), .ZN(net124367) );
  XNOR2_X2 U2540 ( .A(n802), .B(\SUMB[2][18] ), .ZN(\SUMB[3][17] ) );
  NAND2_X4 U2541 ( .A1(n798), .A2(n799), .ZN(n801) );
  INV_X1 U2542 ( .A(\ab[3][17] ), .ZN(n798) );
  NAND2_X2 U2543 ( .A1(\CARRYB[2][17] ), .A2(\ab[3][17] ), .ZN(n800) );
  NOR2_X2 U2544 ( .A1(net88344), .A2(net119855), .ZN(\ab[4][16] ) );
  NAND2_X4 U2545 ( .A1(\SUMB[3][17] ), .A2(\ab[4][16] ), .ZN(net80836) );
  NAND3_X2 U2546 ( .A1(net80668), .A2(net80667), .A3(net149917), .ZN(
        \CARRYB[29][1] ) );
  NAND3_X2 U2547 ( .A1(net80667), .A2(net80668), .A3(net149917), .ZN(net93672)
         );
  NAND2_X4 U2548 ( .A1(net120657), .A2(n804), .ZN(net84208) );
  INV_X4 U2549 ( .A(net84208), .ZN(net87944) );
  INV_X1 U2550 ( .A(\ab[17][9] ), .ZN(net120656) );
  NOR2_X1 U2551 ( .A1(net70452), .A2(net70461), .ZN(\ab[17][9] ) );
  NAND2_X1 U2552 ( .A1(\ab[17][9] ), .A2(\CARRYB[16][9] ), .ZN(net80814) );
  NAND3_X2 U2553 ( .A1(net79980), .A2(net79981), .A3(n805), .ZN(
        \CARRYB[16][9] ) );
  NAND2_X2 U2554 ( .A1(\SUMB[15][10] ), .A2(net121214), .ZN(net79981) );
  CLKBUF_X3 U2555 ( .A(\CARRYB[15][9] ), .Z(net121214) );
  NAND2_X2 U2556 ( .A1(\ab[16][9] ), .A2(\SUMB[15][10] ), .ZN(net79980) );
  NAND3_X4 U2557 ( .A1(net79909), .A2(net79908), .A3(net79907), .ZN(
        \CARRYB[24][4] ) );
  NAND2_X4 U2558 ( .A1(net87941), .A2(net87940), .ZN(net82544) );
  INV_X1 U2559 ( .A(\ab[25][3] ), .ZN(net87939) );
  NAND2_X4 U2560 ( .A1(n3), .A2(\ab[25][3] ), .ZN(net87940) );
  NAND3_X2 U2561 ( .A1(net81007), .A2(net81006), .A3(net87940), .ZN(net123427)
         );
  NAND3_X2 U2562 ( .A1(net81006), .A2(net81007), .A3(net87940), .ZN(
        \CARRYB[25][3] ) );
  NOR2_X4 U2563 ( .A1(net77886), .A2(net70445), .ZN(\ab[25][3] ) );
  INV_X4 U2564 ( .A(A[25]), .ZN(net70445) );
  NAND2_X4 U2565 ( .A1(net86024), .A2(net86023), .ZN(\SUMB[24][4] ) );
  INV_X2 U2566 ( .A(net93813), .ZN(net86022) );
  NAND3_X4 U2567 ( .A1(net80352), .A2(net90996), .A3(net80353), .ZN(
        \CARRYB[10][12] ) );
  NAND2_X2 U2568 ( .A1(\CARRYB[10][12] ), .A2(\ab[11][12] ), .ZN(net83630) );
  NAND2_X2 U2569 ( .A1(\SUMB[10][13] ), .A2(\CARRYB[10][12] ), .ZN(net80251)
         );
  BUF_X4 U2570 ( .A(net80351), .Z(net90996) );
  NAND2_X4 U2571 ( .A1(net89065), .A2(net89982), .ZN(net80353) );
  INV_X1 U2572 ( .A(net84820), .ZN(net89982) );
  INV_X4 U2573 ( .A(\CARRYB[9][12] ), .ZN(net84820) );
  NAND2_X4 U2574 ( .A1(net84819), .A2(net84820), .ZN(net84822) );
  NAND2_X4 U2575 ( .A1(\SUMB[9][13] ), .A2(\ab[10][12] ), .ZN(net80352) );
  NAND2_X2 U2576 ( .A1(\CARRYB[9][12] ), .A2(\ab[10][12] ), .ZN(net80351) );
  NAND2_X4 U2577 ( .A1(net80351), .A2(net84822), .ZN(net80983) );
  XNOR2_X2 U2578 ( .A(net85399), .B(net80346), .ZN(net89065) );
  XNOR2_X2 U2580 ( .A(net85399), .B(net80346), .ZN(\SUMB[9][13] ) );
  NAND2_X1 U2581 ( .A1(\SUMB[9][13] ), .A2(net80983), .ZN(net120653) );
  NOR2_X2 U2582 ( .A1(net83784), .A2(net70475), .ZN(\ab[10][12] ) );
  INV_X1 U2583 ( .A(\ab[10][12] ), .ZN(net84819) );
  NAND2_X2 U2584 ( .A1(n2356), .A2(net86884), .ZN(net80686) );
  NAND3_X4 U2585 ( .A1(net80992), .A2(net80991), .A3(net80990), .ZN(
        \CARRYB[27][1] ) );
  NAND3_X2 U2586 ( .A1(net84678), .A2(net84679), .A3(net84680), .ZN(
        \CARRYB[24][3] ) );
  NAND2_X2 U2587 ( .A1(n565), .A2(\CARRYB[8][13] ), .ZN(net80350) );
  NAND3_X4 U2588 ( .A1(net82022), .A2(net82021), .A3(n806), .ZN(
        \CARRYB[12][11] ) );
  NAND2_X4 U2589 ( .A1(net89670), .A2(n808), .ZN(net82021) );
  INV_X1 U2590 ( .A(n807), .ZN(n808) );
  INV_X4 U2591 ( .A(\CARRYB[11][11] ), .ZN(n807) );
  NAND2_X4 U2592 ( .A1(n807), .A2(net84824), .ZN(net84826) );
  NAND3_X2 U2593 ( .A1(net81166), .A2(net81167), .A3(net81168), .ZN(
        \CARRYB[11][11] ) );
  XNOR2_X2 U2594 ( .A(net90262), .B(net81087), .ZN(net124563) );
  XNOR2_X2 U2595 ( .A(net90262), .B(net81087), .ZN(\SUMB[11][12] ) );
  NAND2_X4 U2596 ( .A1(\SUMB[11][12] ), .A2(\ab[12][11] ), .ZN(net82022) );
  NOR2_X4 U2597 ( .A1(net85716), .A2(net70469), .ZN(\ab[13][11] ) );
  NAND3_X2 U2598 ( .A1(net81166), .A2(net81167), .A3(net81168), .ZN(net90604)
         );
  NAND2_X2 U2599 ( .A1(\ab[11][12] ), .A2(\SUMB[10][13] ), .ZN(net80250) );
  NAND2_X2 U2600 ( .A1(net83866), .A2(\SUMB[11][12] ), .ZN(net85457) );
  NAND3_X4 U2601 ( .A1(net80989), .A2(net80988), .A3(net80987), .ZN(
        \CARRYB[26][2] ) );
  NAND2_X4 U2602 ( .A1(\CARRYB[26][2] ), .A2(\ab[27][2] ), .ZN(net93918) );
  NAND2_X2 U2603 ( .A1(\ab[26][2] ), .A2(\CARRYB[25][2] ), .ZN(net80987) );
  NOR2_X4 U2604 ( .A1(net77878), .A2(net70443), .ZN(\ab[26][2] ) );
  INV_X4 U2605 ( .A(A[26]), .ZN(net70443) );
  NAND3_X4 U2606 ( .A1(net80262), .A2(net80261), .A3(net80263), .ZN(
        \CARRYB[25][2] ) );
  NAND2_X2 U2607 ( .A1(net89453), .A2(net87797), .ZN(net80472) );
  NAND3_X2 U2608 ( .A1(net80686), .A2(n809), .A3(net93918), .ZN(
        \CARRYB[27][2] ) );
  NAND3_X2 U2609 ( .A1(net79991), .A2(net79990), .A3(net79989), .ZN(
        \CARRYB[21][5] ) );
  NAND2_X2 U2610 ( .A1(\SUMB[10][12] ), .A2(net87490), .ZN(net81166) );
  NAND2_X1 U2611 ( .A1(\ab[11][11] ), .A2(net88525), .ZN(net81168) );
  NAND2_X4 U2612 ( .A1(net83630), .A2(net83631), .ZN(net81087) );
  NAND2_X4 U2613 ( .A1(net83628), .A2(net83629), .ZN(net83631) );
  NOR2_X4 U2614 ( .A1(net77920), .A2(net70459), .ZN(\ab[18][8] ) );
  INV_X16 U2615 ( .A(A[18]), .ZN(net70459) );
  NAND3_X4 U2616 ( .A1(n812), .A2(n811), .A3(n810), .ZN(\CARRYB[17][8] ) );
  NAND2_X1 U2617 ( .A1(\ab[17][8] ), .A2(\CARRYB[16][8] ), .ZN(n810) );
  NAND2_X4 U2618 ( .A1(n813), .A2(net87945), .ZN(\SUMB[17][9] ) );
  INV_X8 U2619 ( .A(net85807), .ZN(net85808) );
  NAND2_X4 U2620 ( .A1(net85808), .A2(net89819), .ZN(net80812) );
  NAND2_X2 U2621 ( .A1(net87944), .A2(net85807), .ZN(n813) );
  XNOR2_X2 U2622 ( .A(n390), .B(\ab[17][10] ), .ZN(net85325) );
  NAND2_X1 U2623 ( .A1(\ab[17][10] ), .A2(n390), .ZN(net84746) );
  NAND3_X2 U2624 ( .A1(net82561), .A2(net82560), .A3(net82559), .ZN(
        \CARRYB[15][10] ) );
  NAND2_X2 U2625 ( .A1(\SUMB[14][11] ), .A2(\ab[15][10] ), .ZN(net82560) );
  BUF_X4 U2626 ( .A(\SUMB[13][12] ), .Z(net86801) );
  XNOR2_X2 U2627 ( .A(net86801), .B(net90817), .ZN(net88668) );
  NOR2_X1 U2628 ( .A1(net91660), .A2(net70463), .ZN(\ab[16][10] ) );
  NAND2_X4 U2629 ( .A1(net87688), .A2(n815), .ZN(\SUMB[15][11] ) );
  INV_X4 U2630 ( .A(net81169), .ZN(n814) );
  NAND2_X2 U2631 ( .A1(n816), .A2(net81169), .ZN(net87688) );
  NOR2_X1 U2632 ( .A1(net77892), .A2(net70449), .ZN(\ab[23][4] ) );
  NOR2_X1 U2633 ( .A1(net70452), .A2(net70463), .ZN(\ab[16][9] ) );
  XNOR2_X2 U2634 ( .A(net86799), .B(net88668), .ZN(\SUMB[15][10] ) );
  NAND2_X4 U2635 ( .A1(net119921), .A2(n817), .ZN(net82030) );
  NAND3_X2 U2636 ( .A1(net82030), .A2(net82029), .A3(net82031), .ZN(net123303)
         );
  XNOR2_X2 U2637 ( .A(net81983), .B(n821), .ZN(\SUMB[23][5] ) );
  INV_X8 U2638 ( .A(n823), .ZN(n821) );
  NAND2_X4 U2639 ( .A1(net88860), .A2(n821), .ZN(net79906) );
  NAND2_X4 U2640 ( .A1(n821), .A2(\ab[23][5] ), .ZN(net79905) );
  XNOR2_X2 U2641 ( .A(net81983), .B(n821), .ZN(net93813) );
  XNOR2_X2 U2642 ( .A(\SUMB[21][7] ), .B(n822), .ZN(n823) );
  NAND2_X2 U2643 ( .A1(n824), .A2(\CARRYB[21][6] ), .ZN(n819) );
  INV_X4 U2644 ( .A(\CARRYB[21][6] ), .ZN(n818) );
  NAND2_X2 U2645 ( .A1(\SUMB[21][7] ), .A2(net89008), .ZN(net80942) );
  NAND2_X2 U2646 ( .A1(\ab[22][6] ), .A2(\SUMB[21][7] ), .ZN(net80941) );
  NAND2_X1 U2647 ( .A1(\ab[22][6] ), .A2(\CARRYB[21][6] ), .ZN(net80940) );
  INV_X1 U2649 ( .A(\ab[11][12] ), .ZN(net83628) );
  NAND3_X2 U2650 ( .A1(net80251), .A2(net80250), .A3(net83630), .ZN(
        \CARRYB[11][12] ) );
  NOR2_X2 U2651 ( .A1(net83784), .A2(net70473), .ZN(\ab[11][12] ) );
  NAND2_X4 U2652 ( .A1(net124908), .A2(net120511), .ZN(net88079) );
  NAND2_X1 U2653 ( .A1(\ab[5][15] ), .A2(n93), .ZN(net80838) );
  NOR2_X4 U2654 ( .A1(net81424), .A2(net77948), .ZN(\ab[5][15] ) );
  XNOR2_X2 U2655 ( .A(\CARRYB[18][8] ), .B(\ab[19][8] ), .ZN(net88700) );
  NAND2_X4 U2656 ( .A1(\CARRYB[7][13] ), .A2(\ab[8][13] ), .ZN(net87067) );
  NAND2_X4 U2657 ( .A1(net87067), .A2(net87068), .ZN(net81958) );
  INV_X2 U2658 ( .A(\ab[8][13] ), .ZN(net87065) );
  INV_X4 U2659 ( .A(\ab[13][10] ), .ZN(net84007) );
  NAND2_X2 U2660 ( .A1(net84007), .A2(net124392), .ZN(net84211) );
  INV_X4 U2661 ( .A(\SUMB[12][11] ), .ZN(net85465) );
  NAND3_X2 U2662 ( .A1(net81058), .A2(net81057), .A3(net81056), .ZN(net124392)
         );
  NOR2_X1 U2663 ( .A1(net91660), .A2(net70465), .ZN(\ab[15][10] ) );
  XNOR2_X2 U2664 ( .A(n150), .B(n826), .ZN(net88692) );
  NAND2_X1 U2665 ( .A1(\ab[18][9] ), .A2(\SUMB[17][10] ), .ZN(net80880) );
  NAND3_X4 U2666 ( .A1(n829), .A2(n828), .A3(n827), .ZN(\CARRYB[15][9] ) );
  XNOR2_X2 U2667 ( .A(net84163), .B(net93756), .ZN(\SUMB[14][10] ) );
  INV_X4 U2668 ( .A(net120648), .ZN(net82263) );
  NAND2_X2 U2669 ( .A1(net89255), .A2(\CARRYB[14][9] ), .ZN(n829) );
  XNOR2_X2 U2670 ( .A(net84163), .B(net87942), .ZN(net89255) );
  XNOR2_X2 U2671 ( .A(n832), .B(\SUMB[9][14] ), .ZN(\SUMB[10][13] ) );
  XNOR2_X2 U2672 ( .A(\CARRYB[9][13] ), .B(\ab[10][13] ), .ZN(n832) );
  NAND2_X2 U2673 ( .A1(\ab[10][13] ), .A2(\SUMB[9][14] ), .ZN(net80247) );
  NAND2_X2 U2674 ( .A1(\ab[10][13] ), .A2(\CARRYB[9][13] ), .ZN(net80246) );
  NOR2_X2 U2675 ( .A1(net70460), .A2(net70477), .ZN(\ab[9][13] ) );
  NAND2_X2 U2676 ( .A1(\ab[9][13] ), .A2(\CARRYB[8][13] ), .ZN(net80348) );
  XNOR2_X2 U2677 ( .A(net81995), .B(n833), .ZN(\SUMB[8][14] ) );
  NAND2_X2 U2678 ( .A1(\CARRYB[7][14] ), .A2(\SUMB[7][15] ), .ZN(net80355) );
  NAND2_X2 U2679 ( .A1(\ab[8][14] ), .A2(\CARRYB[7][14] ), .ZN(net80356) );
  XNOR2_X2 U2680 ( .A(net81663), .B(n91), .ZN(\SUMB[26][3] ) );
  NAND2_X1 U2681 ( .A1(\SUMB[25][4] ), .A2(net84891), .ZN(net81053) );
  NAND2_X4 U2682 ( .A1(n834), .A2(n835), .ZN(net92317) );
  INV_X4 U2683 ( .A(net81157), .ZN(net92325) );
  NAND2_X4 U2684 ( .A1(n837), .A2(n836), .ZN(net81157) );
  NAND2_X4 U2685 ( .A1(net87654), .A2(net87655), .ZN(n837) );
  INV_X2 U2686 ( .A(net81548), .ZN(net87655) );
  INV_X4 U2687 ( .A(net93672), .ZN(net87654) );
  XNOR2_X2 U2688 ( .A(\CARRYB[13][11] ), .B(\ab[14][11] ), .ZN(net90817) );
  NAND2_X1 U2689 ( .A1(\CARRYB[13][11] ), .A2(\ab[14][11] ), .ZN(net82556) );
  NOR2_X1 U2690 ( .A1(net70482), .A2(n331), .ZN(n838) );
  NOR2_X1 U2691 ( .A1(net70482), .A2(n331), .ZN(\ab[2][24] ) );
  INV_X2 U2692 ( .A(\SUMB[6][21] ), .ZN(n839) );
  INV_X4 U2693 ( .A(n839), .ZN(n840) );
  XNOR2_X2 U2694 ( .A(n841), .B(n34), .ZN(\SUMB[3][22] ) );
  XNOR2_X2 U2695 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .ZN(n841) );
  NAND2_X2 U2696 ( .A1(\ab[7][22] ), .A2(\CARRYB[6][22] ), .ZN(n877) );
  CLKBUF_X2 U2697 ( .A(\SUMB[10][4] ), .Z(n842) );
  INV_X4 U2698 ( .A(\CARRYB[7][11] ), .ZN(n1659) );
  XNOR2_X2 U2699 ( .A(net87855), .B(net90671), .ZN(n843) );
  NAND2_X4 U2700 ( .A1(n885), .A2(net123509), .ZN(n887) );
  NOR2_X1 U2701 ( .A1(net70452), .A2(net77938), .ZN(\ab[6][9] ) );
  INV_X1 U2702 ( .A(\CARRYB[14][0] ), .ZN(n845) );
  INV_X2 U2703 ( .A(n845), .ZN(n846) );
  NAND3_X2 U2704 ( .A1(net80838), .A2(net80839), .A3(net80840), .ZN(n847) );
  INV_X4 U2705 ( .A(net83134), .ZN(net86702) );
  CLKBUF_X3 U2706 ( .A(\SUMB[14][12] ), .Z(net125062) );
  XNOR2_X2 U2707 ( .A(n2367), .B(n1233), .ZN(n848) );
  NAND2_X2 U2708 ( .A1(\ab[19][9] ), .A2(\CARRYB[18][9] ), .ZN(n935) );
  INV_X4 U2709 ( .A(\SUMB[7][21] ), .ZN(n850) );
  INV_X8 U2710 ( .A(n850), .ZN(n851) );
  NAND2_X4 U2711 ( .A1(n1548), .A2(n1549), .ZN(n2111) );
  NAND2_X2 U2712 ( .A1(\CARRYB[26][3] ), .A2(\ab[27][3] ), .ZN(n1535) );
  INV_X2 U2713 ( .A(net91301), .ZN(net83151) );
  NAND2_X4 U2714 ( .A1(\CARRYB[11][9] ), .A2(\ab[12][9] ), .ZN(net88297) );
  XNOR2_X2 U2715 ( .A(n1880), .B(n1217), .ZN(n853) );
  INV_X4 U2716 ( .A(\CARRYB[21][7] ), .ZN(net83120) );
  NAND2_X2 U2717 ( .A1(net81491), .A2(\CARRYB[21][7] ), .ZN(net83121) );
  NAND3_X2 U2718 ( .A1(n1919), .A2(n1918), .A3(n1917), .ZN(n854) );
  XNOR2_X1 U2719 ( .A(\SUMB[6][22] ), .B(n855), .ZN(\SUMB[7][21] ) );
  XNOR2_X2 U2720 ( .A(\CARRYB[6][21] ), .B(\ab[7][21] ), .ZN(n855) );
  XNOR2_X2 U2721 ( .A(n1663), .B(\SUMB[20][10] ), .ZN(n856) );
  BUF_X8 U2722 ( .A(\SUMB[9][2] ), .Z(net124757) );
  NAND3_X2 U2723 ( .A1(n2219), .A2(n2220), .A3(n2221), .ZN(\CARRYB[10][19] )
         );
  NAND2_X4 U2724 ( .A1(\CARRYB[3][14] ), .A2(\ab[4][14] ), .ZN(net92718) );
  XNOR2_X2 U2725 ( .A(\CARRYB[4][20] ), .B(\ab[5][20] ), .ZN(n1210) );
  NOR2_X1 U2726 ( .A1(net80727), .A2(net77948), .ZN(\ab[5][20] ) );
  NAND3_X2 U2727 ( .A1(n2305), .A2(n2304), .A3(n2306), .ZN(\CARRYB[9][16] ) );
  XNOR2_X2 U2728 ( .A(net82396), .B(\SUMB[19][10] ), .ZN(n859) );
  NAND2_X4 U2729 ( .A1(net81033), .A2(n937), .ZN(net82396) );
  XOR2_X2 U2730 ( .A(\ab[13][17] ), .B(\CARRYB[12][17] ), .Z(n860) );
  NOR2_X4 U2731 ( .A1(net82890), .A2(net70469), .ZN(\ab[13][17] ) );
  NAND2_X2 U2732 ( .A1(n299), .A2(net123142), .ZN(n909) );
  NAND2_X2 U2733 ( .A1(\SUMB[6][17] ), .A2(n1368), .ZN(n2251) );
  NAND3_X2 U2735 ( .A1(n1933), .A2(n1934), .A3(n1935), .ZN(\CARRYB[3][21] ) );
  INV_X4 U2736 ( .A(\CARRYB[3][10] ), .ZN(n888) );
  XNOR2_X2 U2737 ( .A(\SUMB[8][6] ), .B(\ab[9][5] ), .ZN(n1448) );
  XNOR2_X2 U2738 ( .A(n862), .B(n871), .ZN(\SUMB[16][3] ) );
  INV_X4 U2739 ( .A(\CARRYB[11][12] ), .ZN(net120585) );
  INV_X2 U2740 ( .A(\SUMB[2][22] ), .ZN(n865) );
  INV_X4 U2741 ( .A(n865), .ZN(n866) );
  INV_X2 U2742 ( .A(\ab[19][9] ), .ZN(net87133) );
  NAND2_X1 U2743 ( .A1(\ab[8][19] ), .A2(\SUMB[7][20] ), .ZN(net79956) );
  XNOR2_X2 U2744 ( .A(n368), .B(\SUMB[19][9] ), .ZN(n869) );
  NAND3_X2 U2745 ( .A1(net79867), .A2(net79868), .A3(n1062), .ZN(
        \CARRYB[25][5] ) );
  NAND2_X1 U2746 ( .A1(\ab[11][0] ), .A2(\SUMB[10][1] ), .ZN(n1141) );
  XOR2_X1 U2747 ( .A(n1139), .B(\SUMB[10][1] ), .Z(PRODUCT[11]) );
  INV_X2 U2748 ( .A(n2060), .ZN(n1458) );
  NAND3_X2 U2749 ( .A1(n1910), .A2(n1909), .A3(n1908), .ZN(\CARRYB[4][7] ) );
  NAND2_X1 U2750 ( .A1(n1781), .A2(n1782), .ZN(n1784) );
  NAND2_X2 U2751 ( .A1(\CARRYB[11][12] ), .A2(\ab[12][12] ), .ZN(n1019) );
  XNOR2_X2 U2752 ( .A(n1942), .B(n1256), .ZN(net124104) );
  NAND3_X2 U2753 ( .A1(n1969), .A2(n1968), .A3(n1967), .ZN(\CARRYB[14][3] ) );
  NAND2_X4 U2754 ( .A1(net123899), .A2(n872), .ZN(n1456) );
  INV_X2 U2755 ( .A(net82757), .ZN(net123897) );
  NAND2_X1 U2756 ( .A1(\CARRYB[12][13] ), .A2(\SUMB[12][14] ), .ZN(n1575) );
  NAND2_X4 U2757 ( .A1(n1386), .A2(n428), .ZN(n1388) );
  NAND2_X1 U2758 ( .A1(\ab[8][16] ), .A2(\CARRYB[7][16] ), .ZN(n2297) );
  NOR2_X1 U2759 ( .A1(n2354), .A2(n242), .ZN(\ab[1][28] ) );
  NAND2_X4 U2760 ( .A1(net123842), .A2(net123843), .ZN(n874) );
  NAND2_X4 U2761 ( .A1(n874), .A2(n873), .ZN(\SUMB[8][10] ) );
  INV_X2 U2762 ( .A(net120922), .ZN(net123843) );
  NAND2_X4 U2763 ( .A1(\SUMB[8][10] ), .A2(\ab[9][9] ), .ZN(n1620) );
  NAND2_X4 U2764 ( .A1(\SUMB[8][10] ), .A2(\CARRYB[8][9] ), .ZN(n1619) );
  NAND2_X2 U2765 ( .A1(net124104), .A2(n1679), .ZN(n1318) );
  NAND2_X2 U2766 ( .A1(n1504), .A2(\SUMB[1][13] ), .ZN(n886) );
  INV_X4 U2767 ( .A(n1679), .ZN(n1317) );
  NAND2_X2 U2768 ( .A1(\SUMB[13][8] ), .A2(\CARRYB[13][7] ), .ZN(net84998) );
  NAND2_X4 U2769 ( .A1(\ab[3][11] ), .A2(\SUMB[2][12] ), .ZN(n2029) );
  NAND2_X2 U2770 ( .A1(\ab[3][11] ), .A2(\CARRYB[2][11] ), .ZN(n2030) );
  NAND2_X2 U2771 ( .A1(n875), .A2(n876), .ZN(n878) );
  INV_X1 U2773 ( .A(\ab[7][22] ), .ZN(n875) );
  NAND2_X1 U2774 ( .A1(n1606), .A2(\SUMB[18][12] ), .ZN(n881) );
  NAND2_X2 U2775 ( .A1(n879), .A2(n880), .ZN(n882) );
  NAND2_X4 U2776 ( .A1(n881), .A2(n882), .ZN(\SUMB[19][11] ) );
  INV_X4 U2777 ( .A(n1606), .ZN(n879) );
  INV_X1 U2778 ( .A(\SUMB[18][12] ), .ZN(n880) );
  NAND2_X2 U2779 ( .A1(net86864), .A2(net93243), .ZN(n883) );
  NAND2_X4 U2780 ( .A1(net123592), .A2(net123591), .ZN(n884) );
  NAND2_X4 U2781 ( .A1(n883), .A2(n884), .ZN(\SUMB[2][14] ) );
  INV_X4 U2782 ( .A(net93243), .ZN(net123591) );
  INV_X4 U2783 ( .A(net86864), .ZN(net123592) );
  XNOR2_X2 U2784 ( .A(n2303), .B(net88703), .ZN(\SUMB[9][16] ) );
  INV_X4 U2785 ( .A(net88703), .ZN(net88704) );
  XNOR2_X2 U2786 ( .A(\CARRYB[6][6] ), .B(\ab[7][6] ), .ZN(n1309) );
  NAND2_X2 U2787 ( .A1(\ab[15][6] ), .A2(\SUMB[14][7] ), .ZN(n1437) );
  NAND2_X2 U2788 ( .A1(\CARRYB[2][4] ), .A2(\SUMB[2][5] ), .ZN(n1147) );
  NOR2_X4 U2789 ( .A1(net124610), .A2(net70486), .ZN(\ab[0][26] ) );
  NAND3_X2 U2790 ( .A1(net82664), .A2(net82665), .A3(net82666), .ZN(
        \CARRYB[18][11] ) );
  INV_X4 U2791 ( .A(net80517), .ZN(net86407) );
  NAND3_X2 U2792 ( .A1(net80803), .A2(net80802), .A3(net80801), .ZN(
        \CARRYB[9][17] ) );
  NAND2_X4 U2793 ( .A1(net80801), .A2(n928), .ZN(n925) );
  NAND3_X2 U2794 ( .A1(net81954), .A2(net81953), .A3(n935), .ZN(
        \CARRYB[19][9] ) );
  NAND2_X2 U2795 ( .A1(\CARRYB[1][12] ), .A2(\ab[2][12] ), .ZN(n2082) );
  NAND2_X4 U2796 ( .A1(n887), .A2(n886), .ZN(\SUMB[2][12] ) );
  INV_X1 U2797 ( .A(\ab[4][10] ), .ZN(n889) );
  NOR2_X1 U2798 ( .A1(net70482), .A2(net77956), .ZN(\ab[4][24] ) );
  NOR2_X1 U2799 ( .A1(net70482), .A2(net77948), .ZN(\ab[5][24] ) );
  NOR2_X1 U2800 ( .A1(net70482), .A2(net77940), .ZN(\ab[6][24] ) );
  NOR2_X1 U2801 ( .A1(net77930), .A2(net70482), .ZN(\ab[7][24] ) );
  NAND2_X1 U2802 ( .A1(\ab[1][23] ), .A2(\ab[0][24] ), .ZN(net82045) );
  NAND2_X1 U2803 ( .A1(\ab[6][24] ), .A2(\SUMB[5][25] ), .ZN(n905) );
  NAND2_X2 U2804 ( .A1(\ab[4][17] ), .A2(n861), .ZN(n1893) );
  NAND2_X2 U2805 ( .A1(\ab[6][20] ), .A2(\SUMB[5][21] ), .ZN(net79936) );
  NAND3_X2 U2806 ( .A1(n1466), .A2(n1467), .A3(n1468), .ZN(\CARRYB[12][17] )
         );
  INV_X2 U2807 ( .A(\SUMB[12][18] ), .ZN(n993) );
  XOR2_X2 U2808 ( .A(\CARRYB[16][12] ), .B(\ab[17][12] ), .Z(n891) );
  XOR2_X2 U2809 ( .A(\SUMB[16][13] ), .B(n891), .Z(\SUMB[17][12] ) );
  NAND2_X1 U2810 ( .A1(\ab[17][12] ), .A2(\CARRYB[16][12] ), .ZN(n894) );
  NAND3_X4 U2812 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(\CARRYB[16][12] )
         );
  INV_X2 U2813 ( .A(\ab[1][11] ), .ZN(n1023) );
  CLKBUF_X3 U2814 ( .A(\CARRYB[3][20] ), .Z(n1009) );
  INV_X4 U2815 ( .A(net88449), .ZN(net123428) );
  NAND2_X4 U2816 ( .A1(\SUMB[1][13] ), .A2(n588), .ZN(n2081) );
  XNOR2_X2 U2817 ( .A(\ab[21][1] ), .B(\SUMB[20][2] ), .ZN(n1266) );
  INV_X2 U2818 ( .A(\SUMB[4][14] ), .ZN(n1356) );
  NAND2_X4 U2819 ( .A1(n1346), .A2(n1347), .ZN(n1349) );
  NAND2_X4 U2820 ( .A1(n1290), .A2(n1291), .ZN(n1773) );
  NAND2_X4 U2821 ( .A1(n2155), .A2(\ab[24][5] ), .ZN(n2157) );
  XNOR2_X2 U2822 ( .A(\CARRYB[17][10] ), .B(n897), .ZN(net87009) );
  XNOR2_X2 U2823 ( .A(n898), .B(\SUMB[12][16] ), .ZN(\SUMB[13][15] ) );
  XNOR2_X2 U2824 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .ZN(n898) );
  INV_X8 U2825 ( .A(\CARRYB[1][12] ), .ZN(n1044) );
  XOR2_X2 U2826 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .Z(n899) );
  XOR2_X2 U2827 ( .A(n899), .B(n908), .Z(\SUMB[5][25] ) );
  XOR2_X2 U2828 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .Z(n900) );
  XOR2_X2 U2829 ( .A(n900), .B(\SUMB[5][25] ), .Z(\SUMB[6][24] ) );
  NAND2_X1 U2830 ( .A1(\ab[5][25] ), .A2(\CARRYB[4][25] ), .ZN(n901) );
  NAND2_X2 U2831 ( .A1(\ab[5][25] ), .A2(n908), .ZN(n902) );
  NAND2_X2 U2832 ( .A1(\CARRYB[4][25] ), .A2(n908), .ZN(n903) );
  NAND3_X4 U2833 ( .A1(n901), .A2(n902), .A3(n903), .ZN(\CARRYB[5][25] ) );
  NAND2_X1 U2834 ( .A1(\ab[6][24] ), .A2(\CARRYB[5][24] ), .ZN(n904) );
  NAND2_X1 U2835 ( .A1(\CARRYB[5][24] ), .A2(\SUMB[5][25] ), .ZN(n906) );
  NAND3_X4 U2836 ( .A1(n904), .A2(n905), .A3(n906), .ZN(\CARRYB[6][24] ) );
  INV_X2 U2837 ( .A(\SUMB[4][26] ), .ZN(n907) );
  INV_X8 U2838 ( .A(n907), .ZN(n908) );
  NAND2_X4 U2839 ( .A1(n911), .A2(n912), .ZN(\SUMB[4][13] ) );
  NAND2_X4 U2840 ( .A1(n1417), .A2(n1418), .ZN(net82089) );
  NAND2_X4 U2841 ( .A1(\ab[0][12] ), .A2(\ab[1][11] ), .ZN(n2334) );
  NAND2_X2 U2842 ( .A1(\CARRYB[2][11] ), .A2(\ab[3][11] ), .ZN(n915) );
  NAND2_X4 U2843 ( .A1(n913), .A2(n914), .ZN(n916) );
  INV_X2 U2844 ( .A(\ab[3][11] ), .ZN(n914) );
  NAND2_X4 U2845 ( .A1(n2374), .A2(\ab[6][10] ), .ZN(n1590) );
  NAND2_X2 U2846 ( .A1(\ab[1][20] ), .A2(\ab[0][21] ), .ZN(n2341) );
  NAND2_X4 U2847 ( .A1(n1162), .A2(n1161), .ZN(n1942) );
  INV_X8 U2848 ( .A(net81815), .ZN(net84303) );
  XNOR2_X2 U2849 ( .A(\CARRYB[22][2] ), .B(\ab[23][2] ), .ZN(net121523) );
  NAND2_X4 U2850 ( .A1(\CARRYB[4][12] ), .A2(\ab[5][12] ), .ZN(net81204) );
  INV_X4 U2851 ( .A(\CARRYB[2][18] ), .ZN(n1547) );
  OAI21_X4 U2852 ( .B1(n918), .B2(net123019), .A(n919), .ZN(n917) );
  NAND2_X2 U2853 ( .A1(n917), .A2(net123028), .ZN(net80801) );
  NAND2_X2 U2854 ( .A1(n917), .A2(n920), .ZN(net80803) );
  NAND2_X2 U2855 ( .A1(n920), .A2(net123028), .ZN(net80802) );
  NAND2_X2 U2856 ( .A1(n921), .A2(\ab[10][16] ), .ZN(net80805) );
  NAND2_X2 U2857 ( .A1(n921), .A2(\CARRYB[9][16] ), .ZN(net80806) );
  XNOR2_X2 U2858 ( .A(net80366), .B(\SUMB[6][19] ), .ZN(n922) );
  XNOR2_X2 U2859 ( .A(\SUMB[7][19] ), .B(net79939), .ZN(n923) );
  XNOR2_X2 U2860 ( .A(n923), .B(n925), .ZN(n924) );
  INV_X4 U2861 ( .A(net123019), .ZN(net123062) );
  OAI21_X4 U2862 ( .B1(n929), .B2(net123062), .A(\CARRYB[7][17] ), .ZN(n919)
         );
  INV_X4 U2863 ( .A(net123055), .ZN(net123028) );
  INV_X4 U2864 ( .A(n923), .ZN(n920) );
  INV_X4 U2865 ( .A(n924), .ZN(n921) );
  XNOR2_X2 U2866 ( .A(n922), .B(net123019), .ZN(n926) );
  INV_X2 U2867 ( .A(net123072), .ZN(net82890) );
  CLKBUF_X3 U2868 ( .A(n922), .Z(n929) );
  XNOR2_X2 U2869 ( .A(n921), .B(net81945), .ZN(\SUMB[10][16] ) );
  NAND3_X2 U2870 ( .A1(n931), .A2(n932), .A3(n930), .ZN(\CARRYB[7][17] ) );
  NAND2_X1 U2871 ( .A1(\ab[7][17] ), .A2(\CARRYB[6][17] ), .ZN(n930) );
  NAND2_X2 U2872 ( .A1(\ab[7][17] ), .A2(net90702), .ZN(n931) );
  INV_X4 U2873 ( .A(\CARRYB[6][18] ), .ZN(net80658) );
  INV_X1 U2874 ( .A(\ab[7][18] ), .ZN(net80657) );
  XNOR2_X2 U2875 ( .A(net86557), .B(\SUMB[5][20] ), .ZN(\SUMB[6][19] ) );
  XNOR2_X2 U2876 ( .A(net82396), .B(\SUMB[19][10] ), .ZN(\SUMB[20][9] ) );
  NAND2_X2 U2877 ( .A1(net86403), .A2(net86404), .ZN(n937) );
  INV_X4 U2878 ( .A(\CARRYB[19][9] ), .ZN(net86404) );
  INV_X1 U2879 ( .A(\ab[20][9] ), .ZN(net86403) );
  XNOR2_X2 U2880 ( .A(\SUMB[18][11] ), .B(n934), .ZN(\SUMB[19][10] ) );
  NAND2_X1 U2881 ( .A1(\ab[20][9] ), .A2(\SUMB[19][10] ), .ZN(net81034) );
  XNOR2_X2 U2882 ( .A(\CARRYB[18][10] ), .B(\ab[19][10] ), .ZN(n934) );
  BUF_X8 U2883 ( .A(\CARRYB[19][9] ), .Z(net82255) );
  NAND2_X2 U2884 ( .A1(n936), .A2(\ab[19][9] ), .ZN(net81953) );
  XNOR2_X2 U2885 ( .A(net85979), .B(n936), .ZN(\SUMB[19][9] ) );
  XNOR2_X2 U2886 ( .A(net85979), .B(n936), .ZN(net89289) );
  NAND2_X2 U2887 ( .A1(net90802), .A2(n936), .ZN(net81954) );
  INV_X1 U2888 ( .A(net87134), .ZN(net90802) );
  INV_X4 U2889 ( .A(\CARRYB[18][9] ), .ZN(net87134) );
  NAND2_X4 U2890 ( .A1(net87133), .A2(net87134), .ZN(net87136) );
  NOR2_X1 U2891 ( .A1(net70452), .A2(net70455), .ZN(\ab[20][9] ) );
  NAND2_X4 U2892 ( .A1(\SUMB[23][6] ), .A2(n2148), .ZN(n1121) );
  XNOR2_X2 U2893 ( .A(n1820), .B(n1264), .ZN(n938) );
  XNOR2_X2 U2894 ( .A(n1820), .B(n1264), .ZN(n939) );
  NAND3_X2 U2895 ( .A1(n1822), .A2(n1823), .A3(n1824), .ZN(\CARRYB[7][7] ) );
  XNOR2_X2 U2896 ( .A(net124874), .B(\SUMB[24][2] ), .ZN(n940) );
  INV_X4 U2897 ( .A(\CARRYB[17][5] ), .ZN(n1005) );
  NAND2_X2 U2898 ( .A1(n682), .A2(n390), .ZN(n1579) );
  NAND2_X1 U2899 ( .A1(\ab[15][0] ), .A2(\SUMB[14][1] ), .ZN(n1411) );
  CLKBUF_X2 U2900 ( .A(\SUMB[8][5] ), .Z(net121926) );
  XNOR2_X2 U2901 ( .A(n942), .B(\SUMB[13][4] ), .ZN(\SUMB[14][3] ) );
  NAND3_X2 U2902 ( .A1(n1962), .A2(n1961), .A3(n1963), .ZN(n943) );
  NOR2_X2 U2903 ( .A1(net84698), .A2(net77964), .ZN(\ab[3][14] ) );
  INV_X4 U2904 ( .A(\ab[4][14] ), .ZN(net92716) );
  XNOR2_X2 U2905 ( .A(\CARRYB[20][4] ), .B(n945), .ZN(n944) );
  INV_X4 U2906 ( .A(n66), .ZN(n1341) );
  NAND3_X4 U2907 ( .A1(n2117), .A2(net81060), .A3(net81059), .ZN(net85043) );
  INV_X2 U2908 ( .A(\SUMB[3][9] ), .ZN(n947) );
  XNOR2_X2 U2909 ( .A(n856), .B(n1095), .ZN(n949) );
  XNOR2_X2 U2910 ( .A(n2362), .B(n1325), .ZN(n950) );
  NAND2_X2 U2911 ( .A1(\ab[16][5] ), .A2(\SUMB[15][6] ), .ZN(n2072) );
  XOR2_X2 U2912 ( .A(\CARRYB[17][13] ), .B(\ab[18][13] ), .Z(n951) );
  NOR2_X2 U2913 ( .A1(net82890), .A2(net77956), .ZN(\ab[4][17] ) );
  XNOR2_X2 U2914 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .ZN(n952) );
  INV_X4 U2915 ( .A(\ab[16][8] ), .ZN(n2153) );
  NAND2_X1 U2916 ( .A1(n1187), .A2(\CARRYB[15][11] ), .ZN(n2098) );
  NAND2_X1 U2917 ( .A1(\CARRYB[3][18] ), .A2(\SUMB[3][19] ), .ZN(n1722) );
  NAND2_X2 U2918 ( .A1(\ab[6][13] ), .A2(\CARRYB[5][13] ), .ZN(n1161) );
  NAND2_X2 U2919 ( .A1(net83736), .A2(net125375), .ZN(n953) );
  NAND2_X4 U2920 ( .A1(net121606), .A2(net121607), .ZN(n954) );
  NAND2_X4 U2921 ( .A1(n953), .A2(n954), .ZN(\SUMB[9][10] ) );
  INV_X4 U2922 ( .A(net125375), .ZN(net121607) );
  XNOR2_X2 U2923 ( .A(n1742), .B(n852), .ZN(n1242) );
  INV_X8 U2924 ( .A(\CARRYB[14][12] ), .ZN(n1850) );
  NAND2_X4 U2925 ( .A1(\SUMB[1][20] ), .A2(\CARRYB[1][19] ), .ZN(n2143) );
  NAND2_X2 U2926 ( .A1(\CARRYB[3][9] ), .A2(\ab[4][9] ), .ZN(n1961) );
  BUF_X8 U2927 ( .A(\CARRYB[12][7] ), .Z(n1588) );
  NAND2_X2 U2928 ( .A1(\CARRYB[12][7] ), .A2(\ab[13][7] ), .ZN(n2023) );
  NAND2_X2 U2929 ( .A1(\ab[18][0] ), .A2(\SUMB[17][1] ), .ZN(n1810) );
  NAND2_X4 U2930 ( .A1(\ab[18][5] ), .A2(n1719), .ZN(n2231) );
  NAND2_X2 U2931 ( .A1(\SUMB[23][1] ), .A2(\ab[24][0] ), .ZN(n1570) );
  INV_X2 U2932 ( .A(net70476), .ZN(n1118) );
  INV_X8 U2933 ( .A(B[21]), .ZN(net70476) );
  NAND2_X4 U2934 ( .A1(net121453), .A2(net121454), .ZN(n956) );
  NAND2_X4 U2935 ( .A1(net121455), .A2(n956), .ZN(net90731) );
  NAND2_X1 U2936 ( .A1(\CARRYB[4][21] ), .A2(\ab[5][21] ), .ZN(n959) );
  NAND2_X2 U2937 ( .A1(n959), .A2(n960), .ZN(n1435) );
  INV_X4 U2938 ( .A(\CARRYB[4][21] ), .ZN(n957) );
  INV_X2 U2939 ( .A(\ab[5][21] ), .ZN(n958) );
  XOR2_X2 U2940 ( .A(\CARRYB[16][12] ), .B(\ab[17][12] ), .Z(n961) );
  XOR2_X2 U2941 ( .A(net90103), .B(n961), .Z(net88647) );
  NOR2_X2 U2942 ( .A1(net80643), .A2(net77948), .ZN(\ab[5][21] ) );
  NAND2_X2 U2943 ( .A1(\ab[14][14] ), .A2(\SUMB[13][15] ), .ZN(net80479) );
  XNOR2_X1 U2944 ( .A(net90525), .B(net81290), .ZN(net90103) );
  NOR2_X2 U2945 ( .A1(net83784), .A2(net70461), .ZN(\ab[17][12] ) );
  NAND2_X1 U2946 ( .A1(\ab[18][11] ), .A2(net88647), .ZN(net82665) );
  NAND3_X4 U2947 ( .A1(net80255), .A2(net80254), .A3(n2295), .ZN(
        \CARRYB[23][2] ) );
  XOR2_X2 U2948 ( .A(\CARRYB[6][1] ), .B(\ab[7][1] ), .Z(n964) );
  XOR2_X1 U2949 ( .A(\SUMB[6][2] ), .B(n964), .Z(\SUMB[7][1] ) );
  NAND2_X2 U2950 ( .A1(\CARRYB[6][1] ), .A2(\SUMB[6][2] ), .ZN(n965) );
  NAND2_X2 U2951 ( .A1(\ab[7][1] ), .A2(\SUMB[6][2] ), .ZN(n966) );
  NAND2_X1 U2952 ( .A1(\ab[7][1] ), .A2(\CARRYB[6][1] ), .ZN(n967) );
  NAND3_X2 U2953 ( .A1(n965), .A2(n966), .A3(n967), .ZN(\CARRYB[7][1] ) );
  XOR2_X2 U2954 ( .A(\CARRYB[7][1] ), .B(\ab[8][1] ), .Z(n968) );
  XOR2_X2 U2955 ( .A(\SUMB[7][2] ), .B(n968), .Z(\SUMB[8][1] ) );
  NAND2_X1 U2956 ( .A1(\CARRYB[7][1] ), .A2(\SUMB[7][2] ), .ZN(n969) );
  NAND2_X2 U2957 ( .A1(\ab[8][1] ), .A2(\SUMB[7][2] ), .ZN(n970) );
  NAND2_X1 U2958 ( .A1(\ab[8][1] ), .A2(\CARRYB[7][1] ), .ZN(n971) );
  NAND3_X2 U2959 ( .A1(n969), .A2(n970), .A3(n971), .ZN(\CARRYB[8][1] ) );
  NOR2_X1 U2960 ( .A1(net77866), .A2(net77930), .ZN(\ab[7][1] ) );
  NOR2_X1 U2961 ( .A1(net77866), .A2(net77924), .ZN(\ab[8][1] ) );
  NAND2_X4 U2962 ( .A1(n1045), .A2(n1046), .ZN(n1504) );
  NAND2_X4 U2963 ( .A1(net120174), .A2(n1044), .ZN(n1046) );
  NAND2_X2 U2964 ( .A1(n1261), .A2(\CARRYB[8][7] ), .ZN(n2016) );
  NAND2_X4 U2965 ( .A1(net88156), .A2(net88157), .ZN(n1321) );
  NAND2_X4 U2966 ( .A1(n1180), .A2(n1179), .ZN(n2015) );
  NAND2_X4 U2967 ( .A1(n1177), .A2(n1178), .ZN(n1180) );
  INV_X4 U2968 ( .A(\ab[2][12] ), .ZN(net120174) );
  NAND2_X2 U2969 ( .A1(n67), .A2(\SUMB[6][10] ), .ZN(n2003) );
  INV_X2 U2970 ( .A(\SUMB[6][10] ), .ZN(n1263) );
  CLKBUF_X3 U2971 ( .A(\SUMB[5][16] ), .Z(n1119) );
  NAND2_X4 U2972 ( .A1(\SUMB[12][8] ), .A2(\ab[13][7] ), .ZN(n2022) );
  NAND2_X2 U2973 ( .A1(\SUMB[11][4] ), .A2(\ab[12][3] ), .ZN(n1673) );
  NAND2_X4 U2974 ( .A1(net84304), .A2(net84303), .ZN(n1622) );
  NAND2_X2 U2975 ( .A1(n1720), .A2(\SUMB[3][15] ), .ZN(n975) );
  NAND2_X4 U2976 ( .A1(n973), .A2(n974), .ZN(n976) );
  NAND2_X4 U2977 ( .A1(n976), .A2(n975), .ZN(\SUMB[4][14] ) );
  INV_X4 U2978 ( .A(n1720), .ZN(n973) );
  INV_X4 U2979 ( .A(\SUMB[3][15] ), .ZN(n974) );
  INV_X8 U2980 ( .A(\CARRYB[5][13] ), .ZN(n1160) );
  NAND2_X1 U2981 ( .A1(\ab[10][3] ), .A2(\SUMB[9][4] ), .ZN(n1802) );
  NAND2_X4 U2982 ( .A1(net93308), .A2(net93309), .ZN(n1125) );
  NAND3_X4 U2983 ( .A1(n2253), .A2(n2254), .A3(n2252), .ZN(\CARRYB[8][15] ) );
  NAND2_X2 U2984 ( .A1(n977), .A2(n978), .ZN(n980) );
  INV_X4 U2985 ( .A(\CARRYB[5][19] ), .ZN(n977) );
  INV_X1 U2986 ( .A(\ab[6][19] ), .ZN(n978) );
  NOR2_X4 U2987 ( .A1(net86565), .A2(net77940), .ZN(\ab[6][19] ) );
  INV_X2 U2988 ( .A(net123291), .ZN(net121150) );
  NAND2_X4 U2989 ( .A1(net85540), .A2(net88934), .ZN(net85543) );
  NAND2_X2 U2990 ( .A1(\CARRYB[9][14] ), .A2(\ab[10][14] ), .ZN(n1039) );
  NAND2_X4 U2991 ( .A1(n1168), .A2(n1169), .ZN(n1171) );
  NAND3_X2 U2992 ( .A1(n2019), .A2(n2020), .A3(n2021), .ZN(\CARRYB[12][7] ) );
  NOR2_X2 U2993 ( .A1(net86565), .A2(net70491), .ZN(\ab[2][19] ) );
  NAND2_X2 U2994 ( .A1(\SUMB[15][9] ), .A2(\ab[16][8] ), .ZN(n2300) );
  NAND2_X1 U2995 ( .A1(\SUMB[2][22] ), .A2(\CARRYB[2][21] ), .ZN(n1935) );
  NAND2_X2 U2996 ( .A1(n1186), .A2(\ab[3][14] ), .ZN(n1987) );
  NAND3_X2 U2997 ( .A1(n1883), .A2(n1884), .A3(n1885), .ZN(\CARRYB[5][20] ) );
  NAND2_X2 U2998 ( .A1(n57), .A2(n1692), .ZN(n983) );
  NAND2_X4 U2999 ( .A1(n981), .A2(n982), .ZN(n984) );
  NAND2_X4 U3000 ( .A1(n983), .A2(n984), .ZN(\SUMB[2][21] ) );
  INV_X4 U3001 ( .A(n1828), .ZN(n981) );
  INV_X4 U3002 ( .A(n1692), .ZN(n982) );
  INV_X2 U3003 ( .A(\SUMB[2][21] ), .ZN(n1432) );
  XNOR2_X2 U3004 ( .A(n985), .B(\CARRYB[11][3] ), .ZN(\SUMB[12][3] ) );
  NAND2_X2 U3005 ( .A1(\CARRYB[11][2] ), .A2(\SUMB[11][3] ), .ZN(n1995) );
  NAND2_X1 U3006 ( .A1(\CARRYB[6][21] ), .A2(\SUMB[6][22] ), .ZN(n986) );
  NAND2_X1 U3007 ( .A1(\ab[7][21] ), .A2(\CARRYB[6][21] ), .ZN(n988) );
  NAND3_X2 U3008 ( .A1(n986), .A2(n987), .A3(n988), .ZN(\CARRYB[7][21] ) );
  NAND2_X2 U3009 ( .A1(n1088), .A2(n1089), .ZN(n991) );
  NAND2_X4 U3010 ( .A1(n989), .A2(n990), .ZN(n992) );
  NAND2_X4 U3011 ( .A1(n991), .A2(n992), .ZN(\SUMB[4][23] ) );
  INV_X4 U3012 ( .A(n1088), .ZN(n989) );
  INV_X4 U3013 ( .A(n1089), .ZN(n990) );
  NAND2_X2 U3014 ( .A1(\SUMB[12][18] ), .A2(n1571), .ZN(n994) );
  NAND2_X4 U3015 ( .A1(n993), .A2(n860), .ZN(n995) );
  NAND2_X4 U3016 ( .A1(n994), .A2(n995), .ZN(\SUMB[13][17] ) );
  XNOR2_X1 U3017 ( .A(\ab[13][17] ), .B(\CARRYB[12][17] ), .ZN(n1571) );
  XNOR2_X2 U3018 ( .A(\SUMB[22][9] ), .B(n1273), .ZN(\SUMB[23][8] ) );
  XOR2_X2 U3019 ( .A(\CARRYB[9][6] ), .B(\ab[10][6] ), .Z(n996) );
  NAND2_X1 U3020 ( .A1(\CARRYB[9][6] ), .A2(\SUMB[9][7] ), .ZN(n997) );
  NAND2_X2 U3021 ( .A1(\ab[10][6] ), .A2(\SUMB[9][7] ), .ZN(n998) );
  NAND2_X1 U3022 ( .A1(\ab[10][6] ), .A2(\CARRYB[9][6] ), .ZN(n999) );
  NAND3_X2 U3023 ( .A1(n997), .A2(n998), .A3(n999), .ZN(\CARRYB[10][6] ) );
  NAND2_X2 U3024 ( .A1(n1214), .A2(n1994), .ZN(n1002) );
  NAND2_X4 U3025 ( .A1(n1000), .A2(n1001), .ZN(n1003) );
  NAND2_X4 U3026 ( .A1(n1002), .A2(n1003), .ZN(\SUMB[6][8] ) );
  INV_X4 U3027 ( .A(n1214), .ZN(n1000) );
  NAND3_X4 U3028 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(\CARRYB[9][6] ) );
  NOR2_X1 U3029 ( .A1(net77906), .A2(net70475), .ZN(\ab[10][6] ) );
  INV_X8 U3030 ( .A(net84357), .ZN(net84358) );
  INV_X4 U3031 ( .A(\SUMB[24][6] ), .ZN(net84304) );
  NAND2_X2 U3032 ( .A1(n849), .A2(n215), .ZN(n1387) );
  NAND3_X4 U3033 ( .A1(n1793), .A2(n1794), .A3(n1795), .ZN(\CARRYB[12][13] )
         );
  INV_X2 U3034 ( .A(\CARRYB[8][18] ), .ZN(n1050) );
  CLKBUF_X3 U3035 ( .A(n854), .Z(n1379) );
  NAND3_X2 U3036 ( .A1(n1398), .A2(n1397), .A3(n1396), .ZN(\CARRYB[5][9] ) );
  NAND3_X4 U3037 ( .A1(n1676), .A2(n1677), .A3(n1678), .ZN(\CARRYB[13][3] ) );
  NAND2_X4 U3038 ( .A1(net120628), .A2(net120627), .ZN(net83202) );
  INV_X4 U3039 ( .A(n1005), .ZN(n1719) );
  NOR2_X1 U3040 ( .A1(net70452), .A2(net70467), .ZN(\ab[14][9] ) );
  NOR2_X1 U3041 ( .A1(net70452), .A2(net70469), .ZN(\ab[13][9] ) );
  XNOR2_X2 U3042 ( .A(\ab[2][20] ), .B(\CARRYB[1][20] ), .ZN(n1424) );
  NAND3_X4 U3043 ( .A1(net119921), .A2(net119920), .A3(n209), .ZN(net82031) );
  XNOR2_X2 U3044 ( .A(\ab[2][20] ), .B(n2341), .ZN(n1004) );
  NAND2_X1 U3045 ( .A1(\CARRYB[9][18] ), .A2(\SUMB[9][19] ), .ZN(n1876) );
  NAND2_X1 U3046 ( .A1(\ab[5][21] ), .A2(\CARRYB[4][21] ), .ZN(n1117) );
  NAND2_X1 U3047 ( .A1(\CARRYB[17][5] ), .A2(\ab[18][5] ), .ZN(n1007) );
  NAND2_X2 U3048 ( .A1(n1005), .A2(n1006), .ZN(n1008) );
  NAND2_X2 U3049 ( .A1(n1007), .A2(n1008), .ZN(n1718) );
  INV_X1 U3050 ( .A(\ab[18][5] ), .ZN(n1006) );
  INV_X4 U3051 ( .A(n2339), .ZN(\CARRYB[1][19] ) );
  NAND2_X2 U3052 ( .A1(\ab[1][19] ), .A2(\ab[0][20] ), .ZN(n2339) );
  NAND2_X2 U3053 ( .A1(\ab[20][4] ), .A2(\CARRYB[19][4] ), .ZN(n2228) );
  INV_X4 U3054 ( .A(n1426), .ZN(n1427) );
  XNOR2_X2 U3055 ( .A(n1010), .B(\CARRYB[14][3] ), .ZN(\SUMB[15][3] ) );
  NAND2_X2 U3057 ( .A1(\ab[10][3] ), .A2(\CARRYB[9][3] ), .ZN(n1803) );
  NAND3_X4 U3058 ( .A1(n1060), .A2(n1061), .A3(n1059), .ZN(\CARRYB[14][13] )
         );
  NAND2_X2 U3059 ( .A1(net120651), .A2(net120652), .ZN(n1011) );
  INV_X2 U3060 ( .A(net80983), .ZN(net120651) );
  NAND2_X2 U3061 ( .A1(\CARRYB[1][5] ), .A2(\SUMB[1][6] ), .ZN(n1866) );
  NOR2_X2 U3062 ( .A1(net70470), .A2(net77964), .ZN(\ab[3][18] ) );
  NAND2_X4 U3063 ( .A1(n1012), .A2(n1013), .ZN(n1014) );
  NAND2_X4 U3064 ( .A1(n1014), .A2(n2143), .ZN(n1927) );
  INV_X2 U3065 ( .A(\CARRYB[1][19] ), .ZN(n1013) );
  NAND2_X2 U3066 ( .A1(n1927), .A2(\ab[2][19] ), .ZN(n1526) );
  NAND2_X1 U3067 ( .A1(\ab[10][17] ), .A2(n1016), .ZN(n1017) );
  NAND2_X1 U3068 ( .A1(n1015), .A2(\CARRYB[9][17] ), .ZN(n1018) );
  NAND2_X2 U3069 ( .A1(n1017), .A2(n1018), .ZN(net88226) );
  INV_X1 U3070 ( .A(\ab[10][17] ), .ZN(n1015) );
  INV_X2 U3071 ( .A(\CARRYB[9][17] ), .ZN(n1016) );
  NAND2_X2 U3072 ( .A1(n1019), .A2(n1020), .ZN(net89026) );
  INV_X1 U3073 ( .A(\ab[12][12] ), .ZN(net120586) );
  NOR2_X2 U3074 ( .A1(net83784), .A2(net70471), .ZN(\ab[12][12] ) );
  NOR2_X2 U3075 ( .A1(net77914), .A2(net70459), .ZN(\ab[18][7] ) );
  NOR2_X2 U3076 ( .A1(net77914), .A2(net70461), .ZN(\ab[17][7] ) );
  NOR2_X2 U3077 ( .A1(net77914), .A2(net70453), .ZN(\ab[21][7] ) );
  NOR2_X2 U3078 ( .A1(net77912), .A2(net70473), .ZN(\ab[11][7] ) );
  NOR2_X2 U3079 ( .A1(net77912), .A2(net70475), .ZN(\ab[10][7] ) );
  NOR2_X2 U3080 ( .A1(net77912), .A2(net77956), .ZN(\ab[4][7] ) );
  NAND2_X2 U3081 ( .A1(\SUMB[13][8] ), .A2(\ab[14][7] ), .ZN(net84999) );
  NAND2_X2 U3082 ( .A1(\ab[17][7] ), .A2(\CARRYB[16][7] ), .ZN(net81265) );
  INV_X4 U3083 ( .A(\ab[6][7] ), .ZN(n1313) );
  NAND2_X2 U3084 ( .A1(\SUMB[8][8] ), .A2(\ab[9][7] ), .ZN(n2017) );
  INV_X4 U3085 ( .A(\ab[8][7] ), .ZN(n1831) );
  NAND2_X1 U3086 ( .A1(\ab[4][7] ), .A2(\CARRYB[3][7] ), .ZN(n1908) );
  NAND2_X4 U3087 ( .A1(net120513), .A2(net120514), .ZN(n1021) );
  NAND2_X4 U3088 ( .A1(n1021), .A2(net120515), .ZN(\SUMB[10][9] ) );
  NAND2_X4 U3089 ( .A1(net120517), .A2(net120518), .ZN(n1022) );
  NAND2_X4 U3090 ( .A1(net120519), .A2(n1022), .ZN(\SUMB[15][7] ) );
  BUF_X4 U3091 ( .A(\SUMB[10][9] ), .Z(net88928) );
  NAND2_X4 U3092 ( .A1(net86893), .A2(net86894), .ZN(net86896) );
  NOR2_X4 U3093 ( .A1(net70456), .A2(net80409), .ZN(\ab[1][11] ) );
  INV_X8 U3094 ( .A(n1780), .ZN(\SUMB[23][6] ) );
  NAND2_X2 U3095 ( .A1(\SUMB[10][15] ), .A2(\ab[11][14] ), .ZN(n1843) );
  NAND2_X4 U3096 ( .A1(n1846), .A2(n1847), .ZN(n1849) );
  INV_X4 U3097 ( .A(\SUMB[15][12] ), .ZN(n1847) );
  NAND2_X4 U3098 ( .A1(n1321), .A2(n1320), .ZN(net81756) );
  INV_X4 U3099 ( .A(\CARRYB[16][5] ), .ZN(n1380) );
  NAND2_X4 U3100 ( .A1(net120463), .A2(net120464), .ZN(net120466) );
  INV_X4 U3101 ( .A(\CARRYB[10][8] ), .ZN(net120463) );
  NAND2_X2 U3102 ( .A1(net88928), .A2(net86844), .ZN(n1027) );
  NAND2_X4 U3103 ( .A1(net120467), .A2(net120468), .ZN(n1028) );
  NAND2_X4 U3104 ( .A1(n1027), .A2(n1028), .ZN(\SUMB[11][8] ) );
  INV_X4 U3105 ( .A(net88928), .ZN(net120467) );
  NOR2_X4 U3106 ( .A1(net77920), .A2(net70473), .ZN(\ab[11][8] ) );
  XNOR2_X2 U3107 ( .A(net84883), .B(n838), .ZN(net90671) );
  NAND2_X2 U3108 ( .A1(\SUMB[9][5] ), .A2(\CARRYB[9][4] ), .ZN(n1926) );
  XNOR2_X2 U3109 ( .A(n2327), .B(\ab[2][4] ), .ZN(n1135) );
  INV_X2 U3110 ( .A(n2327), .ZN(\CARRYB[1][4] ) );
  NAND2_X4 U3111 ( .A1(n645), .A2(n1372), .ZN(n1374) );
  NAND3_X4 U3112 ( .A1(net82028), .A2(net82027), .A3(n1941), .ZN(
        \CARRYB[2][17] ) );
  NAND2_X2 U3113 ( .A1(n1694), .A2(\CARRYB[5][10] ), .ZN(n1170) );
  INV_X1 U3115 ( .A(\ab[5][10] ), .ZN(n1030) );
  NAND2_X1 U3116 ( .A1(\ab[7][15] ), .A2(\CARRYB[6][15] ), .ZN(n2208) );
  NAND2_X2 U3117 ( .A1(net120359), .A2(net93792), .ZN(n1034) );
  NAND2_X2 U3118 ( .A1(\SUMB[2][15] ), .A2(n1792), .ZN(n1558) );
  NAND2_X2 U3119 ( .A1(net84978), .A2(net84979), .ZN(n1035) );
  NAND2_X2 U3120 ( .A1(n170), .A2(n393), .ZN(n1036) );
  XNOR2_X2 U3121 ( .A(\CARRYB[10][3] ), .B(\ab[11][3] ), .ZN(n1200) );
  BUF_X8 U3122 ( .A(\CARRYB[26][3] ), .Z(n1272) );
  NAND2_X4 U3123 ( .A1(\CARRYB[14][5] ), .A2(n864), .ZN(n1979) );
  NAND2_X4 U3124 ( .A1(\CARRYB[8][11] ), .A2(\ab[9][11] ), .ZN(net86895) );
  NAND2_X4 U3125 ( .A1(n1037), .A2(n1038), .ZN(n1040) );
  NAND2_X4 U3126 ( .A1(n1041), .A2(n1042), .ZN(n1043) );
  NAND2_X4 U3127 ( .A1(n1795), .A2(n1043), .ZN(n1753) );
  INV_X1 U3128 ( .A(\ab[12][13] ), .ZN(n1042) );
  NOR2_X2 U3129 ( .A1(net70460), .A2(net70471), .ZN(\ab[12][13] ) );
  XOR2_X1 U3130 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .Z(n1315) );
  NAND2_X2 U3131 ( .A1(\ab[2][12] ), .A2(\CARRYB[1][12] ), .ZN(n1045) );
  NAND3_X4 U3132 ( .A1(net79935), .A2(net79936), .A3(net79937), .ZN(
        \CARRYB[6][20] ) );
  NAND2_X4 U3133 ( .A1(n1500), .A2(\ab[16][4] ), .ZN(n2105) );
  NAND2_X1 U3134 ( .A1(\ab[22][8] ), .A2(\SUMB[21][9] ), .ZN(net81179) );
  NAND2_X4 U3135 ( .A1(n1788), .A2(n1789), .ZN(n1791) );
  INV_X2 U3136 ( .A(n848), .ZN(n1789) );
  NAND2_X2 U3137 ( .A1(\CARRYB[11][14] ), .A2(\SUMB[11][15] ), .ZN(n1066) );
  NAND3_X2 U3138 ( .A1(n1568), .A2(n1569), .A3(n1570), .ZN(\CARRYB[24][0] ) );
  NAND2_X4 U3139 ( .A1(n2243), .A2(net83151), .ZN(n1757) );
  XNOR2_X2 U3140 ( .A(\CARRYB[17][3] ), .B(\ab[18][3] ), .ZN(n1268) );
  NAND2_X2 U3141 ( .A1(\ab[2][22] ), .A2(\CARRYB[1][22] ), .ZN(n1048) );
  NAND2_X2 U3142 ( .A1(n1047), .A2(n2345), .ZN(n1049) );
  NAND2_X2 U3143 ( .A1(n1048), .A2(n1049), .ZN(n1457) );
  INV_X2 U3144 ( .A(\ab[2][22] ), .ZN(n1047) );
  NAND2_X1 U3145 ( .A1(\CARRYB[8][18] ), .A2(n1051), .ZN(n1052) );
  NAND2_X1 U3146 ( .A1(n1050), .A2(\ab[9][18] ), .ZN(n1053) );
  NAND2_X2 U3147 ( .A1(n1052), .A2(n1053), .ZN(net79950) );
  INV_X1 U3148 ( .A(\ab[9][18] ), .ZN(n1051) );
  NAND2_X2 U3149 ( .A1(\ab[0][23] ), .A2(n2196), .ZN(n2345) );
  NAND2_X2 U3150 ( .A1(\ab[5][13] ), .A2(\CARRYB[4][13] ), .ZN(n1980) );
  NAND2_X4 U3151 ( .A1(\CARRYB[1][10] ), .A2(\SUMB[1][11] ), .ZN(n1654) );
  NAND2_X4 U3152 ( .A1(n1355), .A2(n1262), .ZN(n1358) );
  INV_X8 U3153 ( .A(n2338), .ZN(\SUMB[1][16] ) );
  NAND2_X4 U3154 ( .A1(n2192), .A2(n1740), .ZN(n1765) );
  NAND2_X4 U3155 ( .A1(n1738), .A2(n1739), .ZN(n1740) );
  NAND2_X4 U3156 ( .A1(n1603), .A2(net86601), .ZN(n1605) );
  NAND2_X2 U3157 ( .A1(\ab[4][21] ), .A2(\SUMB[3][22] ), .ZN(n2277) );
  NAND2_X4 U3158 ( .A1(net119979), .A2(n1054), .ZN(net119982) );
  INV_X4 U3159 ( .A(\CARRYB[11][9] ), .ZN(net119979) );
  NOR2_X4 U3160 ( .A1(n1111), .A2(net81673), .ZN(\ab[0][25] ) );
  XNOR2_X2 U3161 ( .A(net121859), .B(net149611), .ZN(net119817) );
  NAND2_X4 U3162 ( .A1(\SUMB[26][2] ), .A2(\CARRYB[26][1] ), .ZN(net80992) );
  XNOR2_X2 U3163 ( .A(\CARRYB[25][2] ), .B(net93792), .ZN(net93791) );
  XNOR2_X2 U3164 ( .A(\CARRYB[14][7] ), .B(\ab[15][7] ), .ZN(net83755) );
  NAND3_X2 U3165 ( .A1(net80257), .A2(n500), .A3(net80258), .ZN(net93840) );
  NAND2_X4 U3166 ( .A1(net86407), .A2(\SUMB[10][17] ), .ZN(n1055) );
  NAND2_X4 U3167 ( .A1(net86409), .A2(n1055), .ZN(\SUMB[11][16] ) );
  INV_X4 U3168 ( .A(net88225), .ZN(\SUMB[10][17] ) );
  NAND2_X1 U3169 ( .A1(\CARRYB[10][16] ), .A2(\SUMB[10][17] ), .ZN(net80523)
         );
  NAND2_X1 U3170 ( .A1(\ab[11][16] ), .A2(\SUMB[10][17] ), .ZN(net80522) );
  XNOR2_X2 U3171 ( .A(net88226), .B(\SUMB[9][18] ), .ZN(net88225) );
  NAND2_X2 U3172 ( .A1(net80517), .A2(net88225), .ZN(net86409) );
  XNOR2_X2 U3173 ( .A(\CARRYB[10][16] ), .B(net81394), .ZN(net80517) );
  INV_X4 U3174 ( .A(\ab[11][16] ), .ZN(net81394) );
  NAND2_X1 U3175 ( .A1(\ab[10][17] ), .A2(n573), .ZN(net80519) );
  NAND2_X1 U3176 ( .A1(\CARRYB[9][17] ), .A2(n573), .ZN(net80520) );
  NAND2_X1 U3177 ( .A1(\ab[10][17] ), .A2(\CARRYB[9][17] ), .ZN(net80518) );
  NAND2_X1 U3178 ( .A1(\ab[11][16] ), .A2(\CARRYB[10][16] ), .ZN(net80521) );
  NAND2_X2 U3179 ( .A1(net81285), .A2(net81284), .ZN(n1056) );
  NAND2_X2 U3180 ( .A1(net80794), .A2(n1056), .ZN(net80825) );
  INV_X1 U3181 ( .A(\ab[5][22] ), .ZN(net81284) );
  INV_X4 U3182 ( .A(\CARRYB[4][22] ), .ZN(net81285) );
  NOR2_X1 U3183 ( .A1(net70478), .A2(net77948), .ZN(\ab[5][22] ) );
  INV_X16 U3184 ( .A(B[22]), .ZN(net70478) );
  NAND2_X1 U3185 ( .A1(\CARRYB[4][22] ), .A2(\SUMB[4][23] ), .ZN(net80796) );
  NAND2_X1 U3186 ( .A1(\ab[4][22] ), .A2(\CARRYB[3][22] ), .ZN(n1057) );
  NAND2_X2 U3187 ( .A1(\CARRYB[3][22] ), .A2(\SUMB[3][23] ), .ZN(net84312) );
  XOR2_X2 U3188 ( .A(\CARRYB[3][22] ), .B(\ab[4][22] ), .Z(net84311) );
  XOR2_X2 U3189 ( .A(\SUMB[3][23] ), .B(net84311), .Z(\SUMB[4][22] ) );
  XNOR2_X2 U3190 ( .A(\CARRYB[13][14] ), .B(\ab[14][14] ), .ZN(net85119) );
  XNOR2_X2 U3191 ( .A(\CARRYB[14][13] ), .B(\ab[15][13] ), .ZN(net93107) );
  NAND2_X1 U3192 ( .A1(\ab[15][13] ), .A2(\CARRYB[14][13] ), .ZN(n1058) );
  NAND2_X1 U3193 ( .A1(\ab[14][13] ), .A2(\CARRYB[13][13] ), .ZN(n1059) );
  NAND2_X2 U3194 ( .A1(\SUMB[13][14] ), .A2(n695), .ZN(n1061) );
  NAND2_X1 U3195 ( .A1(\CARRYB[13][14] ), .A2(\SUMB[13][15] ), .ZN(net80478)
         );
  NAND2_X1 U3196 ( .A1(\ab[14][14] ), .A2(\CARRYB[13][14] ), .ZN(net80480) );
  XNOR2_X2 U3197 ( .A(net89094), .B(net80110), .ZN(net88916) );
  NAND2_X2 U3198 ( .A1(net81815), .A2(net88916), .ZN(net84305) );
  NAND3_X1 U3199 ( .A1(net79969), .A2(net79970), .A3(net79968), .ZN(net86696)
         );
  NAND2_X1 U3200 ( .A1(\ab[25][5] ), .A2(net86696), .ZN(n1062) );
  XNOR2_X2 U3201 ( .A(net80110), .B(\SUMB[23][7] ), .ZN(\SUMB[24][6] ) );
  NAND2_X1 U3202 ( .A1(\ab[24][6] ), .A2(net89094), .ZN(net79864) );
  NAND3_X2 U3203 ( .A1(net79969), .A2(net79968), .A3(net79970), .ZN(
        \CARRYB[24][5] ) );
  NAND3_X2 U3204 ( .A1(net82658), .A2(net82657), .A3(n1063), .ZN(
        \CARRYB[13][14] ) );
  NAND3_X4 U3205 ( .A1(n1066), .A2(n1065), .A3(n1064), .ZN(\CARRYB[12][14] )
         );
  XNOR2_X2 U3206 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .ZN(net84481) );
  NAND2_X1 U3207 ( .A1(\ab[13][14] ), .A2(\CARRYB[12][14] ), .ZN(n1063) );
  NAND2_X1 U3208 ( .A1(\ab[12][14] ), .A2(\CARRYB[11][14] ), .ZN(n1064) );
  NAND2_X2 U3209 ( .A1(\ab[12][14] ), .A2(\SUMB[11][15] ), .ZN(n1065) );
  FA_X1 U3210 ( .A(n111), .B(\ab[12][15] ), .CI(\SUMB[11][16] ), .S(net88756)
         );
  XNOR2_X2 U3211 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .ZN(n1067) );
  XNOR2_X2 U3212 ( .A(net80825), .B(\SUMB[4][23] ), .ZN(\SUMB[5][22] ) );
  NOR2_X1 U3213 ( .A1(net70478), .A2(net77956), .ZN(\ab[4][22] ) );
  NAND2_X2 U3214 ( .A1(\ab[3][22] ), .A2(\SUMB[2][23] ), .ZN(n1069) );
  XNOR2_X2 U3215 ( .A(net87855), .B(net90671), .ZN(\SUMB[3][23] ) );
  XNOR2_X2 U3216 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .ZN(net87855) );
  XNOR2_X2 U3217 ( .A(net84883), .B(\ab[2][24] ), .ZN(\SUMB[2][24] ) );
  NAND2_X1 U3218 ( .A1(n39), .A2(\ab[2][24] ), .ZN(net84299) );
  NAND2_X2 U3219 ( .A1(\SUMB[1][25] ), .A2(n838), .ZN(net84298) );
  NAND2_X1 U3220 ( .A1(\ab[3][23] ), .A2(\CARRYB[2][23] ), .ZN(net84300) );
  NAND2_X2 U3221 ( .A1(\SUMB[2][24] ), .A2(\ab[3][23] ), .ZN(net84301) );
  NOR2_X4 U3222 ( .A1(net77898), .A2(net70445), .ZN(\ab[25][5] ) );
  INV_X1 U3223 ( .A(\ab[25][5] ), .ZN(net86697) );
  NAND2_X2 U3224 ( .A1(\ab[25][5] ), .A2(\CARRYB[24][5] ), .ZN(net86699) );
  NAND2_X1 U3225 ( .A1(n262), .A2(\SUMB[23][7] ), .ZN(net79865) );
  NAND2_X2 U3226 ( .A1(\CARRYB[2][23] ), .A2(\SUMB[2][24] ), .ZN(net84302) );
  NAND3_X4 U3227 ( .A1(n1074), .A2(n1073), .A3(n1072), .ZN(\CARRYB[21][7] ) );
  NAND2_X1 U3228 ( .A1(\CARRYB[21][7] ), .A2(\ab[22][7] ), .ZN(n1071) );
  NAND2_X1 U3229 ( .A1(\ab[21][7] ), .A2(\CARRYB[20][7] ), .ZN(n1072) );
  NAND2_X2 U3230 ( .A1(\SUMB[20][8] ), .A2(\ab[21][7] ), .ZN(n1073) );
  NAND2_X2 U3231 ( .A1(\CARRYB[20][7] ), .A2(\SUMB[20][8] ), .ZN(n1074) );
  XNOR2_X2 U3234 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .ZN(net81113) );
  XNOR2_X2 U3235 ( .A(\CARRYB[20][7] ), .B(\ab[21][7] ), .ZN(net83134) );
  NAND2_X1 U3236 ( .A1(\ab[21][8] ), .A2(\CARRYB[20][8] ), .ZN(net81036) );
  XNOR2_X2 U3237 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .ZN(net90801) );
  NAND3_X2 U3238 ( .A1(net83575), .A2(n1077), .A3(net83576), .ZN(
        \CARRYB[2][23] ) );
  XNOR2_X2 U3239 ( .A(\ab[2][23] ), .B(net82124), .ZN(net88004) );
  NAND2_X1 U3240 ( .A1(\ab[2][23] ), .A2(net82124), .ZN(n1077) );
  NAND2_X2 U3241 ( .A1(net82043), .A2(net82044), .ZN(net82046) );
  INV_X4 U3242 ( .A(\ab[1][23] ), .ZN(net82043) );
  XOR2_X2 U3243 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Z(net83044) );
  XNOR2_X2 U3244 ( .A(net88004), .B(n2357), .ZN(\SUMB[2][23] ) );
  XNOR2_X2 U3245 ( .A(net86937), .B(net92319), .ZN(net92323) );
  XNOR2_X2 U3246 ( .A(\ab[31][0] ), .B(net92320), .ZN(net92319) );
  INV_X4 U3247 ( .A(A[31]), .ZN(n1078) );
  XNOR2_X2 U3248 ( .A(\SUMB[26][5] ), .B(net82807), .ZN(net86937) );
  XOR2_X2 U3249 ( .A(\CARRYB[26][4] ), .B(\ab[27][4] ), .Z(net82807) );
  NOR2_X1 U3250 ( .A1(net70441), .A2(net77892), .ZN(\ab[27][4] ) );
  NAND3_X2 U3251 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(\CARRYB[26][4] ) );
  NAND2_X1 U3252 ( .A1(\ab[26][4] ), .A2(n1082), .ZN(n1081) );
  BUF_X8 U3253 ( .A(\CARRYB[25][4] ), .Z(n1082) );
  NAND2_X1 U3254 ( .A1(n1082), .A2(\SUMB[25][5] ), .ZN(n1079) );
  NOR2_X1 U3255 ( .A1(net70443), .A2(net77898), .ZN(\ab[26][5] ) );
  XNOR2_X2 U3256 ( .A(\CARRYB[24][6] ), .B(net81946), .ZN(n1083) );
  OR2_X2 U3257 ( .A1(net70445), .A2(net77906), .ZN(net81946) );
  NAND3_X2 U3258 ( .A1(net79865), .A2(net79864), .A3(net79863), .ZN(
        \CARRYB[24][6] ) );
  XOR2_X2 U3259 ( .A(\CARRYB[23][7] ), .B(\ab[24][7] ), .Z(n1084) );
  NOR2_X1 U3260 ( .A1(net70447), .A2(net77912), .ZN(\ab[24][7] ) );
  NOR2_X2 U3261 ( .A1(net84358), .A2(net77964), .ZN(\ab[3][23] ) );
  INV_X2 U3262 ( .A(net70480), .ZN(net84357) );
  INV_X8 U3263 ( .A(B[23]), .ZN(net70480) );
  NOR2_X2 U3264 ( .A1(net70480), .A2(net86101), .ZN(\ab[1][23] ) );
  XNOR2_X2 U3265 ( .A(\ab[18][12] ), .B(\CARRYB[17][12] ), .ZN(net88165) );
  NAND2_X1 U3266 ( .A1(\CARRYB[17][12] ), .A2(\SUMB[17][13] ), .ZN(net80451)
         );
  NAND2_X1 U3267 ( .A1(\ab[18][12] ), .A2(\CARRYB[17][12] ), .ZN(net80449) );
  XNOR2_X2 U3268 ( .A(\SUMB[17][12] ), .B(net89353), .ZN(\SUMB[18][11] ) );
  XNOR2_X2 U3269 ( .A(\SUMB[15][14] ), .B(net81290), .ZN(\SUMB[16][13] ) );
  NAND2_X1 U3270 ( .A1(\ab[16][12] ), .A2(\CARRYB[15][12] ), .ZN(n1085) );
  XNOR2_X2 U3271 ( .A(\SUMB[14][15] ), .B(net86054), .ZN(\SUMB[15][14] ) );
  NAND2_X1 U3272 ( .A1(\ab[16][13] ), .A2(\SUMB[15][14] ), .ZN(net80274) );
  XNOR2_X2 U3273 ( .A(\CARRYB[15][13] ), .B(\ab[16][13] ), .ZN(net81290) );
  NAND2_X2 U3274 ( .A1(\ab[16][12] ), .A2(\CARRYB[15][12] ), .ZN(net87005) );
  XNOR2_X2 U3275 ( .A(net82641), .B(\SUMB[15][13] ), .ZN(\SUMB[16][12] ) );
  INV_X1 U3276 ( .A(\ab[16][12] ), .ZN(net87003) );
  NAND2_X1 U3277 ( .A1(\ab[15][14] ), .A2(\SUMB[14][15] ), .ZN(net84309) );
  NAND2_X1 U3278 ( .A1(\CARRYB[14][14] ), .A2(\SUMB[14][15] ), .ZN(net84308)
         );
  NAND2_X1 U3279 ( .A1(\CARRYB[15][13] ), .A2(net90525), .ZN(net80273) );
  NAND2_X1 U3280 ( .A1(\ab[16][13] ), .A2(\CARRYB[15][13] ), .ZN(net80275) );
  NOR2_X1 U3281 ( .A1(net84698), .A2(net70467), .ZN(\ab[14][14] ) );
  INV_X16 U3282 ( .A(B[24]), .ZN(net70482) );
  XNOR2_X2 U3283 ( .A(\CARRYB[3][23] ), .B(\ab[4][23] ), .ZN(n1088) );
  NAND2_X2 U3284 ( .A1(\ab[4][23] ), .A2(\SUMB[3][24] ), .ZN(net80793) );
  NAND2_X2 U3285 ( .A1(\CARRYB[3][23] ), .A2(\SUMB[3][24] ), .ZN(net80792) );
  NAND2_X2 U3286 ( .A1(\CARRYB[3][23] ), .A2(\ab[4][23] ), .ZN(net80791) );
  NAND2_X4 U3287 ( .A1(net83116), .A2(net83115), .ZN(n1090) );
  INV_X4 U3288 ( .A(\CARRYB[23][6] ), .ZN(net83116) );
  INV_X2 U3289 ( .A(\ab[24][6] ), .ZN(net83115) );
  XNOR2_X2 U3290 ( .A(n949), .B(n867), .ZN(net89094) );
  NAND2_X2 U3291 ( .A1(\ab[24][6] ), .A2(\CARRYB[23][6] ), .ZN(net79863) );
  XNOR2_X2 U3292 ( .A(\SUMB[22][8] ), .B(net88961), .ZN(\SUMB[23][7] ) );
  NAND2_X1 U3293 ( .A1(\SUMB[22][8] ), .A2(\CARRYB[22][7] ), .ZN(net86412) );
  NAND3_X2 U3294 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(\CARRYB[11][15] )
         );
  NAND2_X1 U3295 ( .A1(\ab[11][15] ), .A2(\CARRYB[10][15] ), .ZN(n1093) );
  NAND2_X2 U3296 ( .A1(\ab[11][15] ), .A2(\SUMB[10][16] ), .ZN(n1092) );
  NOR2_X2 U3297 ( .A1(net81424), .A2(net70471), .ZN(\ab[12][15] ) );
  XNOR2_X2 U3298 ( .A(\CARRYB[10][15] ), .B(\ab[11][15] ), .ZN(n1094) );
  NOR2_X1 U3299 ( .A1(net70460), .A2(net70465), .ZN(\ab[15][13] ) );
  NAND2_X1 U3300 ( .A1(\ab[23][7] ), .A2(\CARRYB[22][7] ), .ZN(net86414) );
  INV_X1 U3301 ( .A(\ab[22][7] ), .ZN(net81491) );
  NOR2_X1 U3302 ( .A1(net84698), .A2(net70469), .ZN(\ab[13][14] ) );
  XNOR2_X2 U3303 ( .A(n1095), .B(\SUMB[21][9] ), .ZN(\SUMB[22][8] ) );
  NAND2_X4 U3304 ( .A1(n1098), .A2(n1099), .ZN(n1095) );
  NAND2_X4 U3305 ( .A1(n1096), .A2(n1097), .ZN(n1099) );
  INV_X1 U3306 ( .A(\ab[22][8] ), .ZN(n1097) );
  INV_X4 U3307 ( .A(\CARRYB[21][8] ), .ZN(n1096) );
  NAND2_X2 U3308 ( .A1(\CARRYB[21][8] ), .A2(\ab[22][8] ), .ZN(n1098) );
  NAND2_X1 U3309 ( .A1(n856), .A2(\CARRYB[21][8] ), .ZN(net81178) );
  NAND2_X1 U3310 ( .A1(\ab[22][8] ), .A2(\CARRYB[21][8] ), .ZN(net81180) );
  NOR2_X4 U3311 ( .A1(net77920), .A2(net70453), .ZN(\ab[21][8] ) );
  NAND3_X4 U3312 ( .A1(n1100), .A2(net81956), .A3(net81955), .ZN(
        \CARRYB[20][8] ) );
  NAND2_X2 U3313 ( .A1(net89467), .A2(net89289), .ZN(n1100) );
  XOR2_X2 U3314 ( .A(n32), .B(net79950), .Z(\SUMB[9][18] ) );
  NAND2_X1 U3315 ( .A1(\ab[9][18] ), .A2(\SUMB[8][19] ), .ZN(net79952) );
  NAND2_X1 U3316 ( .A1(\CARRYB[8][18] ), .A2(n32), .ZN(net79951) );
  NAND2_X1 U3317 ( .A1(\ab[9][18] ), .A2(\CARRYB[8][18] ), .ZN(net79953) );
  XNOR2_X2 U3318 ( .A(\SUMB[7][20] ), .B(net86231), .ZN(\SUMB[8][19] ) );
  XNOR2_X2 U3319 ( .A(\CARRYB[7][19] ), .B(\ab[8][19] ), .ZN(net86231) );
  NAND2_X1 U3320 ( .A1(\CARRYB[7][19] ), .A2(\SUMB[7][20] ), .ZN(net79955) );
  NAND3_X4 U3321 ( .A1(n1103), .A2(n1102), .A3(n1101), .ZN(\CARRYB[7][19] ) );
  NAND2_X2 U3322 ( .A1(\ab[8][19] ), .A2(\CARRYB[7][19] ), .ZN(net79957) );
  NAND2_X1 U3323 ( .A1(\ab[7][19] ), .A2(\CARRYB[6][19] ), .ZN(n1101) );
  NAND2_X2 U3324 ( .A1(\ab[7][19] ), .A2(\SUMB[6][20] ), .ZN(n1102) );
  NOR2_X1 U3325 ( .A1(net86565), .A2(net77926), .ZN(\ab[8][19] ) );
  INV_X8 U3326 ( .A(B[19]), .ZN(net86565) );
  NAND2_X2 U3327 ( .A1(\ab[7][20] ), .A2(n840), .ZN(net79960) );
  NAND2_X1 U3328 ( .A1(\CARRYB[6][20] ), .A2(n840), .ZN(net79959) );
  NAND2_X1 U3329 ( .A1(\ab[7][20] ), .A2(\CARRYB[6][20] ), .ZN(net79961) );
  XNOR2_X2 U3330 ( .A(\CARRYB[6][19] ), .B(\ab[7][19] ), .ZN(n1104) );
  XNOR2_X2 U3331 ( .A(n1104), .B(\SUMB[6][20] ), .ZN(\SUMB[7][19] ) );
  NAND2_X1 U3332 ( .A1(\ab[19][10] ), .A2(\SUMB[18][11] ), .ZN(net82669) );
  NAND2_X1 U3333 ( .A1(\SUMB[18][11] ), .A2(\CARRYB[18][10] ), .ZN(net82668)
         );
  XNOR2_X2 U3334 ( .A(\ab[18][11] ), .B(\CARRYB[17][11] ), .ZN(net89353) );
  NOR2_X1 U3335 ( .A1(net85716), .A2(net70459), .ZN(\ab[18][11] ) );
  NAND2_X1 U3336 ( .A1(\ab[18][11] ), .A2(\CARRYB[17][11] ), .ZN(net82664) );
  NAND3_X4 U3337 ( .A1(net87011), .A2(net87010), .A3(net87012), .ZN(
        \CARRYB[17][11] ) );
  NOR2_X1 U3338 ( .A1(net70460), .A2(net70463), .ZN(\ab[16][13] ) );
  NAND2_X1 U3339 ( .A1(\ab[13][15] ), .A2(\SUMB[12][16] ), .ZN(net79892) );
  NAND2_X1 U3340 ( .A1(net93674), .A2(\SUMB[12][16] ), .ZN(net79893) );
  NAND2_X1 U3341 ( .A1(\ab[13][15] ), .A2(net93674), .ZN(net79891) );
  CLKBUF_X2 U3342 ( .A(\CARRYB[12][15] ), .Z(net93674) );
  NAND2_X2 U3343 ( .A1(\SUMB[7][19] ), .A2(n1109), .ZN(n1107) );
  INV_X4 U3344 ( .A(n1108), .ZN(n1109) );
  INV_X4 U3345 ( .A(\CARRYB[7][18] ), .ZN(n1108) );
  XNOR2_X2 U3346 ( .A(\ab[8][18] ), .B(n1108), .ZN(net79939) );
  NAND3_X2 U3347 ( .A1(n1110), .A2(net80303), .A3(net80302), .ZN(
        \CARRYB[7][18] ) );
  NAND2_X1 U3348 ( .A1(\SUMB[6][19] ), .A2(\CARRYB[6][18] ), .ZN(n1110) );
  NAND2_X2 U3349 ( .A1(\SUMB[7][19] ), .A2(\ab[8][18] ), .ZN(n1106) );
  NOR2_X1 U3350 ( .A1(n182), .A2(net70477), .ZN(\ab[9][18] ) );
  NAND2_X2 U3351 ( .A1(\ab[7][18] ), .A2(\CARRYB[6][18] ), .ZN(net80302) );
  INV_X8 U3352 ( .A(B[25]), .ZN(n1111) );
  NOR2_X2 U3353 ( .A1(n1111), .A2(net80409), .ZN(\ab[1][25] ) );
  NAND3_X4 U3354 ( .A1(n1114), .A2(n1113), .A3(n1112), .ZN(\CARRYB[18][10] )
         );
  NAND2_X1 U3355 ( .A1(\CARRYB[18][10] ), .A2(\ab[19][10] ), .ZN(net82667) );
  NAND2_X2 U3356 ( .A1(\ab[18][10] ), .A2(\SUMB[17][11] ), .ZN(n1114) );
  NAND2_X2 U3357 ( .A1(\CARRYB[17][10] ), .A2(\SUMB[17][11] ), .ZN(n1113) );
  NAND2_X1 U3358 ( .A1(\CARRYB[17][10] ), .A2(\ab[18][10] ), .ZN(n1112) );
  NOR2_X1 U3359 ( .A1(net91660), .A2(net70457), .ZN(\ab[19][10] ) );
  XNOR2_X2 U3360 ( .A(\SUMB[1][25] ), .B(n39), .ZN(net84883) );
  NAND2_X2 U3361 ( .A1(\SUMB[1][25] ), .A2(n39), .ZN(net84297) );
  XNOR2_X2 U3362 ( .A(\ab[0][26] ), .B(\ab[1][25] ), .ZN(
        \*UDW_*112644/net78437 ) );
  INV_X16 U3363 ( .A(B[26]), .ZN(net70486) );
  NOR2_X1 U3364 ( .A1(net80643), .A2(net77940), .ZN(\ab[6][21] ) );
  NAND3_X2 U3365 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(\CARRYB[5][21] ) );
  NAND2_X1 U3366 ( .A1(\SUMB[4][22] ), .A2(\CARRYB[4][21] ), .ZN(n1115) );
  XNOR2_X2 U3367 ( .A(net93880), .B(\SUMB[24][2] ), .ZN(\SUMB[25][1] ) );
  INV_X8 U3368 ( .A(B[20]), .ZN(net70474) );
  XNOR2_X2 U3369 ( .A(net124618), .B(\SUMB[1][14] ), .ZN(n1120) );
  NAND2_X2 U3370 ( .A1(\SUMB[6][16] ), .A2(n676), .ZN(n2210) );
  INV_X1 U3371 ( .A(net83850), .ZN(net93747) );
  XNOR2_X2 U3372 ( .A(net93713), .B(net83358), .ZN(\SUMB[23][1] ) );
  XNOR2_X2 U3373 ( .A(\CARRYB[15][8] ), .B(n2153), .ZN(n1279) );
  XNOR2_X2 U3374 ( .A(n1122), .B(n1389), .ZN(\SUMB[5][7] ) );
  NOR2_X2 U3375 ( .A1(net70452), .A2(net77946), .ZN(\ab[5][9] ) );
  NOR2_X2 U3376 ( .A1(net70452), .A2(net77924), .ZN(\ab[8][9] ) );
  NAND2_X2 U3377 ( .A1(\SUMB[7][10] ), .A2(\ab[8][9] ), .ZN(n2084) );
  NAND2_X1 U3378 ( .A1(\ab[18][9] ), .A2(\CARRYB[17][9] ), .ZN(n2154) );
  NAND2_X2 U3380 ( .A1(n596), .A2(\SUMB[20][3] ), .ZN(n2185) );
  NAND3_X2 U3382 ( .A1(net80817), .A2(net80818), .A3(net80816), .ZN(n1184) );
  INV_X8 U3383 ( .A(net86661), .ZN(net86662) );
  NAND2_X4 U3384 ( .A1(\ab[3][7] ), .A2(net85036), .ZN(n1648) );
  NAND2_X4 U3385 ( .A1(net86662), .A2(n1719), .ZN(n2233) );
  NAND2_X4 U3387 ( .A1(n1125), .A2(n1124), .ZN(\SUMB[12][8] ) );
  INV_X4 U3388 ( .A(net82548), .ZN(net93308) );
  NAND2_X4 U3389 ( .A1(\SUMB[15][5] ), .A2(\ab[16][4] ), .ZN(n2104) );
  NAND3_X2 U3390 ( .A1(n2307), .A2(n2308), .A3(n2309), .ZN(\CARRYB[12][16] )
         );
  XNOR2_X2 U3391 ( .A(n1539), .B(\SUMB[3][26] ), .ZN(n1185) );
  NAND2_X4 U3392 ( .A1(n288), .A2(n1157), .ZN(n2057) );
  NAND2_X2 U3393 ( .A1(n1193), .A2(\SUMB[11][7] ), .ZN(n1919) );
  NAND2_X4 U3394 ( .A1(n1500), .A2(\SUMB[15][5] ), .ZN(n2103) );
  NAND3_X4 U3397 ( .A1(n1813), .A2(n1814), .A3(n1815), .ZN(\CARRYB[19][0] ) );
  NAND2_X2 U3398 ( .A1(\SUMB[9][4] ), .A2(\CARRYB[9][3] ), .ZN(n1804) );
  NAND2_X2 U3399 ( .A1(\CARRYB[1][18] ), .A2(\ab[2][18] ), .ZN(n1711) );
  NAND2_X2 U3400 ( .A1(n1732), .A2(n1588), .ZN(n1446) );
  NAND2_X2 U3401 ( .A1(\ab[16][3] ), .A2(\SUMB[15][4] ), .ZN(n1130) );
  NAND3_X4 U3402 ( .A1(n1990), .A2(n1991), .A3(n1992), .ZN(\CARRYB[15][3] ) );
  XNOR2_X2 U3403 ( .A(n1132), .B(n1133), .ZN(n1312) );
  XNOR2_X2 U3404 ( .A(n2066), .B(\SUMB[14][17] ), .ZN(n1132) );
  XNOR2_X2 U3405 ( .A(\CARRYB[15][15] ), .B(\ab[16][15] ), .ZN(n1133) );
  XNOR2_X2 U3406 ( .A(\CARRYB[18][3] ), .B(\ab[19][3] ), .ZN(n2110) );
  XNOR2_X2 U3407 ( .A(n558), .B(n1869), .ZN(n1229) );
  NOR2_X1 U3408 ( .A1(net70486), .A2(net77956), .ZN(\ab[4][26] ) );
  INV_X8 U3409 ( .A(B[27]), .ZN(n2355) );
  NAND2_X4 U3410 ( .A1(n1523), .A2(n1522), .ZN(net91088) );
  NAND2_X2 U3411 ( .A1(\CARRYB[8][6] ), .A2(\SUMB[8][7] ), .ZN(n1292) );
  NAND2_X2 U3412 ( .A1(\CARRYB[10][3] ), .A2(\SUMB[10][4] ), .ZN(n1672) );
  NAND2_X4 U3413 ( .A1(net88166), .A2(n1317), .ZN(n1319) );
  NAND2_X4 U3414 ( .A1(\CARRYB[19][6] ), .A2(n1190), .ZN(n2211) );
  NOR2_X1 U3415 ( .A1(net70482), .A2(net77966), .ZN(\ab[3][24] ) );
  XOR2_X2 U3416 ( .A(\SUMB[1][5] ), .B(n1135), .Z(\SUMB[2][4] ) );
  NAND2_X1 U3417 ( .A1(\CARRYB[1][4] ), .A2(\SUMB[1][5] ), .ZN(n1136) );
  NAND2_X2 U3418 ( .A1(\ab[2][4] ), .A2(\SUMB[1][5] ), .ZN(n1137) );
  NAND2_X1 U3419 ( .A1(\ab[2][4] ), .A2(\CARRYB[1][4] ), .ZN(n1138) );
  NAND3_X2 U3420 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(\CARRYB[2][4] ) );
  NAND3_X2 U3421 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(\CARRYB[11][0] ) );
  XOR2_X1 U3422 ( .A(\ab[12][0] ), .B(\SUMB[11][1] ), .Z(n1143) );
  XOR2_X2 U3423 ( .A(n1143), .B(\CARRYB[11][0] ), .Z(PRODUCT[12]) );
  NAND2_X2 U3424 ( .A1(\ab[12][0] ), .A2(\CARRYB[11][0] ), .ZN(n1145) );
  NAND3_X2 U3425 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(\CARRYB[12][0] ) );
  NAND2_X2 U3426 ( .A1(\ab[3][4] ), .A2(\SUMB[2][5] ), .ZN(n1148) );
  NAND2_X1 U3427 ( .A1(\ab[3][4] ), .A2(\CARRYB[2][4] ), .ZN(n1149) );
  NAND3_X2 U3428 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(\CARRYB[3][4] ) );
  NOR2_X2 U3429 ( .A1(net77892), .A2(net77970), .ZN(\ab[2][4] ) );
  NOR2_X1 U3430 ( .A1(net77892), .A2(net77966), .ZN(\ab[3][4] ) );
  NAND2_X2 U3431 ( .A1(n2244), .A2(net148233), .ZN(n1364) );
  NAND3_X4 U3432 ( .A1(n1620), .A2(n1619), .A3(n1621), .ZN(\CARRYB[9][9] ) );
  NAND2_X1 U3433 ( .A1(\ab[5][20] ), .A2(\CARRYB[4][20] ), .ZN(n1885) );
  NAND2_X2 U3434 ( .A1(n1783), .A2(n1784), .ZN(n2060) );
  NAND2_X2 U3435 ( .A1(\CARRYB[9][1] ), .A2(\ab[10][1] ), .ZN(n1471) );
  NAND3_X4 U3436 ( .A1(n2229), .A2(n2230), .A3(n2228), .ZN(\CARRYB[20][4] ) );
  NAND2_X4 U3437 ( .A1(n1150), .A2(n1151), .ZN(n1153) );
  NAND2_X4 U3438 ( .A1(n1153), .A2(n1152), .ZN(\SUMB[15][5] ) );
  INV_X4 U3439 ( .A(n1721), .ZN(n1150) );
  NAND2_X2 U3440 ( .A1(\ab[9][6] ), .A2(\CARRYB[8][6] ), .ZN(n1294) );
  XNOR2_X2 U3441 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .ZN(n1204) );
  XNOR2_X1 U3442 ( .A(\CARRYB[2][11] ), .B(\ab[3][11] ), .ZN(n1869) );
  NAND2_X2 U3443 ( .A1(\CARRYB[6][6] ), .A2(\SUMB[6][7] ), .ZN(n1335) );
  NAND2_X2 U3444 ( .A1(\ab[2][10] ), .A2(n2332), .ZN(n1155) );
  INV_X4 U3445 ( .A(\ab[2][10] ), .ZN(n1154) );
  INV_X8 U3446 ( .A(n2335), .ZN(\SUMB[1][11] ) );
  NAND2_X4 U3447 ( .A1(net92716), .A2(net92717), .ZN(n1158) );
  NAND2_X4 U3448 ( .A1(n1158), .A2(net92718), .ZN(n1720) );
  INV_X4 U3449 ( .A(\CARRYB[3][14] ), .ZN(net92717) );
  INV_X1 U3450 ( .A(\ab[6][13] ), .ZN(n1159) );
  NAND2_X4 U3451 ( .A1(n1984), .A2(n1163), .ZN(n1361) );
  INV_X2 U3452 ( .A(\ab[2][15] ), .ZN(net92724) );
  NOR2_X2 U3453 ( .A1(net84698), .A2(net119855), .ZN(\ab[4][14] ) );
  NAND3_X4 U3454 ( .A1(n1988), .A2(n1987), .A3(n1989), .ZN(\CARRYB[3][14] ) );
  NOR2_X4 U3455 ( .A1(net70460), .A2(net77940), .ZN(\ab[6][13] ) );
  NAND2_X2 U3456 ( .A1(n1361), .A2(\SUMB[1][16] ), .ZN(n1353) );
  INV_X4 U3457 ( .A(n1361), .ZN(n1351) );
  NAND2_X4 U3458 ( .A1(net85455), .A2(net85456), .ZN(n1505) );
  OR2_X1 U3459 ( .A1(net70451), .A2(net70452), .ZN(n1929) );
  NOR2_X1 U3460 ( .A1(net70452), .A2(net70453), .ZN(\ab[21][9] ) );
  NOR2_X1 U3461 ( .A1(net70452), .A2(net70457), .ZN(\ab[19][9] ) );
  NAND2_X2 U3462 ( .A1(n1837), .A2(n1260), .ZN(n1166) );
  NAND2_X4 U3463 ( .A1(n1164), .A2(n1165), .ZN(n1167) );
  NAND2_X4 U3464 ( .A1(n1166), .A2(n1167), .ZN(\SUMB[13][5] ) );
  INV_X4 U3465 ( .A(n1837), .ZN(n1164) );
  INV_X4 U3466 ( .A(n1260), .ZN(n1165) );
  NAND2_X4 U3467 ( .A1(n1170), .A2(n1171), .ZN(\SUMB[6][10] ) );
  INV_X4 U3468 ( .A(n1694), .ZN(n1168) );
  INV_X1 U3469 ( .A(\CARRYB[5][10] ), .ZN(n1169) );
  NAND3_X4 U3470 ( .A1(n2080), .A2(n2081), .A3(n2082), .ZN(n1207) );
  NAND2_X2 U3471 ( .A1(n1563), .A2(\CARRYB[8][9] ), .ZN(n1174) );
  NAND2_X4 U3472 ( .A1(n1172), .A2(n1173), .ZN(n1175) );
  INV_X4 U3473 ( .A(n1563), .ZN(n1173) );
  INV_X2 U3474 ( .A(\ab[9][9] ), .ZN(n1563) );
  NAND2_X4 U3475 ( .A1(n1345), .A2(\ab[14][12] ), .ZN(n1488) );
  NAND2_X4 U3476 ( .A1(\SUMB[7][12] ), .A2(\ab[8][11] ), .ZN(n2127) );
  XNOR2_X2 U3477 ( .A(n1176), .B(n946), .ZN(\SUMB[9][7] ) );
  INV_X4 U3478 ( .A(n2243), .ZN(n1755) );
  NAND2_X2 U3479 ( .A1(\CARRYB[8][8] ), .A2(\ab[9][8] ), .ZN(n1179) );
  INV_X1 U3480 ( .A(\ab[9][8] ), .ZN(n1178) );
  NAND2_X2 U3481 ( .A1(\CARRYB[6][13] ), .A2(\ab[7][13] ), .ZN(n1320) );
  INV_X4 U3482 ( .A(net88702), .ZN(net85469) );
  NAND2_X4 U3483 ( .A1(n1373), .A2(n1374), .ZN(n1730) );
  NAND3_X1 U3484 ( .A1(net80355), .A2(net80356), .A3(n2272), .ZN(n1235) );
  NAND2_X4 U3485 ( .A1(n1195), .A2(n176), .ZN(n2076) );
  NAND2_X4 U3486 ( .A1(\SUMB[16][5] ), .A2(\ab[17][4] ), .ZN(n2075) );
  NAND2_X4 U3487 ( .A1(n1275), .A2(\ab[12][5] ), .ZN(n1637) );
  INV_X4 U3488 ( .A(\SUMB[15][9] ), .ZN(n1449) );
  NAND2_X2 U3489 ( .A1(\ab[12][3] ), .A2(\CARRYB[11][3] ), .ZN(n1674) );
  NAND2_X4 U3490 ( .A1(n1201), .A2(\ab[17][5] ), .ZN(n1382) );
  NAND2_X2 U3491 ( .A1(\CARRYB[6][6] ), .A2(\ab[7][6] ), .ZN(n1333) );
  NAND2_X4 U3492 ( .A1(\ab[24][2] ), .A2(\CARRYB[23][2] ), .ZN(net80258) );
  NAND3_X2 U3493 ( .A1(n1670), .A2(n1671), .A3(n1672), .ZN(\CARRYB[11][3] ) );
  NAND2_X2 U3494 ( .A1(\SUMB[4][9] ), .A2(\CARRYB[4][8] ), .ZN(n1966) );
  CLKBUF_X3 U3495 ( .A(\SUMB[4][9] ), .Z(n1217) );
  NAND2_X2 U3496 ( .A1(\SUMB[22][1] ), .A2(\ab[23][0] ), .ZN(n1799) );
  NOR2_X1 U3497 ( .A1(net70452), .A2(net77966), .ZN(\ab[3][9] ) );
  NAND3_X4 U3498 ( .A1(net80920), .A2(net80922), .A3(net80921), .ZN(
        \CARRYB[24][1] ) );
  NAND2_X4 U3499 ( .A1(n1544), .A2(net85254), .ZN(n1679) );
  XNOR2_X2 U3500 ( .A(net92378), .B(n284), .ZN(PRODUCT[28]) );
  NAND3_X4 U3501 ( .A1(net84116), .A2(n1648), .A3(net84118), .ZN(
        \CARRYB[3][7] ) );
  NAND3_X1 U3502 ( .A1(n2011), .A2(n2376), .A3(n2012), .ZN(net91001) );
  NAND3_X2 U3503 ( .A1(n1796), .A2(n1797), .A3(n1798), .ZN(\CARRYB[22][0] ) );
  NAND3_X4 U3504 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(\CARRYB[10][14] )
         );
  NAND2_X4 U3505 ( .A1(n176), .A2(\ab[17][4] ), .ZN(n2074) );
  XNOR2_X2 U3506 ( .A(n1182), .B(n1183), .ZN(net92322) );
  XNOR2_X2 U3507 ( .A(n1184), .B(net92341), .ZN(n1183) );
  NAND2_X4 U3508 ( .A1(\ab[15][4] ), .A2(n1211), .ZN(n1705) );
  NAND2_X4 U3509 ( .A1(\ab[3][20] ), .A2(\CARRYB[2][20] ), .ZN(n2192) );
  XNOR2_X2 U3510 ( .A(n2065), .B(\SUMB[14][13] ), .ZN(n1187) );
  XNOR2_X2 U3511 ( .A(n1821), .B(\SUMB[6][8] ), .ZN(n1188) );
  INV_X4 U3512 ( .A(n1188), .ZN(\SUMB[7][7] ) );
  CLKBUF_X3 U3513 ( .A(\SUMB[16][6] ), .Z(n1270) );
  NAND3_X2 U3514 ( .A1(n2279), .A2(n2280), .A3(n2281), .ZN(\CARRYB[6][19] ) );
  XNOR2_X2 U3515 ( .A(\CARRYB[10][13] ), .B(\ab[11][13] ), .ZN(n1221) );
  INV_X4 U3516 ( .A(n1192), .ZN(n1193) );
  INV_X2 U3517 ( .A(n1298), .ZN(n1194) );
  XNOR2_X2 U3518 ( .A(n1585), .B(n1236), .ZN(n1195) );
  NAND2_X4 U3519 ( .A1(net87310), .A2(n1367), .ZN(net85212) );
  NAND2_X1 U3521 ( .A1(\CARRYB[14][12] ), .A2(\SUMB[14][13] ), .ZN(n2198) );
  NAND3_X2 U3522 ( .A1(n2198), .A2(n2199), .A3(n2200), .ZN(\CARRYB[15][12] )
         );
  INV_X4 U3523 ( .A(\SUMB[2][27] ), .ZN(n1196) );
  XNOR2_X2 U3524 ( .A(n1198), .B(\SUMB[8][7] ), .ZN(\SUMB[9][6] ) );
  NAND2_X4 U3525 ( .A1(\CARRYB[18][5] ), .A2(\ab[19][5] ), .ZN(net84708) );
  NAND2_X4 U3526 ( .A1(net85373), .A2(net85732), .ZN(n1523) );
  XNOR2_X2 U3527 ( .A(n1200), .B(n842), .ZN(\SUMB[11][3] ) );
  NAND3_X2 U3528 ( .A1(n2071), .A2(n2072), .A3(n2073), .ZN(n1201) );
  NAND2_X4 U3529 ( .A1(n1617), .A2(net91243), .ZN(n1522) );
  NAND3_X2 U3530 ( .A1(n1652), .A2(n1653), .A3(n1654), .ZN(n1203) );
  XNOR2_X2 U3531 ( .A(n1204), .B(\SUMB[19][11] ), .ZN(\SUMB[20][10] ) );
  NAND3_X2 U3532 ( .A1(n1958), .A2(n1959), .A3(n1960), .ZN(\CARRYB[5][23] ) );
  NAND3_X2 U3533 ( .A1(net81365), .A2(net81367), .A3(n2035), .ZN(
        \CARRYB[7][14] ) );
  INV_X2 U3534 ( .A(n1767), .ZN(n1768) );
  NOR2_X2 U3535 ( .A1(net70460), .A2(net70475), .ZN(\ab[10][13] ) );
  NAND3_X2 U3538 ( .A1(n1409), .A2(n1410), .A3(n1411), .ZN(\CARRYB[15][0] ) );
  XNOR2_X2 U3539 ( .A(n1210), .B(\SUMB[4][21] ), .ZN(\SUMB[5][20] ) );
  CLKBUF_X3 U3540 ( .A(\SUMB[15][6] ), .Z(n1236) );
  NAND3_X2 U3541 ( .A1(n2150), .A2(n2151), .A3(n2152), .ZN(n1211) );
  CLKBUF_X3 U3542 ( .A(\SUMB[13][5] ), .Z(n1253) );
  NAND2_X2 U3543 ( .A1(n943), .A2(\ab[5][9] ), .ZN(n1396) );
  XNOR2_X2 U3544 ( .A(\SUMB[5][19] ), .B(n1212), .ZN(net90702) );
  XNOR2_X2 U3545 ( .A(\CARRYB[5][18] ), .B(\ab[6][18] ), .ZN(n1212) );
  CLKBUF_X2 U3546 ( .A(\SUMB[6][24] ), .Z(n1213) );
  INV_X4 U3547 ( .A(\CARRYB[4][13] ), .ZN(n1541) );
  XNOR2_X2 U3550 ( .A(n1215), .B(\SUMB[11][17] ), .ZN(\SUMB[12][16] ) );
  XNOR2_X2 U3551 ( .A(\ab[12][16] ), .B(\CARRYB[11][16] ), .ZN(n1215) );
  XNOR2_X2 U3552 ( .A(n1216), .B(n1220), .ZN(\SUMB[10][15] ) );
  XNOR2_X2 U3553 ( .A(\CARRYB[9][15] ), .B(n1624), .ZN(n1216) );
  NAND2_X2 U3554 ( .A1(n1943), .A2(\SUMB[18][8] ), .ZN(n1510) );
  INV_X2 U3555 ( .A(\SUMB[2][26] ), .ZN(n1218) );
  XNOR2_X2 U3556 ( .A(n1221), .B(\SUMB[10][14] ), .ZN(\SUMB[11][13] ) );
  NAND3_X2 U3557 ( .A1(n1437), .A2(n1436), .A3(n1438), .ZN(net90347) );
  XNOR2_X2 U3558 ( .A(n1993), .B(n1253), .ZN(n1222) );
  XNOR2_X2 U3559 ( .A(n1223), .B(\SUMB[11][18] ), .ZN(\SUMB[12][17] ) );
  XNOR2_X2 U3560 ( .A(\CARRYB[11][17] ), .B(\ab[12][17] ), .ZN(n1223) );
  XNOR2_X2 U3561 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .ZN(n1226) );
  XNOR2_X2 U3562 ( .A(n1227), .B(n367), .ZN(\SUMB[10][14] ) );
  NAND2_X2 U3563 ( .A1(net91088), .A2(\CARRYB[11][9] ), .ZN(net88295) );
  FA_X1 U3564 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .CI(n844), .S(n1231) );
  XNOR2_X2 U3565 ( .A(n1232), .B(n20), .ZN(\SUMB[20][2] ) );
  XNOR2_X2 U3566 ( .A(\CARRYB[20][2] ), .B(\ab[21][2] ), .ZN(n2171) );
  NAND2_X2 U3567 ( .A1(\ab[7][6] ), .A2(\SUMB[6][7] ), .ZN(n1334) );
  NAND2_X2 U3568 ( .A1(n1627), .A2(n1628), .ZN(n1630) );
  XNOR2_X2 U3569 ( .A(\CARRYB[22][6] ), .B(n1234), .ZN(n2282) );
  NAND3_X2 U3570 ( .A1(n2102), .A2(n2101), .A3(n2100), .ZN(n1237) );
  NAND2_X2 U3571 ( .A1(n1121), .A2(n2149), .ZN(n1301) );
  XOR2_X2 U3572 ( .A(\SUMB[9][20] ), .B(n2215), .Z(\SUMB[10][19] ) );
  XNOR2_X2 U3573 ( .A(n1238), .B(\SUMB[3][2] ), .ZN(\SUMB[4][1] ) );
  XNOR2_X2 U3574 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .ZN(n1238) );
  XNOR2_X2 U3575 ( .A(n1371), .B(net88800), .ZN(net89876) );
  XNOR2_X2 U3576 ( .A(\SUMB[16][12] ), .B(n1239), .ZN(\SUMB[17][11] ) );
  XNOR2_X2 U3577 ( .A(\CARRYB[16][11] ), .B(\ab[17][11] ), .ZN(n1239) );
  XNOR2_X2 U3578 ( .A(\SUMB[11][5] ), .B(n1243), .ZN(\SUMB[12][4] ) );
  XNOR2_X2 U3579 ( .A(n1244), .B(\SUMB[1][26] ), .ZN(\SUMB[2][25] ) );
  XNOR2_X2 U3580 ( .A(\ab[2][25] ), .B(n349), .ZN(n1244) );
  INV_X4 U3581 ( .A(n1245), .ZN(n1246) );
  NAND3_X2 U3582 ( .A1(n2241), .A2(n2240), .A3(n2242), .ZN(\CARRYB[5][19] ) );
  XNOR2_X2 U3583 ( .A(\SUMB[5][21] ), .B(n1247), .ZN(\SUMB[6][20] ) );
  XNOR2_X2 U3584 ( .A(\CARRYB[5][20] ), .B(\ab[6][20] ), .ZN(n1247) );
  NAND2_X2 U3586 ( .A1(\CARRYB[14][12] ), .A2(\ab[15][12] ), .ZN(n1852) );
  NOR2_X2 U3587 ( .A1(net81424), .A2(net70465), .ZN(\ab[15][15] ) );
  INV_X2 U3588 ( .A(n615), .ZN(n1250) );
  NAND3_X2 U3589 ( .A1(net79906), .A2(net79905), .A3(net79904), .ZN(n1251) );
  NAND2_X2 U3590 ( .A1(\ab[13][3] ), .A2(\CARRYB[12][3] ), .ZN(n1678) );
  NAND3_X2 U3591 ( .A1(n1673), .A2(n1674), .A3(n1675), .ZN(\CARRYB[12][3] ) );
  NAND2_X4 U3592 ( .A1(net86662), .A2(\ab[18][5] ), .ZN(n2232) );
  XNOR2_X2 U3593 ( .A(n1254), .B(n24), .ZN(\SUMB[19][2] ) );
  NAND2_X4 U3594 ( .A1(\SUMB[9][12] ), .A2(net82678), .ZN(net80956) );
  NAND3_X2 U3595 ( .A1(n2091), .A2(n2090), .A3(n2089), .ZN(n1255) );
  NOR2_X2 U3596 ( .A1(net83784), .A2(net77956), .ZN(\ab[4][12] ) );
  NAND3_X2 U3597 ( .A1(net79906), .A2(net79905), .A3(net79904), .ZN(
        \CARRYB[23][5] ) );
  NAND2_X1 U3598 ( .A1(\CARRYB[6][23] ), .A2(n1213), .ZN(n2268) );
  NAND2_X1 U3599 ( .A1(\ab[7][23] ), .A2(n1213), .ZN(n2267) );
  XNOR2_X2 U3600 ( .A(\SUMB[8][20] ), .B(n1257), .ZN(\SUMB[9][19] ) );
  XNOR2_X2 U3601 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .ZN(n1257) );
  NAND2_X4 U3604 ( .A1(\CARRYB[18][7] ), .A2(\ab[19][7] ), .ZN(n2010) );
  INV_X4 U3605 ( .A(n1730), .ZN(n1627) );
  INV_X4 U3606 ( .A(net124563), .ZN(net85456) );
  INV_X4 U3607 ( .A(n1263), .ZN(n1264) );
  XNOR2_X2 U3608 ( .A(n1903), .B(\CARRYB[9][4] ), .ZN(\SUMB[10][4] ) );
  XNOR2_X2 U3609 ( .A(\ab[10][4] ), .B(\SUMB[9][5] ), .ZN(n1903) );
  XNOR2_X2 U3610 ( .A(n1267), .B(\SUMB[12][3] ), .ZN(\SUMB[13][2] ) );
  XNOR2_X2 U3611 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .ZN(n1267) );
  XNOR2_X2 U3612 ( .A(n1268), .B(n1241), .ZN(\SUMB[18][3] ) );
  INV_X2 U3613 ( .A(net88867), .ZN(net88868) );
  INV_X2 U3614 ( .A(net88859), .ZN(net88860) );
  FA_X1 U3615 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), 
        .S(n1269) );
  INV_X4 U3616 ( .A(n1781), .ZN(n1271) );
  INV_X4 U3617 ( .A(\CARRYB[10][5] ), .ZN(n1781) );
  NAND3_X2 U3618 ( .A1(n1575), .A2(n1574), .A3(n1573), .ZN(\CARRYB[13][13] )
         );
  XNOR2_X2 U3619 ( .A(\CARRYB[22][8] ), .B(\ab[23][8] ), .ZN(n1273) );
  XNOR2_X2 U3620 ( .A(\CARRYB[25][4] ), .B(\ab[26][4] ), .ZN(n1310) );
  NAND2_X1 U3621 ( .A1(\ab[13][17] ), .A2(n1240), .ZN(n2223) );
  NAND2_X1 U3622 ( .A1(\CARRYB[12][17] ), .A2(n1240), .ZN(n2224) );
  XNOR2_X2 U3623 ( .A(\CARRYB[10][4] ), .B(\ab[11][4] ), .ZN(n1276) );
  INV_X2 U3624 ( .A(\SUMB[8][21] ), .ZN(n1277) );
  XNOR2_X2 U3626 ( .A(net86427), .B(net88656), .ZN(n1281) );
  INV_X2 U3627 ( .A(net88655), .ZN(net88656) );
  INV_X4 U3628 ( .A(n1449), .ZN(n1282) );
  XNOR2_X2 U3629 ( .A(\CARRYB[19][11] ), .B(n1283), .ZN(n2142) );
  OR2_X1 U3630 ( .A1(net70455), .A2(net85716), .ZN(n1283) );
  NAND2_X2 U3631 ( .A1(\SUMB[13][10] ), .A2(net85043), .ZN(n1940) );
  NAND2_X2 U3632 ( .A1(\ab[3][10] ), .A2(n1203), .ZN(n1645) );
  NAND3_X2 U3633 ( .A1(net80957), .A2(net80956), .A3(net80958), .ZN(net88525)
         );
  NAND2_X2 U3634 ( .A1(\CARRYB[4][19] ), .A2(\SUMB[4][20] ), .ZN(n2242) );
  NAND2_X4 U3635 ( .A1(n1286), .A2(n1285), .ZN(n1287) );
  NAND2_X4 U3636 ( .A1(n1287), .A2(n2019), .ZN(n1902) );
  INV_X2 U3637 ( .A(\ab[12][7] ), .ZN(n1285) );
  NAND2_X2 U3638 ( .A1(\CARRYB[9][8] ), .A2(n1503), .ZN(n1290) );
  NAND2_X4 U3639 ( .A1(n1288), .A2(n1289), .ZN(n1291) );
  INV_X8 U3640 ( .A(n1503), .ZN(n1288) );
  NOR2_X2 U3641 ( .A1(net77914), .A2(net70471), .ZN(\ab[12][7] ) );
  INV_X1 U3642 ( .A(\ab[10][8] ), .ZN(n1503) );
  NAND2_X4 U3643 ( .A1(n1430), .A2(\ab[7][8] ), .ZN(n2058) );
  NAND2_X4 U3644 ( .A1(\SUMB[26][1] ), .A2(\ab[27][0] ), .ZN(net80768) );
  NAND2_X4 U3645 ( .A1(\CARRYB[26][0] ), .A2(n1281), .ZN(net80769) );
  NAND2_X4 U3646 ( .A1(n1755), .A2(net87573), .ZN(n1756) );
  NAND2_X4 U3647 ( .A1(n1377), .A2(n1378), .ZN(\SUMB[7][15] ) );
  NAND2_X2 U3648 ( .A1(n1375), .A2(n2204), .ZN(n1378) );
  NAND2_X2 U3649 ( .A1(\ab[9][6] ), .A2(\SUMB[8][7] ), .ZN(n1293) );
  NAND2_X2 U3650 ( .A1(n1635), .A2(n1298), .ZN(n1299) );
  NAND2_X2 U3651 ( .A1(n1297), .A2(n1194), .ZN(n1300) );
  NAND2_X4 U3652 ( .A1(n1299), .A2(n1300), .ZN(\SUMB[13][4] ) );
  INV_X4 U3653 ( .A(n1635), .ZN(n1297) );
  INV_X1 U3654 ( .A(\SUMB[12][5] ), .ZN(n1298) );
  NAND3_X4 U3655 ( .A1(n1826), .A2(n1827), .A3(n1825), .ZN(\CARRYB[8][6] ) );
  NAND2_X2 U3656 ( .A1(\CARRYB[6][7] ), .A2(\SUMB[6][8] ), .ZN(n1824) );
  NAND2_X2 U3657 ( .A1(\SUMB[6][8] ), .A2(\ab[7][7] ), .ZN(n1823) );
  NAND2_X2 U3658 ( .A1(\CARRYB[12][4] ), .A2(\SUMB[12][5] ), .ZN(n1641) );
  NAND2_X2 U3659 ( .A1(\ab[13][4] ), .A2(\CARRYB[12][4] ), .ZN(n1639) );
  NAND3_X2 U3660 ( .A1(n2061), .A2(n2062), .A3(n2063), .ZN(\CARRYB[11][5] ) );
  INV_X1 U3661 ( .A(net88157), .ZN(net88444) );
  INV_X8 U3662 ( .A(\CARRYB[6][13] ), .ZN(net88157) );
  NAND2_X2 U3663 ( .A1(\SUMB[9][15] ), .A2(\ab[10][14] ), .ZN(n1303) );
  NAND2_X2 U3664 ( .A1(\SUMB[9][15] ), .A2(\CARRYB[9][14] ), .ZN(n1304) );
  NAND2_X1 U3665 ( .A1(\CARRYB[10][13] ), .A2(\ab[11][13] ), .ZN(n1305) );
  NAND2_X2 U3666 ( .A1(\SUMB[10][14] ), .A2(\CARRYB[10][13] ), .ZN(n1306) );
  NAND2_X2 U3667 ( .A1(\SUMB[10][14] ), .A2(\ab[11][13] ), .ZN(n1307) );
  NAND3_X4 U3668 ( .A1(n1307), .A2(n1306), .A3(n1305), .ZN(\CARRYB[11][13] )
         );
  NAND2_X4 U3669 ( .A1(n1780), .A2(n896), .ZN(n2149) );
  NAND3_X4 U3670 ( .A1(n1832), .A2(n1833), .A3(n1834), .ZN(\CARRYB[11][4] ) );
  XNOR2_X2 U3671 ( .A(n1973), .B(n1308), .ZN(\SUMB[14][6] ) );
  XNOR2_X2 U3673 ( .A(\SUMB[25][5] ), .B(n1310), .ZN(\SUMB[26][4] ) );
  NAND3_X2 U3674 ( .A1(net80676), .A2(net80675), .A3(net80674), .ZN(
        \CARRYB[21][6] ) );
  NAND3_X2 U3675 ( .A1(n2011), .A2(n2012), .A3(n2376), .ZN(\CARRYB[19][7] ) );
  NOR2_X1 U3676 ( .A1(net91660), .A2(net70455), .ZN(\ab[20][10] ) );
  NOR2_X1 U3677 ( .A1(net70454), .A2(net77946), .ZN(\ab[5][10] ) );
  INV_X4 U3679 ( .A(\ab[3][18] ), .ZN(n1546) );
  NAND2_X4 U3680 ( .A1(\SUMB[3][21] ), .A2(n1009), .ZN(n2239) );
  XNOR2_X2 U3681 ( .A(net121785), .B(n1311), .ZN(\SUMB[4][11] ) );
  XNOR2_X2 U3682 ( .A(\CARRYB[3][11] ), .B(\ab[4][11] ), .ZN(n1311) );
  XNOR2_X2 U3683 ( .A(n1312), .B(n1369), .ZN(\SUMB[17][14] ) );
  INV_X2 U3684 ( .A(net70474), .ZN(net81080) );
  INV_X4 U3685 ( .A(net85465), .ZN(net87064) );
  NOR2_X2 U3686 ( .A1(net88344), .A2(net77940), .ZN(\ab[6][16] ) );
  NOR2_X1 U3687 ( .A1(net124723), .A2(net70467), .ZN(\ab[14][16] ) );
  XNOR2_X2 U3688 ( .A(n1314), .B(\SUMB[8][22] ), .ZN(\SUMB[9][21] ) );
  XNOR2_X2 U3689 ( .A(\ab[9][21] ), .B(\CARRYB[8][21] ), .ZN(n1314) );
  NAND2_X4 U3690 ( .A1(\ab[3][8] ), .A2(n1427), .ZN(n1906) );
  NAND2_X1 U3691 ( .A1(\ab[9][21] ), .A2(\SUMB[8][22] ), .ZN(n1687) );
  INV_X4 U3692 ( .A(\CARRYB[26][3] ), .ZN(n1533) );
  NAND2_X2 U3693 ( .A1(\CARRYB[8][16] ), .A2(n1600), .ZN(n1601) );
  INV_X4 U3694 ( .A(\CARRYB[14][11] ), .ZN(n1770) );
  NAND2_X4 U3695 ( .A1(n952), .A2(n1282), .ZN(n1451) );
  NAND3_X2 U3696 ( .A1(n2091), .A2(n2090), .A3(n2089), .ZN(\CARRYB[4][13] ) );
  XOR2_X2 U3697 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .Z(n1316) );
  XOR2_X2 U3698 ( .A(n1316), .B(\SUMB[6][4] ), .Z(\SUMB[7][3] ) );
  NAND3_X2 U3699 ( .A1(net88206), .A2(net88207), .A3(net88208), .ZN(
        \CARRYB[4][6] ) );
  NAND3_X4 U3700 ( .A1(net88209), .A2(net88210), .A3(net88211), .ZN(
        \CARRYB[5][5] ) );
  NAND2_X1 U3701 ( .A1(\ab[20][8] ), .A2(\CARRYB[19][8] ), .ZN(net81955) );
  NAND3_X2 U3702 ( .A1(net82557), .A2(net82558), .A3(net82556), .ZN(
        \CARRYB[14][11] ) );
  NAND2_X2 U3703 ( .A1(n2095), .A2(n1733), .ZN(n1727) );
  NAND2_X4 U3704 ( .A1(n1318), .A2(n1319), .ZN(\SUMB[7][12] ) );
  XNOR2_X2 U3705 ( .A(net88165), .B(\SUMB[17][13] ), .ZN(\SUMB[18][12] ) );
  NAND2_X2 U3706 ( .A1(n1246), .A2(\ab[3][9] ), .ZN(n1655) );
  INV_X1 U3707 ( .A(\ab[7][13] ), .ZN(net88156) );
  NOR2_X4 U3708 ( .A1(net70460), .A2(net77932), .ZN(\ab[7][13] ) );
  NAND3_X2 U3709 ( .A1(net82099), .A2(n1923), .A3(net82101), .ZN(
        \CARRYB[9][4] ) );
  XNOR2_X2 U3710 ( .A(n1219), .B(n1322), .ZN(\SUMB[3][25] ) );
  XNOR2_X2 U3711 ( .A(\ab[3][25] ), .B(\CARRYB[2][25] ), .ZN(n1322) );
  NAND2_X4 U3712 ( .A1(n1541), .A2(n1540), .ZN(n1543) );
  NAND2_X4 U3713 ( .A1(\SUMB[1][20] ), .A2(\ab[2][19] ), .ZN(n2144) );
  INV_X8 U3714 ( .A(\CARRYB[17][9] ), .ZN(net83850) );
  NAND3_X2 U3715 ( .A1(n1715), .A2(n1714), .A3(n1716), .ZN(\CARRYB[3][17] ) );
  NAND2_X2 U3716 ( .A1(\ab[6][17] ), .A2(\SUMB[5][18] ), .ZN(n2246) );
  NAND2_X4 U3717 ( .A1(net83120), .A2(\ab[22][7] ), .ZN(n1759) );
  XNOR2_X2 U3718 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .ZN(n1323) );
  XNOR2_X2 U3719 ( .A(\CARRYB[4][9] ), .B(\ab[5][9] ), .ZN(n1350) );
  NAND2_X4 U3720 ( .A1(net84948), .A2(net84947), .ZN(n1901) );
  NOR2_X1 U3721 ( .A1(net124723), .A2(net70473), .ZN(\ab[11][16] ) );
  NAND2_X2 U3722 ( .A1(\SUMB[8][15] ), .A2(n1235), .ZN(n2292) );
  NAND2_X4 U3723 ( .A1(n1662), .A2(n1661), .ZN(net80993) );
  NAND3_X4 U3724 ( .A1(n2028), .A2(n2029), .A3(n2030), .ZN(\CARRYB[3][11] ) );
  NAND2_X2 U3725 ( .A1(n1326), .A2(n1327), .ZN(n1328) );
  INV_X4 U3726 ( .A(\ab[4][8] ), .ZN(n1326) );
  INV_X4 U3727 ( .A(\CARRYB[3][8] ), .ZN(n1327) );
  XOR2_X2 U3728 ( .A(n1329), .B(n853), .Z(\SUMB[6][7] ) );
  NAND2_X1 U3729 ( .A1(\CARRYB[5][7] ), .A2(\ab[6][7] ), .ZN(n1330) );
  NAND2_X2 U3731 ( .A1(n29), .A2(\SUMB[5][8] ), .ZN(n1332) );
  NAND3_X4 U3732 ( .A1(n1335), .A2(n1334), .A3(n1333), .ZN(\CARRYB[7][6] ) );
  NAND2_X2 U3733 ( .A1(\ab[9][16] ), .A2(net88704), .ZN(n2305) );
  NOR2_X1 U3734 ( .A1(net70460), .A2(net77948), .ZN(\ab[5][13] ) );
  INV_X4 U3735 ( .A(n621), .ZN(n1761) );
  NAND2_X4 U3736 ( .A1(\ab[21][1] ), .A2(\CARRYB[20][1] ), .ZN(n2162) );
  NAND3_X4 U3737 ( .A1(net80565), .A2(net83296), .A3(net80566), .ZN(
        \CARRYB[16][7] ) );
  NAND2_X4 U3739 ( .A1(n1336), .A2(n1337), .ZN(\SUMB[21][4] ) );
  NAND2_X4 U3740 ( .A1(n2044), .A2(n2045), .ZN(n2047) );
  NAND2_X4 U3741 ( .A1(n1790), .A2(n1791), .ZN(\SUMB[5][19] ) );
  XNOR2_X2 U3742 ( .A(\CARRYB[16][14] ), .B(n1338), .ZN(n1369) );
  OR2_X1 U3743 ( .A1(net70461), .A2(net84698), .ZN(n1338) );
  XNOR2_X2 U3744 ( .A(n1339), .B(n1229), .ZN(\SUMB[4][10] ) );
  NAND3_X2 U3745 ( .A1(n1746), .A2(n1745), .A3(n1744), .ZN(\CARRYB[5][10] ) );
  NAND2_X4 U3746 ( .A1(\ab[2][20] ), .A2(\SUMB[1][21] ), .ZN(n2052) );
  NAND2_X2 U3747 ( .A1(n2197), .A2(n848), .ZN(n1790) );
  XNOR2_X2 U3748 ( .A(\CARRYB[5][15] ), .B(\ab[6][15] ), .ZN(n1695) );
  XNOR2_X2 U3749 ( .A(\CARRYB[8][14] ), .B(\ab[9][14] ), .ZN(n1587) );
  XNOR2_X2 U3750 ( .A(n1340), .B(n1864), .ZN(\SUMB[8][7] ) );
  XNOR2_X2 U3751 ( .A(n165), .B(n1831), .ZN(n1340) );
  INV_X2 U3752 ( .A(\CARRYB[6][9] ), .ZN(n1699) );
  NAND2_X2 U3753 ( .A1(net88704), .A2(\CARRYB[8][16] ), .ZN(n2304) );
  NAND2_X1 U3754 ( .A1(\ab[13][12] ), .A2(\CARRYB[12][12] ), .ZN(n2125) );
  NAND2_X2 U3755 ( .A1(net87683), .A2(\ab[2][17] ), .ZN(n1941) );
  XNOR2_X2 U3756 ( .A(n1342), .B(\SUMB[2][25] ), .ZN(\SUMB[3][24] ) );
  XNOR2_X2 U3757 ( .A(\ab[3][24] ), .B(\CARRYB[2][24] ), .ZN(n1342) );
  INV_X2 U3758 ( .A(\ab[2][17] ), .ZN(net87682) );
  INV_X4 U3759 ( .A(n2109), .ZN(n1346) );
  NAND2_X4 U3760 ( .A1(n1455), .A2(n2071), .ZN(n1585) );
  INV_X4 U3761 ( .A(net93878), .ZN(net85540) );
  XNOR2_X2 U3762 ( .A(n1258), .B(n1350), .ZN(\SUMB[5][9] ) );
  NAND3_X2 U3763 ( .A1(net84297), .A2(net84298), .A3(net84299), .ZN(
        \CARRYB[2][24] ) );
  NAND2_X4 U3764 ( .A1(n1351), .A2(n1352), .ZN(n1354) );
  NAND2_X4 U3765 ( .A1(n1353), .A2(n1354), .ZN(\SUMB[2][15] ) );
  NAND2_X2 U3766 ( .A1(n362), .A2(n1356), .ZN(n1357) );
  NAND2_X4 U3767 ( .A1(n1357), .A2(n1358), .ZN(\SUMB[5][13] ) );
  INV_X4 U3768 ( .A(n362), .ZN(n1355) );
  NAND2_X4 U3769 ( .A1(\SUMB[7][12] ), .A2(\CARRYB[7][11] ), .ZN(n2126) );
  INV_X2 U3770 ( .A(net83151), .ZN(net87573) );
  XNOR2_X2 U3771 ( .A(\SUMB[5][24] ), .B(n1359), .ZN(\SUMB[6][23] ) );
  XNOR2_X2 U3772 ( .A(\ab[6][23] ), .B(\CARRYB[5][23] ), .ZN(n1359) );
  NOR2_X2 U3773 ( .A1(net77868), .A2(n242), .ZN(\ab[1][1] ) );
  XNOR2_X2 U3774 ( .A(n1360), .B(\SUMB[6][24] ), .ZN(\SUMB[7][23] ) );
  XNOR2_X2 U3775 ( .A(\ab[7][23] ), .B(\CARRYB[6][23] ), .ZN(n1360) );
  NAND2_X1 U3776 ( .A1(\CARRYB[13][16] ), .A2(n1250), .ZN(n2227) );
  NAND3_X2 U3777 ( .A1(net80478), .A2(net80479), .A3(net80480), .ZN(
        \CARRYB[14][14] ) );
  NAND2_X1 U3778 ( .A1(\ab[12][16] ), .A2(\SUMB[11][17] ), .ZN(n2308) );
  NAND2_X1 U3779 ( .A1(\CARRYB[11][16] ), .A2(\SUMB[11][17] ), .ZN(n2309) );
  NAND3_X2 U3780 ( .A1(n2056), .A2(n2055), .A3(n2054), .ZN(\CARRYB[3][19] ) );
  INV_X4 U3781 ( .A(n1439), .ZN(n1362) );
  NAND3_X2 U3782 ( .A1(net81205), .A2(net81204), .A3(net81206), .ZN(n1439) );
  NAND2_X4 U3783 ( .A1(net84706), .A2(net84707), .ZN(n1582) );
  NAND2_X4 U3784 ( .A1(net87064), .A2(n1506), .ZN(n1508) );
  INV_X1 U3785 ( .A(\ab[5][12] ), .ZN(net87464) );
  NOR2_X2 U3786 ( .A1(net83784), .A2(net77948), .ZN(\ab[5][12] ) );
  NAND2_X4 U3787 ( .A1(n1364), .A2(n1365), .ZN(\SUMB[21][3] ) );
  INV_X4 U3788 ( .A(n2244), .ZN(n1363) );
  NAND3_X4 U3789 ( .A1(n1801), .A2(n1800), .A3(n1799), .ZN(\CARRYB[23][0] ) );
  NAND2_X2 U3790 ( .A1(\ab[12][2] ), .A2(\CARRYB[11][2] ), .ZN(n1997) );
  NAND3_X4 U3791 ( .A1(n1707), .A2(n1706), .A3(n1705), .ZN(n1500) );
  NAND3_X4 U3792 ( .A1(n1702), .A2(n1704), .A3(n1703), .ZN(\CARRYB[14][5] ) );
  NAND3_X2 U3793 ( .A1(n2037), .A2(n2038), .A3(n2039), .ZN(\CARRYB[17][5] ) );
  NAND3_X4 U3794 ( .A1(n2302), .A2(net79993), .A3(net79992), .ZN(
        \CARRYB[22][4] ) );
  NAND2_X1 U3795 ( .A1(\ab[27][3] ), .A2(n1272), .ZN(net80818) );
  NAND2_X1 U3796 ( .A1(\ab[5][17] ), .A2(\CARRYB[4][17] ), .ZN(n2203) );
  NAND2_X4 U3797 ( .A1(net87309), .A2(net87308), .ZN(n1367) );
  XNOR2_X2 U3798 ( .A(n1370), .B(n1123), .ZN(\SUMB[15][6] ) );
  XNOR2_X2 U3799 ( .A(\CARRYB[14][6] ), .B(\ab[15][6] ), .ZN(n1370) );
  XNOR2_X2 U3800 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .ZN(n1371) );
  NAND2_X4 U3801 ( .A1(n935), .A2(net87136), .ZN(net85979) );
  INV_X2 U3802 ( .A(\ab[13][12] ), .ZN(n1372) );
  INV_X4 U3803 ( .A(n2204), .ZN(n1376) );
  NOR2_X2 U3804 ( .A1(net83784), .A2(net70469), .ZN(\ab[13][12] ) );
  XNOR2_X2 U3805 ( .A(n1936), .B(n863), .ZN(\SUMB[17][4] ) );
  NAND2_X2 U3806 ( .A1(\ab[14][7] ), .A2(\CARRYB[13][7] ), .ZN(net85000) );
  NAND2_X2 U3807 ( .A1(\SUMB[7][16] ), .A2(n858), .ZN(n2254) );
  NAND2_X4 U3808 ( .A1(n1380), .A2(n1381), .ZN(n1383) );
  INV_X4 U3809 ( .A(\ab[17][5] ), .ZN(n1381) );
  NAND2_X4 U3810 ( .A1(\SUMB[20][2] ), .A2(\CARRYB[20][1] ), .ZN(n2163) );
  XNOR2_X2 U3811 ( .A(\CARRYB[5][6] ), .B(\ab[6][6] ), .ZN(n1552) );
  NAND2_X2 U3812 ( .A1(\CARRYB[18][3] ), .A2(n1209), .ZN(n2273) );
  NAND2_X2 U3813 ( .A1(\ab[1][10] ), .A2(\ab[0][11] ), .ZN(n2332) );
  XNOR2_X2 U3814 ( .A(n1384), .B(n1189), .ZN(\SUMB[18][4] ) );
  XNOR2_X2 U3815 ( .A(\CARRYB[17][4] ), .B(\ab[18][4] ), .ZN(n1384) );
  NAND3_X2 U3816 ( .A1(net84926), .A2(net84925), .A3(net84924), .ZN(
        \CARRYB[3][6] ) );
  NAND2_X2 U3817 ( .A1(net87003), .A2(net87004), .ZN(n1385) );
  NAND2_X1 U3818 ( .A1(\CARRYB[16][11] ), .A2(\ab[17][11] ), .ZN(net87010) );
  NAND2_X2 U3819 ( .A1(\ab[17][11] ), .A2(\SUMB[16][12] ), .ZN(net87012) );
  INV_X4 U3820 ( .A(n1608), .ZN(n1386) );
  NOR2_X2 U3821 ( .A1(net83784), .A2(net70463), .ZN(\ab[16][12] ) );
  NAND2_X4 U3822 ( .A1(n2046), .A2(n2047), .ZN(n2112) );
  NAND2_X4 U3823 ( .A1(net83121), .A2(n1759), .ZN(net80264) );
  NAND2_X4 U3824 ( .A1(n1515), .A2(n1964), .ZN(n1880) );
  NAND2_X2 U3825 ( .A1(n1453), .A2(n1454), .ZN(n1455) );
  NOR2_X1 U3826 ( .A1(net124723), .A2(net77932), .ZN(\ab[7][16] ) );
  NOR2_X4 U3827 ( .A1(net124723), .A2(net77926), .ZN(\ab[8][16] ) );
  NOR2_X4 U3828 ( .A1(net124723), .A2(net70471), .ZN(\ab[12][16] ) );
  NAND2_X4 U3829 ( .A1(n1859), .A2(n1860), .ZN(n2109) );
  NAND2_X2 U3830 ( .A1(\ab[3][8] ), .A2(\CARRYB[2][8] ), .ZN(n1905) );
  XNOR2_X2 U3831 ( .A(\CARRYB[2][8] ), .B(\ab[3][8] ), .ZN(n1452) );
  NAND3_X4 U3832 ( .A1(net80805), .A2(net80806), .A3(n2164), .ZN(
        \CARRYB[10][16] ) );
  NAND2_X4 U3833 ( .A1(\CARRYB[26][0] ), .A2(\ab[27][0] ), .ZN(net80767) );
  NAND3_X4 U3834 ( .A1(n2027), .A2(net81535), .A3(net81533), .ZN(
        \CARRYB[26][0] ) );
  NAND3_X4 U3835 ( .A1(n2127), .A2(n2126), .A3(n2128), .ZN(\CARRYB[8][11] ) );
  NAND3_X4 U3836 ( .A1(n1982), .A2(n1981), .A3(n1980), .ZN(\CARRYB[5][13] ) );
  NAND2_X1 U3837 ( .A1(\ab[19][8] ), .A2(\CARRYB[18][8] ), .ZN(n1392) );
  NAND3_X4 U3838 ( .A1(n1395), .A2(n1394), .A3(n1393), .ZN(\CARRYB[4][10] ) );
  NAND2_X2 U3839 ( .A1(n572), .A2(\ab[5][9] ), .ZN(n1397) );
  NAND3_X2 U3840 ( .A1(n2077), .A2(n2078), .A3(n2079), .ZN(n1425) );
  XNOR2_X2 U3841 ( .A(n128), .B(n1399), .ZN(\SUMB[3][10] ) );
  NAND2_X2 U3842 ( .A1(\ab[3][21] ), .A2(\SUMB[2][22] ), .ZN(n1934) );
  NAND2_X2 U3843 ( .A1(n6), .A2(\SUMB[16][8] ), .ZN(net81267) );
  NAND2_X4 U3844 ( .A1(net86697), .A2(net86698), .ZN(n1400) );
  NAND2_X4 U3845 ( .A1(net86699), .A2(n1400), .ZN(net81815) );
  INV_X4 U3846 ( .A(\CARRYB[24][5] ), .ZN(net86698) );
  NAND2_X4 U3847 ( .A1(net86704), .A2(n1401), .ZN(\SUMB[21][7] ) );
  NAND2_X2 U3848 ( .A1(\ab[12][6] ), .A2(\SUMB[11][7] ), .ZN(n1918) );
  XOR2_X2 U3849 ( .A(\CARRYB[5][1] ), .B(\ab[6][1] ), .Z(n1402) );
  XOR2_X2 U3850 ( .A(\SUMB[5][2] ), .B(n1402), .Z(\SUMB[6][1] ) );
  NAND2_X2 U3851 ( .A1(\CARRYB[5][1] ), .A2(\SUMB[5][2] ), .ZN(n1403) );
  NAND2_X2 U3852 ( .A1(\ab[6][1] ), .A2(\SUMB[5][2] ), .ZN(n1404) );
  NAND2_X2 U3853 ( .A1(\ab[6][1] ), .A2(\CARRYB[5][1] ), .ZN(n1405) );
  NAND3_X2 U3854 ( .A1(n1403), .A2(n1404), .A3(n1405), .ZN(\CARRYB[6][1] ) );
  XOR2_X1 U3855 ( .A(\CARRYB[15][0] ), .B(\ab[16][0] ), .Z(net86649) );
  NAND2_X2 U3856 ( .A1(\ab[16][0] ), .A2(\CARRYB[15][0] ), .ZN(n1406) );
  XOR2_X1 U3857 ( .A(net86653), .B(\CARRYB[16][0] ), .Z(PRODUCT[17]) );
  NAND2_X2 U3858 ( .A1(\ab[17][0] ), .A2(\CARRYB[16][0] ), .ZN(n1407) );
  NAND3_X2 U3859 ( .A1(net86654), .A2(n1407), .A3(net86656), .ZN(
        \CARRYB[17][0] ) );
  XOR2_X1 U3860 ( .A(\SUMB[14][1] ), .B(\ab[15][0] ), .Z(n1408) );
  XOR2_X2 U3861 ( .A(n846), .B(n1408), .Z(PRODUCT[15]) );
  NAND2_X2 U3862 ( .A1(\CARRYB[14][0] ), .A2(\ab[15][0] ), .ZN(n1410) );
  NOR2_X1 U3863 ( .A1(net77866), .A2(net77938), .ZN(\ab[6][1] ) );
  NOR2_X2 U3864 ( .A1(net77860), .A2(net70465), .ZN(\ab[15][0] ) );
  NAND3_X4 U3865 ( .A1(n2211), .A2(n2212), .A3(n2213), .ZN(\CARRYB[20][6] ) );
  NAND2_X2 U3866 ( .A1(\ab[20][6] ), .A2(\CARRYB[19][6] ), .ZN(n2213) );
  NAND3_X4 U3867 ( .A1(n2160), .A2(net80852), .A3(net80850), .ZN(
        \CARRYB[20][1] ) );
  NAND3_X2 U3868 ( .A1(n2209), .A2(n2210), .A3(n2208), .ZN(\CARRYB[7][15] ) );
  NAND2_X4 U3869 ( .A1(net86630), .A2(n1412), .ZN(\SUMB[14][13] ) );
  NOR2_X2 U3870 ( .A1(net77900), .A2(n242), .ZN(\ab[1][5] ) );
  NOR2_X2 U3871 ( .A1(net70436), .A2(net83263), .ZN(\ab[1][0] ) );
  NAND2_X1 U3872 ( .A1(\ab[3][19] ), .A2(\CARRYB[2][19] ), .ZN(n2054) );
  NAND2_X4 U3873 ( .A1(n1488), .A2(n1489), .ZN(net83535) );
  XNOR2_X2 U3874 ( .A(n1413), .B(n2142), .ZN(\SUMB[20][11] ) );
  NAND2_X4 U3875 ( .A1(\ab[0][5] ), .A2(\ab[1][4] ), .ZN(n2327) );
  NAND2_X1 U3876 ( .A1(\CARRYB[8][21] ), .A2(\SUMB[8][22] ), .ZN(n1688) );
  NAND3_X4 U3877 ( .A1(n2293), .A2(n2292), .A3(n2294), .ZN(\CARRYB[9][14] ) );
  NAND3_X4 U3878 ( .A1(net80247), .A2(net80248), .A3(net80246), .ZN(
        \CARRYB[10][13] ) );
  NOR2_X2 U3879 ( .A1(net77886), .A2(net70459), .ZN(\ab[18][3] ) );
  NAND3_X4 U3880 ( .A1(n2106), .A2(n2108), .A3(n2107), .ZN(\CARRYB[17][3] ) );
  NAND2_X2 U3881 ( .A1(\ab[6][12] ), .A2(\CARRYB[5][12] ), .ZN(n1983) );
  INV_X1 U3882 ( .A(\ab[6][12] ), .ZN(net86440) );
  NOR2_X2 U3883 ( .A1(net83784), .A2(net77940), .ZN(\ab[6][12] ) );
  INV_X4 U3884 ( .A(n1732), .ZN(n1444) );
  NAND2_X4 U3885 ( .A1(n1190), .A2(\ab[20][6] ), .ZN(n2212) );
  INV_X8 U3886 ( .A(\CARRYB[24][4] ), .ZN(net82551) );
  XNOR2_X2 U3887 ( .A(net86427), .B(net88656), .ZN(\SUMB[26][1] ) );
  NAND2_X4 U3888 ( .A1(\CARRYB[24][4] ), .A2(\ab[25][4] ), .ZN(n1854) );
  NAND3_X2 U3889 ( .A1(net86412), .A2(net86413), .A3(net86414), .ZN(
        \CARRYB[23][7] ) );
  NAND2_X2 U3890 ( .A1(n2135), .A2(n1420), .ZN(n1421) );
  NAND2_X4 U3891 ( .A1(n1421), .A2(n1422), .ZN(\SUMB[4][19] ) );
  INV_X4 U3892 ( .A(n2135), .ZN(n1419) );
  NAND2_X2 U3893 ( .A1(n708), .A2(\SUMB[4][19] ), .ZN(n1577) );
  INV_X4 U3894 ( .A(\SUMB[4][19] ), .ZN(n1576) );
  NAND3_X4 U3895 ( .A1(n2085), .A2(n2084), .A3(n2083), .ZN(\CARRYB[8][9] ) );
  NOR2_X4 U3896 ( .A1(net70472), .A2(net80409), .ZN(\ab[1][19] ) );
  NOR2_X4 U3897 ( .A1(net86565), .A2(net77948), .ZN(\ab[5][19] ) );
  INV_X8 U3898 ( .A(net81080), .ZN(net80727) );
  NOR2_X4 U3899 ( .A1(net70472), .A2(net82149), .ZN(net81354) );
  XNOR2_X2 U3900 ( .A(\SUMB[16][14] ), .B(n1423), .ZN(\SUMB[17][13] ) );
  XNOR2_X2 U3901 ( .A(\ab[17][13] ), .B(\CARRYB[16][13] ), .ZN(n1423) );
  NOR2_X2 U3902 ( .A1(net70452), .A2(net77970), .ZN(\ab[2][9] ) );
  NAND2_X2 U3903 ( .A1(\ab[8][9] ), .A2(\CARRYB[7][9] ), .ZN(n2083) );
  NOR2_X4 U3904 ( .A1(net123000), .A2(net70491), .ZN(\ab[2][17] ) );
  XOR2_X1 U3905 ( .A(\CARRYB[17][0] ), .B(\ab[18][0] ), .Z(n1808) );
  NAND3_X2 U3906 ( .A1(n2150), .A2(n2151), .A3(n2152), .ZN(\CARRYB[14][4] ) );
  NAND2_X2 U3907 ( .A1(\CARRYB[15][5] ), .A2(\SUMB[15][6] ), .ZN(n2073) );
  INV_X2 U3908 ( .A(\SUMB[2][9] ), .ZN(n1426) );
  XNOR2_X2 U3909 ( .A(n1428), .B(\SUMB[2][10] ), .ZN(\SUMB[3][9] ) );
  XNOR2_X2 U3910 ( .A(n1246), .B(\ab[3][9] ), .ZN(n1428) );
  NAND3_X4 U3911 ( .A1(net81513), .A2(net81514), .A3(net81515), .ZN(
        \CARRYB[3][13] ) );
  NAND3_X2 U3912 ( .A1(net86158), .A2(net86159), .A3(n1019), .ZN(
        \CARRYB[12][12] ) );
  NAND2_X4 U3913 ( .A1(n1433), .A2(n1434), .ZN(\SUMB[3][20] ) );
  INV_X4 U3914 ( .A(n1765), .ZN(n1431) );
  NAND2_X4 U3915 ( .A1(\ab[4][19] ), .A2(\SUMB[3][20] ), .ZN(n2137) );
  NAND3_X4 U3916 ( .A1(n2237), .A2(n2239), .A3(n2238), .ZN(\CARRYB[4][20] ) );
  XNOR2_X2 U3917 ( .A(\SUMB[4][22] ), .B(n1435), .ZN(\SUMB[5][21] ) );
  NAND3_X2 U3918 ( .A1(n1964), .A2(n1966), .A3(n1965), .ZN(\CARRYB[5][8] ) );
  NAND2_X2 U3919 ( .A1(\CARRYB[14][6] ), .A2(\SUMB[14][7] ), .ZN(n1436) );
  NAND3_X2 U3920 ( .A1(n1437), .A2(n1436), .A3(n1438), .ZN(\CARRYB[15][6] ) );
  NAND3_X2 U3921 ( .A1(net86170), .A2(net86171), .A3(net86172), .ZN(
        \CARRYB[2][14] ) );
  NAND3_X4 U3922 ( .A1(n1974), .A2(n1976), .A3(n1975), .ZN(\CARRYB[14][6] ) );
  NOR2_X2 U3923 ( .A1(net77908), .A2(net70465), .ZN(\ab[15][6] ) );
  NOR2_X4 U3924 ( .A1(net84698), .A2(net70491), .ZN(\ab[2][14] ) );
  NAND2_X4 U3925 ( .A1(n1460), .A2(n1459), .ZN(\SUMB[11][5] ) );
  NAND2_X2 U3926 ( .A1(\CARRYB[4][7] ), .A2(\SUMB[4][8] ), .ZN(n1948) );
  NAND2_X2 U3927 ( .A1(\ab[5][7] ), .A2(\SUMB[4][8] ), .ZN(n1947) );
  NAND2_X4 U3928 ( .A1(n1858), .A2(n1857), .ZN(n1860) );
  NAND3_X2 U3929 ( .A1(n1839), .A2(n1840), .A3(n1841), .ZN(\CARRYB[10][15] )
         );
  NAND2_X1 U3930 ( .A1(\SUMB[5][6] ), .A2(\CARRYB[5][5] ), .ZN(n1440) );
  NAND2_X1 U3931 ( .A1(\SUMB[5][6] ), .A2(\ab[6][5] ), .ZN(n1441) );
  NAND2_X1 U3932 ( .A1(\ab[6][5] ), .A2(\CARRYB[5][5] ), .ZN(n1442) );
  NAND3_X2 U3933 ( .A1(n1440), .A2(n1441), .A3(n1442), .ZN(\CARRYB[6][5] ) );
  NOR2_X1 U3934 ( .A1(net77898), .A2(net77938), .ZN(\ab[6][5] ) );
  NAND2_X4 U3935 ( .A1(n1763), .A2(n1762), .ZN(n2001) );
  INV_X1 U3937 ( .A(\ab[7][7] ), .ZN(n1499) );
  NAND2_X4 U3938 ( .A1(n1556), .A2(n1557), .ZN(n1559) );
  NAND2_X4 U3939 ( .A1(n1444), .A2(n1445), .ZN(n1447) );
  NAND2_X4 U3940 ( .A1(n1447), .A2(n1446), .ZN(\SUMB[13][7] ) );
  XNOR2_X2 U3941 ( .A(\CARRYB[14][14] ), .B(\ab[15][14] ), .ZN(net86054) );
  NAND2_X4 U3942 ( .A1(\ab[21][0] ), .A2(n1237), .ZN(n1807) );
  NAND2_X2 U3943 ( .A1(\CARRYB[17][0] ), .A2(\SUMB[17][1] ), .ZN(n1811) );
  NAND2_X2 U3944 ( .A1(\ab[18][0] ), .A2(\CARRYB[17][0] ), .ZN(n1809) );
  XOR2_X2 U3945 ( .A(\SUMB[4][2] ), .B(\ab[5][1] ), .Z(n1481) );
  XNOR2_X2 U3946 ( .A(n1448), .B(n1206), .ZN(\SUMB[9][5] ) );
  NAND2_X2 U3947 ( .A1(n194), .A2(n2060), .ZN(n1459) );
  NAND2_X2 U3948 ( .A1(n1279), .A2(n1449), .ZN(n1450) );
  NAND2_X4 U3949 ( .A1(n1450), .A2(n1451), .ZN(\SUMB[16][8] ) );
  XNOR2_X2 U3950 ( .A(n1452), .B(n1427), .ZN(\SUMB[3][8] ) );
  NAND2_X2 U3951 ( .A1(n1514), .A2(n1513), .ZN(n1515) );
  INV_X1 U3952 ( .A(\ab[16][5] ), .ZN(n1453) );
  NAND2_X2 U3953 ( .A1(\ab[4][9] ), .A2(\SUMB[3][10] ), .ZN(n1962) );
  NAND3_X2 U3954 ( .A1(net81034), .A2(net81035), .A3(net81033), .ZN(
        \CARRYB[20][9] ) );
  NAND2_X2 U3955 ( .A1(\CARRYB[17][9] ), .A2(\ab[18][9] ), .ZN(n1554) );
  XNOR2_X2 U3956 ( .A(n1457), .B(\SUMB[1][23] ), .ZN(\SUMB[2][22] ) );
  NOR2_X2 U3957 ( .A1(net70491), .A2(net70478), .ZN(\ab[2][22] ) );
  NAND2_X2 U3958 ( .A1(\SUMB[23][6] ), .A2(n1251), .ZN(net79968) );
  INV_X4 U3959 ( .A(\CARRYB[23][5] ), .ZN(n2155) );
  NAND2_X4 U3960 ( .A1(\SUMB[1][12] ), .A2(\CARRYB[1][11] ), .ZN(n1644) );
  NAND3_X4 U3961 ( .A1(n1777), .A2(n1779), .A3(n1778), .ZN(\CARRYB[11][7] ) );
  XNOR2_X2 U3962 ( .A(n1461), .B(n1259), .ZN(\SUMB[4][9] ) );
  XNOR2_X2 U3963 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .ZN(n1461) );
  NAND2_X2 U3964 ( .A1(n173), .A2(\ab[11][7] ), .ZN(n1777) );
  XOR2_X2 U3965 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .Z(n1462) );
  XOR2_X2 U3966 ( .A(n1462), .B(\SUMB[10][19] ), .Z(\SUMB[11][18] ) );
  NAND2_X1 U3967 ( .A1(\ab[11][18] ), .A2(\CARRYB[10][18] ), .ZN(n1463) );
  NAND2_X1 U3968 ( .A1(\ab[11][18] ), .A2(\SUMB[10][19] ), .ZN(n1464) );
  NAND2_X1 U3969 ( .A1(\CARRYB[10][18] ), .A2(\SUMB[10][19] ), .ZN(n1465) );
  NAND3_X2 U3970 ( .A1(n1463), .A2(n1464), .A3(n1465), .ZN(\CARRYB[11][18] )
         );
  NAND2_X1 U3971 ( .A1(\CARRYB[11][17] ), .A2(\ab[12][17] ), .ZN(n1466) );
  NAND2_X1 U3972 ( .A1(\CARRYB[11][17] ), .A2(\SUMB[11][18] ), .ZN(n1467) );
  XNOR2_X2 U3973 ( .A(n1469), .B(\SUMB[3][25] ), .ZN(\SUMB[4][24] ) );
  XNOR2_X2 U3974 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .ZN(n1469) );
  NAND2_X2 U3975 ( .A1(\ab[11][4] ), .A2(n2370), .ZN(n1834) );
  NAND2_X2 U3976 ( .A1(\SUMB[9][2] ), .A2(\ab[10][1] ), .ZN(n1472) );
  NAND2_X2 U3977 ( .A1(\SUMB[9][2] ), .A2(\CARRYB[9][1] ), .ZN(n1473) );
  NAND3_X2 U3978 ( .A1(n2289), .A2(n2290), .A3(n2291), .ZN(\CARRYB[9][19] ) );
  NAND3_X2 U3979 ( .A1(n2072), .A2(n2073), .A3(n2071), .ZN(\CARRYB[16][5] ) );
  NOR2_X1 U3980 ( .A1(net70454), .A2(net119855), .ZN(\ab[4][10] ) );
  NAND2_X1 U3981 ( .A1(\ab[5][23] ), .A2(\SUMB[4][24] ), .ZN(n1959) );
  XOR2_X2 U3982 ( .A(\CARRYB[1][3] ), .B(\ab[2][3] ), .Z(n1474) );
  XOR2_X2 U3983 ( .A(\SUMB[1][4] ), .B(n1474), .Z(\SUMB[2][3] ) );
  NAND2_X1 U3984 ( .A1(\CARRYB[1][3] ), .A2(\SUMB[1][4] ), .ZN(n1475) );
  NAND2_X2 U3985 ( .A1(\ab[2][3] ), .A2(\SUMB[1][4] ), .ZN(n1476) );
  NAND2_X1 U3986 ( .A1(\ab[2][3] ), .A2(\CARRYB[1][3] ), .ZN(n1477) );
  NAND3_X2 U3987 ( .A1(n1475), .A2(n1476), .A3(n1477), .ZN(\CARRYB[2][3] ) );
  NAND2_X1 U3988 ( .A1(\ab[4][1] ), .A2(\CARRYB[3][1] ), .ZN(n1478) );
  NAND2_X2 U3989 ( .A1(\ab[4][1] ), .A2(\SUMB[3][2] ), .ZN(n1479) );
  NAND2_X1 U3990 ( .A1(\CARRYB[3][1] ), .A2(\SUMB[3][2] ), .ZN(n1480) );
  NAND3_X2 U3991 ( .A1(n1478), .A2(n1479), .A3(n1480), .ZN(\CARRYB[4][1] ) );
  XOR2_X2 U3992 ( .A(n1481), .B(\CARRYB[4][1] ), .Z(\SUMB[5][1] ) );
  NAND2_X1 U3993 ( .A1(\ab[5][1] ), .A2(\SUMB[4][2] ), .ZN(n1482) );
  NAND2_X2 U3994 ( .A1(\ab[5][1] ), .A2(\CARRYB[4][1] ), .ZN(n1483) );
  NAND2_X1 U3995 ( .A1(\SUMB[4][2] ), .A2(\CARRYB[4][1] ), .ZN(n1484) );
  NAND3_X2 U3996 ( .A1(n1482), .A2(n1483), .A3(n1484), .ZN(\CARRYB[5][1] ) );
  NOR2_X2 U3997 ( .A1(net77882), .A2(net77970), .ZN(\ab[2][3] ) );
  XNOR2_X2 U3998 ( .A(net85734), .B(net85036), .ZN(\SUMB[3][7] ) );
  NAND3_X4 U3999 ( .A1(n1999), .A2(n1998), .A3(n2000), .ZN(\CARRYB[13][6] ) );
  XNOR2_X2 U4000 ( .A(n1485), .B(\SUMB[1][12] ), .ZN(\SUMB[2][11] ) );
  NAND2_X2 U4001 ( .A1(\CARRYB[8][5] ), .A2(\SUMB[8][6] ), .ZN(n1785) );
  INV_X2 U4002 ( .A(\ab[14][12] ), .ZN(n1487) );
  NOR2_X2 U4003 ( .A1(net83784), .A2(net70467), .ZN(\ab[14][12] ) );
  NAND2_X4 U4004 ( .A1(n2116), .A2(n1696), .ZN(net81663) );
  NAND3_X2 U4005 ( .A1(n2201), .A2(n2202), .A3(n2203), .ZN(n1490) );
  NAND2_X2 U4006 ( .A1(\CARRYB[3][18] ), .A2(n1693), .ZN(n1493) );
  NAND2_X4 U4007 ( .A1(n1491), .A2(n1492), .ZN(n1494) );
  NAND2_X4 U4008 ( .A1(n1493), .A2(n1494), .ZN(\SUMB[4][18] ) );
  INV_X4 U4009 ( .A(n1693), .ZN(n1491) );
  INV_X2 U4010 ( .A(\CARRYB[3][18] ), .ZN(n1492) );
  NOR2_X4 U4011 ( .A1(net77920), .A2(net70451), .ZN(\ab[22][8] ) );
  XNOR2_X2 U4012 ( .A(\SUMB[5][4] ), .B(n1495), .ZN(\SUMB[6][3] ) );
  XNOR2_X2 U4013 ( .A(\CARRYB[5][3] ), .B(\ab[6][3] ), .ZN(n1495) );
  NAND2_X4 U4014 ( .A1(n1496), .A2(n1497), .ZN(\SUMB[6][16] ) );
  NAND2_X2 U4015 ( .A1(n397), .A2(\SUMB[1][19] ), .ZN(net85602) );
  NAND2_X4 U4016 ( .A1(n287), .A2(n1498), .ZN(net85603) );
  NAND3_X2 U4017 ( .A1(n1922), .A2(n1921), .A3(n1920), .ZN(n1501) );
  XNOR2_X2 U4018 ( .A(n1502), .B(\SUMB[15][15] ), .ZN(\SUMB[16][14] ) );
  XNOR2_X2 U4019 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .ZN(n1502) );
  NAND2_X4 U4020 ( .A1(n1816), .A2(n1817), .ZN(n1819) );
  NAND2_X2 U4021 ( .A1(\SUMB[12][5] ), .A2(\ab[13][4] ), .ZN(n1640) );
  NAND2_X2 U4022 ( .A1(\ab[8][6] ), .A2(\CARRYB[7][6] ), .ZN(n1825) );
  XNOR2_X2 U4023 ( .A(\CARRYB[14][4] ), .B(\ab[15][4] ), .ZN(n1581) );
  NAND3_X4 U4024 ( .A1(n2042), .A2(n2041), .A3(n2040), .ZN(\CARRYB[18][4] ) );
  NAND2_X4 U4025 ( .A1(net85457), .A2(n1505), .ZN(\SUMB[12][11] ) );
  NAND2_X2 U4026 ( .A1(n1937), .A2(net85465), .ZN(n1507) );
  NAND2_X4 U4027 ( .A1(n1509), .A2(net85469), .ZN(n1511) );
  INV_X4 U4028 ( .A(n1943), .ZN(n1509) );
  NAND2_X4 U4029 ( .A1(net84825), .A2(net84826), .ZN(net83866) );
  XNOR2_X2 U4030 ( .A(\SUMB[21][10] ), .B(n1512), .ZN(\SUMB[22][9] ) );
  XOR2_X2 U4031 ( .A(\CARRYB[21][9] ), .B(n1929), .Z(n1512) );
  NAND2_X2 U4032 ( .A1(\ab[2][20] ), .A2(\CARRYB[1][20] ), .ZN(n2051) );
  INV_X2 U4033 ( .A(\ab[5][8] ), .ZN(n1513) );
  NAND3_X4 U4034 ( .A1(n2076), .A2(n2075), .A3(n2074), .ZN(\CARRYB[17][4] ) );
  NOR2_X4 U4035 ( .A1(net70452), .A2(net86101), .ZN(\ab[1][9] ) );
  NAND2_X2 U4036 ( .A1(n1518), .A2(n1517), .ZN(n2331) );
  INV_X4 U4037 ( .A(\ab[1][9] ), .ZN(n1516) );
  NAND2_X2 U4038 ( .A1(\ab[7][5] ), .A2(\CARRYB[6][5] ), .ZN(n1520) );
  NAND3_X2 U4039 ( .A1(n1519), .A2(n1520), .A3(n1521), .ZN(\CARRYB[7][5] ) );
  NOR2_X1 U4040 ( .A1(net77898), .A2(net77930), .ZN(\ab[7][5] ) );
  NAND2_X4 U4041 ( .A1(n1523), .A2(n1522), .ZN(\SUMB[11][10] ) );
  NAND2_X4 U4042 ( .A1(\SUMB[12][12] ), .A2(net121285), .ZN(net82159) );
  NAND2_X1 U4043 ( .A1(\ab[14][12] ), .A2(\CARRYB[13][12] ), .ZN(n2122) );
  NAND3_X2 U4044 ( .A1(n2201), .A2(n2202), .A3(n2203), .ZN(\CARRYB[5][17] ) );
  NAND2_X4 U4045 ( .A1(n1524), .A2(n1525), .ZN(n1527) );
  NAND2_X4 U4046 ( .A1(n1527), .A2(n1526), .ZN(\SUMB[2][19] ) );
  INV_X1 U4047 ( .A(\ab[2][19] ), .ZN(n1525) );
  INV_X4 U4048 ( .A(n1528), .ZN(n1529) );
  XNOR2_X2 U4049 ( .A(n1530), .B(\CARRYB[12][4] ), .ZN(n1635) );
  XOR2_X2 U4050 ( .A(\CARRYB[8][22] ), .B(\ab[9][22] ), .Z(n1531) );
  XOR2_X2 U4051 ( .A(\SUMB[8][23] ), .B(n1531), .Z(\SUMB[9][22] ) );
  XOR2_X2 U4052 ( .A(\SUMB[13][18] ), .B(n1532), .Z(\SUMB[14][17] ) );
  INV_X1 U4053 ( .A(\ab[27][3] ), .ZN(n1534) );
  NAND2_X2 U4054 ( .A1(net81052), .A2(n2116), .ZN(n1537) );
  NAND2_X4 U4055 ( .A1(n1538), .A2(net81053), .ZN(\CARRYB[26][3] ) );
  INV_X4 U4056 ( .A(n1537), .ZN(n1538) );
  NOR2_X4 U4057 ( .A1(net77886), .A2(net70441), .ZN(\ab[27][3] ) );
  INV_X2 U4058 ( .A(n2345), .ZN(\CARRYB[1][22] ) );
  XNOR2_X2 U4059 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .ZN(n1539) );
  INV_X4 U4060 ( .A(n1845), .ZN(n1540) );
  NAND2_X2 U4061 ( .A1(\CARRYB[6][12] ), .A2(\ab[7][12] ), .ZN(n1544) );
  INV_X2 U4062 ( .A(\ab[5][13] ), .ZN(n1845) );
  INV_X1 U4063 ( .A(n1770), .ZN(n1545) );
  NAND2_X2 U4064 ( .A1(\ab[3][18] ), .A2(\CARRYB[2][18] ), .ZN(n1548) );
  NAND2_X2 U4065 ( .A1(n1546), .A2(n1547), .ZN(n1549) );
  NAND3_X4 U4066 ( .A1(n1713), .A2(n1712), .A3(n1711), .ZN(\CARRYB[2][18] ) );
  NAND2_X2 U4067 ( .A1(\ab[19][4] ), .A2(\CARRYB[18][4] ), .ZN(n2234) );
  NAND3_X2 U4068 ( .A1(net80796), .A2(net80795), .A3(net80794), .ZN(
        \CARRYB[5][22] ) );
  INV_X4 U4069 ( .A(n1792), .ZN(n1556) );
  NAND2_X2 U4070 ( .A1(n1301), .A2(net90433), .ZN(n2115) );
  NAND2_X2 U4071 ( .A1(n1501), .A2(\SUMB[13][6] ), .ZN(n1704) );
  NAND2_X2 U4072 ( .A1(\ab[11][7] ), .A2(\SUMB[10][8] ), .ZN(n1778) );
  NAND2_X2 U4073 ( .A1(\CARRYB[2][8] ), .A2(n1427), .ZN(n1907) );
  NAND2_X2 U4074 ( .A1(\CARRYB[2][24] ), .A2(\SUMB[2][25] ), .ZN(n2170) );
  XNOR2_X2 U4075 ( .A(n1550), .B(\SUMB[9][21] ), .ZN(\SUMB[10][20] ) );
  XNOR2_X2 U4076 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .ZN(n1550) );
  NAND2_X2 U4077 ( .A1(\ab[16][8] ), .A2(\CARRYB[15][8] ), .ZN(n2299) );
  NAND2_X4 U4078 ( .A1(n1616), .A2(n2010), .ZN(n1943) );
  NOR2_X4 U4079 ( .A1(net70454), .A2(net77970), .ZN(\ab[2][10] ) );
  NAND2_X2 U4080 ( .A1(\SUMB[4][9] ), .A2(\ab[5][8] ), .ZN(n1965) );
  NOR2_X4 U4081 ( .A1(net70456), .A2(net77970), .ZN(\ab[2][11] ) );
  NAND2_X4 U4082 ( .A1(\SUMB[1][12] ), .A2(n289), .ZN(n1643) );
  NAND2_X2 U4083 ( .A1(\SUMB[3][9] ), .A2(\CARRYB[3][8] ), .ZN(n1946) );
  XOR2_X2 U4084 ( .A(\SUMB[9][22] ), .B(n2321), .Z(\SUMB[10][21] ) );
  NAND3_X4 U4085 ( .A1(n1643), .A2(n1644), .A3(n1642), .ZN(\CARRYB[2][11] ) );
  NAND2_X2 U4086 ( .A1(n1501), .A2(\ab[14][5] ), .ZN(n1702) );
  NAND3_X2 U4087 ( .A1(n2266), .A2(n2267), .A3(n2268), .ZN(\CARRYB[7][23] ) );
  NAND3_X2 U4088 ( .A1(n2276), .A2(n2277), .A3(n2278), .ZN(\CARRYB[4][21] ) );
  NAND2_X2 U4089 ( .A1(\ab[5][20] ), .A2(\SUMB[4][21] ), .ZN(n1884) );
  NAND3_X4 U4090 ( .A1(n2232), .A2(n2233), .A3(n2231), .ZN(\CARRYB[18][5] ) );
  NAND2_X4 U4091 ( .A1(n1818), .A2(n1819), .ZN(n2135) );
  NAND2_X4 U4092 ( .A1(n1554), .A2(n1555), .ZN(net81782) );
  XNOR2_X2 U4093 ( .A(\CARRYB[13][7] ), .B(\ab[14][7] ), .ZN(n1553) );
  NOR2_X1 U4094 ( .A1(net70452), .A2(net77956), .ZN(\ab[4][9] ) );
  NOR2_X1 U4095 ( .A1(net85716), .A2(net70465), .ZN(\ab[15][11] ) );
  NAND2_X4 U4096 ( .A1(net83850), .A2(net85017), .ZN(n1555) );
  INV_X1 U4097 ( .A(\ab[18][9] ), .ZN(net85017) );
  NAND3_X4 U4098 ( .A1(net80813), .A2(net80812), .A3(net80814), .ZN(
        \CARRYB[17][9] ) );
  INV_X4 U4099 ( .A(n2343), .ZN(\CARRYB[1][21] ) );
  NAND3_X2 U4100 ( .A1(net85000), .A2(net84999), .A3(net84998), .ZN(
        \CARRYB[14][7] ) );
  NOR2_X1 U4101 ( .A1(net77914), .A2(net70467), .ZN(\ab[14][7] ) );
  NAND3_X4 U4102 ( .A1(n2024), .A2(n2023), .A3(n2022), .ZN(\CARRYB[13][7] ) );
  NAND2_X4 U4103 ( .A1(n1558), .A2(n1559), .ZN(\SUMB[3][14] ) );
  XNOR2_X2 U4104 ( .A(\CARRYB[13][5] ), .B(\ab[14][5] ), .ZN(n1584) );
  NAND2_X2 U4105 ( .A1(\CARRYB[13][6] ), .A2(\ab[14][6] ), .ZN(n1974) );
  NAND2_X2 U4106 ( .A1(\CARRYB[7][8] ), .A2(\ab[8][8] ), .ZN(n2004) );
  XOR2_X2 U4107 ( .A(\CARRYB[5][25] ), .B(\ab[6][25] ), .Z(n1560) );
  XOR2_X2 U4108 ( .A(\SUMB[5][26] ), .B(n1560), .Z(\SUMB[6][25] ) );
  XOR2_X2 U4109 ( .A(\CARRYB[4][26] ), .B(\ab[5][26] ), .Z(n1561) );
  XOR2_X2 U4110 ( .A(\SUMB[4][27] ), .B(n1561), .Z(\SUMB[5][26] ) );
  NOR2_X1 U4111 ( .A1(net77940), .A2(net82239), .ZN(\ab[6][25] ) );
  NOR2_X1 U4112 ( .A1(net77948), .A2(net70486), .ZN(\ab[5][26] ) );
  NAND2_X4 U4113 ( .A1(net84212), .A2(net84211), .ZN(n1937) );
  XNOR2_X2 U4114 ( .A(n1649), .B(\SUMB[3][8] ), .ZN(\SUMB[4][7] ) );
  NAND3_X4 U4115 ( .A1(net81069), .A2(net81068), .A3(net81067), .ZN(
        \CARRYB[19][6] ) );
  NAND2_X2 U4116 ( .A1(\ab[6][3] ), .A2(\SUMB[5][4] ), .ZN(n1565) );
  NAND2_X2 U4117 ( .A1(\CARRYB[23][0] ), .A2(n23), .ZN(n1568) );
  NOR2_X1 U4118 ( .A1(net77886), .A2(net77938), .ZN(\ab[6][3] ) );
  NOR2_X2 U4119 ( .A1(net77858), .A2(net70447), .ZN(\ab[24][0] ) );
  NOR2_X2 U4120 ( .A1(net70492), .A2(net83263), .ZN(\ab[1][29] ) );
  NAND2_X2 U4121 ( .A1(\ab[0][22] ), .A2(\ab[1][21] ), .ZN(n2343) );
  NAND2_X2 U4122 ( .A1(\ab[22][0] ), .A2(\CARRYB[21][0] ), .ZN(n1796) );
  XNOR2_X2 U4123 ( .A(\CARRYB[12][5] ), .B(\ab[13][5] ), .ZN(n1837) );
  NOR2_X4 U4124 ( .A1(net70478), .A2(net82149), .ZN(\ab[0][22] ) );
  NAND2_X2 U4125 ( .A1(n1769), .A2(\CARRYB[14][11] ), .ZN(n1772) );
  NAND2_X4 U4126 ( .A1(net83796), .A2(net83797), .ZN(n1696) );
  XNOR2_X2 U4127 ( .A(n1572), .B(\SUMB[2][28] ), .ZN(\SUMB[3][27] ) );
  XNOR2_X2 U4128 ( .A(\ab[3][27] ), .B(\CARRYB[2][27] ), .ZN(n1572) );
  XOR2_X1 U4129 ( .A(n2099), .B(\SUMB[19][1] ), .Z(PRODUCT[20]) );
  NAND2_X4 U4130 ( .A1(n1771), .A2(n1772), .ZN(net81169) );
  NAND3_X4 U4131 ( .A1(net82408), .A2(net82407), .A3(n1882), .ZN(
        \CARRYB[21][4] ) );
  NAND2_X2 U4132 ( .A1(\ab[18][7] ), .A2(net87619), .ZN(n2118) );
  NAND2_X1 U4133 ( .A1(\ab[13][13] ), .A2(\CARRYB[12][13] ), .ZN(n1573) );
  NAND2_X4 U4134 ( .A1(n1577), .A2(n1578), .ZN(\SUMB[5][18] ) );
  NOR2_X1 U4135 ( .A1(net91660), .A2(net70461), .ZN(\ab[17][10] ) );
  XNOR2_X2 U4136 ( .A(n1581), .B(n1225), .ZN(\SUMB[15][4] ) );
  NAND2_X2 U4137 ( .A1(\SUMB[8][15] ), .A2(\ab[9][14] ), .ZN(n2293) );
  INV_X1 U4138 ( .A(\ab[19][5] ), .ZN(net84706) );
  NAND2_X4 U4139 ( .A1(net84710), .A2(net84711), .ZN(n1583) );
  NAND2_X4 U4140 ( .A1(net84712), .A2(n1583), .ZN(n2243) );
  INV_X4 U4141 ( .A(net80694), .ZN(net84711) );
  XNOR2_X2 U4142 ( .A(n1584), .B(n1202), .ZN(\SUMB[14][5] ) );
  XNOR2_X2 U4143 ( .A(\CARRYB[19][6] ), .B(\ab[20][6] ), .ZN(net84348) );
  XNOR2_X2 U4144 ( .A(n1585), .B(n1236), .ZN(\SUMB[16][5] ) );
  XNOR2_X2 U4145 ( .A(n1586), .B(n1275), .ZN(\SUMB[12][5] ) );
  XNOR2_X2 U4146 ( .A(\CARRYB[11][5] ), .B(\ab[12][5] ), .ZN(n1586) );
  NAND2_X2 U4147 ( .A1(\CARRYB[1][22] ), .A2(\SUMB[1][23] ), .ZN(n1932) );
  NAND2_X2 U4148 ( .A1(\ab[2][22] ), .A2(\SUMB[1][23] ), .ZN(n1931) );
  XOR2_X1 U4149 ( .A(n1812), .B(\CARRYB[18][0] ), .Z(PRODUCT[19]) );
  NAND2_X2 U4150 ( .A1(\SUMB[18][1] ), .A2(\CARRYB[18][0] ), .ZN(n1815) );
  NAND2_X2 U4151 ( .A1(\ab[2][21] ), .A2(n1692), .ZN(n2190) );
  XNOR2_X2 U4152 ( .A(n1587), .B(\SUMB[8][15] ), .ZN(\SUMB[9][14] ) );
  INV_X1 U4153 ( .A(\ab[6][10] ), .ZN(n1589) );
  NAND2_X2 U4154 ( .A1(\ab[0][13] ), .A2(n237), .ZN(n2336) );
  NAND2_X4 U4155 ( .A1(n1594), .A2(n1595), .ZN(\SUMB[7][16] ) );
  NAND3_X4 U4156 ( .A1(n2218), .A2(n2217), .A3(n2216), .ZN(\CARRYB[9][20] ) );
  NAND2_X2 U4157 ( .A1(\CARRYB[8][20] ), .A2(n1278), .ZN(n2218) );
  NAND2_X2 U4158 ( .A1(n1301), .A2(n145), .ZN(n1597) );
  NAND2_X4 U4159 ( .A1(n340), .A2(n1596), .ZN(n1598) );
  NAND2_X4 U4160 ( .A1(n1597), .A2(n1598), .ZN(\SUMB[25][4] ) );
  INV_X4 U4161 ( .A(n1766), .ZN(n1603) );
  XNOR2_X2 U4162 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .ZN(n1606) );
  NAND2_X4 U4163 ( .A1(n1612), .A2(n1613), .ZN(n2248) );
  XNOR2_X2 U4164 ( .A(\SUMB[12][15] ), .B(net84481), .ZN(\SUMB[13][14] ) );
  INV_X8 U4165 ( .A(n2342), .ZN(\SUMB[1][20] ) );
  NAND2_X1 U4166 ( .A1(\ab[5][16] ), .A2(\CARRYB[4][16] ), .ZN(n1896) );
  XNOR2_X2 U4167 ( .A(\CARRYB[13][6] ), .B(n1607), .ZN(n1973) );
  XNOR2_X2 U4168 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .ZN(n1608) );
  XNOR2_X2 U4169 ( .A(n557), .B(n866), .ZN(\SUMB[3][21] ) );
  XNOR2_X2 U4170 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .ZN(n1609) );
  NAND2_X2 U4171 ( .A1(n1900), .A2(\CARRYB[6][16] ), .ZN(n1612) );
  NAND2_X4 U4172 ( .A1(n1611), .A2(n1610), .ZN(n1613) );
  INV_X4 U4173 ( .A(n1900), .ZN(n1610) );
  INV_X4 U4174 ( .A(\CARRYB[6][16] ), .ZN(n1611) );
  INV_X1 U4175 ( .A(\ab[7][16] ), .ZN(n1900) );
  NAND2_X2 U4176 ( .A1(n1424), .A2(\SUMB[1][21] ), .ZN(n1684) );
  NAND2_X2 U4177 ( .A1(\CARRYB[13][3] ), .A2(\SUMB[13][4] ), .ZN(n1969) );
  NAND2_X2 U4178 ( .A1(\CARRYB[18][7] ), .A2(\SUMB[18][8] ), .ZN(n2012) );
  NAND3_X4 U4179 ( .A1(n2158), .A2(net80836), .A3(net80835), .ZN(
        \CARRYB[4][16] ) );
  INV_X1 U4180 ( .A(\ab[19][7] ), .ZN(n1614) );
  NAND3_X4 U4181 ( .A1(net81066), .A2(net81065), .A3(n2118), .ZN(
        \CARRYB[18][7] ) );
  NAND2_X4 U4182 ( .A1(n1756), .A2(n1757), .ZN(\SUMB[13][8] ) );
  NOR2_X1 U4183 ( .A1(net70452), .A2(net70477), .ZN(\ab[9][9] ) );
  NAND3_X4 U4184 ( .A1(net80350), .A2(net80348), .A3(net80349), .ZN(
        \CARRYB[9][13] ) );
  XNOR2_X2 U4185 ( .A(\CARRYB[7][9] ), .B(\ab[8][9] ), .ZN(n1836) );
  XNOR2_X2 U4186 ( .A(n1207), .B(\ab[3][12] ), .ZN(n1928) );
  NAND3_X4 U4187 ( .A1(net84302), .A2(net84301), .A3(net84300), .ZN(
        \CARRYB[3][23] ) );
  NAND2_X4 U4188 ( .A1(net84305), .A2(n1622), .ZN(\SUMB[25][5] ) );
  NAND2_X1 U4189 ( .A1(\ab[15][14] ), .A2(\CARRYB[14][14] ), .ZN(n1623) );
  NAND3_X4 U4190 ( .A1(net84308), .A2(net84309), .A3(n1623), .ZN(
        \CARRYB[15][14] ) );
  NAND2_X2 U4191 ( .A1(\ab[16][14] ), .A2(\CARRYB[15][14] ), .ZN(n1952) );
  NAND3_X2 U4192 ( .A1(net80838), .A2(net80839), .A3(net80840), .ZN(
        \CARRYB[5][15] ) );
  XNOR2_X2 U4193 ( .A(\SUMB[4][24] ), .B(n1625), .ZN(\SUMB[5][23] ) );
  XNOR2_X2 U4194 ( .A(\CARRYB[4][23] ), .B(\ab[5][23] ), .ZN(n1625) );
  XNOR2_X2 U4195 ( .A(\SUMB[6][23] ), .B(n1626), .ZN(\SUMB[7][22] ) );
  NAND2_X1 U4196 ( .A1(\ab[18][12] ), .A2(\SUMB[17][13] ), .ZN(n2255) );
  XOR2_X2 U4197 ( .A(net82532), .B(\SUMB[16][2] ), .Z(\SUMB[17][1] ) );
  NAND2_X4 U4198 ( .A1(n1630), .A2(n1629), .ZN(\SUMB[13][12] ) );
  NAND2_X2 U4199 ( .A1(n1187), .A2(n1881), .ZN(n1848) );
  NAND2_X2 U4200 ( .A1(\ab[6][15] ), .A2(n847), .ZN(n2032) );
  INV_X1 U4201 ( .A(\ab[14][4] ), .ZN(n1632) );
  NAND2_X2 U4202 ( .A1(n1275), .A2(\CARRYB[11][5] ), .ZN(n1638) );
  NAND3_X4 U4203 ( .A1(n1638), .A2(n1637), .A3(n1636), .ZN(\CARRYB[12][5] ) );
  NAND2_X2 U4204 ( .A1(\SUMB[2][11] ), .A2(\ab[3][10] ), .ZN(n1646) );
  NAND2_X2 U4205 ( .A1(\SUMB[2][11] ), .A2(n1203), .ZN(n1647) );
  NAND3_X4 U4206 ( .A1(n1647), .A2(n1646), .A3(n1645), .ZN(\CARRYB[3][10] ) );
  NOR2_X4 U4207 ( .A1(net77892), .A2(net70467), .ZN(\ab[14][4] ) );
  INV_X4 U4208 ( .A(\CARRYB[25][3] ), .ZN(net83796) );
  NOR2_X2 U4209 ( .A1(net77912), .A2(net77966), .ZN(\ab[3][7] ) );
  NAND2_X4 U4210 ( .A1(n1700), .A2(n1701), .ZN(n1820) );
  XNOR2_X2 U4211 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .ZN(n1649) );
  NOR2_X4 U4212 ( .A1(n392), .A2(net70452), .ZN(\ab[0][9] ) );
  XOR2_X2 U4213 ( .A(n1651), .B(\SUMB[1][11] ), .Z(\SUMB[2][10] ) );
  NAND3_X2 U4214 ( .A1(n1652), .A2(n1653), .A3(n1654), .ZN(\CARRYB[2][10] ) );
  NAND2_X2 U4215 ( .A1(n1246), .A2(\SUMB[2][10] ), .ZN(n1656) );
  NAND2_X2 U4216 ( .A1(\ab[3][9] ), .A2(\SUMB[2][10] ), .ZN(n1657) );
  NAND3_X4 U4217 ( .A1(n1657), .A2(n1656), .A3(n1655), .ZN(\CARRYB[3][9] ) );
  NAND2_X2 U4218 ( .A1(\CARRYB[7][11] ), .A2(n1838), .ZN(n1661) );
  NAND2_X4 U4219 ( .A1(n1659), .A2(n1660), .ZN(n1662) );
  INV_X4 U4220 ( .A(n1838), .ZN(n1660) );
  INV_X4 U4221 ( .A(\ab[8][11] ), .ZN(n1838) );
  NAND3_X4 U4222 ( .A1(n1895), .A2(n1894), .A3(n1893), .ZN(\CARRYB[4][17] ) );
  XNOR2_X2 U4223 ( .A(n1663), .B(n568), .ZN(\SUMB[21][9] ) );
  XNOR2_X2 U4224 ( .A(\CARRYB[20][9] ), .B(\ab[21][9] ), .ZN(n1663) );
  XNOR2_X2 U4225 ( .A(\SUMB[3][19] ), .B(\ab[4][18] ), .ZN(n1693) );
  NAND2_X2 U4226 ( .A1(\ab[16][2] ), .A2(\CARRYB[15][2] ), .ZN(n1664) );
  NAND2_X2 U4227 ( .A1(\ab[16][2] ), .A2(\SUMB[15][3] ), .ZN(n1665) );
  NAND2_X2 U4228 ( .A1(\CARRYB[15][2] ), .A2(\SUMB[15][3] ), .ZN(n1666) );
  NAND3_X4 U4229 ( .A1(n1666), .A2(n1665), .A3(n1664), .ZN(\CARRYB[16][2] ) );
  NAND2_X2 U4230 ( .A1(\ab[17][2] ), .A2(\SUMB[16][3] ), .ZN(n1667) );
  NAND3_X4 U4231 ( .A1(n1668), .A2(n1669), .A3(n1667), .ZN(\CARRYB[17][2] ) );
  NAND2_X1 U4232 ( .A1(\ab[11][3] ), .A2(\CARRYB[10][3] ), .ZN(n1670) );
  NAND2_X2 U4233 ( .A1(\ab[11][3] ), .A2(\SUMB[10][4] ), .ZN(n1671) );
  NAND2_X2 U4234 ( .A1(\CARRYB[12][3] ), .A2(\SUMB[12][4] ), .ZN(n1676) );
  NAND2_X2 U4235 ( .A1(\ab[13][3] ), .A2(\SUMB[12][4] ), .ZN(n1677) );
  NOR2_X2 U4236 ( .A1(net77866), .A2(net70443), .ZN(\ab[26][1] ) );
  NOR2_X1 U4237 ( .A1(net77886), .A2(net70469), .ZN(\ab[13][3] ) );
  NAND2_X2 U4238 ( .A1(\CARRYB[6][9] ), .A2(\ab[7][9] ), .ZN(n1700) );
  NAND2_X2 U4239 ( .A1(\CARRYB[12][6] ), .A2(\SUMB[12][7] ), .ZN(n1998) );
  NAND2_X2 U4240 ( .A1(n854), .A2(\ab[13][6] ), .ZN(n1999) );
  NAND3_X2 U4241 ( .A1(n1919), .A2(n1918), .A3(n1917), .ZN(\CARRYB[12][6] ) );
  NAND3_X4 U4242 ( .A1(n2121), .A2(n2120), .A3(n2122), .ZN(\CARRYB[14][12] )
         );
  NAND2_X2 U4243 ( .A1(\CARRYB[5][18] ), .A2(\SUMB[5][19] ), .ZN(n1680) );
  NAND2_X2 U4244 ( .A1(\ab[6][18] ), .A2(\CARRYB[5][18] ), .ZN(n1682) );
  NAND3_X4 U4245 ( .A1(n1680), .A2(n1681), .A3(n1682), .ZN(\CARRYB[6][18] ) );
  NAND3_X4 U4246 ( .A1(n2140), .A2(n2141), .A3(n2139), .ZN(\CARRYB[5][18] ) );
  NAND2_X1 U4247 ( .A1(\ab[9][21] ), .A2(\CARRYB[8][21] ), .ZN(n1686) );
  NAND3_X2 U4248 ( .A1(n1686), .A2(n1687), .A3(n1688), .ZN(\CARRYB[9][21] ) );
  NAND2_X1 U4249 ( .A1(\ab[10][20] ), .A2(\CARRYB[9][20] ), .ZN(n1689) );
  NAND2_X1 U4250 ( .A1(\ab[10][20] ), .A2(\SUMB[9][21] ), .ZN(n1690) );
  NAND2_X1 U4251 ( .A1(\CARRYB[9][20] ), .A2(\SUMB[9][21] ), .ZN(n1691) );
  NAND3_X2 U4252 ( .A1(n1689), .A2(n1690), .A3(n1691), .ZN(\CARRYB[10][20] )
         );
  NOR2_X2 U4253 ( .A1(net84358), .A2(net77940), .ZN(\ab[6][23] ) );
  NAND2_X1 U4254 ( .A1(\ab[6][23] ), .A2(n1231), .ZN(n2180) );
  XNOR2_X2 U4255 ( .A(n1695), .B(n1119), .ZN(\SUMB[6][15] ) );
  INV_X1 U4256 ( .A(\ab[26][3] ), .ZN(net83797) );
  XNOR2_X2 U4257 ( .A(\SUMB[13][16] ), .B(n1697), .ZN(\SUMB[14][15] ) );
  XNOR2_X2 U4258 ( .A(\CARRYB[13][15] ), .B(\ab[14][15] ), .ZN(n1697) );
  NAND2_X1 U4259 ( .A1(\CARRYB[18][11] ), .A2(\SUMB[18][12] ), .ZN(n2258) );
  NAND3_X4 U4260 ( .A1(n2088), .A2(n2087), .A3(n2086), .ZN(\CARRYB[9][8] ) );
  NAND2_X2 U4261 ( .A1(n1222), .A2(\CARRYB[14][3] ), .ZN(n1990) );
  NAND3_X4 U4262 ( .A1(n1977), .A2(n1979), .A3(n1978), .ZN(\CARRYB[15][5] ) );
  NAND2_X1 U4263 ( .A1(\ab[27][3] ), .A2(\SUMB[26][4] ), .ZN(net80817) );
  INV_X1 U4264 ( .A(\ab[7][9] ), .ZN(n1698) );
  NAND2_X2 U4265 ( .A1(\ab[14][5] ), .A2(\SUMB[13][6] ), .ZN(n1703) );
  NAND2_X2 U4266 ( .A1(\SUMB[17][5] ), .A2(\ab[18][4] ), .ZN(n2041) );
  NAND2_X2 U4267 ( .A1(\SUMB[8][6] ), .A2(\ab[9][5] ), .ZN(n1787) );
  XNOR2_X2 U4268 ( .A(n1500), .B(\ab[16][4] ), .ZN(n1731) );
  XNOR2_X2 U4269 ( .A(\CARRYB[14][5] ), .B(\ab[15][5] ), .ZN(n1721) );
  NAND2_X2 U4270 ( .A1(\CARRYB[17][4] ), .A2(\SUMB[17][5] ), .ZN(n2042) );
  NAND2_X2 U4271 ( .A1(\ab[13][6] ), .A2(n553), .ZN(n2000) );
  NAND2_X2 U4272 ( .A1(\CARRYB[4][17] ), .A2(\SUMB[4][18] ), .ZN(n2201) );
  NOR2_X1 U4273 ( .A1(net81424), .A2(net70473), .ZN(\ab[11][15] ) );
  NAND2_X1 U4274 ( .A1(\ab[10][18] ), .A2(\SUMB[9][19] ), .ZN(n1875) );
  NAND2_X2 U4275 ( .A1(\ab[5][18] ), .A2(n1768), .ZN(n2139) );
  INV_X1 U4276 ( .A(\ab[9][15] ), .ZN(n1708) );
  NAND2_X2 U4277 ( .A1(\ab[3][17] ), .A2(\SUMB[2][18] ), .ZN(n1715) );
  XNOR2_X2 U4278 ( .A(n1717), .B(n1249), .ZN(\SUMB[11][7] ) );
  NOR2_X1 U4279 ( .A1(net77926), .A2(net84358), .ZN(\ab[8][23] ) );
  NOR2_X1 U4280 ( .A1(net84358), .A2(net77932), .ZN(\ab[7][23] ) );
  NOR2_X1 U4281 ( .A1(net84358), .A2(net77956), .ZN(\ab[4][23] ) );
  NAND2_X2 U4282 ( .A1(n1888), .A2(\CARRYB[3][19] ), .ZN(n1818) );
  INV_X2 U4283 ( .A(\ab[4][19] ), .ZN(n1888) );
  NAND2_X2 U4284 ( .A1(\CARRYB[18][4] ), .A2(\ab[19][4] ), .ZN(n1859) );
  NAND2_X2 U4285 ( .A1(\ab[4][18] ), .A2(\CARRYB[3][18] ), .ZN(n1723) );
  NAND3_X2 U4286 ( .A1(n1722), .A2(n1723), .A3(n1724), .ZN(\CARRYB[4][18] ) );
  NAND2_X4 U4287 ( .A1(n1725), .A2(n1726), .ZN(n1728) );
  INV_X2 U4288 ( .A(n1733), .ZN(n1726) );
  NAND2_X4 U4289 ( .A1(n1848), .A2(n1849), .ZN(n2095) );
  NAND2_X2 U4290 ( .A1(\ab[17][5] ), .A2(n1201), .ZN(n2037) );
  XNOR2_X2 U4291 ( .A(\SUMB[4][18] ), .B(n1729), .ZN(\SUMB[5][17] ) );
  XNOR2_X2 U4292 ( .A(\CARRYB[4][17] ), .B(\ab[5][17] ), .ZN(n1729) );
  XNOR2_X2 U4293 ( .A(\SUMB[13][13] ), .B(net83535), .ZN(\SUMB[14][12] ) );
  NAND2_X2 U4294 ( .A1(\SUMB[12][8] ), .A2(\CARRYB[12][7] ), .ZN(n2024) );
  NAND2_X2 U4295 ( .A1(\SUMB[12][6] ), .A2(\CARRYB[12][5] ), .ZN(n1922) );
  NAND2_X2 U4296 ( .A1(\ab[7][9] ), .A2(\SUMB[6][10] ), .ZN(n2002) );
  NAND2_X1 U4297 ( .A1(\ab[7][16] ), .A2(\CARRYB[6][16] ), .ZN(n2249) );
  XNOR2_X2 U4298 ( .A(n1193), .B(\ab[12][6] ), .ZN(n1764) );
  XNOR2_X2 U4299 ( .A(n288), .B(n2014), .ZN(\SUMB[7][8] ) );
  NAND2_X4 U4300 ( .A1(n1735), .A2(net82760), .ZN(\CARRYB[4][12] ) );
  INV_X4 U4301 ( .A(n1734), .ZN(n1735) );
  NAND3_X4 U4302 ( .A1(n1913), .A2(n1912), .A3(n1911), .ZN(\CARRYB[19][2] ) );
  INV_X4 U4303 ( .A(\CARRYB[3][19] ), .ZN(n1817) );
  NAND2_X4 U4304 ( .A1(\ab[6][16] ), .A2(\CARRYB[5][16] ), .ZN(n2205) );
  XNOR2_X2 U4305 ( .A(n1736), .B(\SUMB[7][16] ), .ZN(\SUMB[8][15] ) );
  XNOR2_X2 U4306 ( .A(n1737), .B(\SUMB[3][21] ), .ZN(\SUMB[4][20] ) );
  XNOR2_X2 U4307 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .ZN(n1737) );
  INV_X4 U4308 ( .A(\ab[3][20] ), .ZN(n1738) );
  INV_X4 U4309 ( .A(\CARRYB[2][20] ), .ZN(n1739) );
  NOR2_X2 U4310 ( .A1(net80727), .A2(net77964), .ZN(\ab[3][20] ) );
  INV_X2 U4311 ( .A(net83357), .ZN(net83358) );
  NAND2_X1 U4312 ( .A1(\ab[3][21] ), .A2(\CARRYB[2][21] ), .ZN(n1933) );
  XNOR2_X2 U4313 ( .A(n1741), .B(\SUMB[4][17] ), .ZN(\SUMB[5][16] ) );
  XNOR2_X2 U4314 ( .A(n1743), .B(net89255), .ZN(\SUMB[15][9] ) );
  NAND2_X2 U4315 ( .A1(\ab[9][14] ), .A2(n1235), .ZN(n2294) );
  NAND2_X1 U4316 ( .A1(\ab[5][10] ), .A2(\CARRYB[4][10] ), .ZN(n1744) );
  NAND2_X2 U4317 ( .A1(\ab[6][10] ), .A2(\CARRYB[5][10] ), .ZN(n1747) );
  NOR2_X1 U4318 ( .A1(net70459), .A2(net70460), .ZN(\ab[18][13] ) );
  NOR2_X1 U4319 ( .A1(net70460), .A2(net70461), .ZN(\ab[17][13] ) );
  NOR2_X1 U4320 ( .A1(net70460), .A2(net70467), .ZN(\ab[14][13] ) );
  NOR2_X1 U4321 ( .A1(net70460), .A2(net70469), .ZN(\ab[13][13] ) );
  NAND2_X2 U4322 ( .A1(n2043), .A2(\CARRYB[6][15] ), .ZN(n1751) );
  NAND2_X4 U4323 ( .A1(n1750), .A2(n1749), .ZN(n1752) );
  NAND2_X4 U4324 ( .A1(n1751), .A2(n1752), .ZN(n2204) );
  INV_X8 U4325 ( .A(\CARRYB[6][15] ), .ZN(n1750) );
  INV_X1 U4326 ( .A(\ab[7][15] ), .ZN(n2043) );
  NAND3_X2 U4327 ( .A1(n2003), .A2(n2002), .A3(n1700), .ZN(\CARRYB[7][9] ) );
  XNOR2_X2 U4328 ( .A(\SUMB[11][14] ), .B(n1753), .ZN(\SUMB[12][13] ) );
  XNOR2_X2 U4329 ( .A(\CARRYB[2][14] ), .B(\ab[3][14] ), .ZN(n1792) );
  XNOR2_X2 U4330 ( .A(n1754), .B(net89289), .ZN(\SUMB[20][8] ) );
  XNOR2_X2 U4331 ( .A(\CARRYB[19][8] ), .B(\ab[20][8] ), .ZN(n1754) );
  INV_X4 U4332 ( .A(net82834), .ZN(net83172) );
  NAND2_X4 U4333 ( .A1(n1853), .A2(n1852), .ZN(n2065) );
  NAND3_X4 U4334 ( .A1(n2006), .A2(n2004), .A3(n2005), .ZN(\CARRYB[8][8] ) );
  NAND2_X2 U4335 ( .A1(\CARRYB[11][7] ), .A2(\SUMB[11][8] ), .ZN(n2021) );
  XNOR2_X2 U4336 ( .A(n2171), .B(net122087), .ZN(\SUMB[21][2] ) );
  NAND3_X2 U4337 ( .A1(n2283), .A2(n2284), .A3(n2285), .ZN(\CARRYB[23][6] ) );
  NAND2_X2 U4339 ( .A1(n621), .A2(n1830), .ZN(n1762) );
  NAND2_X4 U4340 ( .A1(n1761), .A2(n1760), .ZN(n1763) );
  INV_X4 U4341 ( .A(\ab[8][8] ), .ZN(n1830) );
  NAND2_X4 U4342 ( .A1(n1850), .A2(n1851), .ZN(n1853) );
  XNOR2_X2 U4343 ( .A(\CARRYB[6][17] ), .B(\ab[7][17] ), .ZN(n1766) );
  NAND3_X2 U4344 ( .A1(net80879), .A2(net80880), .A3(n2154), .ZN(
        \CARRYB[18][9] ) );
  NAND3_X4 U4345 ( .A1(net80561), .A2(net80562), .A3(net80563), .ZN(
        \CARRYB[15][8] ) );
  NAND2_X4 U4346 ( .A1(n1770), .A2(\ab[15][11] ), .ZN(n1771) );
  INV_X1 U4347 ( .A(\ab[15][11] ), .ZN(n1769) );
  NOR2_X2 U4348 ( .A1(net70460), .A2(net70473), .ZN(\ab[11][13] ) );
  NAND2_X2 U4349 ( .A1(\SUMB[18][5] ), .A2(\CARRYB[18][4] ), .ZN(n2236) );
  XNOR2_X2 U4350 ( .A(\CARRYB[15][6] ), .B(\ab[16][6] ), .ZN(n1856) );
  NAND3_X2 U4351 ( .A1(n1776), .A2(n1775), .A3(n1774), .ZN(\CARRYB[10][8] ) );
  NAND2_X2 U4352 ( .A1(n173), .A2(\SUMB[10][8] ), .ZN(n1779) );
  NAND2_X4 U4353 ( .A1(n1121), .A2(n2149), .ZN(\SUMB[24][5] ) );
  NOR2_X1 U4354 ( .A1(net70477), .A2(net70478), .ZN(\ab[9][22] ) );
  NOR2_X1 U4355 ( .A1(net70478), .A2(net77926), .ZN(\ab[8][22] ) );
  NOR2_X1 U4356 ( .A1(net70478), .A2(net77932), .ZN(\ab[7][22] ) );
  NOR2_X1 U4357 ( .A1(net70478), .A2(net77940), .ZN(\ab[6][22] ) );
  NOR2_X2 U4358 ( .A1(net80643), .A2(net77964), .ZN(\ab[3][21] ) );
  NAND2_X2 U4359 ( .A1(n1891), .A2(n1890), .ZN(n1892) );
  INV_X4 U4360 ( .A(n1835), .ZN(n1782) );
  NAND3_X2 U4361 ( .A1(n1786), .A2(n1785), .A3(n1787), .ZN(\CARRYB[9][5] ) );
  INV_X1 U4362 ( .A(\ab[11][5] ), .ZN(n1835) );
  NOR2_X1 U4363 ( .A1(net77898), .A2(net70477), .ZN(\ab[9][5] ) );
  NAND2_X2 U4364 ( .A1(n2373), .A2(n868), .ZN(n1913) );
  INV_X4 U4365 ( .A(\CARRYB[5][16] ), .ZN(n1891) );
  NAND2_X2 U4366 ( .A1(\ab[12][13] ), .A2(\SUMB[11][14] ), .ZN(n1794) );
  NAND2_X2 U4367 ( .A1(\ab[23][0] ), .A2(\CARRYB[22][0] ), .ZN(n1800) );
  NAND2_X2 U4368 ( .A1(n36), .A2(\SUMB[22][1] ), .ZN(n1801) );
  NAND3_X2 U4369 ( .A1(net82848), .A2(net82849), .A3(net82850), .ZN(
        \CARRYB[9][3] ) );
  NAND3_X2 U4370 ( .A1(n1802), .A2(n1803), .A3(n1804), .ZN(\CARRYB[10][3] ) );
  NAND3_X4 U4371 ( .A1(n1805), .A2(n1807), .A3(n1806), .ZN(\CARRYB[21][0] ) );
  NAND3_X2 U4372 ( .A1(n1809), .A2(n1810), .A3(n1811), .ZN(\CARRYB[18][0] ) );
  NAND2_X2 U4374 ( .A1(\ab[19][0] ), .A2(\SUMB[18][1] ), .ZN(n1813) );
  NAND2_X2 U4375 ( .A1(\ab[19][0] ), .A2(\CARRYB[18][0] ), .ZN(n1814) );
  NOR2_X1 U4376 ( .A1(net77858), .A2(net70453), .ZN(\ab[21][0] ) );
  NAND2_X1 U4377 ( .A1(\ab[15][11] ), .A2(net125062), .ZN(n2093) );
  INV_X8 U4378 ( .A(n1888), .ZN(n1816) );
  XNOR2_X2 U4379 ( .A(n1820), .B(n1264), .ZN(\SUMB[7][9] ) );
  NAND3_X4 U4380 ( .A1(n2189), .A2(n2190), .A3(n2191), .ZN(\CARRYB[2][21] ) );
  XNOR2_X2 U4381 ( .A(\ab[2][21] ), .B(\CARRYB[1][21] ), .ZN(n1828) );
  NAND2_X2 U4382 ( .A1(\ab[11][5] ), .A2(\SUMB[10][6] ), .ZN(n2062) );
  NOR2_X1 U4383 ( .A1(net77892), .A2(net70473), .ZN(\ab[11][4] ) );
  XNOR2_X2 U4384 ( .A(n1836), .B(n1325), .ZN(\SUMB[8][9] ) );
  XNOR2_X2 U4385 ( .A(n11), .B(n1270), .ZN(\SUMB[17][5] ) );
  NAND2_X1 U4386 ( .A1(\ab[10][15] ), .A2(\CARRYB[9][15] ), .ZN(n1839) );
  NAND2_X1 U4387 ( .A1(\ab[11][14] ), .A2(\CARRYB[10][14] ), .ZN(n1842) );
  XNOR2_X2 U4388 ( .A(net82601), .B(net121926), .ZN(\SUMB[9][4] ) );
  INV_X4 U4389 ( .A(n1881), .ZN(n1846) );
  INV_X1 U4390 ( .A(\ab[15][12] ), .ZN(n1851) );
  INV_X1 U4391 ( .A(\ab[16][11] ), .ZN(n1881) );
  NOR2_X4 U4392 ( .A1(net83784), .A2(net70465), .ZN(\ab[15][12] ) );
  NAND2_X4 U4393 ( .A1(net82551), .A2(net82550), .ZN(n1855) );
  INV_X2 U4394 ( .A(\ab[25][4] ), .ZN(net82550) );
  NAND3_X2 U4395 ( .A1(n2025), .A2(net81530), .A3(net81531), .ZN(
        \CARRYB[25][0] ) );
  NAND2_X1 U4396 ( .A1(\ab[24][5] ), .A2(\CARRYB[23][5] ), .ZN(net79970) );
  NAND2_X4 U4397 ( .A1(n1892), .A2(n2205), .ZN(n2064) );
  NAND2_X2 U4398 ( .A1(\ab[17][1] ), .A2(\SUMB[16][2] ), .ZN(net82534) );
  NOR2_X1 U4399 ( .A1(net77868), .A2(net70451), .ZN(\ab[22][1] ) );
  NAND3_X4 U4400 ( .A1(n2161), .A2(n2162), .A3(n2163), .ZN(\CARRYB[21][1] ) );
  XNOR2_X2 U4401 ( .A(\SUMB[12][17] ), .B(n2296), .ZN(\SUMB[13][16] ) );
  NAND2_X2 U4402 ( .A1(\SUMB[7][17] ), .A2(\CARRYB[7][16] ), .ZN(n2298) );
  XNOR2_X2 U4403 ( .A(n1904), .B(\SUMB[3][22] ), .ZN(\SUMB[4][21] ) );
  INV_X1 U4404 ( .A(\ab[19][4] ), .ZN(n1857) );
  NOR2_X2 U4405 ( .A1(net77892), .A2(net70457), .ZN(\ab[19][4] ) );
  NOR2_X1 U4406 ( .A1(net91660), .A2(net70459), .ZN(\ab[18][10] ) );
  NAND2_X2 U4407 ( .A1(n1251), .A2(n2195), .ZN(n2156) );
  NOR2_X1 U4408 ( .A1(net84698), .A2(net70473), .ZN(\ab[11][14] ) );
  NAND2_X2 U4409 ( .A1(\SUMB[5][17] ), .A2(\CARRYB[5][16] ), .ZN(n2207) );
  NOR2_X1 U4410 ( .A1(net77912), .A2(net77924), .ZN(\ab[8][7] ) );
  XOR2_X2 U4411 ( .A(\CARRYB[1][5] ), .B(\ab[2][5] ), .Z(n1865) );
  XOR2_X2 U4412 ( .A(\SUMB[1][6] ), .B(n1865), .Z(\SUMB[2][5] ) );
  NAND2_X2 U4413 ( .A1(\ab[2][5] ), .A2(\SUMB[1][6] ), .ZN(n1867) );
  NAND2_X1 U4414 ( .A1(\ab[2][5] ), .A2(\CARRYB[1][5] ), .ZN(n1868) );
  NAND3_X2 U4415 ( .A1(n1866), .A2(n1867), .A3(n1868), .ZN(\CARRYB[2][5] ) );
  NOR2_X2 U4416 ( .A1(net77898), .A2(net77970), .ZN(\ab[2][5] ) );
  NOR2_X1 U4417 ( .A1(net77898), .A2(net77966), .ZN(\ab[3][5] ) );
  NAND2_X2 U4418 ( .A1(\ab[3][18] ), .A2(\SUMB[2][19] ), .ZN(n2146) );
  NAND2_X1 U4419 ( .A1(\CARRYB[13][15] ), .A2(\SUMB[13][16] ), .ZN(n1870) );
  NAND2_X1 U4420 ( .A1(\ab[14][15] ), .A2(\CARRYB[13][15] ), .ZN(n1872) );
  XOR2_X2 U4421 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .Z(n1873) );
  XOR2_X2 U4422 ( .A(n1873), .B(\SUMB[10][18] ), .Z(\SUMB[11][17] ) );
  NAND2_X1 U4423 ( .A1(\ab[10][18] ), .A2(\CARRYB[9][18] ), .ZN(n1874) );
  NAND2_X1 U4424 ( .A1(\ab[11][17] ), .A2(\CARRYB[10][17] ), .ZN(n1877) );
  NAND2_X1 U4425 ( .A1(\ab[11][17] ), .A2(\SUMB[10][18] ), .ZN(n1878) );
  NAND2_X1 U4426 ( .A1(\CARRYB[10][17] ), .A2(\SUMB[10][18] ), .ZN(n1879) );
  NAND3_X2 U4427 ( .A1(n1877), .A2(n1878), .A3(n1879), .ZN(\CARRYB[11][17] )
         );
  NOR2_X1 U4428 ( .A1(net81424), .A2(net70467), .ZN(\ab[14][15] ) );
  NOR2_X1 U4429 ( .A1(net70449), .A2(net77920), .ZN(\ab[23][8] ) );
  NAND3_X4 U4430 ( .A1(n2286), .A2(n2287), .A3(n2288), .ZN(\CARRYB[8][20] ) );
  XNOR2_X2 U4431 ( .A(n1880), .B(n1217), .ZN(\SUMB[5][8] ) );
  NAND3_X4 U4432 ( .A1(n2053), .A2(n2052), .A3(n2051), .ZN(\CARRYB[2][20] ) );
  NAND2_X2 U4433 ( .A1(\ab[6][20] ), .A2(\CARRYB[5][20] ), .ZN(net79937) );
  NAND2_X2 U4434 ( .A1(\CARRYB[2][18] ), .A2(\SUMB[2][19] ), .ZN(n2147) );
  XNOR2_X2 U4435 ( .A(n1886), .B(\CARRYB[9][19] ), .ZN(n2215) );
  XNOR2_X2 U4436 ( .A(n1887), .B(\SUMB[2][20] ), .ZN(\SUMB[3][19] ) );
  XNOR2_X2 U4437 ( .A(\CARRYB[2][19] ), .B(\ab[3][19] ), .ZN(n1887) );
  XNOR2_X2 U4438 ( .A(n1889), .B(\CARRYB[8][20] ), .ZN(n2214) );
  INV_X1 U4439 ( .A(\ab[6][16] ), .ZN(n1890) );
  NAND2_X2 U4440 ( .A1(\SUMB[3][18] ), .A2(\ab[4][17] ), .ZN(n1894) );
  NAND2_X2 U4441 ( .A1(n861), .A2(\SUMB[3][18] ), .ZN(n1895) );
  NAND2_X2 U4442 ( .A1(n1242), .A2(\CARRYB[4][16] ), .ZN(n1898) );
  NAND3_X4 U4443 ( .A1(n1898), .A2(n1897), .A3(n1896), .ZN(\CARRYB[5][16] ) );
  XNOR2_X2 U4444 ( .A(\CARRYB[12][16] ), .B(\ab[13][16] ), .ZN(n2296) );
  INV_X4 U4445 ( .A(n2341), .ZN(\CARRYB[1][20] ) );
  NAND2_X2 U4446 ( .A1(\SUMB[3][20] ), .A2(\CARRYB[3][19] ), .ZN(n2138) );
  XNOR2_X2 U4447 ( .A(n1899), .B(n1379), .ZN(\SUMB[13][6] ) );
  XNOR2_X2 U4448 ( .A(n1902), .B(n1248), .ZN(\SUMB[12][7] ) );
  NAND2_X2 U4449 ( .A1(\CARRYB[16][3] ), .A2(\ab[17][3] ), .ZN(n2106) );
  NAND2_X1 U4450 ( .A1(\ab[3][24] ), .A2(\CARRYB[2][24] ), .ZN(n2168) );
  NAND3_X2 U4451 ( .A1(n2245), .A2(n2246), .A3(n2247), .ZN(\CARRYB[6][17] ) );
  NOR2_X1 U4452 ( .A1(net84698), .A2(net70463), .ZN(\ab[16][14] ) );
  NOR2_X1 U4453 ( .A1(net84698), .A2(net70465), .ZN(\ab[15][14] ) );
  NOR2_X1 U4454 ( .A1(net84698), .A2(net70471), .ZN(\ab[12][14] ) );
  XOR2_X1 U4455 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .Z(n2099) );
  XNOR2_X2 U4456 ( .A(\CARRYB[3][21] ), .B(\ab[4][21] ), .ZN(n1904) );
  NAND3_X4 U4457 ( .A1(n1907), .A2(n1906), .A3(n1905), .ZN(\CARRYB[3][8] ) );
  NAND3_X2 U4458 ( .A1(n1914), .A2(n1916), .A3(n1915), .ZN(\CARRYB[20][2] ) );
  NOR2_X2 U4459 ( .A1(net82239), .A2(net77946), .ZN(\ab[5][25] ) );
  NOR2_X2 U4460 ( .A1(net82239), .A2(net77956), .ZN(\ab[4][25] ) );
  NOR2_X1 U4461 ( .A1(net82239), .A2(net77966), .ZN(\ab[3][25] ) );
  XNOR2_X2 U4462 ( .A(net82154), .B(net90731), .ZN(\SUMB[6][11] ) );
  NAND3_X2 U4463 ( .A1(n1946), .A2(n1945), .A3(n1944), .ZN(\CARRYB[4][8] ) );
  NAND3_X2 U4464 ( .A1(n1922), .A2(n1921), .A3(n1920), .ZN(\CARRYB[13][5] ) );
  NAND2_X2 U4465 ( .A1(\ab[9][4] ), .A2(\SUMB[8][5] ), .ZN(n1923) );
  NAND2_X2 U4467 ( .A1(\CARRYB[9][4] ), .A2(\ab[10][4] ), .ZN(n1925) );
  NAND3_X2 U4468 ( .A1(n1926), .A2(n1925), .A3(n1924), .ZN(\CARRYB[10][4] ) );
  NAND2_X2 U4469 ( .A1(net82045), .A2(net82046), .ZN(n2347) );
  NAND2_X1 U4470 ( .A1(\ab[2][22] ), .A2(\CARRYB[1][22] ), .ZN(n1930) );
  XNOR2_X2 U4471 ( .A(n176), .B(\ab[17][4] ), .ZN(n1936) );
  NAND3_X4 U4472 ( .A1(n1940), .A2(n1939), .A3(n1938), .ZN(\CARRYB[14][9] ) );
  NAND2_X2 U4473 ( .A1(\ab[7][15] ), .A2(\SUMB[6][16] ), .ZN(n2209) );
  XNOR2_X2 U4474 ( .A(n1256), .B(n1942), .ZN(\SUMB[6][13] ) );
  NOR2_X1 U4475 ( .A1(net70470), .A2(net77940), .ZN(\ab[6][18] ) );
  NOR2_X1 U4476 ( .A1(net70470), .A2(net77948), .ZN(\ab[5][18] ) );
  NOR2_X1 U4477 ( .A1(net70470), .A2(net119855), .ZN(\ab[4][18] ) );
  NAND3_X2 U4478 ( .A1(n1949), .A2(n1950), .A3(n1951), .ZN(\CARRYB[6][6] ) );
  NOR2_X1 U4479 ( .A1(net77906), .A2(net77938), .ZN(\ab[6][6] ) );
  NAND2_X2 U4480 ( .A1(\SUMB[19][9] ), .A2(\ab[20][8] ), .ZN(net81956) );
  XNOR2_X2 U4481 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .ZN(net81945) );
  NAND2_X2 U4482 ( .A1(\ab[16][14] ), .A2(n1269), .ZN(n1953) );
  NAND2_X2 U4483 ( .A1(\CARRYB[15][14] ), .A2(n1269), .ZN(n1954) );
  NAND2_X1 U4484 ( .A1(\ab[17][13] ), .A2(\CARRYB[16][13] ), .ZN(n1955) );
  NAND2_X1 U4485 ( .A1(\ab[17][13] ), .A2(\SUMB[16][14] ), .ZN(n1956) );
  NAND2_X1 U4486 ( .A1(\CARRYB[16][13] ), .A2(\SUMB[16][14] ), .ZN(n1957) );
  NAND3_X2 U4487 ( .A1(n1955), .A2(n1956), .A3(n1957), .ZN(\CARRYB[17][13] )
         );
  NAND2_X1 U4488 ( .A1(\CARRYB[4][23] ), .A2(\SUMB[4][24] ), .ZN(n1958) );
  NAND2_X1 U4489 ( .A1(\ab[5][23] ), .A2(\CARRYB[4][23] ), .ZN(n1960) );
  NOR2_X1 U4490 ( .A1(net84358), .A2(net77948), .ZN(\ab[5][23] ) );
  NAND3_X4 U4491 ( .A1(net80791), .A2(net80792), .A3(net80793), .ZN(
        \CARRYB[4][23] ) );
  NAND2_X1 U4492 ( .A1(\CARRYB[5][23] ), .A2(n1231), .ZN(n2181) );
  NAND2_X2 U4493 ( .A1(\ab[6][23] ), .A2(\CARRYB[5][23] ), .ZN(n2179) );
  NAND3_X2 U4494 ( .A1(n1962), .A2(n1961), .A3(n1963), .ZN(\CARRYB[4][9] ) );
  NAND2_X2 U4495 ( .A1(\ab[15][2] ), .A2(\SUMB[14][3] ), .ZN(n1971) );
  NAND2_X2 U4496 ( .A1(\CARRYB[14][2] ), .A2(\SUMB[14][3] ), .ZN(n1972) );
  NOR2_X2 U4497 ( .A1(net91660), .A2(net70469), .ZN(\ab[13][10] ) );
  NAND2_X1 U4498 ( .A1(\ab[20][10] ), .A2(\SUMB[19][11] ), .ZN(n2130) );
  NAND2_X1 U4499 ( .A1(\ab[2][25] ), .A2(n349), .ZN(n2165) );
  NAND2_X1 U4500 ( .A1(\ab[2][25] ), .A2(\SUMB[1][26] ), .ZN(n2166) );
  NAND3_X4 U4501 ( .A1(net80845), .A2(net80844), .A3(n2159), .ZN(
        \CARRYB[7][13] ) );
  NAND2_X2 U4502 ( .A1(\ab[14][6] ), .A2(\SUMB[13][7] ), .ZN(n1975) );
  NAND2_X2 U4504 ( .A1(\SUMB[4][14] ), .A2(n1255), .ZN(n1982) );
  NAND3_X4 U4505 ( .A1(net81713), .A2(net81714), .A3(n1983), .ZN(
        \CARRYB[6][12] ) );
  NAND3_X2 U4506 ( .A1(n1986), .A2(n1985), .A3(n1984), .ZN(\CARRYB[2][15] ) );
  NAND2_X2 U4507 ( .A1(n17), .A2(\ab[15][3] ), .ZN(n1991) );
  NOR2_X1 U4508 ( .A1(net77886), .A2(net70465), .ZN(\ab[15][3] ) );
  NAND2_X2 U4509 ( .A1(\CARRYB[8][8] ), .A2(\SUMB[8][9] ), .ZN(n2088) );
  NAND2_X2 U4510 ( .A1(\SUMB[8][9] ), .A2(\ab[9][8] ), .ZN(n2087) );
  NAND2_X2 U4511 ( .A1(\ab[25][4] ), .A2(\SUMB[24][5] ), .ZN(n2114) );
  XNOR2_X2 U4512 ( .A(n1993), .B(n1253), .ZN(\SUMB[14][4] ) );
  NAND2_X2 U4513 ( .A1(\ab[12][2] ), .A2(\SUMB[11][3] ), .ZN(n1996) );
  NAND3_X2 U4514 ( .A1(n1995), .A2(n1996), .A3(n1997), .ZN(\CARRYB[12][2] ) );
  NOR2_X1 U4515 ( .A1(net77878), .A2(net70471), .ZN(\ab[12][2] ) );
  NOR2_X1 U4516 ( .A1(net85716), .A2(net70457), .ZN(\ab[19][11] ) );
  NOR2_X1 U4517 ( .A1(net85716), .A2(net70461), .ZN(\ab[17][11] ) );
  NOR2_X1 U4518 ( .A1(net85716), .A2(net70463), .ZN(\ab[16][11] ) );
  NOR2_X1 U4519 ( .A1(net83784), .A2(net70459), .ZN(\ab[18][12] ) );
  XNOR2_X2 U4520 ( .A(net149004), .B(net81586), .ZN(\SUMB[7][10] ) );
  NAND2_X2 U4521 ( .A1(n938), .A2(\CARRYB[7][8] ), .ZN(n2006) );
  NAND2_X2 U4522 ( .A1(net88702), .A2(\ab[19][7] ), .ZN(n2011) );
  XNOR2_X2 U4523 ( .A(n1425), .B(\ab[7][8] ), .ZN(n2014) );
  NAND3_X4 U4524 ( .A1(n2069), .A2(n2070), .A3(n2068), .ZN(\CARRYB[6][13] ) );
  NOR2_X1 U4525 ( .A1(net77892), .A2(net70443), .ZN(\ab[26][4] ) );
  NAND2_X2 U4526 ( .A1(\SUMB[2][21] ), .A2(\CARRYB[2][20] ), .ZN(n2194) );
  NAND2_X2 U4527 ( .A1(\ab[3][20] ), .A2(\SUMB[2][21] ), .ZN(n2193) );
  NAND3_X2 U4528 ( .A1(n2016), .A2(n2017), .A3(n2018), .ZN(\CARRYB[9][7] ) );
  NAND2_X2 U4529 ( .A1(\ab[12][7] ), .A2(\SUMB[11][8] ), .ZN(n2020) );
  NAND2_X2 U4530 ( .A1(\CARRYB[24][0] ), .A2(\ab[25][0] ), .ZN(n2025) );
  NOR2_X1 U4531 ( .A1(net77912), .A2(net70477), .ZN(\ab[9][7] ) );
  XNOR2_X2 U4532 ( .A(net81493), .B(net88868), .ZN(\SUMB[22][3] ) );
  XNOR2_X2 U4533 ( .A(n2031), .B(\SUMB[8][16] ), .ZN(\SUMB[9][15] ) );
  NOR2_X2 U4534 ( .A1(net86565), .A2(net119855), .ZN(\ab[4][19] ) );
  NOR2_X2 U4535 ( .A1(net86565), .A2(net77932), .ZN(\ab[7][19] ) );
  NOR2_X2 U4536 ( .A1(net86565), .A2(net70477), .ZN(\ab[9][19] ) );
  NOR2_X2 U4537 ( .A1(net86565), .A2(net70475), .ZN(\ab[10][19] ) );
  NOR2_X2 U4538 ( .A1(net86565), .A2(net70473), .ZN(\ab[11][19] ) );
  NOR2_X2 U4539 ( .A1(net70471), .A2(net86565), .ZN(\ab[12][19] ) );
  NAND2_X2 U4540 ( .A1(\ab[6][15] ), .A2(\SUMB[5][16] ), .ZN(n2033) );
  NAND2_X2 U4541 ( .A1(\SUMB[5][16] ), .A2(n847), .ZN(n2034) );
  NAND3_X4 U4542 ( .A1(n2033), .A2(n2034), .A3(n2032), .ZN(\CARRYB[6][15] ) );
  NAND2_X2 U4543 ( .A1(\ab[7][14] ), .A2(\SUMB[6][15] ), .ZN(n2035) );
  NOR2_X1 U4544 ( .A1(net70457), .A2(net83784), .ZN(\ab[19][12] ) );
  XNOR2_X2 U4545 ( .A(n851), .B(n2036), .ZN(\SUMB[8][20] ) );
  XNOR2_X2 U4546 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .ZN(n2036) );
  NAND2_X2 U4547 ( .A1(\ab[17][5] ), .A2(\SUMB[16][6] ), .ZN(n2038) );
  NAND2_X2 U4548 ( .A1(\SUMB[16][6] ), .A2(\CARRYB[16][5] ), .ZN(n2039) );
  NAND2_X2 U4549 ( .A1(\ab[24][5] ), .A2(\SUMB[23][6] ), .ZN(net79969) );
  NAND2_X1 U4550 ( .A1(\SUMB[9][20] ), .A2(\ab[10][19] ), .ZN(n2220) );
  NAND2_X1 U4551 ( .A1(\SUMB[9][20] ), .A2(\CARRYB[9][19] ), .ZN(n2221) );
  NAND2_X1 U4552 ( .A1(\ab[19][11] ), .A2(\SUMB[18][12] ), .ZN(n2257) );
  INV_X4 U4553 ( .A(\CARRYB[5][17] ), .ZN(n2044) );
  NAND2_X1 U4554 ( .A1(\ab[9][15] ), .A2(\CARRYB[8][15] ), .ZN(n2050) );
  NAND2_X1 U4555 ( .A1(\ab[11][5] ), .A2(\CARRYB[10][5] ), .ZN(n2063) );
  NOR2_X1 U4556 ( .A1(net77920), .A2(net77930), .ZN(\ab[7][8] ) );
  NOR2_X1 U4557 ( .A1(net77898), .A2(net70473), .ZN(\ab[11][5] ) );
  XNOR2_X2 U4558 ( .A(n2065), .B(\SUMB[14][13] ), .ZN(\SUMB[15][12] ) );
  XOR2_X2 U4559 ( .A(\CARRYB[14][16] ), .B(\ab[15][16] ), .Z(n2066) );
  NOR2_X1 U4560 ( .A1(net70465), .A2(net124723), .ZN(\ab[15][16] ) );
  NAND2_X1 U4561 ( .A1(\CARRYB[19][10] ), .A2(\SUMB[19][11] ), .ZN(n2131) );
  NOR2_X1 U4562 ( .A1(net70469), .A2(n182), .ZN(\ab[13][18] ) );
  NOR2_X1 U4563 ( .A1(n182), .A2(net70471), .ZN(\ab[12][18] ) );
  NOR2_X1 U4564 ( .A1(n182), .A2(net70473), .ZN(\ab[11][18] ) );
  NOR2_X1 U4565 ( .A1(n182), .A2(net70475), .ZN(\ab[10][18] ) );
  NOR2_X1 U4566 ( .A1(net70470), .A2(net77926), .ZN(\ab[8][18] ) );
  NAND2_X1 U4567 ( .A1(\CARRYB[8][11] ), .A2(\ab[9][11] ), .ZN(n2067) );
  NAND3_X4 U4568 ( .A1(net81258), .A2(net81259), .A3(n2067), .ZN(
        \CARRYB[9][11] ) );
  NAND3_X4 U4569 ( .A1(net81262), .A2(net81261), .A3(net81260), .ZN(
        \CARRYB[10][10] ) );
  NAND2_X1 U4570 ( .A1(\ab[6][13] ), .A2(\CARRYB[5][13] ), .ZN(n2068) );
  NAND2_X2 U4571 ( .A1(\SUMB[5][9] ), .A2(\ab[6][8] ), .ZN(n2078) );
  NAND3_X4 U4572 ( .A1(net81212), .A2(net81213), .A3(net81211), .ZN(
        \CARRYB[7][11] ) );
  NAND2_X2 U4573 ( .A1(\SUMB[7][10] ), .A2(\CARRYB[7][9] ), .ZN(n2085) );
  NAND3_X2 U4574 ( .A1(net81205), .A2(net81204), .A3(net81206), .ZN(
        \CARRYB[5][12] ) );
  NOR2_X1 U4575 ( .A1(net91660), .A2(net77930), .ZN(\ab[7][10] ) );
  NAND3_X4 U4576 ( .A1(n2168), .A2(n2169), .A3(n2170), .ZN(\CARRYB[3][24] ) );
  NAND2_X2 U4577 ( .A1(\ab[3][24] ), .A2(\SUMB[2][25] ), .ZN(n2169) );
  NAND2_X1 U4578 ( .A1(\ab[15][11] ), .A2(n1545), .ZN(n2092) );
  NAND2_X1 U4579 ( .A1(n1545), .A2(net125062), .ZN(n2094) );
  NAND3_X2 U4580 ( .A1(n2092), .A2(n2093), .A3(n2094), .ZN(\CARRYB[15][11] )
         );
  NAND2_X1 U4581 ( .A1(\ab[16][11] ), .A2(n1187), .ZN(n2096) );
  NAND3_X2 U4582 ( .A1(n2096), .A2(n2098), .A3(n2097), .ZN(\CARRYB[16][11] )
         );
  NAND3_X2 U4583 ( .A1(net81178), .A2(net81179), .A3(net81180), .ZN(
        \CARRYB[22][8] ) );
  NOR2_X1 U4584 ( .A1(net85716), .A2(net70473), .ZN(\ab[11][11] ) );
  NOR2_X1 U4585 ( .A1(net70486), .A2(n331), .ZN(\ab[2][26] ) );
  NAND2_X2 U4586 ( .A1(\ab[20][0] ), .A2(\SUMB[19][1] ), .ZN(n2101) );
  NAND3_X2 U4587 ( .A1(n2101), .A2(n2102), .A3(n2100), .ZN(\CARRYB[20][0] ) );
  NOR2_X1 U4588 ( .A1(net77892), .A2(net70463), .ZN(\ab[16][4] ) );
  XNOR2_X2 U4589 ( .A(n2110), .B(n1209), .ZN(\SUMB[19][3] ) );
  XNOR2_X2 U4590 ( .A(n2111), .B(\SUMB[2][19] ), .ZN(\SUMB[3][18] ) );
  XNOR2_X2 U4591 ( .A(n2112), .B(\SUMB[5][18] ), .ZN(\SUMB[6][17] ) );
  XNOR2_X2 U4592 ( .A(n2119), .B(\CARRYB[20][10] ), .ZN(\SUMB[21][10] ) );
  XNOR2_X2 U4593 ( .A(\SUMB[20][11] ), .B(\ab[21][10] ), .ZN(n2119) );
  NAND2_X2 U4594 ( .A1(\ab[14][12] ), .A2(\SUMB[13][13] ), .ZN(n2121) );
  NAND2_X2 U4595 ( .A1(\ab[13][12] ), .A2(\SUMB[12][13] ), .ZN(n2124) );
  NOR2_X1 U4596 ( .A1(net70456), .A2(net77924), .ZN(\ab[8][11] ) );
  NAND2_X1 U4597 ( .A1(\ab[20][10] ), .A2(\CARRYB[19][10] ), .ZN(n2129) );
  NAND3_X2 U4598 ( .A1(n2129), .A2(n2130), .A3(n2131), .ZN(\CARRYB[20][10] )
         );
  NAND2_X1 U4599 ( .A1(\ab[21][9] ), .A2(n370), .ZN(n2132) );
  NAND2_X1 U4600 ( .A1(\ab[21][9] ), .A2(n568), .ZN(n2133) );
  NAND2_X1 U4601 ( .A1(\SUMB[20][10] ), .A2(n370), .ZN(n2134) );
  NAND3_X2 U4602 ( .A1(n2132), .A2(n2133), .A3(n2134), .ZN(\CARRYB[21][9] ) );
  NAND2_X2 U4603 ( .A1(\ab[4][19] ), .A2(\CARRYB[3][19] ), .ZN(n2136) );
  NAND3_X4 U4604 ( .A1(n2138), .A2(n2137), .A3(n2136), .ZN(\CARRYB[4][19] ) );
  NAND3_X2 U4605 ( .A1(n2256), .A2(n2257), .A3(n2258), .ZN(\CARRYB[19][11] )
         );
  NOR2_X1 U4606 ( .A1(net70453), .A2(net91660), .ZN(\ab[21][10] ) );
  NAND2_X2 U4607 ( .A1(\CARRYB[1][19] ), .A2(\ab[2][19] ), .ZN(n2145) );
  NAND3_X4 U4608 ( .A1(n2143), .A2(n2144), .A3(n2145), .ZN(\CARRYB[2][19] ) );
  INV_X4 U4609 ( .A(n896), .ZN(n2148) );
  NOR2_X1 U4610 ( .A1(net77878), .A2(net70451), .ZN(\ab[22][2] ) );
  NOR2_X1 U4611 ( .A1(net70452), .A2(net70459), .ZN(\ab[18][9] ) );
  NAND2_X1 U4612 ( .A1(\ab[7][13] ), .A2(\CARRYB[6][13] ), .ZN(n2159) );
  NAND2_X2 U4613 ( .A1(\ab[20][1] ), .A2(\SUMB[19][2] ), .ZN(n2160) );
  NAND2_X2 U4614 ( .A1(n349), .A2(\SUMB[1][26] ), .ZN(n2167) );
  XOR2_X2 U4615 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .Z(n2172) );
  XOR2_X2 U4616 ( .A(n2172), .B(n1197), .Z(\SUMB[3][26] ) );
  NAND2_X1 U4617 ( .A1(\ab[3][26] ), .A2(\CARRYB[2][26] ), .ZN(n2173) );
  NAND2_X2 U4618 ( .A1(\ab[3][26] ), .A2(n1197), .ZN(n2174) );
  NAND2_X2 U4619 ( .A1(\CARRYB[2][26] ), .A2(n1197), .ZN(n2175) );
  NAND3_X2 U4620 ( .A1(n2173), .A2(n2174), .A3(n2175), .ZN(\CARRYB[3][26] ) );
  NAND2_X1 U4621 ( .A1(\ab[4][25] ), .A2(\CARRYB[3][25] ), .ZN(n2176) );
  NAND2_X1 U4622 ( .A1(\ab[4][25] ), .A2(\SUMB[3][26] ), .ZN(n2177) );
  NAND2_X1 U4623 ( .A1(\CARRYB[3][25] ), .A2(\SUMB[3][26] ), .ZN(n2178) );
  NAND3_X2 U4624 ( .A1(n2176), .A2(n2177), .A3(n2178), .ZN(\CARRYB[4][25] ) );
  NAND3_X2 U4625 ( .A1(n2179), .A2(n2180), .A3(n2181), .ZN(\CARRYB[6][23] ) );
  NAND2_X1 U4626 ( .A1(\ab[7][22] ), .A2(\SUMB[6][23] ), .ZN(n2182) );
  NAND2_X1 U4627 ( .A1(\CARRYB[6][22] ), .A2(\SUMB[6][23] ), .ZN(n2183) );
  NAND3_X2 U4628 ( .A1(n877), .A2(n2182), .A3(n2183), .ZN(\CARRYB[7][22] ) );
  XNOR2_X2 U4629 ( .A(n2184), .B(\SUMB[7][23] ), .ZN(\SUMB[8][22] ) );
  XNOR2_X2 U4630 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .ZN(n2184) );
  NOR2_X1 U4631 ( .A1(net123000), .A2(net70471), .ZN(\ab[12][17] ) );
  NOR2_X1 U4632 ( .A1(net123000), .A2(net70473), .ZN(\ab[11][17] ) );
  NAND3_X4 U4633 ( .A1(n2301), .A2(n2300), .A3(n2299), .ZN(\CARRYB[16][8] ) );
  NAND2_X2 U4634 ( .A1(\SUMB[20][3] ), .A2(\ab[21][2] ), .ZN(n2186) );
  NAND3_X2 U4635 ( .A1(n2185), .A2(n2186), .A3(n2187), .ZN(\CARRYB[21][2] ) );
  NOR2_X2 U4636 ( .A1(net77878), .A2(net70453), .ZN(\ab[21][2] ) );
  XNOR2_X2 U4637 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .ZN(n2188) );
  NAND2_X2 U4638 ( .A1(\SUMB[15][9] ), .A2(\CARRYB[15][8] ), .ZN(n2301) );
  NAND2_X2 U4639 ( .A1(\CARRYB[1][21] ), .A2(n1692), .ZN(n2191) );
  NAND3_X4 U4640 ( .A1(n2193), .A2(n2194), .A3(n2192), .ZN(\CARRYB[3][20] ) );
  NOR2_X1 U4641 ( .A1(net70470), .A2(net77932), .ZN(\ab[7][18] ) );
  NOR2_X1 U4642 ( .A1(net80643), .A2(net70477), .ZN(\ab[9][21] ) );
  NOR2_X1 U4643 ( .A1(net80643), .A2(net77926), .ZN(\ab[8][21] ) );
  NOR2_X1 U4644 ( .A1(net80643), .A2(net77932), .ZN(\ab[7][21] ) );
  XNOR2_X2 U4645 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .ZN(n2197) );
  NAND2_X2 U4646 ( .A1(\ab[6][16] ), .A2(\SUMB[5][17] ), .ZN(n2206) );
  NOR2_X2 U4647 ( .A1(net123000), .A2(net77948), .ZN(\ab[5][17] ) );
  NOR2_X1 U4648 ( .A1(net77908), .A2(net70455), .ZN(\ab[20][6] ) );
  XOR2_X2 U4649 ( .A(n2214), .B(n1278), .Z(\SUMB[9][20] ) );
  NAND2_X1 U4650 ( .A1(\ab[9][20] ), .A2(\CARRYB[8][20] ), .ZN(n2216) );
  NAND2_X2 U4651 ( .A1(\ab[9][20] ), .A2(n1278), .ZN(n2217) );
  NAND2_X2 U4652 ( .A1(\ab[10][19] ), .A2(\CARRYB[9][19] ), .ZN(n2219) );
  NAND2_X2 U4653 ( .A1(\ab[13][17] ), .A2(\CARRYB[12][17] ), .ZN(n2222) );
  NAND3_X2 U4654 ( .A1(n2222), .A2(n2223), .A3(n2224), .ZN(\CARRYB[13][17] )
         );
  NAND2_X1 U4655 ( .A1(\ab[14][16] ), .A2(\CARRYB[13][16] ), .ZN(n2225) );
  NAND2_X1 U4656 ( .A1(\ab[14][16] ), .A2(n1250), .ZN(n2226) );
  NAND3_X2 U4657 ( .A1(n2225), .A2(n2226), .A3(n2227), .ZN(\CARRYB[14][16] )
         );
  NAND3_X2 U4658 ( .A1(net80518), .A2(net80519), .A3(net80520), .ZN(
        \CARRYB[10][17] ) );
  NAND3_X2 U4659 ( .A1(net80521), .A2(net80522), .A3(net80523), .ZN(
        \CARRYB[11][16] ) );
  NAND2_X1 U4660 ( .A1(\ab[4][20] ), .A2(\CARRYB[3][20] ), .ZN(n2237) );
  NAND2_X1 U4661 ( .A1(\ab[5][19] ), .A2(\CARRYB[4][19] ), .ZN(n2240) );
  NAND3_X4 U4662 ( .A1(n2251), .A2(n2250), .A3(n2249), .ZN(\CARRYB[7][16] ) );
  NAND2_X2 U4663 ( .A1(\ab[8][15] ), .A2(\SUMB[7][16] ), .ZN(n2253) );
  NAND3_X2 U4664 ( .A1(net80449), .A2(n2255), .A3(net80451), .ZN(
        \CARRYB[18][12] ) );
  NAND2_X1 U4665 ( .A1(\ab[19][11] ), .A2(\CARRYB[18][11] ), .ZN(n2256) );
  XOR2_X2 U4666 ( .A(\ab[2][28] ), .B(n347), .Z(n2259) );
  XOR2_X2 U4667 ( .A(n2259), .B(\SUMB[1][29] ), .Z(\SUMB[2][28] ) );
  NAND2_X2 U4668 ( .A1(\ab[2][28] ), .A2(n347), .ZN(n2260) );
  NAND2_X2 U4669 ( .A1(\ab[2][28] ), .A2(\SUMB[1][29] ), .ZN(n2261) );
  NAND2_X2 U4670 ( .A1(n347), .A2(\SUMB[1][29] ), .ZN(n2262) );
  NAND2_X1 U4671 ( .A1(\ab[3][27] ), .A2(\CARRYB[2][27] ), .ZN(n2263) );
  NAND2_X1 U4672 ( .A1(\ab[3][27] ), .A2(\SUMB[2][28] ), .ZN(n2264) );
  NAND2_X1 U4673 ( .A1(\CARRYB[2][27] ), .A2(\SUMB[2][28] ), .ZN(n2265) );
  NAND3_X2 U4674 ( .A1(n2263), .A2(n2264), .A3(n2265), .ZN(\CARRYB[3][27] ) );
  NAND2_X1 U4675 ( .A1(\ab[7][23] ), .A2(\CARRYB[6][23] ), .ZN(n2266) );
  NAND2_X1 U4676 ( .A1(\ab[8][22] ), .A2(\CARRYB[7][22] ), .ZN(n2269) );
  NAND2_X1 U4677 ( .A1(\ab[8][22] ), .A2(\SUMB[7][23] ), .ZN(n2270) );
  NAND2_X1 U4678 ( .A1(\CARRYB[7][22] ), .A2(\SUMB[7][23] ), .ZN(n2271) );
  NAND3_X2 U4679 ( .A1(n2269), .A2(n2270), .A3(n2271), .ZN(\CARRYB[8][22] ) );
  NOR2_X1 U4680 ( .A1(n242), .A2(n2353), .ZN(\ab[1][30] ) );
  INV_X8 U4681 ( .A(B[28]), .ZN(n2354) );
  NAND3_X2 U4682 ( .A1(n2272), .A2(net80356), .A3(net80355), .ZN(
        \CARRYB[8][14] ) );
  NAND2_X2 U4683 ( .A1(\SUMB[18][4] ), .A2(\ab[19][3] ), .ZN(n2274) );
  NAND3_X2 U4684 ( .A1(n2273), .A2(n2274), .A3(n2275), .ZN(\CARRYB[19][3] ) );
  NOR2_X1 U4685 ( .A1(net77886), .A2(net70457), .ZN(\ab[19][3] ) );
  NOR2_X1 U4686 ( .A1(n2355), .A2(net77966), .ZN(\ab[3][27] ) );
  NOR2_X2 U4687 ( .A1(net77966), .A2(n2354), .ZN(\ab[3][28] ) );
  INV_X8 U4688 ( .A(B[29]), .ZN(net70492) );
  NAND2_X1 U4689 ( .A1(\ab[4][21] ), .A2(\CARRYB[3][21] ), .ZN(n2278) );
  NAND2_X1 U4690 ( .A1(\ab[6][19] ), .A2(n56), .ZN(n2279) );
  NOR2_X1 U4691 ( .A1(n955), .A2(net77956), .ZN(\ab[4][21] ) );
  NAND2_X1 U4692 ( .A1(\ab[23][6] ), .A2(n351), .ZN(n2283) );
  NAND3_X2 U4693 ( .A1(net80273), .A2(net80274), .A3(net80275), .ZN(
        \CARRYB[16][13] ) );
  NAND2_X1 U4694 ( .A1(\ab[8][20] ), .A2(\CARRYB[7][20] ), .ZN(n2286) );
  NAND2_X2 U4695 ( .A1(n851), .A2(\ab[8][20] ), .ZN(n2287) );
  NAND2_X2 U4696 ( .A1(n851), .A2(\CARRYB[7][20] ), .ZN(n2288) );
  NAND2_X1 U4697 ( .A1(\ab[9][19] ), .A2(\CARRYB[8][19] ), .ZN(n2289) );
  NAND2_X2 U4698 ( .A1(\CARRYB[8][19] ), .A2(\SUMB[8][20] ), .ZN(n2291) );
  NOR2_X1 U4699 ( .A1(net84698), .A2(net70477), .ZN(\ab[9][14] ) );
  XNOR2_X2 U4700 ( .A(\ab[1][27] ), .B(\ab[0][28] ), .ZN(n2350) );
  NOR2_X1 U4701 ( .A1(n175), .A2(net70492), .ZN(\ab[2][29] ) );
  NAND2_X1 U4702 ( .A1(\ab[9][16] ), .A2(\CARRYB[8][16] ), .ZN(n2306) );
  NAND3_X2 U4703 ( .A1(net79951), .A2(net79952), .A3(net79953), .ZN(
        \CARRYB[9][18] ) );
  NAND3_X2 U4704 ( .A1(net79955), .A2(net79956), .A3(net79957), .ZN(
        \CARRYB[8][19] ) );
  NAND3_X2 U4705 ( .A1(net79959), .A2(net79960), .A3(net79961), .ZN(
        \CARRYB[7][20] ) );
  NOR2_X1 U4706 ( .A1(net80727), .A2(net77932), .ZN(\ab[7][20] ) );
  NOR2_X1 U4707 ( .A1(net80727), .A2(net77940), .ZN(\ab[6][20] ) );
  NAND2_X1 U4708 ( .A1(\ab[12][16] ), .A2(\CARRYB[11][16] ), .ZN(n2307) );
  NAND2_X1 U4709 ( .A1(\ab[3][25] ), .A2(\CARRYB[2][25] ), .ZN(n2310) );
  NAND2_X2 U4710 ( .A1(n1219), .A2(\ab[3][25] ), .ZN(n2311) );
  NAND2_X2 U4711 ( .A1(n1219), .A2(\CARRYB[2][25] ), .ZN(n2312) );
  NAND3_X2 U4712 ( .A1(n2310), .A2(n2311), .A3(n2312), .ZN(\CARRYB[3][25] ) );
  NAND2_X1 U4713 ( .A1(\ab[4][24] ), .A2(\CARRYB[3][24] ), .ZN(n2313) );
  NAND2_X1 U4714 ( .A1(\ab[4][24] ), .A2(\SUMB[3][25] ), .ZN(n2314) );
  NAND2_X1 U4715 ( .A1(\CARRYB[3][24] ), .A2(\SUMB[3][25] ), .ZN(n2315) );
  NAND3_X2 U4716 ( .A1(n2313), .A2(n2314), .A3(n2315), .ZN(\CARRYB[4][24] ) );
  NAND2_X1 U4717 ( .A1(\CARRYB[12][16] ), .A2(\SUMB[12][17] ), .ZN(n2316) );
  NAND2_X1 U4718 ( .A1(\ab[13][16] ), .A2(\CARRYB[12][16] ), .ZN(n2318) );
  NAND3_X2 U4719 ( .A1(n2316), .A2(n2317), .A3(n2318), .ZN(\CARRYB[13][16] )
         );
  NOR2_X1 U4720 ( .A1(net124723), .A2(net70469), .ZN(\ab[13][16] ) );
  XOR2_X2 U4721 ( .A(\CARRYB[10][20] ), .B(\ab[11][20] ), .Z(n2319) );
  XOR2_X2 U4722 ( .A(\SUMB[10][21] ), .B(n2319), .Z(\SUMB[11][20] ) );
  XOR2_X2 U4723 ( .A(\CARRYB[3][27] ), .B(\ab[4][27] ), .Z(n2320) );
  XOR2_X2 U4724 ( .A(\SUMB[3][28] ), .B(n2320), .Z(\SUMB[4][27] ) );
  XOR2_X2 U4725 ( .A(\CARRYB[9][21] ), .B(\ab[10][21] ), .Z(n2321) );
  NOR2_X1 U4726 ( .A1(net70473), .A2(net80727), .ZN(\ab[11][20] ) );
  NOR2_X1 U4727 ( .A1(net70463), .A2(net81424), .ZN(\ab[16][15] ) );
  NOR2_X1 U4728 ( .A1(net77956), .A2(n2355), .ZN(\ab[4][27] ) );
  NOR2_X1 U4729 ( .A1(net70475), .A2(net80643), .ZN(\ab[10][21] ) );
  NAND2_X2 U4730 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .ZN(n2322) );
  INV_X4 U4731 ( .A(n2322), .ZN(\CARRYB[1][0] ) );
  NAND2_X2 U4732 ( .A1(\ab[0][3] ), .A2(\ab[1][2] ), .ZN(n2323) );
  INV_X4 U4733 ( .A(n2323), .ZN(\CARRYB[1][2] ) );
  INV_X4 U4734 ( .A(n2324), .ZN(\SUMB[1][2] ) );
  NAND2_X2 U4735 ( .A1(n870), .A2(\ab[1][3] ), .ZN(n2325) );
  XNOR2_X2 U4736 ( .A(\ab[1][3] ), .B(n870), .ZN(n2326) );
  INV_X4 U4737 ( .A(n2326), .ZN(\SUMB[1][3] ) );
  INV_X4 U4738 ( .A(n2328), .ZN(\SUMB[1][4] ) );
  XNOR2_X2 U4739 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .ZN(n2330) );
  INV_X4 U4740 ( .A(n2330), .ZN(\SUMB[1][5] ) );
  INV_X4 U4741 ( .A(\*UDW_*112739/net78703 ), .ZN(\SUMB[1][6] ) );
  INV_X4 U4742 ( .A(n1517), .ZN(\CARRYB[1][9] ) );
  INV_X4 U4743 ( .A(n2331), .ZN(\SUMB[1][9] ) );
  XNOR2_X2 U4744 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .ZN(n2333) );
  INV_X4 U4745 ( .A(n2333), .ZN(\SUMB[1][10] ) );
  INV_X4 U4746 ( .A(n2336), .ZN(\CARRYB[1][12] ) );
  XNOR2_X2 U4747 ( .A(n237), .B(\ab[0][13] ), .ZN(n2337) );
  XNOR2_X2 U4748 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .ZN(n2340) );
  XNOR2_X2 U4749 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .ZN(n2342) );
  XNOR2_X2 U4750 ( .A(\ab[0][22] ), .B(\ab[1][21] ), .ZN(n2344) );
  XNOR2_X2 U4751 ( .A(n2196), .B(\ab[0][23] ), .ZN(n2346) );
  INV_X4 U4752 ( .A(n2347), .ZN(\SUMB[1][23] ) );
  NAND2_X2 U4753 ( .A1(\ab[0][27] ), .A2(\ab[1][26] ), .ZN(n2348) );
  INV_X4 U4754 ( .A(n2348), .ZN(\CARRYB[1][26] ) );
  XNOR2_X2 U4755 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .ZN(n2349) );
  INV_X4 U4756 ( .A(n2349), .ZN(\SUMB[1][26] ) );
  INV_X4 U4757 ( .A(n2350), .ZN(\SUMB[1][27] ) );
  XNOR2_X2 U4758 ( .A(\ab[1][28] ), .B(\ab[0][29] ), .ZN(n2351) );
  INV_X4 U4759 ( .A(n2351), .ZN(\SUMB[1][28] ) );
  XNOR2_X2 U4760 ( .A(\ab[1][29] ), .B(\ab[0][30] ), .ZN(n2352) );
  INV_X4 U4761 ( .A(n2352), .ZN(\SUMB[1][29] ) );
  AND2_X2 U4762 ( .A1(B[31]), .A2(net80392), .ZN(\ab[0][31] ) );
  NOR2_X4 U4763 ( .A1(net70476), .A2(net82149), .ZN(\ab[0][21] ) );
  NOR2_X4 U4764 ( .A1(net81673), .A2(net77898), .ZN(\ab[0][5] ) );
  NOR2_X4 U4765 ( .A1(net77892), .A2(net83263), .ZN(\ab[1][4] ) );
  NOR2_X4 U4766 ( .A1(net77882), .A2(net83263), .ZN(\ab[1][3] ) );
  NOR2_X4 U4767 ( .A1(net81673), .A2(net77878), .ZN(\ab[0][2] ) );
  NOR2_X4 U4768 ( .A1(net77920), .A2(net77970), .ZN(\ab[2][8] ) );
  NOR2_X4 U4769 ( .A1(net82890), .A2(net77964), .ZN(\ab[3][17] ) );
  NOR2_X4 U4770 ( .A1(net77920), .A2(net77966), .ZN(\ab[3][8] ) );
  NOR2_X4 U4771 ( .A1(net77906), .A2(net77966), .ZN(\ab[3][6] ) );
  NOR2_X4 U4772 ( .A1(net77920), .A2(net119855), .ZN(\ab[4][8] ) );
  NOR2_X4 U4773 ( .A1(net77906), .A2(net119855), .ZN(\ab[4][6] ) );
  NOR2_X4 U4774 ( .A1(net77886), .A2(net77956), .ZN(\ab[4][3] ) );
  NOR2_X4 U4775 ( .A1(net77878), .A2(net119855), .ZN(\ab[4][2] ) );
  NOR2_X4 U4776 ( .A1(net77920), .A2(net77946), .ZN(\ab[5][8] ) );
  NOR2_X4 U4777 ( .A1(net77866), .A2(net77946), .ZN(\ab[5][1] ) );
  NOR2_X4 U4778 ( .A1(net81424), .A2(net77940), .ZN(\ab[6][15] ) );
  NOR2_X4 U4779 ( .A1(net77912), .A2(net77938), .ZN(\ab[6][7] ) );
  NOR2_X4 U4780 ( .A1(net77892), .A2(net77938), .ZN(\ab[6][4] ) );
  NOR2_X4 U4781 ( .A1(net77878), .A2(net77938), .ZN(\ab[6][2] ) );
  NOR2_X4 U4782 ( .A1(net77860), .A2(net77938), .ZN(\ab[6][0] ) );
  NOR2_X4 U4783 ( .A1(net123000), .A2(net77932), .ZN(\ab[7][17] ) );
  NOR2_X4 U4784 ( .A1(net70452), .A2(net77930), .ZN(\ab[7][9] ) );
  NOR2_X4 U4785 ( .A1(net77912), .A2(net77930), .ZN(\ab[7][7] ) );
  NOR2_X4 U4786 ( .A1(net77906), .A2(net77930), .ZN(\ab[7][6] ) );
  NOR2_X4 U4787 ( .A1(net77886), .A2(net77930), .ZN(\ab[7][3] ) );
  NOR2_X4 U4788 ( .A1(net80727), .A2(net77926), .ZN(\ab[8][20] ) );
  NOR2_X4 U4789 ( .A1(net70460), .A2(net77926), .ZN(\ab[8][13] ) );
  NOR2_X4 U4790 ( .A1(net77920), .A2(net77924), .ZN(\ab[8][8] ) );
  NOR2_X4 U4791 ( .A1(net80727), .A2(net70477), .ZN(\ab[9][20] ) );
  NOR2_X4 U4792 ( .A1(net77920), .A2(net70477), .ZN(\ab[9][8] ) );
  NOR2_X4 U4793 ( .A1(net77892), .A2(net70477), .ZN(\ab[9][4] ) );
  NOR2_X4 U4794 ( .A1(net77886), .A2(net70477), .ZN(\ab[9][3] ) );
  NOR2_X4 U4795 ( .A1(net77878), .A2(net70477), .ZN(\ab[9][2] ) );
  NOR2_X4 U4796 ( .A1(net80727), .A2(net70475), .ZN(\ab[10][20] ) );
  NOR2_X4 U4797 ( .A1(net81424), .A2(net70475), .ZN(\ab[10][15] ) );
  NOR2_X4 U4798 ( .A1(net77892), .A2(net70475), .ZN(\ab[10][4] ) );
  NOR2_X4 U4799 ( .A1(net77886), .A2(net70475), .ZN(\ab[10][3] ) );
  NOR2_X4 U4800 ( .A1(net77866), .A2(net70475), .ZN(\ab[10][1] ) );
  NOR2_X4 U4801 ( .A1(net77886), .A2(net70473), .ZN(\ab[11][3] ) );
  NOR2_X4 U4802 ( .A1(net77860), .A2(net70473), .ZN(\ab[11][0] ) );
  NOR2_X4 U4803 ( .A1(net77908), .A2(net70471), .ZN(\ab[12][6] ) );
  NOR2_X4 U4804 ( .A1(net77900), .A2(net70471), .ZN(\ab[12][5] ) );
  NOR2_X4 U4805 ( .A1(net77886), .A2(net70471), .ZN(\ab[12][3] ) );
  NOR2_X4 U4806 ( .A1(net77860), .A2(net70471), .ZN(\ab[12][0] ) );
  NOR2_X4 U4807 ( .A1(net77900), .A2(net70469), .ZN(\ab[13][5] ) );
  NOR2_X4 U4808 ( .A1(net77900), .A2(net70467), .ZN(\ab[14][5] ) );
  NOR2_X4 U4809 ( .A1(net77886), .A2(net70467), .ZN(\ab[14][3] ) );
  NOR2_X4 U4810 ( .A1(net77868), .A2(net70467), .ZN(\ab[14][1] ) );
  NOR2_X4 U4811 ( .A1(net77920), .A2(net70465), .ZN(\ab[15][8] ) );
  NOR2_X4 U4812 ( .A1(net77914), .A2(net70465), .ZN(\ab[15][7] ) );
  NOR2_X4 U4813 ( .A1(net77900), .A2(net70465), .ZN(\ab[15][5] ) );
  NOR2_X4 U4814 ( .A1(net77892), .A2(net70465), .ZN(\ab[15][4] ) );
  NOR2_X4 U4815 ( .A1(net77878), .A2(net70465), .ZN(\ab[15][2] ) );
  NOR2_X4 U4816 ( .A1(net77920), .A2(net70463), .ZN(\ab[16][8] ) );
  NOR2_X4 U4817 ( .A1(net77908), .A2(net70463), .ZN(\ab[16][6] ) );
  NOR2_X4 U4818 ( .A1(net77900), .A2(net70463), .ZN(\ab[16][5] ) );
  NOR2_X4 U4819 ( .A1(net77886), .A2(net70463), .ZN(\ab[16][3] ) );
  NOR2_X4 U4820 ( .A1(net77878), .A2(net70463), .ZN(\ab[16][2] ) );
  NOR2_X4 U4821 ( .A1(net77860), .A2(net70463), .ZN(\ab[16][0] ) );
  NOR2_X4 U4822 ( .A1(net77920), .A2(net70461), .ZN(\ab[17][8] ) );
  NOR2_X4 U4823 ( .A1(net77900), .A2(net70461), .ZN(\ab[17][5] ) );
  NOR2_X4 U4824 ( .A1(net77892), .A2(net70461), .ZN(\ab[17][4] ) );
  NOR2_X4 U4825 ( .A1(net77886), .A2(net70461), .ZN(\ab[17][3] ) );
  NOR2_X4 U4826 ( .A1(net77878), .A2(net70461), .ZN(\ab[17][2] ) );
  NOR2_X4 U4827 ( .A1(net77868), .A2(net70461), .ZN(\ab[17][1] ) );
  NOR2_X4 U4828 ( .A1(net77860), .A2(net70461), .ZN(\ab[17][0] ) );
  NOR2_X4 U4829 ( .A1(net77900), .A2(net70459), .ZN(\ab[18][5] ) );
  NOR2_X4 U4830 ( .A1(net77892), .A2(net70459), .ZN(\ab[18][4] ) );
  NOR2_X4 U4831 ( .A1(net77878), .A2(net70459), .ZN(\ab[18][2] ) );
  NOR2_X4 U4832 ( .A1(net77868), .A2(net70459), .ZN(\ab[18][1] ) );
  NOR2_X4 U4833 ( .A1(net77860), .A2(net70459), .ZN(\ab[18][0] ) );
  NOR2_X4 U4834 ( .A1(net77914), .A2(net70457), .ZN(\ab[19][7] ) );
  NOR2_X4 U4835 ( .A1(net77900), .A2(net70457), .ZN(\ab[19][5] ) );
  NOR2_X4 U4836 ( .A1(net77878), .A2(net70457), .ZN(\ab[19][2] ) );
  NOR2_X4 U4837 ( .A1(net77858), .A2(net70457), .ZN(\ab[19][0] ) );
  NOR2_X4 U4838 ( .A1(net77920), .A2(net70455), .ZN(\ab[20][8] ) );
  NOR2_X4 U4839 ( .A1(net77914), .A2(net70455), .ZN(\ab[20][7] ) );
  NOR2_X4 U4840 ( .A1(net77892), .A2(net70455), .ZN(\ab[20][4] ) );
  NOR2_X4 U4841 ( .A1(net77878), .A2(net70455), .ZN(\ab[20][2] ) );
  NOR2_X4 U4842 ( .A1(net77868), .A2(net70455), .ZN(\ab[20][1] ) );
  NOR2_X4 U4843 ( .A1(net77858), .A2(net70455), .ZN(\ab[20][0] ) );
  NOR2_X4 U4844 ( .A1(net77892), .A2(net70453), .ZN(\ab[21][4] ) );
  NOR2_X4 U4845 ( .A1(net77886), .A2(net70453), .ZN(\ab[21][3] ) );
  NOR2_X4 U4846 ( .A1(net77868), .A2(net70453), .ZN(\ab[21][1] ) );
  NOR2_X4 U4847 ( .A1(net77908), .A2(net70451), .ZN(\ab[22][6] ) );
  NOR2_X4 U4848 ( .A1(net77892), .A2(net70451), .ZN(\ab[22][4] ) );
  NOR2_X4 U4849 ( .A1(net77858), .A2(net70451), .ZN(\ab[22][0] ) );
  NOR2_X4 U4850 ( .A1(net77908), .A2(net70449), .ZN(\ab[23][6] ) );
  NOR2_X4 U4851 ( .A1(net77900), .A2(net70449), .ZN(\ab[23][5] ) );
  NOR2_X4 U4852 ( .A1(net77878), .A2(net70449), .ZN(\ab[23][2] ) );
  NOR2_X4 U4853 ( .A1(net77858), .A2(net70449), .ZN(\ab[23][0] ) );
  NOR2_X4 U4854 ( .A1(net77906), .A2(net70447), .ZN(\ab[24][6] ) );
  NOR2_X4 U4855 ( .A1(net77878), .A2(net70447), .ZN(\ab[24][2] ) );
  NOR2_X4 U4856 ( .A1(net77886), .A2(net70443), .ZN(\ab[26][3] ) );
  INV_X4 U4857 ( .A(net70435), .ZN(PRODUCT[0]) );
  NOR2_X1 U15 ( .A1(n348), .A2(net92311), .ZN(n1181) );
  NAND2_X2 U17 ( .A1(n581), .A2(n582), .ZN(n584) );
  NAND2_X2 U29 ( .A1(net119817), .A2(\CARRYB[3][14] ), .ZN(n529) );
  NAND3_X4 U30 ( .A1(net80673), .A2(net80672), .A3(net80671), .ZN(
        \CARRYB[20][7] ) );
  NAND2_X2 U35 ( .A1(net91001), .A2(net88699), .ZN(net80673) );
  INV_X2 U40 ( .A(net83054), .ZN(n2356) );
  NAND2_X2 U65 ( .A1(net123363), .A2(\ab[28][1] ), .ZN(net79880) );
  INV_X4 U67 ( .A(n476), .ZN(n12) );
  INV_X2 U105 ( .A(net89104), .ZN(n582) );
  XNOR2_X2 U140 ( .A(n2001), .B(n221), .ZN(n1261) );
  INV_X4 U148 ( .A(n939), .ZN(n221) );
  INV_X2 U160 ( .A(\SUMB[3][14] ), .ZN(n910) );
  NAND2_X4 U177 ( .A1(n214), .A2(n213), .ZN(n857) );
  NAND2_X2 U178 ( .A1(\CARRYB[3][13] ), .A2(n212), .ZN(n213) );
  INV_X8 U217 ( .A(\CARRYB[26][2] ), .ZN(net83054) );
  NAND2_X2 U236 ( .A1(\CARRYB[27][2] ), .A2(\ab[28][2] ), .ZN(n115) );
  XOR2_X2 U253 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Z(n2357) );
  NAND2_X2 U262 ( .A1(net121452), .A2(net121451), .ZN(n193) );
  INV_X2 U287 ( .A(n565), .ZN(net85399) );
  INV_X1 U290 ( .A(\CARRYB[1][16] ), .ZN(n2358) );
  INV_X2 U309 ( .A(n2358), .ZN(n2359) );
  NAND2_X2 U330 ( .A1(net85044), .A2(net88455), .ZN(n2117) );
  NAND2_X2 U350 ( .A1(net81070), .A2(n193), .ZN(n486) );
  INV_X4 U402 ( .A(\CARRYB[8][12] ), .ZN(net84868) );
  NAND2_X2 U428 ( .A1(\CARRYB[8][12] ), .A2(\ab[9][12] ), .ZN(net81373) );
  NAND2_X4 U430 ( .A1(net85461), .A2(n517), .ZN(n2360) );
  NAND2_X2 U443 ( .A1(net85461), .A2(n517), .ZN(\SUMB[8][13] ) );
  INV_X2 U444 ( .A(net92790), .ZN(net92568) );
  NAND2_X2 U446 ( .A1(n9), .A2(net92568), .ZN(n499) );
  NAND2_X4 U448 ( .A1(n817), .A2(net87363), .ZN(net82029) );
  NAND2_X4 U455 ( .A1(\CARRYB[21][3] ), .A2(\ab[22][3] ), .ZN(n502) );
  INV_X2 U465 ( .A(n280), .ZN(n2361) );
  INV_X4 U467 ( .A(\ab[2][16] ), .ZN(n280) );
  NAND2_X2 U485 ( .A1(\CARRYB[5][6] ), .A2(\ab[6][6] ), .ZN(n1951) );
  NAND2_X2 U505 ( .A1(\CARRYB[5][6] ), .A2(\SUMB[5][7] ), .ZN(n1949) );
  XNOR2_X2 U569 ( .A(\CARRYB[7][9] ), .B(\ab[8][9] ), .ZN(n2362) );
  NAND3_X2 U579 ( .A1(n892), .A2(n893), .A3(n894), .ZN(\CARRYB[17][12] ) );
  INV_X2 U617 ( .A(n544), .ZN(n547) );
  NAND2_X4 U628 ( .A1(n60), .A2(n61), .ZN(n933) );
  NAND2_X4 U633 ( .A1(n1431), .A2(n1432), .ZN(n1434) );
  NAND2_X4 U637 ( .A1(n58), .A2(n59), .ZN(n61) );
  NAND2_X4 U639 ( .A1(net79863), .A2(n1090), .ZN(net80110) );
  NAND3_X4 U658 ( .A1(net80941), .A2(net80942), .A3(net80940), .ZN(
        \CARRYB[22][6] ) );
  NAND2_X1 U672 ( .A1(\ab[3][17] ), .A2(\CARRYB[2][17] ), .ZN(n1714) );
  NAND2_X2 U682 ( .A1(\SUMB[2][13] ), .A2(\ab[3][12] ), .ZN(n2008) );
  NAND2_X2 U684 ( .A1(\SUMB[2][13] ), .A2(n1324), .ZN(n2007) );
  BUF_X2 U693 ( .A(\SUMB[6][7] ), .Z(n1208) );
  NAND2_X2 U703 ( .A1(\ab[16][1] ), .A2(\CARRYB[15][1] ), .ZN(n648) );
  NAND2_X2 U704 ( .A1(\ab[15][1] ), .A2(\CARRYB[14][1] ), .ZN(n653) );
  NAND2_X4 U716 ( .A1(n2370), .A2(n563), .ZN(n1832) );
  NAND2_X4 U804 ( .A1(n1029), .A2(n1030), .ZN(n1032) );
  INV_X16 U808 ( .A(net70491), .ZN(n26) );
  INV_X2 U828 ( .A(\SUMB[11][6] ), .ZN(n1274) );
  INV_X2 U832 ( .A(net86662), .ZN(net148235) );
  INV_X4 U837 ( .A(n1718), .ZN(n634) );
  XNOR2_X2 U884 ( .A(net86519), .B(net121380), .ZN(n2363) );
  XNOR2_X2 U886 ( .A(net86519), .B(n2365), .ZN(n2364) );
  INV_X32 U899 ( .A(net121380), .ZN(n2365) );
  NAND2_X4 U938 ( .A1(n2363), .A2(n334), .ZN(net147939) );
  NAND2_X2 U961 ( .A1(n1033), .A2(n1034), .ZN(net81070) );
  INV_X4 U995 ( .A(\CARRYB[24][2] ), .ZN(n129) );
  XOR2_X2 U997 ( .A(\CARRYB[2][13] ), .B(\ab[3][13] ), .Z(n2366) );
  NAND2_X2 U1126 ( .A1(\CARRYB[24][2] ), .A2(\ab[25][2] ), .ZN(n131) );
  NAND2_X4 U1153 ( .A1(n597), .A2(\ab[25][0] ), .ZN(net81531) );
  INV_X4 U1156 ( .A(n541), .ZN(n542) );
  NAND2_X2 U1165 ( .A1(n224), .A2(n225), .ZN(n227) );
  INV_X4 U1178 ( .A(n1274), .ZN(n1275) );
  BUF_X4 U1181 ( .A(\CARRYB[21][6] ), .Z(net89008) );
  NAND2_X2 U1214 ( .A1(n372), .A2(\ab[22][2] ), .ZN(net80926) );
  NAND2_X4 U1215 ( .A1(\SUMB[6][17] ), .A2(\ab[7][16] ), .ZN(n2250) );
  NAND2_X2 U1275 ( .A1(n1554), .A2(n1555), .ZN(n150) );
  NAND2_X4 U1527 ( .A1(n877), .A2(n878), .ZN(n1626) );
  INV_X2 U1629 ( .A(\SUMB[14][9] ), .ZN(net88934) );
  NAND2_X4 U1738 ( .A1(net84070), .A2(net81256), .ZN(net84071) );
  XNOR2_X2 U1767 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .ZN(n2367) );
  NAND2_X4 U1772 ( .A1(\SUMB[1][16] ), .A2(\ab[2][15] ), .ZN(n1985) );
  XOR2_X2 U1774 ( .A(\CARRYB[9][1] ), .B(\ab[10][1] ), .Z(n1470) );
  XNOR2_X2 U1869 ( .A(\SUMB[14][2] ), .B(n2368), .ZN(\SUMB[15][1] ) );
  XNOR2_X1 U1973 ( .A(\CARRYB[14][1] ), .B(\ab[15][1] ), .ZN(n2368) );
  XOR2_X2 U1995 ( .A(\ab[19][0] ), .B(\SUMB[18][1] ), .Z(n1812) );
  XNOR2_X2 U2002 ( .A(n396), .B(\CARRYB[17][1] ), .ZN(\SUMB[18][1] ) );
  XNOR2_X2 U2086 ( .A(n566), .B(n2369), .ZN(net85734) );
  INV_X32 U2093 ( .A(\ab[3][7] ), .ZN(n2369) );
  NAND3_X2 U2159 ( .A1(n1926), .A2(n1925), .A3(n1924), .ZN(n2370) );
  XNOR2_X2 U2160 ( .A(n2371), .B(\SUMB[3][6] ), .ZN(\SUMB[4][5] ) );
  XNOR2_X2 U2193 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .ZN(n2371) );
  NAND2_X2 U2194 ( .A1(\ab[14][3] ), .A2(\CARRYB[13][3] ), .ZN(n1967) );
  NAND2_X2 U2252 ( .A1(\SUMB[9][5] ), .A2(\ab[10][4] ), .ZN(n1924) );
  XNOR2_X2 U2254 ( .A(n23), .B(\ab[24][0] ), .ZN(n2372) );
  XNOR2_X2 U2335 ( .A(n2372), .B(\CARRYB[23][0] ), .ZN(PRODUCT[24]) );
  NAND3_X2 U2338 ( .A1(net81110), .A2(net81111), .A3(net81112), .ZN(n2373) );
  CLKBUF_X3 U2379 ( .A(\SUMB[15][4] ), .Z(n871) );
  NAND2_X4 U2452 ( .A1(\ab[22][1] ), .A2(\CARRYB[21][1] ), .ZN(net82542) );
  NAND2_X2 U2526 ( .A1(\ab[21][1] ), .A2(\SUMB[20][2] ), .ZN(n2161) );
  CLKBUF_X3 U2579 ( .A(\SUMB[21][1] ), .Z(n1280) );
  NAND2_X4 U2648 ( .A1(n1383), .A2(n1382), .ZN(n11) );
  NAND2_X2 U2734 ( .A1(\SUMB[8][13] ), .A2(net89149), .ZN(net81375) );
  INV_X4 U2772 ( .A(n1456), .ZN(n2374) );
  INV_X2 U2811 ( .A(n1456), .ZN(\SUMB[5][11] ) );
  INV_X2 U3056 ( .A(n585), .ZN(n289) );
  INV_X2 U3114 ( .A(\CARRYB[23][2] ), .ZN(net147938) );
  NAND2_X4 U3232 ( .A1(n1582), .A2(net84708), .ZN(net92542) );
  INV_X2 U3233 ( .A(net88887), .ZN(net88800) );
  INV_X4 U3379 ( .A(\CARRYB[21][4] ), .ZN(n73) );
  OR2_X2 U3381 ( .A1(net81424), .A2(net77964), .ZN(n353) );
  INV_X16 U3386 ( .A(n90), .ZN(net81424) );
  NAND2_X2 U3395 ( .A1(net88303), .A2(\CARRYB[11][10] ), .ZN(net92552) );
  XNOR2_X2 U3396 ( .A(n1309), .B(n1208), .ZN(n2375) );
  NAND2_X4 U3520 ( .A1(\ab[6][7] ), .A2(n853), .ZN(n1331) );
  NAND2_X2 U3536 ( .A1(\CARRYB[6][7] ), .A2(n1499), .ZN(n1443) );
  INV_X4 U3537 ( .A(\SUMB[12][8] ), .ZN(n313) );
  INV_X8 U3548 ( .A(n1277), .ZN(n1278) );
  NAND2_X2 U3549 ( .A1(net82548), .A2(net149580), .ZN(n1124) );
  CLKBUF_X3 U3585 ( .A(n152), .Z(n290) );
  NAND2_X2 U3602 ( .A1(n1730), .A2(n1191), .ZN(n1629) );
  NAND2_X1 U3603 ( .A1(\ab[10][16] ), .A2(\CARRYB[9][16] ), .ZN(n2164) );
  CLKBUF_X2 U3625 ( .A(n2010), .Z(n2376) );
  BUF_X4 U3672 ( .A(\SUMB[5][9] ), .Z(n1214) );
  NAND3_X2 U3678 ( .A1(n1964), .A2(n1966), .A3(n1965), .ZN(n2377) );
  NAND3_X2 U3730 ( .A1(net81216), .A2(n461), .A3(net81215), .ZN(n2378) );
  BUF_X8 U3738 ( .A(\SUMB[18][2] ), .Z(n359) );
  NAND2_X2 U3936 ( .A1(\CARRYB[18][1] ), .A2(\SUMB[18][2] ), .ZN(net81097) );
  INV_X2 U4338 ( .A(net123000), .ZN(net123072) );
  NAND2_X4 U4373 ( .A1(n805), .A2(n660), .ZN(net81992) );
  NAND2_X4 U4466 ( .A1(\CARRYB[4][14] ), .A2(\ab[5][14] ), .ZN(n480) );
  NAND2_X4 U4503 ( .A1(net83919), .A2(\ab[5][14] ), .ZN(n479) );
  NOR2_X1 U4858 ( .A1(net123000), .A2(net70475), .ZN(\ab[10][17] ) );
  XNOR2_X2 U4859 ( .A(n173), .B(\ab[11][7] ), .ZN(n1717) );
  NAND2_X4 U4860 ( .A1(\CARRYB[13][6] ), .A2(\SUMB[13][7] ), .ZN(n1976) );
  NAND2_X4 U4861 ( .A1(\ab[23][2] ), .A2(n394), .ZN(n2295) );
  CLKBUF_X3 U4862 ( .A(\SUMB[9][10] ), .Z(net91419) );
  NAND3_X2 U4863 ( .A1(net119921), .A2(n490), .A3(net82029), .ZN(n123) );
endmodule


module single_cycle ( clk, reset, instructionAddr_out, instruction, 
        dmem_addr_out, dmem_write_out, dmem_read_in, dmem_writeEnable_out, 
        dmem_dsize );
  output [0:31] instructionAddr_out;
  input [0:31] instruction;
  output [0:31] dmem_addr_out;
  output [0:31] dmem_write_out;
  input [0:31] dmem_read_in;
  output [0:1] dmem_dsize;
  input clk, reset;
  output dmem_writeEnable_out;
  wire   n10944, \REGFILE/reg_out[31][31] , \REGFILE/reg_out[31][30] ,
         \REGFILE/reg_out[31][29] , \REGFILE/reg_out[31][28] ,
         \REGFILE/reg_out[31][27] , \REGFILE/reg_out[31][26] ,
         \REGFILE/reg_out[31][25] , \REGFILE/reg_out[31][24] ,
         \REGFILE/reg_out[31][23] , \REGFILE/reg_out[31][22] ,
         \REGFILE/reg_out[31][21] , \REGFILE/reg_out[31][20] ,
         \REGFILE/reg_out[31][19] , \REGFILE/reg_out[31][18] ,
         \REGFILE/reg_out[31][17] , \REGFILE/reg_out[31][16] ,
         \REGFILE/reg_out[31][15] , \REGFILE/reg_out[31][14] ,
         \REGFILE/reg_out[31][13] , \REGFILE/reg_out[31][12] ,
         \REGFILE/reg_out[31][11] , \REGFILE/reg_out[31][10] ,
         \REGFILE/reg_out[31][9] , \REGFILE/reg_out[31][8] ,
         \REGFILE/reg_out[31][7] , \REGFILE/reg_out[31][6] ,
         \REGFILE/reg_out[31][5] , \REGFILE/reg_out[31][4] ,
         \REGFILE/reg_out[31][3] , \REGFILE/reg_out[31][2] ,
         \REGFILE/reg_out[31][1] , \REGFILE/reg_out[31][0] ,
         \REGFILE/reg_out[30][31] , \REGFILE/reg_out[30][30] ,
         \REGFILE/reg_out[30][29] , \REGFILE/reg_out[30][28] ,
         \REGFILE/reg_out[30][27] , \REGFILE/reg_out[30][26] ,
         \REGFILE/reg_out[30][25] , \REGFILE/reg_out[30][24] ,
         \REGFILE/reg_out[30][23] , \REGFILE/reg_out[30][22] ,
         \REGFILE/reg_out[30][21] , \REGFILE/reg_out[30][20] ,
         \REGFILE/reg_out[30][19] , \REGFILE/reg_out[30][18] ,
         \REGFILE/reg_out[30][17] , \REGFILE/reg_out[30][16] ,
         \REGFILE/reg_out[30][15] , \REGFILE/reg_out[30][14] ,
         \REGFILE/reg_out[30][13] , \REGFILE/reg_out[30][12] ,
         \REGFILE/reg_out[30][11] , \REGFILE/reg_out[30][10] ,
         \REGFILE/reg_out[30][9] , \REGFILE/reg_out[30][8] ,
         \REGFILE/reg_out[30][7] , \REGFILE/reg_out[30][6] ,
         \REGFILE/reg_out[30][5] , \REGFILE/reg_out[30][4] ,
         \REGFILE/reg_out[30][3] , \REGFILE/reg_out[30][2] ,
         \REGFILE/reg_out[30][1] , \REGFILE/reg_out[30][0] ,
         \REGFILE/reg_out[29][31] , \REGFILE/reg_out[29][30] ,
         \REGFILE/reg_out[29][29] , \REGFILE/reg_out[29][28] ,
         \REGFILE/reg_out[29][27] , \REGFILE/reg_out[29][26] ,
         \REGFILE/reg_out[29][25] , \REGFILE/reg_out[29][24] ,
         \REGFILE/reg_out[29][23] , \REGFILE/reg_out[29][22] ,
         \REGFILE/reg_out[29][21] , \REGFILE/reg_out[29][20] ,
         \REGFILE/reg_out[29][19] , \REGFILE/reg_out[29][18] ,
         \REGFILE/reg_out[29][17] , \REGFILE/reg_out[29][16] ,
         \REGFILE/reg_out[29][15] , \REGFILE/reg_out[29][14] ,
         \REGFILE/reg_out[29][13] , \REGFILE/reg_out[29][12] ,
         \REGFILE/reg_out[29][11] , \REGFILE/reg_out[29][10] ,
         \REGFILE/reg_out[29][9] , \REGFILE/reg_out[29][8] ,
         \REGFILE/reg_out[29][7] , \REGFILE/reg_out[29][6] ,
         \REGFILE/reg_out[29][5] , \REGFILE/reg_out[29][4] ,
         \REGFILE/reg_out[29][3] , \REGFILE/reg_out[29][2] ,
         \REGFILE/reg_out[29][1] , \REGFILE/reg_out[29][0] ,
         \REGFILE/reg_out[28][31] , \REGFILE/reg_out[28][30] ,
         \REGFILE/reg_out[28][29] , \REGFILE/reg_out[28][28] ,
         \REGFILE/reg_out[28][27] , \REGFILE/reg_out[28][26] ,
         \REGFILE/reg_out[28][25] , \REGFILE/reg_out[28][24] ,
         \REGFILE/reg_out[28][23] , \REGFILE/reg_out[28][22] ,
         \REGFILE/reg_out[28][21] , \REGFILE/reg_out[28][20] ,
         \REGFILE/reg_out[28][19] , \REGFILE/reg_out[28][18] ,
         \REGFILE/reg_out[28][17] , \REGFILE/reg_out[28][16] ,
         \REGFILE/reg_out[28][15] , \REGFILE/reg_out[28][14] ,
         \REGFILE/reg_out[28][13] , \REGFILE/reg_out[28][12] ,
         \REGFILE/reg_out[28][11] , \REGFILE/reg_out[28][10] ,
         \REGFILE/reg_out[28][9] , \REGFILE/reg_out[28][8] ,
         \REGFILE/reg_out[28][7] , \REGFILE/reg_out[28][6] ,
         \REGFILE/reg_out[28][5] , \REGFILE/reg_out[28][4] ,
         \REGFILE/reg_out[28][3] , \REGFILE/reg_out[28][2] ,
         \REGFILE/reg_out[28][1] , \REGFILE/reg_out[28][0] ,
         \REGFILE/reg_out[27][31] , \REGFILE/reg_out[27][30] ,
         \REGFILE/reg_out[27][29] , \REGFILE/reg_out[27][28] ,
         \REGFILE/reg_out[27][27] , \REGFILE/reg_out[27][26] ,
         \REGFILE/reg_out[27][25] , \REGFILE/reg_out[27][24] ,
         \REGFILE/reg_out[27][23] , \REGFILE/reg_out[27][22] ,
         \REGFILE/reg_out[27][21] , \REGFILE/reg_out[27][20] ,
         \REGFILE/reg_out[27][19] , \REGFILE/reg_out[27][18] ,
         \REGFILE/reg_out[27][17] , \REGFILE/reg_out[27][16] ,
         \REGFILE/reg_out[27][15] , \REGFILE/reg_out[27][14] ,
         \REGFILE/reg_out[27][13] , \REGFILE/reg_out[27][12] ,
         \REGFILE/reg_out[27][11] , \REGFILE/reg_out[27][10] ,
         \REGFILE/reg_out[27][9] , \REGFILE/reg_out[27][8] ,
         \REGFILE/reg_out[27][7] , \REGFILE/reg_out[27][6] ,
         \REGFILE/reg_out[27][5] , \REGFILE/reg_out[27][4] ,
         \REGFILE/reg_out[27][3] , \REGFILE/reg_out[27][2] ,
         \REGFILE/reg_out[27][1] , \REGFILE/reg_out[27][0] ,
         \REGFILE/reg_out[26][31] , \REGFILE/reg_out[26][30] ,
         \REGFILE/reg_out[26][29] , \REGFILE/reg_out[26][28] ,
         \REGFILE/reg_out[26][27] , \REGFILE/reg_out[26][26] ,
         \REGFILE/reg_out[26][25] , \REGFILE/reg_out[26][24] ,
         \REGFILE/reg_out[26][23] , \REGFILE/reg_out[26][22] ,
         \REGFILE/reg_out[26][21] , \REGFILE/reg_out[26][20] ,
         \REGFILE/reg_out[26][19] , \REGFILE/reg_out[26][18] ,
         \REGFILE/reg_out[26][17] , \REGFILE/reg_out[26][16] ,
         \REGFILE/reg_out[26][15] , \REGFILE/reg_out[26][14] ,
         \REGFILE/reg_out[26][13] , \REGFILE/reg_out[26][12] ,
         \REGFILE/reg_out[26][11] , \REGFILE/reg_out[26][10] ,
         \REGFILE/reg_out[26][9] , \REGFILE/reg_out[26][8] ,
         \REGFILE/reg_out[26][7] , \REGFILE/reg_out[26][6] ,
         \REGFILE/reg_out[26][5] , \REGFILE/reg_out[26][4] ,
         \REGFILE/reg_out[26][3] , \REGFILE/reg_out[26][2] ,
         \REGFILE/reg_out[26][1] , \REGFILE/reg_out[26][0] ,
         \REGFILE/reg_out[25][31] , \REGFILE/reg_out[25][30] ,
         \REGFILE/reg_out[25][29] , \REGFILE/reg_out[25][28] ,
         \REGFILE/reg_out[25][27] , \REGFILE/reg_out[25][26] ,
         \REGFILE/reg_out[25][25] , \REGFILE/reg_out[25][24] ,
         \REGFILE/reg_out[25][23] , \REGFILE/reg_out[25][22] ,
         \REGFILE/reg_out[25][21] , \REGFILE/reg_out[25][20] ,
         \REGFILE/reg_out[25][19] , \REGFILE/reg_out[25][18] ,
         \REGFILE/reg_out[25][17] , \REGFILE/reg_out[25][16] ,
         \REGFILE/reg_out[25][15] , \REGFILE/reg_out[25][14] ,
         \REGFILE/reg_out[25][13] , \REGFILE/reg_out[25][12] ,
         \REGFILE/reg_out[25][11] , \REGFILE/reg_out[25][10] ,
         \REGFILE/reg_out[25][9] , \REGFILE/reg_out[25][8] ,
         \REGFILE/reg_out[25][7] , \REGFILE/reg_out[25][5] ,
         \REGFILE/reg_out[25][4] , \REGFILE/reg_out[25][3] ,
         \REGFILE/reg_out[25][2] , \REGFILE/reg_out[25][1] ,
         \REGFILE/reg_out[25][0] , \REGFILE/reg_out[24][31] ,
         \REGFILE/reg_out[24][30] , \REGFILE/reg_out[24][29] ,
         \REGFILE/reg_out[24][28] , \REGFILE/reg_out[24][27] ,
         \REGFILE/reg_out[24][26] , \REGFILE/reg_out[24][25] ,
         \REGFILE/reg_out[24][24] , \REGFILE/reg_out[24][23] ,
         \REGFILE/reg_out[24][22] , \REGFILE/reg_out[24][21] ,
         \REGFILE/reg_out[24][20] , \REGFILE/reg_out[24][19] ,
         \REGFILE/reg_out[24][18] , \REGFILE/reg_out[24][17] ,
         \REGFILE/reg_out[24][16] , \REGFILE/reg_out[24][15] ,
         \REGFILE/reg_out[24][14] , \REGFILE/reg_out[24][13] ,
         \REGFILE/reg_out[24][12] , \REGFILE/reg_out[24][11] ,
         \REGFILE/reg_out[24][10] , \REGFILE/reg_out[24][9] ,
         \REGFILE/reg_out[24][8] , \REGFILE/reg_out[24][7] ,
         \REGFILE/reg_out[24][6] , \REGFILE/reg_out[24][5] ,
         \REGFILE/reg_out[24][4] , \REGFILE/reg_out[24][3] ,
         \REGFILE/reg_out[24][2] , \REGFILE/reg_out[24][1] ,
         \REGFILE/reg_out[24][0] , \REGFILE/reg_out[23][31] ,
         \REGFILE/reg_out[23][30] , \REGFILE/reg_out[23][29] ,
         \REGFILE/reg_out[23][28] , \REGFILE/reg_out[23][27] ,
         \REGFILE/reg_out[23][26] , \REGFILE/reg_out[23][25] ,
         \REGFILE/reg_out[23][24] , \REGFILE/reg_out[23][23] ,
         \REGFILE/reg_out[23][22] , \REGFILE/reg_out[23][21] ,
         \REGFILE/reg_out[23][20] , \REGFILE/reg_out[23][19] ,
         \REGFILE/reg_out[23][18] , \REGFILE/reg_out[23][17] ,
         \REGFILE/reg_out[23][16] , \REGFILE/reg_out[23][15] ,
         \REGFILE/reg_out[23][14] , \REGFILE/reg_out[23][13] ,
         \REGFILE/reg_out[23][12] , \REGFILE/reg_out[23][11] ,
         \REGFILE/reg_out[23][10] , \REGFILE/reg_out[23][9] ,
         \REGFILE/reg_out[23][8] , \REGFILE/reg_out[23][7] ,
         \REGFILE/reg_out[23][6] , \REGFILE/reg_out[23][5] ,
         \REGFILE/reg_out[23][4] , \REGFILE/reg_out[23][3] ,
         \REGFILE/reg_out[23][2] , \REGFILE/reg_out[23][1] ,
         \REGFILE/reg_out[23][0] , \REGFILE/reg_out[22][31] ,
         \REGFILE/reg_out[22][30] , \REGFILE/reg_out[22][29] ,
         \REGFILE/reg_out[22][28] , \REGFILE/reg_out[22][27] ,
         \REGFILE/reg_out[22][26] , \REGFILE/reg_out[22][25] ,
         \REGFILE/reg_out[22][24] , \REGFILE/reg_out[22][23] ,
         \REGFILE/reg_out[22][22] , \REGFILE/reg_out[22][21] ,
         \REGFILE/reg_out[22][20] , \REGFILE/reg_out[22][19] ,
         \REGFILE/reg_out[22][18] , \REGFILE/reg_out[22][17] ,
         \REGFILE/reg_out[22][16] , \REGFILE/reg_out[22][15] ,
         \REGFILE/reg_out[22][14] , \REGFILE/reg_out[22][13] ,
         \REGFILE/reg_out[22][12] , \REGFILE/reg_out[22][11] ,
         \REGFILE/reg_out[22][10] , \REGFILE/reg_out[22][9] ,
         \REGFILE/reg_out[22][8] , \REGFILE/reg_out[22][7] ,
         \REGFILE/reg_out[22][6] , \REGFILE/reg_out[22][5] ,
         \REGFILE/reg_out[22][4] , \REGFILE/reg_out[22][3] ,
         \REGFILE/reg_out[22][2] , \REGFILE/reg_out[22][1] ,
         \REGFILE/reg_out[22][0] , \REGFILE/reg_out[21][31] ,
         \REGFILE/reg_out[21][30] , \REGFILE/reg_out[21][29] ,
         \REGFILE/reg_out[21][28] , \REGFILE/reg_out[21][27] ,
         \REGFILE/reg_out[21][26] , \REGFILE/reg_out[21][25] ,
         \REGFILE/reg_out[21][24] , \REGFILE/reg_out[21][23] ,
         \REGFILE/reg_out[21][22] , \REGFILE/reg_out[21][21] ,
         \REGFILE/reg_out[21][20] , \REGFILE/reg_out[21][19] ,
         \REGFILE/reg_out[21][18] , \REGFILE/reg_out[21][17] ,
         \REGFILE/reg_out[21][16] , \REGFILE/reg_out[21][15] ,
         \REGFILE/reg_out[21][14] , \REGFILE/reg_out[21][13] ,
         \REGFILE/reg_out[21][12] , \REGFILE/reg_out[21][11] ,
         \REGFILE/reg_out[21][10] , \REGFILE/reg_out[21][9] ,
         \REGFILE/reg_out[21][8] , \REGFILE/reg_out[21][7] ,
         \REGFILE/reg_out[21][6] , \REGFILE/reg_out[21][5] ,
         \REGFILE/reg_out[21][4] , \REGFILE/reg_out[21][3] ,
         \REGFILE/reg_out[21][2] , \REGFILE/reg_out[21][1] ,
         \REGFILE/reg_out[21][0] , \REGFILE/reg_out[20][31] ,
         \REGFILE/reg_out[20][30] , \REGFILE/reg_out[20][29] ,
         \REGFILE/reg_out[20][28] , \REGFILE/reg_out[20][27] ,
         \REGFILE/reg_out[20][26] , \REGFILE/reg_out[20][25] ,
         \REGFILE/reg_out[20][24] , \REGFILE/reg_out[20][23] ,
         \REGFILE/reg_out[20][22] , \REGFILE/reg_out[20][21] ,
         \REGFILE/reg_out[20][20] , \REGFILE/reg_out[20][19] ,
         \REGFILE/reg_out[20][18] , \REGFILE/reg_out[20][17] ,
         \REGFILE/reg_out[20][16] , \REGFILE/reg_out[20][15] ,
         \REGFILE/reg_out[20][14] , \REGFILE/reg_out[20][13] ,
         \REGFILE/reg_out[20][12] , \REGFILE/reg_out[20][11] ,
         \REGFILE/reg_out[20][10] , \REGFILE/reg_out[20][9] ,
         \REGFILE/reg_out[20][8] , \REGFILE/reg_out[20][7] ,
         \REGFILE/reg_out[20][6] , \REGFILE/reg_out[20][5] ,
         \REGFILE/reg_out[20][4] , \REGFILE/reg_out[20][3] ,
         \REGFILE/reg_out[20][2] , \REGFILE/reg_out[20][1] ,
         \REGFILE/reg_out[20][0] , \REGFILE/reg_out[19][31] ,
         \REGFILE/reg_out[19][30] , \REGFILE/reg_out[19][29] ,
         \REGFILE/reg_out[19][28] , \REGFILE/reg_out[19][27] ,
         \REGFILE/reg_out[19][26] , \REGFILE/reg_out[19][25] ,
         \REGFILE/reg_out[19][24] , \REGFILE/reg_out[19][23] ,
         \REGFILE/reg_out[19][22] , \REGFILE/reg_out[19][21] ,
         \REGFILE/reg_out[19][20] , \REGFILE/reg_out[19][19] ,
         \REGFILE/reg_out[19][18] , \REGFILE/reg_out[19][17] ,
         \REGFILE/reg_out[19][16] , \REGFILE/reg_out[19][15] ,
         \REGFILE/reg_out[19][14] , \REGFILE/reg_out[19][13] ,
         \REGFILE/reg_out[19][12] , \REGFILE/reg_out[19][11] ,
         \REGFILE/reg_out[19][10] , \REGFILE/reg_out[19][9] ,
         \REGFILE/reg_out[19][8] , \REGFILE/reg_out[19][7] ,
         \REGFILE/reg_out[19][6] , \REGFILE/reg_out[19][5] ,
         \REGFILE/reg_out[19][4] , \REGFILE/reg_out[19][3] ,
         \REGFILE/reg_out[19][2] , \REGFILE/reg_out[19][1] ,
         \REGFILE/reg_out[19][0] , \REGFILE/reg_out[18][31] ,
         \REGFILE/reg_out[18][30] , \REGFILE/reg_out[18][29] ,
         \REGFILE/reg_out[18][28] , \REGFILE/reg_out[18][27] ,
         \REGFILE/reg_out[18][26] , \REGFILE/reg_out[18][25] ,
         \REGFILE/reg_out[18][24] , \REGFILE/reg_out[18][23] ,
         \REGFILE/reg_out[18][22] , \REGFILE/reg_out[18][21] ,
         \REGFILE/reg_out[18][20] , \REGFILE/reg_out[18][19] ,
         \REGFILE/reg_out[18][18] , \REGFILE/reg_out[18][17] ,
         \REGFILE/reg_out[18][16] , \REGFILE/reg_out[18][15] ,
         \REGFILE/reg_out[18][14] , \REGFILE/reg_out[18][13] ,
         \REGFILE/reg_out[18][12] , \REGFILE/reg_out[18][11] ,
         \REGFILE/reg_out[18][10] , \REGFILE/reg_out[18][9] ,
         \REGFILE/reg_out[18][8] , \REGFILE/reg_out[18][7] ,
         \REGFILE/reg_out[18][6] , \REGFILE/reg_out[18][5] ,
         \REGFILE/reg_out[18][4] , \REGFILE/reg_out[18][3] ,
         \REGFILE/reg_out[18][2] , \REGFILE/reg_out[18][1] ,
         \REGFILE/reg_out[18][0] , \REGFILE/reg_out[17][31] ,
         \REGFILE/reg_out[17][30] , \REGFILE/reg_out[17][29] ,
         \REGFILE/reg_out[17][28] , \REGFILE/reg_out[17][27] ,
         \REGFILE/reg_out[17][26] , \REGFILE/reg_out[17][25] ,
         \REGFILE/reg_out[17][24] , \REGFILE/reg_out[17][23] ,
         \REGFILE/reg_out[17][22] , \REGFILE/reg_out[17][21] ,
         \REGFILE/reg_out[17][20] , \REGFILE/reg_out[17][19] ,
         \REGFILE/reg_out[17][18] , \REGFILE/reg_out[17][17] ,
         \REGFILE/reg_out[17][16] , \REGFILE/reg_out[17][15] ,
         \REGFILE/reg_out[17][14] , \REGFILE/reg_out[17][13] ,
         \REGFILE/reg_out[17][12] , \REGFILE/reg_out[17][11] ,
         \REGFILE/reg_out[17][10] , \REGFILE/reg_out[17][9] ,
         \REGFILE/reg_out[17][8] , \REGFILE/reg_out[17][7] ,
         \REGFILE/reg_out[17][6] , \REGFILE/reg_out[17][5] ,
         \REGFILE/reg_out[17][4] , \REGFILE/reg_out[17][3] ,
         \REGFILE/reg_out[17][2] , \REGFILE/reg_out[17][1] ,
         \REGFILE/reg_out[17][0] , \REGFILE/reg_out[16][31] ,
         \REGFILE/reg_out[16][30] , \REGFILE/reg_out[16][29] ,
         \REGFILE/reg_out[16][28] , \REGFILE/reg_out[16][27] ,
         \REGFILE/reg_out[16][26] , \REGFILE/reg_out[16][25] ,
         \REGFILE/reg_out[16][24] , \REGFILE/reg_out[16][23] ,
         \REGFILE/reg_out[16][22] , \REGFILE/reg_out[16][21] ,
         \REGFILE/reg_out[16][20] , \REGFILE/reg_out[16][19] ,
         \REGFILE/reg_out[16][18] , \REGFILE/reg_out[16][17] ,
         \REGFILE/reg_out[16][16] , \REGFILE/reg_out[16][15] ,
         \REGFILE/reg_out[16][14] , \REGFILE/reg_out[16][13] ,
         \REGFILE/reg_out[16][12] , \REGFILE/reg_out[16][11] ,
         \REGFILE/reg_out[16][10] , \REGFILE/reg_out[16][9] ,
         \REGFILE/reg_out[16][8] , \REGFILE/reg_out[16][7] ,
         \REGFILE/reg_out[16][6] , \REGFILE/reg_out[16][5] ,
         \REGFILE/reg_out[16][4] , \REGFILE/reg_out[16][3] ,
         \REGFILE/reg_out[16][2] , \REGFILE/reg_out[16][1] ,
         \REGFILE/reg_out[16][0] , \REGFILE/reg_out[15][31] ,
         \REGFILE/reg_out[15][30] , \REGFILE/reg_out[15][29] ,
         \REGFILE/reg_out[15][28] , \REGFILE/reg_out[15][27] ,
         \REGFILE/reg_out[15][26] , \REGFILE/reg_out[15][25] ,
         \REGFILE/reg_out[15][24] , \REGFILE/reg_out[15][23] ,
         \REGFILE/reg_out[15][22] , \REGFILE/reg_out[15][21] ,
         \REGFILE/reg_out[15][20] , \REGFILE/reg_out[15][19] ,
         \REGFILE/reg_out[15][18] , \REGFILE/reg_out[15][17] ,
         \REGFILE/reg_out[15][16] , \REGFILE/reg_out[15][15] ,
         \REGFILE/reg_out[15][14] , \REGFILE/reg_out[15][13] ,
         \REGFILE/reg_out[15][12] , \REGFILE/reg_out[15][11] ,
         \REGFILE/reg_out[15][10] , \REGFILE/reg_out[15][9] ,
         \REGFILE/reg_out[15][8] , \REGFILE/reg_out[15][7] ,
         \REGFILE/reg_out[15][6] , \REGFILE/reg_out[15][5] ,
         \REGFILE/reg_out[15][4] , \REGFILE/reg_out[15][3] ,
         \REGFILE/reg_out[15][2] , \REGFILE/reg_out[15][1] ,
         \REGFILE/reg_out[15][0] , \REGFILE/reg_out[14][31] ,
         \REGFILE/reg_out[14][30] , \REGFILE/reg_out[14][29] ,
         \REGFILE/reg_out[14][28] , \REGFILE/reg_out[14][27] ,
         \REGFILE/reg_out[14][26] , \REGFILE/reg_out[14][25] ,
         \REGFILE/reg_out[14][24] , \REGFILE/reg_out[14][23] ,
         \REGFILE/reg_out[14][22] , \REGFILE/reg_out[14][21] ,
         \REGFILE/reg_out[14][20] , \REGFILE/reg_out[14][19] ,
         \REGFILE/reg_out[14][18] , \REGFILE/reg_out[14][17] ,
         \REGFILE/reg_out[14][16] , \REGFILE/reg_out[14][15] ,
         \REGFILE/reg_out[14][14] , \REGFILE/reg_out[14][13] ,
         \REGFILE/reg_out[14][12] , \REGFILE/reg_out[14][11] ,
         \REGFILE/reg_out[14][10] , \REGFILE/reg_out[14][9] ,
         \REGFILE/reg_out[14][8] , \REGFILE/reg_out[14][7] ,
         \REGFILE/reg_out[14][6] , \REGFILE/reg_out[14][5] ,
         \REGFILE/reg_out[14][4] , \REGFILE/reg_out[14][3] ,
         \REGFILE/reg_out[14][2] , \REGFILE/reg_out[14][1] ,
         \REGFILE/reg_out[14][0] , \REGFILE/reg_out[13][31] ,
         \REGFILE/reg_out[13][30] , \REGFILE/reg_out[13][29] ,
         \REGFILE/reg_out[13][28] , \REGFILE/reg_out[13][27] ,
         \REGFILE/reg_out[13][26] , \REGFILE/reg_out[13][25] ,
         \REGFILE/reg_out[13][24] , \REGFILE/reg_out[13][23] ,
         \REGFILE/reg_out[13][22] , \REGFILE/reg_out[13][21] ,
         \REGFILE/reg_out[13][20] , \REGFILE/reg_out[13][19] ,
         \REGFILE/reg_out[13][18] , \REGFILE/reg_out[13][17] ,
         \REGFILE/reg_out[13][16] , \REGFILE/reg_out[13][15] ,
         \REGFILE/reg_out[13][14] , \REGFILE/reg_out[13][13] ,
         \REGFILE/reg_out[13][12] , \REGFILE/reg_out[13][11] ,
         \REGFILE/reg_out[13][10] , \REGFILE/reg_out[13][9] ,
         \REGFILE/reg_out[13][8] , \REGFILE/reg_out[13][7] ,
         \REGFILE/reg_out[13][6] , \REGFILE/reg_out[13][5] ,
         \REGFILE/reg_out[13][4] , \REGFILE/reg_out[13][3] ,
         \REGFILE/reg_out[13][2] , \REGFILE/reg_out[13][1] ,
         \REGFILE/reg_out[13][0] , \REGFILE/reg_out[12][31] ,
         \REGFILE/reg_out[12][30] , \REGFILE/reg_out[12][29] ,
         \REGFILE/reg_out[12][28] , \REGFILE/reg_out[12][27] ,
         \REGFILE/reg_out[12][26] , \REGFILE/reg_out[12][25] ,
         \REGFILE/reg_out[12][24] , \REGFILE/reg_out[12][23] ,
         \REGFILE/reg_out[12][22] , \REGFILE/reg_out[12][21] ,
         \REGFILE/reg_out[12][20] , \REGFILE/reg_out[12][19] ,
         \REGFILE/reg_out[12][18] , \REGFILE/reg_out[12][17] ,
         \REGFILE/reg_out[12][16] , \REGFILE/reg_out[12][15] ,
         \REGFILE/reg_out[12][13] , \REGFILE/reg_out[12][12] ,
         \REGFILE/reg_out[12][11] , \REGFILE/reg_out[12][10] ,
         \REGFILE/reg_out[12][9] , \REGFILE/reg_out[12][8] ,
         \REGFILE/reg_out[12][7] , \REGFILE/reg_out[12][6] ,
         \REGFILE/reg_out[12][5] , \REGFILE/reg_out[12][4] ,
         \REGFILE/reg_out[12][3] , \REGFILE/reg_out[12][2] ,
         \REGFILE/reg_out[12][1] , \REGFILE/reg_out[12][0] ,
         \REGFILE/reg_out[11][31] , \REGFILE/reg_out[11][30] ,
         \REGFILE/reg_out[11][29] , \REGFILE/reg_out[11][28] ,
         \REGFILE/reg_out[11][27] , \REGFILE/reg_out[11][26] ,
         \REGFILE/reg_out[11][25] , \REGFILE/reg_out[11][24] ,
         \REGFILE/reg_out[11][23] , \REGFILE/reg_out[11][22] ,
         \REGFILE/reg_out[11][21] , \REGFILE/reg_out[11][20] ,
         \REGFILE/reg_out[11][19] , \REGFILE/reg_out[11][18] ,
         \REGFILE/reg_out[11][17] , \REGFILE/reg_out[11][16] ,
         \REGFILE/reg_out[11][15] , \REGFILE/reg_out[11][14] ,
         \REGFILE/reg_out[11][13] , \REGFILE/reg_out[11][12] ,
         \REGFILE/reg_out[11][11] , \REGFILE/reg_out[11][10] ,
         \REGFILE/reg_out[11][9] , \REGFILE/reg_out[11][8] ,
         \REGFILE/reg_out[11][7] , \REGFILE/reg_out[11][6] ,
         \REGFILE/reg_out[11][5] , \REGFILE/reg_out[11][4] ,
         \REGFILE/reg_out[11][3] , \REGFILE/reg_out[11][2] ,
         \REGFILE/reg_out[11][1] , \REGFILE/reg_out[11][0] ,
         \REGFILE/reg_out[10][31] , \REGFILE/reg_out[10][30] ,
         \REGFILE/reg_out[10][29] , \REGFILE/reg_out[10][28] ,
         \REGFILE/reg_out[10][27] , \REGFILE/reg_out[10][26] ,
         \REGFILE/reg_out[10][25] , \REGFILE/reg_out[10][24] ,
         \REGFILE/reg_out[10][23] , \REGFILE/reg_out[10][22] ,
         \REGFILE/reg_out[10][21] , \REGFILE/reg_out[10][20] ,
         \REGFILE/reg_out[10][19] , \REGFILE/reg_out[10][18] ,
         \REGFILE/reg_out[10][17] , \REGFILE/reg_out[10][16] ,
         \REGFILE/reg_out[10][15] , \REGFILE/reg_out[10][14] ,
         \REGFILE/reg_out[10][13] , \REGFILE/reg_out[10][12] ,
         \REGFILE/reg_out[10][11] , \REGFILE/reg_out[10][10] ,
         \REGFILE/reg_out[10][9] , \REGFILE/reg_out[10][8] ,
         \REGFILE/reg_out[10][7] , \REGFILE/reg_out[10][5] ,
         \REGFILE/reg_out[10][4] , \REGFILE/reg_out[10][3] ,
         \REGFILE/reg_out[10][2] , \REGFILE/reg_out[10][1] ,
         \REGFILE/reg_out[10][0] , \REGFILE/reg_out[9][31] ,
         \REGFILE/reg_out[9][30] , \REGFILE/reg_out[9][29] ,
         \REGFILE/reg_out[9][28] , \REGFILE/reg_out[9][27] ,
         \REGFILE/reg_out[9][26] , \REGFILE/reg_out[9][25] ,
         \REGFILE/reg_out[9][24] , \REGFILE/reg_out[9][23] ,
         \REGFILE/reg_out[9][22] , \REGFILE/reg_out[9][21] ,
         \REGFILE/reg_out[9][20] , \REGFILE/reg_out[9][19] ,
         \REGFILE/reg_out[9][18] , \REGFILE/reg_out[9][17] ,
         \REGFILE/reg_out[9][16] , \REGFILE/reg_out[9][15] ,
         \REGFILE/reg_out[9][14] , \REGFILE/reg_out[9][13] ,
         \REGFILE/reg_out[9][12] , \REGFILE/reg_out[9][11] ,
         \REGFILE/reg_out[9][10] , \REGFILE/reg_out[9][9] ,
         \REGFILE/reg_out[9][8] , \REGFILE/reg_out[9][7] ,
         \REGFILE/reg_out[9][6] , \REGFILE/reg_out[9][5] ,
         \REGFILE/reg_out[9][4] , \REGFILE/reg_out[9][3] ,
         \REGFILE/reg_out[9][2] , \REGFILE/reg_out[9][1] ,
         \REGFILE/reg_out[9][0] , \REGFILE/reg_out[8][31] ,
         \REGFILE/reg_out[8][30] , \REGFILE/reg_out[8][29] ,
         \REGFILE/reg_out[8][28] , \REGFILE/reg_out[8][27] ,
         \REGFILE/reg_out[8][26] , \REGFILE/reg_out[8][25] ,
         \REGFILE/reg_out[8][24] , \REGFILE/reg_out[8][23] ,
         \REGFILE/reg_out[8][22] , \REGFILE/reg_out[8][21] ,
         \REGFILE/reg_out[8][20] , \REGFILE/reg_out[8][19] ,
         \REGFILE/reg_out[8][18] , \REGFILE/reg_out[8][17] ,
         \REGFILE/reg_out[8][16] , \REGFILE/reg_out[8][15] ,
         \REGFILE/reg_out[8][14] , \REGFILE/reg_out[8][13] ,
         \REGFILE/reg_out[8][12] , \REGFILE/reg_out[8][11] ,
         \REGFILE/reg_out[8][10] , \REGFILE/reg_out[8][9] ,
         \REGFILE/reg_out[8][8] , \REGFILE/reg_out[8][7] ,
         \REGFILE/reg_out[8][6] , \REGFILE/reg_out[8][5] ,
         \REGFILE/reg_out[8][4] , \REGFILE/reg_out[8][3] ,
         \REGFILE/reg_out[8][2] , \REGFILE/reg_out[8][1] ,
         \REGFILE/reg_out[8][0] , \REGFILE/reg_out[7][31] ,
         \REGFILE/reg_out[7][30] , \REGFILE/reg_out[7][29] ,
         \REGFILE/reg_out[7][28] , \REGFILE/reg_out[7][27] ,
         \REGFILE/reg_out[7][26] , \REGFILE/reg_out[7][25] ,
         \REGFILE/reg_out[7][24] , \REGFILE/reg_out[7][23] ,
         \REGFILE/reg_out[7][22] , \REGFILE/reg_out[7][21] ,
         \REGFILE/reg_out[7][20] , \REGFILE/reg_out[7][19] ,
         \REGFILE/reg_out[7][18] , \REGFILE/reg_out[7][17] ,
         \REGFILE/reg_out[7][16] , \REGFILE/reg_out[7][15] ,
         \REGFILE/reg_out[7][14] , \REGFILE/reg_out[7][13] ,
         \REGFILE/reg_out[7][12] , \REGFILE/reg_out[7][11] ,
         \REGFILE/reg_out[7][10] , \REGFILE/reg_out[7][9] ,
         \REGFILE/reg_out[7][8] , \REGFILE/reg_out[7][7] ,
         \REGFILE/reg_out[7][6] , \REGFILE/reg_out[7][5] ,
         \REGFILE/reg_out[7][4] , \REGFILE/reg_out[7][3] ,
         \REGFILE/reg_out[7][2] , \REGFILE/reg_out[7][1] ,
         \REGFILE/reg_out[7][0] , \REGFILE/reg_out[6][31] ,
         \REGFILE/reg_out[6][30] , \REGFILE/reg_out[6][29] ,
         \REGFILE/reg_out[6][28] , \REGFILE/reg_out[6][27] ,
         \REGFILE/reg_out[6][26] , \REGFILE/reg_out[6][25] ,
         \REGFILE/reg_out[6][24] , \REGFILE/reg_out[6][23] ,
         \REGFILE/reg_out[6][22] , \REGFILE/reg_out[6][21] ,
         \REGFILE/reg_out[6][20] , \REGFILE/reg_out[6][19] ,
         \REGFILE/reg_out[6][18] , \REGFILE/reg_out[6][17] ,
         \REGFILE/reg_out[6][16] , \REGFILE/reg_out[6][15] ,
         \REGFILE/reg_out[6][14] , \REGFILE/reg_out[6][13] ,
         \REGFILE/reg_out[6][12] , \REGFILE/reg_out[6][11] ,
         \REGFILE/reg_out[6][10] , \REGFILE/reg_out[6][9] ,
         \REGFILE/reg_out[6][8] , \REGFILE/reg_out[6][7] ,
         \REGFILE/reg_out[6][6] , \REGFILE/reg_out[6][5] ,
         \REGFILE/reg_out[6][4] , \REGFILE/reg_out[6][3] ,
         \REGFILE/reg_out[6][2] , \REGFILE/reg_out[6][1] ,
         \REGFILE/reg_out[6][0] , \REGFILE/reg_out[5][31] ,
         \REGFILE/reg_out[5][30] , \REGFILE/reg_out[5][29] ,
         \REGFILE/reg_out[5][28] , \REGFILE/reg_out[5][27] ,
         \REGFILE/reg_out[5][26] , \REGFILE/reg_out[5][25] ,
         \REGFILE/reg_out[5][24] , \REGFILE/reg_out[5][23] ,
         \REGFILE/reg_out[5][22] , \REGFILE/reg_out[5][21] ,
         \REGFILE/reg_out[5][20] , \REGFILE/reg_out[5][19] ,
         \REGFILE/reg_out[5][18] , \REGFILE/reg_out[5][17] ,
         \REGFILE/reg_out[5][16] , \REGFILE/reg_out[5][15] ,
         \REGFILE/reg_out[5][14] , \REGFILE/reg_out[5][13] ,
         \REGFILE/reg_out[5][12] , \REGFILE/reg_out[5][11] ,
         \REGFILE/reg_out[5][10] , \REGFILE/reg_out[5][9] ,
         \REGFILE/reg_out[5][8] , \REGFILE/reg_out[5][7] ,
         \REGFILE/reg_out[5][6] , \REGFILE/reg_out[5][5] ,
         \REGFILE/reg_out[5][4] , \REGFILE/reg_out[5][3] ,
         \REGFILE/reg_out[5][2] , \REGFILE/reg_out[5][1] ,
         \REGFILE/reg_out[5][0] , \REGFILE/reg_out[4][31] ,
         \REGFILE/reg_out[4][30] , \REGFILE/reg_out[4][29] ,
         \REGFILE/reg_out[4][28] , \REGFILE/reg_out[4][27] ,
         \REGFILE/reg_out[4][26] , \REGFILE/reg_out[4][25] ,
         \REGFILE/reg_out[4][24] , \REGFILE/reg_out[4][23] ,
         \REGFILE/reg_out[4][22] , \REGFILE/reg_out[4][21] ,
         \REGFILE/reg_out[4][20] , \REGFILE/reg_out[4][19] ,
         \REGFILE/reg_out[4][18] , \REGFILE/reg_out[4][17] ,
         \REGFILE/reg_out[4][16] , \REGFILE/reg_out[4][15] ,
         \REGFILE/reg_out[4][14] , \REGFILE/reg_out[4][13] ,
         \REGFILE/reg_out[4][12] , \REGFILE/reg_out[4][11] ,
         \REGFILE/reg_out[4][10] , \REGFILE/reg_out[4][9] ,
         \REGFILE/reg_out[4][8] , \REGFILE/reg_out[4][7] ,
         \REGFILE/reg_out[4][6] , \REGFILE/reg_out[4][5] ,
         \REGFILE/reg_out[4][4] , \REGFILE/reg_out[4][3] ,
         \REGFILE/reg_out[4][2] , \REGFILE/reg_out[4][1] ,
         \REGFILE/reg_out[4][0] , \REGFILE/reg_out[3][31] ,
         \REGFILE/reg_out[3][30] , \REGFILE/reg_out[3][29] ,
         \REGFILE/reg_out[3][28] , \REGFILE/reg_out[3][27] ,
         \REGFILE/reg_out[3][26] , \REGFILE/reg_out[3][25] ,
         \REGFILE/reg_out[3][24] , \REGFILE/reg_out[3][23] ,
         \REGFILE/reg_out[3][22] , \REGFILE/reg_out[3][21] ,
         \REGFILE/reg_out[3][20] , \REGFILE/reg_out[3][19] ,
         \REGFILE/reg_out[3][18] , \REGFILE/reg_out[3][17] ,
         \REGFILE/reg_out[3][16] , \REGFILE/reg_out[3][15] ,
         \REGFILE/reg_out[3][14] , \REGFILE/reg_out[3][13] ,
         \REGFILE/reg_out[3][12] , \REGFILE/reg_out[3][11] ,
         \REGFILE/reg_out[3][10] , \REGFILE/reg_out[3][9] ,
         \REGFILE/reg_out[3][8] , \REGFILE/reg_out[3][7] ,
         \REGFILE/reg_out[3][6] , \REGFILE/reg_out[3][5] ,
         \REGFILE/reg_out[3][3] , \REGFILE/reg_out[3][2] ,
         \REGFILE/reg_out[3][1] , \REGFILE/reg_out[3][0] ,
         \REGFILE/reg_out[2][31] , \REGFILE/reg_out[2][30] ,
         \REGFILE/reg_out[2][29] , \REGFILE/reg_out[2][28] ,
         \REGFILE/reg_out[2][27] , \REGFILE/reg_out[2][26] ,
         \REGFILE/reg_out[2][25] , \REGFILE/reg_out[2][24] ,
         \REGFILE/reg_out[2][23] , \REGFILE/reg_out[2][22] ,
         \REGFILE/reg_out[2][21] , \REGFILE/reg_out[2][20] ,
         \REGFILE/reg_out[2][19] , \REGFILE/reg_out[2][18] ,
         \REGFILE/reg_out[2][17] , \REGFILE/reg_out[2][16] ,
         \REGFILE/reg_out[2][15] , \REGFILE/reg_out[2][14] ,
         \REGFILE/reg_out[2][13] , \REGFILE/reg_out[2][12] ,
         \REGFILE/reg_out[2][11] , \REGFILE/reg_out[2][10] ,
         \REGFILE/reg_out[2][9] , \REGFILE/reg_out[2][8] ,
         \REGFILE/reg_out[2][7] , \REGFILE/reg_out[2][6] ,
         \REGFILE/reg_out[2][5] , \REGFILE/reg_out[2][4] ,
         \REGFILE/reg_out[2][3] , \REGFILE/reg_out[2][2] ,
         \REGFILE/reg_out[2][1] , \REGFILE/reg_out[2][0] ,
         \REGFILE/reg_out[1][31] , \REGFILE/reg_out[1][30] ,
         \REGFILE/reg_out[1][29] , \REGFILE/reg_out[1][28] ,
         \REGFILE/reg_out[1][27] , \REGFILE/reg_out[1][26] ,
         \REGFILE/reg_out[1][25] , \REGFILE/reg_out[1][24] ,
         \REGFILE/reg_out[1][23] , \REGFILE/reg_out[1][22] ,
         \REGFILE/reg_out[1][21] , \REGFILE/reg_out[1][20] ,
         \REGFILE/reg_out[1][19] , \REGFILE/reg_out[1][18] ,
         \REGFILE/reg_out[1][17] , \REGFILE/reg_out[1][16] ,
         \REGFILE/reg_out[1][15] , \REGFILE/reg_out[1][14] ,
         \REGFILE/reg_out[1][13] , \REGFILE/reg_out[1][12] ,
         \REGFILE/reg_out[1][11] , \REGFILE/reg_out[1][10] ,
         \REGFILE/reg_out[1][9] , \REGFILE/reg_out[1][8] ,
         \REGFILE/reg_out[1][7] , \REGFILE/reg_out[1][6] ,
         \REGFILE/reg_out[1][5] , \REGFILE/reg_out[1][4] ,
         \REGFILE/reg_out[1][3] , \REGFILE/reg_out[1][2] ,
         \REGFILE/reg_out[1][1] , \REGFILE/reg_out[1][0] ,
         \REGFILE/reg_out[0][31] , \REGFILE/reg_out[0][30] ,
         \REGFILE/reg_out[0][29] , \REGFILE/reg_out[0][28] ,
         \REGFILE/reg_out[0][27] , \REGFILE/reg_out[0][26] ,
         \REGFILE/reg_out[0][25] , \REGFILE/reg_out[0][24] ,
         \REGFILE/reg_out[0][23] , \REGFILE/reg_out[0][22] ,
         \REGFILE/reg_out[0][21] , \REGFILE/reg_out[0][20] ,
         \REGFILE/reg_out[0][19] , \REGFILE/reg_out[0][18] ,
         \REGFILE/reg_out[0][17] , \REGFILE/reg_out[0][16] ,
         \REGFILE/reg_out[0][15] , \REGFILE/reg_out[0][14] ,
         \REGFILE/reg_out[0][13] , \REGFILE/reg_out[0][12] ,
         \REGFILE/reg_out[0][11] , \REGFILE/reg_out[0][10] ,
         \REGFILE/reg_out[0][9] , \REGFILE/reg_out[0][8] ,
         \REGFILE/reg_out[0][7] , \REGFILE/reg_out[0][6] ,
         \REGFILE/reg_out[0][5] , \REGFILE/reg_out[0][4] ,
         \REGFILE/reg_out[0][3] , \REGFILE/reg_out[0][2] ,
         \REGFILE/reg_out[0][1] , \REGFILE/reg_out[0][0] ,
         \PCLOGIC/PC_REG/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \PCLOGIC/PC_REG/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ,
         \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ,
         \WIRE_ALU_A/MUX2TO1_32BIT[1].MUX/N1 ,
         \WIRE_ALU_A/MUX2TO1_32BIT[2].MUX/N1 ,
         \WIRE_ALU_A/MUX2TO1_32BIT[3].MUX/N1 ,
         \WIRE_ALU_A/MUX2TO1_32BIT[4].MUX/N1 ,
         \WIRE_ALU_A/MUX2TO1_32BIT[5].MUX/N1 ,
         \WIRE_ALU_A/MUX2TO1_32BIT[6].MUX/N1 ,
         \WIRE_ALU_A/MUX2TO1_32BIT[7].MUX/N1 ,
         \WIRE_ALU_A/MUX2TO1_32BIT[8].MUX/N1 ,
         \WIRE_ALU_A/MUX2TO1_32BIT[9].MUX/N1 ,
         \WIRE_ALU_A/MUX2TO1_32BIT[10].MUX/N1 ,
         \WIRE_ALU_A/MUX2TO1_32BIT[11].MUX/N1 ,
         \WIRE_ALU_A/MUX2TO1_32BIT[12].MUX/N1 ,
         \WIRE_ALU_A/MUX2TO1_32BIT[13].MUX/N1 ,
         \WIRE_ALU_A/MUX2TO1_32BIT[14].MUX/N1 ,
         \WIRE_ALU_A/MUX2TO1_32BIT[15].MUX/N1 , net36391, net36463, net36466,
         net36470, net36479, net36488, net70506, net70507, net70509, net70529,
         net70531, net70534, net70535, net70537, net70541, net70574, net70684,
         net70685, net70687, net70696, net70697, net70701, net70703, net70706,
         net70709, net70710, net70713, net70714, net70717, net70718, net70719,
         net70720, net70727, net70731, net70734, net70735, net70737, net70738,
         net70740, net70750, net70752, net70755, net70757, net70758, net70761,
         net70780, net70811, net70821, net70826, net70837, net70838, net70845,
         net70866, net70868, net70921, net71026, net71027, net71078, net71085,
         net71092, net71094, net71271, net71273, net71277, net71280, net71299,
         net71300, net71394, net71396, net71824, net71906, net71934, net71936,
         net72163, net72312, net72876, net72947, net72962, net73166, net73167,
         net73170, net73394, net73395, net73400, net73416, net73421, net73423,
         net73429, net73434, net73436, net73439, net73443, net73468, net73494,
         net73495, net73496, net73498, net73499, net73503, net73504, net73509,
         net73510, net73512, net73519, net73527, net73529, net73532, net73541,
         net73543, net73608, net73611, net73612, net73613, net73615, net73616,
         net73619, net73620, net73622, net73629, net73630, net73637, net73638,
         net73646, net73652, net73653, net73670, net73684, net73694, net73695,
         net73696, net73697, net73708, net73771, net73778, net73780, net73831,
         net73836, net73837, net73838, net73842, net73848, net73850, net73851,
         net73855, net73858, net73877, net73878, net73879, net73900, net73902,
         net73908, net73938, net73974, net73987, net73988, net73997, net74009,
         net74011, net74051, net74359, net74361, net74799, net74808, net75367,
         net75368, net75397, net75401, net75418, net75419, net75424, net75425,
         net75427, net75437, net75438, net75439, net75440, net75441, net75442,
         net75443, net75451, net75452, net75453, net75454, net75455, net75456,
         net75464, net75466, net75468, net75469, net75475, net75478, net75479,
         net75481, net75482, net75615, net75619, net75620, net75624, net75748,
         net75759, net75761, net75764, net75791, net75792, net75793, net75843,
         net75844, net75847, net75849, net75857, net75859, net75861, net75995,
         net76025, net76031, net76032, net76034, net76154, net76195, net76199,
         net76201, net76202, net76203, net76204, net76205, net76208, net76209,
         net76211, net76217, net76220, net76222, net76234, net76238, net76239,
         net76241, net76242, net76248, net76249, net76255, net76257, net76258,
         net76259, net76260, net76261, net76278, net76274, net76270, net76320,
         net76318, net76452, net76468, net76464, net76480, net76488, net76508,
         net76506, net76502, net76514, net76510, net76550, net76548, net76616,
         net76614, net76650, net76646, net76660, net76658, net76694, net76692,
         net76702, net76708, net76706, net76716, net76866, net76864, net76862,
         net77030, net77042, net77040, net77038, net77086, net77084, net77106,
         net77104, net77102, net77100, net77116, net77114, net77276, net77272,
         net77292, net77290, net77324, net77320, net77318, net77316, net77314,
         net77312, net77310, net77308, net77306, net77304, net77302, net77300,
         net77298, net77328, net77360, net77358, net77348, net77346, net77344,
         net77342, net77338, net77336, net77396, net77394, net77392, net77388,
         net77386, net77384, net77382, net77380, net77376, net77400, net77432,
         net77430, net77428, net77426, net77424, net77422, net77420, net77418,
         net77416, net77414, net77410, net77406, net77440, net77436, net77464,
         net77462, net77460, net77458, net77456, net77454, net77452, net77444,
         net77474, net77506, net77504, net77502, net77500, net77498, net77496,
         net77494, net77492, net77490, net77488, net77484, net77482, net77480,
         net77478, net77508, net77542, net77540, net77538, net77532, net77530,
         net77528, net77526, net77524, net77522, net77520, net77518, net77516,
         net77514, net77548, net77544, net77576, net77574, net77568, net77566,
         net77564, net77562, net77560, net77558, net77556, net77554, net77550,
         net77588, net77608, net77602, net77616, net77614, net77610, net77624,
         net77620, net77618, net77632, net77630, net77626, net77640, net77638,
         net77634, net77656, net77652, net77650, net77670, net77668, net77666,
         net77676, net77704, net77702, net77700, net77698, net77720, net77716,
         net77714, net77744, net77750, net77748, net77746, net77764, net77762,
         net77776, net77774, net77784, net77780, net77778, net77800, net77798,
         net77796, net77794, net77814, net77812, net77810, net77832, net77828,
         net77826, net77836, net77834, net77848, net77846, net77844, net77842,
         net77856, net77854, net77852, net77850, net77999, net78003, net78014,
         net78042, net78051, net78056, net78055, net78109, net78108, net78107,
         net78128, net78127, net78235, net80189, net80208, net80211, net80390,
         net80440, net80443, net81764, net81810, net82342, net82500, net82499,
         net82515, net82613, net82631, net82739, net83168, net83167, net83203,
         net83260, net84475, net84518, net84663, net84754, net84761, net85047,
         net85371, net86238, net86304, net86794, net86793, net87098, net87489,
         net87506, net87633, net88131, net88253, net89184, net90830, net90864,
         net91311, net91561, net91646, net92392, net92447, net93763, net105361,
         net105360, net105352, net105349, net87820, net85731, net76219,
         net75626, net75625, net75617, net72015, net87495, net76252, net76196,
         net76194, net75621, net75618, net75616, net83210, net82738, net81164,
         net80797, net76256, net76224, net76206, net75623, net120684,
         net121496, net121580, net123282, net123932, net124970, net77296,
         net82513, net78126, net77512, net77326, net75417, net75416, net75414,
         net74050, net73849, net123931, net76181, net75396, net75395, net74029,
         net78050, net77280, net73665, net70693, net36414, net105376,
         net105318, net87097, net78105, net75422, net75415, net70732, net70730,
         net70729, net70692, net70690, net70689, net70497, net78104, net75423,
         net73989, net89734, net88102, net87806, net82932, net77816, net76253,
         net75477, net148091, net148116, net148736, net148735, net83261,
         net72414, net91643, net76262, net73533, net77752, net76254, net76235,
         net75763, net75760, net75747, net75465, net73528, net122022, net73585,
         net92782, net81874, net81873, net70691, net70504, net70503, net70502,
         net73500, net71302, net71269, net71266, net73465, net73427, net71227,
         net71228, net75842, net81974, net76251, net76233, net75862, net73511,
         net83408, net82618, net82598, net81601, net77768, net76237, net76236,
         net76198, net75860, net75858, net75845, net75467, net148494,
         net123382, net92446, net87982, net87981, net84760, net84277, net82933,
         net80161, net76197, net75846, n10943, n4797, n4798, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4849, n4850, n4851, n4852, n4853, n4854,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5576,
         n5577, n5578, n5579, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5748, n5749, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5982, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10953, n11001;
  wire   [16:31] aluA;
  wire   [0:31] multOut;
  wire   [6:15] \PCLOGIC/imm26_32 ;
  wire   [16:31] \PCLOGIC/imm16_32 ;
  wire   [16:31] \SELECT_CORRECT_SEGMENTS/selHalf ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31;
  assign \PCLOGIC/imm26_32  [6] = instruction[6];
  assign \PCLOGIC/imm26_32  [7] = instruction[7];
  assign \PCLOGIC/imm26_32  [8] = instruction[8];
  assign \PCLOGIC/imm26_32  [9] = instruction[9];
  assign \PCLOGIC/imm26_32  [10] = instruction[10];
  assign \PCLOGIC/imm26_32  [11] = instruction[11];
  assign \PCLOGIC/imm26_32  [12] = instruction[12];
  assign \PCLOGIC/imm26_32  [13] = instruction[13];
  assign \PCLOGIC/imm26_32  [14] = instruction[14];
  assign \PCLOGIC/imm26_32  [15] = instruction[15];
  assign \PCLOGIC/imm16_32  [16] = instruction[16];
  assign \PCLOGIC/imm16_32  [17] = instruction[17];
  assign \PCLOGIC/imm16_32  [18] = instruction[18];
  assign \PCLOGIC/imm16_32  [19] = instruction[19];
  assign \PCLOGIC/imm16_32  [20] = instruction[20];
  assign \PCLOGIC/imm16_32  [21] = instruction[21];
  assign \PCLOGIC/imm16_32  [22] = instruction[22];
  assign \PCLOGIC/imm16_32  [23] = instruction[23];
  assign \PCLOGIC/imm16_32  [24] = instruction[24];
  assign \PCLOGIC/imm16_32  [25] = instruction[25];
  assign \PCLOGIC/imm16_32  [26] = instruction[26];
  assign \PCLOGIC/imm16_32  [27] = instruction[27];
  assign \PCLOGIC/imm16_32  [28] = instruction[28];
  assign \PCLOGIC/imm16_32  [29] = instruction[29];
  assign \PCLOGIC/imm16_32  [30] = instruction[30];
  assign \PCLOGIC/imm16_32  [31] = instruction[31];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [16] = dmem_read_in[0];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [17] = dmem_read_in[1];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [18] = dmem_read_in[2];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [19] = dmem_read_in[3];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [20] = dmem_read_in[4];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [21] = dmem_read_in[5];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [22] = dmem_read_in[6];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [23] = dmem_read_in[7];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [24] = dmem_read_in[8];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [25] = dmem_read_in[9];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [26] = dmem_read_in[10];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [27] = dmem_read_in[11];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [28] = dmem_read_in[12];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [29] = dmem_read_in[13];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [30] = dmem_read_in[14];
  assign \SELECT_CORRECT_SEGMENTS/selHalf  [31] = dmem_read_in[15];
  assign dmem_dsize[0] = net76468;
  assign dmem_write_out[17] = net121580;

  OAI22_X2 U181 ( .A1(n6223), .A2(n6219), .B1(n10936), .B2(n6217), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U183 ( .A1(n6222), .A2(n6219), .B1(n4940), .B2(n6217), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U184 ( .A1(n6221), .A2(n6219), .B1(n4950), .B2(n6217), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U216 ( .A1(n6223), .A2(net76318), .B1(n4938), .B2(n6215), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U218 ( .A1(n6222), .A2(net76318), .B1(n4957), .B2(n6215), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U219 ( .A1(n6221), .A2(net76318), .B1(n4952), .B2(n6215), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U386 ( .A1(n6223), .A2(n6213), .B1(n10937), .B2(n6176), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U388 ( .A1(n6222), .A2(n6213), .B1(n10934), .B2(n6176), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U389 ( .A1(n6221), .A2(n6214), .B1(n5543), .B2(n6176), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U421 ( .A1(n6223), .A2(n6211), .B1(n10938), .B2(n6209), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U423 ( .A1(n6222), .A2(n6211), .B1(n4937), .B2(n6209), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U424 ( .A1(n6221), .A2(n6211), .B1(n4958), .B2(n6209), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U660 ( .A1(n6223), .A2(n6207), .B1(n10939), .B2(n6205), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U662 ( .A1(n6222), .A2(n6207), .B1(n10935), .B2(n6205), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U663 ( .A1(n6221), .A2(n6207), .B1(n4951), .B2(n6205), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U729 ( .A1(n6223), .A2(n6203), .B1(n5898), .B2(n6202), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U731 ( .A1(n6222), .A2(n6203), .B1(n5397), .B2(n6202), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U732 ( .A1(n6221), .A2(n6203), .B1(n5433), .B2(n6202), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U969 ( .A1(n6223), .A2(n6198), .B1(n10940), .B2(n6196), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U971 ( .A1(n6222), .A2(n6198), .B1(n4956), .B2(n6197), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U972 ( .A1(n6221), .A2(n6198), .B1(n4961), .B2(n6196), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1005 ( .A1(n6223), .A2(n6194), .B1(n10941), .B2(n6192), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1007 ( .A1(n6222), .A2(n6194), .B1(n4959), .B2(n6192), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U1008 ( .A1(n6221), .A2(n6194), .B1(n4960), .B2(n6192), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][31] ), .QN(n5948) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[31]) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][31] ), .QN(n5792) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][31] ), .QN(n5891) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][31] ), .QN(net78127) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][31] ), .QN(net78128) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][31] ), .QN(net80211) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][31] ), .QN(net80440) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][31] ), .QN(net82515) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][31] ), .QN(n5949) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][31] ), .QN(net80208) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][31] ), .QN(net78108) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][31] ), .QN(net78109) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][31] ), .QN(n6002) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][31] ), .QN(n6003) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][31] ), .QN(n5823) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][31] ), .QN(n5999) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][31] ), .QN(n5717) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][31] ), .QN(n4939) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][31] ), .QN(n5765) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][31] ), .QN(net82499) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][31] ), .QN(n5026) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][31] ), .QN(n5790) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][31] ), .QN(n4917) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][31] ), .QN(n5778) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][31] ), .QN(n5788) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][31] ), .QN(n5895) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][31] ), .QN(n5811) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][31] ), .QN(n5893) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][31] ), .QN(n5824) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][31] ), .QN(n5827) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][31] ), .QN(net78235) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][15] ), .QN(n4935) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][15] ), .QN(n4927) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][15] ), .QN(n4945) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][15] ), .QN(n4948) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][15] ), .QN(n5396) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][15] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][15] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][15] ), .QN(n5917) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][15] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][15] ), .QN(n10950) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][15] ), .QN(n4944) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][15] ), .QN(n5784) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][15] ), .QN(n5251) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][15] ), .QN(n4934) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][15] ), .QN(n4919) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][15] ), .QN(n4943) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][15] ), .QN(n5431) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][15] ), .QN(n5122) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][15] ), .QN(n4942) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][15] ), .QN(n5866) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][15] ), .QN(n4941) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][15] ), .QN(n5714) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][15] ), .QN(n5856) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][15] ), .QN(n5121) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][15] ), .QN(n5852) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][15] ), .QN(n5250) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][14] ), .QN(n4933) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][14] ), .QN(n4918) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][14] ), .QN(n4932) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][14] ), .QN(n4926) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][14] ), .QN(n5395) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][14] ), .QN(n4981) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][14] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][14] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][14] ), .QN(n5838) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][14] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][14] ), .QN(n4831) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][14] ), .QN(n5839) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][14] ), .QN(n4936) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][14] ), .QN(n5879) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][14] ), .QN(n5662) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][14] ), .QN(n4931) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][14] ), .QN(n5837) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][14] ), .QN(n4930) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][14] ), .QN(n5841) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][14] ), .QN(n5394) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][14] ), .QN(n5842) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][14] ), .QN(n4929) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][14] ), .QN(n5819) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][14] ), .QN(n5883) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][14] ), .QN(n4928) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][14] ), .QN(n5843) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][14] ), .QN(n5844) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][10] ), .QN(n5249) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][10] ), .QN(n5350) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][10] ), .QN(n5248) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][10] ), .QN(n5349) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][10] ), .QN(n5083) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][10] ), .QN(n5120) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][10] ), .QN(n5114) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][10] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][10] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][10] ), .QN(n5773) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][10] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][10] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][10] ), .QN(n5877) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][10] ), .QN(n5247) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][10] ), .QN(n5025) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][10] ), .QN(n5110) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][10] ), .QN(n5109) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][10] ), .QN(n5082) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][10] ), .QN(n5246) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][10] ), .QN(n5430) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][10] ), .QN(n4979) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][10] ), .QN(n5393) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][10] ), .QN(n5774) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][10] ), .QN(n5108) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][10] ), .QN(n5245) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][10] ), .QN(n5614) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][10] ), .QN(n5107) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][10] ), .QN(n5024) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][10] ), .QN(n5775) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][10] ), .QN(n5119) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][10] ), .QN(n5875) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][10] ), .QN(n5106) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][2] ), .QN(n4987) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][2] ), .QN(n5244) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][2] ), .QN(n5243) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][2] ), .QN(n5242) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][2] ), .QN(n4986) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][2] ), .QN(n5392) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][2] ), .QN(n5241) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][20] ), .QN(n5240) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][20] ), .QN(n5346) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][20] ), .QN(n5239) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][20] ), .QN(n5345) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][20] ), .QN(n5344) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][20] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][20] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][20] ), .QN(n5023) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][20] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][20] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][20] ), .QN(n5681) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][20] ), .QN(n5238) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][20] ), .QN(n5661) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][20] ), .QN(n5237) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][20] ), .QN(n5236) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][20] ), .QN(n5343) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][20] ), .QN(n5235) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][20] ), .QN(n5342) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][20] ), .QN(n5391) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][20] ), .QN(n5341) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][20] ), .QN(n5234) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][20] ), .QN(n5105) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][20] ), .QN(n5081) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][20] ), .QN(n5233) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][20] ), .QN(n5340) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][20] ), .QN(n5682) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][20] ), .QN(n5390) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][20] ), .QN(n5821) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][20] ), .QN(n5232) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][3] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][3] ), .QN(n5429) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][3] ), .QN(n5428) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][3] ), .QN(n5389) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][19] ), .QN(n5227) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][19] ), .QN(n5337) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][19] ), .QN(n5226) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][19] ), .QN(n5336) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][19] ), .QN(n5335) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][19] ), .QN(n5388) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][19] ), .QN(n5426) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][19] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][19] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][19] ), .QN(n5651) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][19] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][19] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][19] ), .QN(n5225) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][19] ), .QN(n4973) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][19] ), .QN(n5104) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][19] ), .QN(n5224) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][19] ), .QN(n5334) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][19] ), .QN(n5223) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][19] ), .QN(n5425) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][19] ), .QN(n5080) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][19] ), .QN(n5118) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][19] ), .QN(n5333) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][19] ), .QN(n5222) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][19] ), .QN(n5221) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][19] ), .QN(n4978) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][19] ), .QN(n5220) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][19] ), .QN(n5332) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][19] ), .QN(n5387) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][19] ), .QN(n5219) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][4] ), .QN(n5218) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][4] ), .QN(n5386) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][4] ), .QN(n5217) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][4] ), .QN(n5216) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][4] ), .QN(n5215) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][11] ), .QN(n5873) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][11] ), .QN(n5858) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][11] ), .QN(n5881) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][11] ), .QN(n5908) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][11] ), .QN(n5871) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][11] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][29] ), .QN(n5987) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][29] ), .QN(n5125) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][29] ), .QN(n4940) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][29] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][29] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][29] ), .QN(n5989) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][29] ), .QN(n5985) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][29] ), .QN(n4937) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][29] ), .QN(n5214) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][29] ), .QN(n4974) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][29] ), .QN(n5123) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][29] ), .QN(net87633) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][29] ), .QN(n5988) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][29] ), .QN(n4977) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][29] ), .QN(n5397) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][29] ), .QN(n5126) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][29] ), .QN(n5213) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][29] ), .QN(n5914) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][29] ), .QN(n5991) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][29] ), .QN(n5328) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][26] ), .QN(n5422) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][26] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][26] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][26] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][26] ), .QN(n5421) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][26] ), .QN(n5212) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][26] ), .QN(n5327) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][26] ), .QN(n5211) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][26] ), .QN(n5210) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][26] ), .QN(n5326) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][26] ), .QN(n5209) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][26] ), .QN(n5420) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][26] ), .QN(n5325) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][26] ), .QN(n5385) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][26] ), .QN(n5208) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][26] ), .QN(n5324) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][26] ), .QN(n5207) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][26] ), .QN(n5323) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][7] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][6] ), .QN(n5206) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][6] ), .QN(n5322) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][6] ), .QN(n5205) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][6] ), .QN(n5321) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][6] ), .QN(n5320) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][6] ), .QN(n5384) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][6] ), .QN(n5419) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][6] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][6] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][6] ), .QN(n5319) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][6] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][6] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][6] ), .QN(n5113) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][6] ), .QN(n5103) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][6] ), .QN(n5204) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][6] ), .QN(n5203) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][6] ), .QN(n5318) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][6] ), .QN(n5202) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][6] ), .QN(n5418) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][6] ), .QN(n5317) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][6] ), .QN(n5383) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][6] ), .QN(n5316) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][6] ), .QN(n5201) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][6] ), .QN(n5200) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][6] ), .QN(n5315) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][6] ), .QN(n5417) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][6] ), .QN(n5382) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][6] ), .QN(n5437) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][5] ), .QN(n5199) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][5] ), .QN(n5314) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][5] ), .QN(n4985) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][5] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][5] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][5] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][5] ), .QN(n5416) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][5] ), .QN(n5313) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][5] ), .QN(n5198) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][5] ), .QN(n5197) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][5] ), .QN(n5381) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][5] ), .QN(n5196) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][5] ), .QN(n5195) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][5] ), .QN(n5309) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][5] ), .QN(n5308) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][21] ), .QN(n5194) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][21] ), .QN(n5307) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][21] ), .QN(n5193) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][21] ), .QN(n5306) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][21] ), .QN(n5305) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][21] ), .QN(n5414) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][21] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][21] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][21] ), .QN(n5304) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][21] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][21] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][21] ), .QN(n5192) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][21] ), .QN(n5191) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][21] ), .QN(n5190) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][21] ), .QN(n5303) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][21] ), .QN(n5189) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][21] ), .QN(n5302) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][21] ), .QN(n5380) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][21] ), .QN(n5301) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][21] ), .QN(n5188) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][21] ), .QN(n5187) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][21] ), .QN(n5300) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][21] ), .QN(n5186) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][21] ), .QN(n5299) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][21] ), .QN(n5810) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][21] ), .QN(n5379) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][21] ), .QN(n5808) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][21] ), .QN(n5185) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[21]), .QN(n5085) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][8] ), .QN(n5102) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][8] ), .QN(n4972) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][8] ), .QN(n5101) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][8] ), .QN(n5079) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][8] ), .QN(n5686) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][8] ), .QN(n5378) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][8] ), .QN(n5028) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][8] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][8] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][8] ), .QN(n5911) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][8] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][8] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][8] ), .QN(n5978) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][8] ), .QN(n5184) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][8] ), .QN(n5183) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][8] ), .QN(n5182) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][8] ), .QN(n5298) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][8] ), .QN(n5181) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][8] ), .QN(n5413) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][8] ), .QN(n5297) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][8] ), .QN(n5377) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][8] ), .QN(n5296) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][8] ), .QN(n5180) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][8] ), .QN(n5179) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][8] ), .QN(n5910) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][8] ), .QN(n5178) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][8] ), .QN(n5295) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][8] ), .QN(n5950) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][8] ), .QN(n5376) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][8] ), .QN(n5977) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][8] ), .QN(n5127) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][13] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][13] ), .QN(n5715) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][13] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][13] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][13] ), .QN(n5816) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][13] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][13] ), .QN(n5801) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][13] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][13] ), .QN(n5835) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][13] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][13] ), .QN(n5767) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][13] ), .QN(n5937) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][13] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][13] ), .QN(n5939) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][13] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][13] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][13] ), .QN(n5799) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][13] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][13] ), .QN(n5719) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][13] ), .QN(n4850) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][13] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][13] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][13] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][13] ), .QN(n4845) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][13] ), .QN(net83260) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][13] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][13] ), .QN(n5803) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][13] ), .QN(net84518) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][13] ), .QN(n5813) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][13] ) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[13]) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[10].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[10]) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][9] ), .QN(n5177) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][9] ), .QN(n5294) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][9] ), .QN(n5176) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][9] ), .QN(n5293) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][9] ), .QN(n5292) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][9] ), .QN(n5375) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][9] ), .QN(n5112) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][9] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][9] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][9] ), .QN(n5022) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][9] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][9] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][9] ), .QN(n5412) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][9] ), .QN(n5175) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][9] ), .QN(n5021) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][9] ), .QN(n5100) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][9] ), .QN(n5174) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][9] ), .QN(n5291) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][9] ), .QN(n5173) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][9] ), .QN(n5411) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][9] ), .QN(n5290) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][9] ), .QN(n5374) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][9] ), .QN(n5289) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][9] ), .QN(n5172) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][9] ), .QN(n5171) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][9] ), .QN(n4976) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][9] ), .QN(n5170) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][9] ), .QN(n5288) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][9] ), .QN(n5653) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][9] ), .QN(n5373) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][9] ), .QN(n5616) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][9] ), .QN(n5169) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][23] ), .QN(n5168) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][23] ), .QN(n5287) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][23] ), .QN(n5286) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][23] ), .QN(n5372) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][23] ), .QN(n5410) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][23] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][23] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][23] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][23] ), .QN(n5409) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][23] ), .QN(n5167) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][23] ), .QN(n5166) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][23] ), .QN(n5285) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][23] ), .QN(n5165) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][23] ), .QN(n5408) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][23] ), .QN(n5284) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][23] ), .QN(n5371) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][23] ), .QN(n5164) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][23] ), .QN(n5283) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][23] ), .QN(n5163) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][23] ), .QN(n5282) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[23]), .QN(n5086) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[20]) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[19]), .QN(n5063) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][16] ), .QN(n5667) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][16] ), .QN(n4859) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][16] ), .QN(n5755) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][16] ), .QN(n5676) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][16] ), .QN(n5786) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][16] ), .QN(n5612) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][16] ), .QN(n5665) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][16] ), .QN(n5610) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][16] ), .QN(n5617) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][16] ), .QN(n5771) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][16] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][12] ), .QN(n5862) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][12] ), .QN(n5860) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][12] ), .QN(n5864) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][12] ), .QN(n4825) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][12] ), .QN(n5673) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][12] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][17] ), .QN(n5099) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][17] ), .QN(n5078) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][17] ), .QN(n5098) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][17] ), .QN(n5077) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][17] ), .QN(n5076) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][17] ), .QN(n5117) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][17] ), .QN(n5111) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][17] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][17] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][17] ), .QN(n5020) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][17] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][17] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][17] ), .QN(n5027) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][17] ), .QN(n5097) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][17] ), .QN(n5019) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][17] ), .QN(n5096) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][17] ), .QN(n5162) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][17] ), .QN(n5281) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][17] ), .QN(n5161) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][17] ), .QN(n5407) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][17] ), .QN(n5075) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][17] ), .QN(n5116) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][17] ), .QN(n5074) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][17] ), .QN(n5095) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][17] ), .QN(n5094) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][17] ), .QN(n5018) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][17] ), .QN(n5160) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][17] ), .QN(n5280) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][17] ), .QN(n5620) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][17] ), .QN(n5370) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][17] ), .QN(n5073) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][17] ), .QN(n5093) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][25] ), .QN(n5279) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][25] ), .QN(n5369) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][25] ), .QN(n5406) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][25] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][25] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][25] ), .QN(n5405) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][25] ), .QN(n5159) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][25] ), .QN(n5278) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][25] ), .QN(n5158) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][25] ), .QN(n5157) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][25] ), .QN(n5277) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][25] ), .QN(n5156) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][25] ), .QN(n5404) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][25] ), .QN(n5155) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][25] ), .QN(n5276) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][25] ), .QN(n5154) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][25] ), .QN(n5275) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][25] ), .QN(n5274) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][25] ), .QN(n5153) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[25]), .QN(n5087) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[22]) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][22] ), .QN(n5152) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][22] ), .QN(n5273) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][22] ), .QN(n5151) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][22] ), .QN(n5272) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][22] ), .QN(n5271) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][22] ), .QN(n5403) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][22] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][22] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][22] ), .QN(n5270) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][22] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][22] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][22] ), .QN(n5402) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][22] ), .QN(n5150) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][22] ), .QN(n5269) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][22] ), .QN(n5149) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][22] ), .QN(n5148) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][22] ), .QN(n5268) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][22] ), .QN(n5147) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][22] ), .QN(n5267) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][22] ), .QN(n5368) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][22] ), .QN(n5266) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][22] ), .QN(n5146) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][22] ), .QN(n5092) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][22] ), .QN(n5017) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][22] ), .QN(n5145) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][22] ), .QN(n5265) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][22] ), .QN(n5621) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][22] ), .QN(n5367) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][22] ), .QN(n5144) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][27] ), .QN(n5356) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][27] ), .QN(n5362) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][27] ), .QN(n5436) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][27] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][27] ), .QN(n5361) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][27] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][27] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][27] ), .QN(n5435) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][27] ), .QN(n5355) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][27] ), .QN(n5360) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][27] ), .QN(n5354) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][27] ), .QN(n5353) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][27] ), .QN(n5352) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][27] ), .QN(n5434) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][27] ), .QN(n5359) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][27] ), .QN(n5432) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][27] ), .QN(n4949) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][18] ), .QN(n5091) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][18] ), .QN(n5072) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][18] ), .QN(n5143) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][18] ), .QN(n5264) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][18] ), .QN(n5366) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][18] ), .QN(n5685) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][18] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][18] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][18] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][18] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][18] ), .QN(n5913) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][18] ), .QN(n5142) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][18] ), .QN(n5857) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][18] ), .QN(n5141) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][18] ), .QN(n5090) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][18] ), .QN(n5071) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][18] ), .QN(n5140) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][18] ), .QN(n5401) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][18] ), .QN(n5263) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][18] ), .QN(n5365) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][18] ), .QN(n5262) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][18] ), .QN(n5139) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][18] ), .QN(n5138) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][18] ), .QN(n5878) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][18] ), .QN(n5089) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][18] ), .QN(n4925) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][18] ), .QN(n4980) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][18] ), .QN(n5115) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][18] ), .QN(n5886) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][18] ), .QN(n5088) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[18]) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[17].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[17]), .QN(n5084) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][28] ), .QN(n5358) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][28] ), .QN(n4950) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][28] ), .QN(n4952) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][28] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][28] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][28] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][28] ), .QN(n5351) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][28] ), .QN(n5069) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][28] ), .QN(n4951) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][28] ), .QN(n5357) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][28] ), .QN(n5433) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][30] ), .QN(n5927) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][30] ), .QN(n5961) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][30] ), .QN(n5070) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][30] ), .QN(n4938) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][30] ), .QN(n5794) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][30] ), .QN(n5925) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][30] ), .QN(n5680) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][30] ), .QN(n5833) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][30] ), .QN(n5963) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][30] ), .QN(n5920) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][30] ), .QN(n5967) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][30] ), .QN(n5924) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][30] ), .QN(n5969) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][30] ), .QN(n5934) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][30] ), .QN(n5973) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][30] ), .QN(n5922) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][30] ), .QN(n5965) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][30] ), .QN(n5124) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][30] ), .QN(n5898) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][30] ), .QN(n5971) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][30] ), .QN(n5854) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][30] ), .QN(n5929) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][30] ), .QN(n5918) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][30] ), .QN(n5992) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][30] ), .QN(n5958) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][30] ), .QN(n5994) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][30] ), .QN(n5959) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][30] ), .QN(n5996) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][30] ), .QN(n4975) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[28]) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[26]) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][24] ), .QN(n5137) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][24] ), .QN(n5261) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][24] ), .QN(n5136) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][24] ), .QN(n5260) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][24] ), .QN(n5259) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][24] ), .QN(n5364) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][24] ), .QN(n5400) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][24] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][24] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][24] ), .QN(n5258) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][24] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][24] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][24] ), .QN(n5399) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][24] ), .QN(n5135) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][24] ), .QN(n5257) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][24] ), .QN(n5134) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][24] ), .QN(n5133) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][24] ), .QN(n5256) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][24] ), .QN(n5132) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][24] ), .QN(n5398) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][24] ), .QN(n5255) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][24] ), .QN(n5363) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][24] ), .QN(n5254) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][24] ), .QN(n5131) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][24] ), .QN(n5130) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][24] ), .QN(n4947) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][24] ), .QN(n5129) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][24] ), .QN(n4946) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][24] ), .QN(n5253) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][24] ), .QN(n5128) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[24]) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[16]) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[14]) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[9].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[9]) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[6]) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[5]) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[3]) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[1]) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][3] ), .QN(n5956) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][11] ), .QN(n5906) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][16] ), .QN(n5903) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][1] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][8] ), .QN(n5869) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][13] ), .QN(n5849) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][14] ), .QN(n5831) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .QN(n5845) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][21] ), .QN(n5807) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][14] ), .QN(n5780) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][14] ), .QN(n5776) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][4] ), .QN(n5770) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][1] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][30] ), .QN(n5671) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][5] ), .QN(n5660) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][15] ), .QN(n5656) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][13] ), .QN(net148735) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][28] ), .QN(n5569) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][28] ), .QN(n5568) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][27] ), .QN(n5567) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][27] ), .QN(n5566) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][28] ), .QN(n5565) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][24] ), .QN(n5564) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][24] ), .QN(n5563) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][27] ), .QN(n5562) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][3] ), .QN(n5559) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][26] ), .QN(n5556) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][26] ), .QN(n5555) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][5] ), .QN(n5554) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][23] ), .QN(n5553) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][25] ), .QN(n5551) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][27] ), .QN(n5550) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][27] ), .QN(n5549) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][27] ), .QN(n5548) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][28] ), .QN(n5547) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][28] ), .QN(n5546) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][28] ), .QN(n5545) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][28] ), .QN(n5544) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][28] ), .QN(n5543) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][27] ), .QN(n5542) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][3] ), .QN(n5534) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][3] ), .QN(n5533) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][3] ), .QN(n5530) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][29] ), .QN(n5523) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][29] ), .QN(n5522) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][26] ), .QN(n5521) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][26] ), .QN(n5518) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][6] ), .QN(n5517) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][5] ), .QN(n5516) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][5] ), .QN(n5515) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][23] ), .QN(n5514) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][23] ), .QN(n5513) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][25] ), .QN(n5508) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][30] ), .QN(n5507) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][20] ), .QN(n5506) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][21] ), .QN(n5505) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][22] ), .QN(n5504) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][26] ), .QN(n5503) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][23] ), .QN(n5502) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][25] ), .QN(n5501) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][20] ), .QN(n5500) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][21] ), .QN(n5499) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][22] ), .QN(n5498) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][27] ), .QN(n5497) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][27] ), .QN(n5496) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][28] ), .QN(n5495) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][28] ), .QN(n5494) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][27] ), .QN(n5493) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][28] ), .QN(n5491) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][27] ), .QN(n5490) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][27] ), .QN(n5489) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][28] ), .QN(n5488) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][28] ), .QN(n5487) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][28] ), .QN(n5486) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][28] ), .QN(n5485) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][28] ), .QN(n5484) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][3] ), .QN(n5476) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][3] ), .QN(n5475) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][3] ), .QN(n5474) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][4] ), .QN(n5468) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][4] ), .QN(n5464) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][29] ), .QN(n5463) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][29] ), .QN(n5462) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][29] ), .QN(n5461) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][29] ), .QN(n5460) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][29] ), .QN(n5459) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][29] ), .QN(n5458) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][26] ), .QN(n5457) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][26] ), .QN(n5456) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][26] ), .QN(n5455) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][26] ), .QN(n5454) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][26] ), .QN(n5453) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][26] ), .QN(n5452) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][5] ), .QN(n5451) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][23] ), .QN(n5450) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][23] ), .QN(n5449) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][23] ), .QN(n5448) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][23] ), .QN(n5447) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][23] ), .QN(n5446) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][25] ), .QN(n5445) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][25] ), .QN(n5444) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][25] ), .QN(n5443) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][25] ), .QN(n5442) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][25] ), .QN(n5441) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][30] ), .QN(n5440) );
  DFF_X1 \PCLOGIC/PC_REG/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[0]), .QN(n5439) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][5] ), .QN(n5310) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][3] ), .QN(n5231) );
  DFF_X1 \PCLOGIC/PC_REG/REG_32BIT[7].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[7]), .QN(n5059) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][28] ), .QN(n5047) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][3] ), .QN(n5046) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][3] ), .QN(n5045) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][5] ), .QN(n5044) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][5] ), .QN(n5043) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][15] ), .QN(n5038) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][20] ), .QN(n5037) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][19] ), .QN(n5036) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][19] ), .QN(n5035) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][21] ), .QN(n5034) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][4] ), .QN(n5033) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][28] ), .QN(n5032) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][18] ), .QN(n5030) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][14] ), .QN(n5029) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][29] ), .QN(n4988) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][5] ), .QN(n4984) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][22] ), .QN(n4983) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][6] ), .QN(n4982) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][28] ), .QN(n4961) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][28] ), .QN(n4960) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][29] ), .QN(n4959) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][28] ), .QN(n4958) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][29] ), .QN(n4957) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][29] ), .QN(n4956) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][27] ), .QN(n4955) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][15] ), .QN(n4954) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][31] ), .QN(n4953) );
  DFF_X1 \PCLOGIC/PC_REG/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[4]), .QN(n4924) );
  DFF_X1 \PCLOGIC/PC_REG/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[2]), .QN(n4923) );
  DFF_X1 \PCLOGIC/PC_REG/REG_32BIT[8].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[8]), .QN(n4909) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][15] ), .QN(n4902) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][1] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][15] ), .QN(n5683) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][19] ), .QN(n5031) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][15] ), .QN(n4901) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][18] ), .QN(n5785) );
  INV_X2 U4891 ( .A(net77744), .ZN(net81764) );
  INV_X2 U4893 ( .A(net88131), .ZN(n4797) );
  INV_X4 U4894 ( .A(net76242), .ZN(n5587) );
  INV_X4 U4895 ( .A(n5083), .ZN(n4798) );
  AOI22_X4 U4896 ( .A1(\REGFILE/reg_out[16][12] ), .A2(net77764), .B1(
        \REGFILE/reg_out[15][12] ), .B2(net75468), .ZN(n6650) );
  AOI22_X2 U4897 ( .A1(\REGFILE/reg_out[19][8] ), .A2(net77810), .B1(
        \REGFILE/reg_out[1][8] ), .B2(net75478), .ZN(n6733) );
  OAI21_X2 U4898 ( .B1(net76502), .B2(n10581), .A(n10580), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U4899 ( .B1(net76506), .B2(n10593), .A(n10592), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  INV_X1 U4902 ( .A(n10141), .ZN(dmem_addr_out[10]) );
  OAI211_X4 U4903 ( .C1(n10141), .C2(net76646), .A(net70740), .B(n10140), .ZN(
        n10142) );
  NAND4_X4 U4904 ( .A1(n9370), .A2(n9371), .A3(n9372), .A4(n9369), .ZN(
        dmem_addr_out[9]) );
  NAND2_X4 U4905 ( .A1(multOut[9]), .A2(net92392), .ZN(n9370) );
  OAI211_X4 U4906 ( .C1(n9377), .C2(net76646), .A(net70740), .B(n9376), .ZN(
        n9378) );
  INV_X8 U4907 ( .A(net77436), .ZN(net77430) );
  INV_X16 U4908 ( .A(net77436), .ZN(net77428) );
  INV_X8 U4909 ( .A(net77430), .ZN(net77416) );
  INV_X8 U4910 ( .A(net77430), .ZN(net77418) );
  INV_X8 U4911 ( .A(net77430), .ZN(net77420) );
  NAND4_X4 U4912 ( .A1(n6543), .A2(n6542), .A3(n6541), .A4(n6540), .ZN(n6549)
         );
  AOI22_X1 U4913 ( .A1(\REGFILE/reg_out[14][28] ), .A2(net77780), .B1(
        \REGFILE/reg_out[13][28] ), .B2(n5663), .ZN(n6304) );
  AOI22_X2 U4915 ( .A1(\REGFILE/reg_out[14][17] ), .A2(net77780), .B1(
        \REGFILE/reg_out[13][17] ), .B2(n5663), .ZN(net75859) );
  AOI22_X2 U4916 ( .A1(\REGFILE/reg_out[14][13] ), .A2(net77780), .B1(n5804), 
        .B2(n5664), .ZN(net75761) );
  INV_X16 U4918 ( .A(n9528), .ZN(n6050) );
  NAND4_X4 U4919 ( .A1(n9698), .A2(n9697), .A3(n9696), .A4(n9695), .ZN(
        dmem_addr_out[7]) );
  NAND2_X4 U4920 ( .A1(net76650), .A2(dmem_addr_out[7]), .ZN(n9702) );
  NAND3_X4 U4921 ( .A1(n9702), .A2(net70740), .A3(n9701), .ZN(n9703) );
  INV_X16 U4922 ( .A(n6058), .ZN(n4802) );
  INV_X16 U4923 ( .A(n6069), .ZN(n4803) );
  INV_X16 U4924 ( .A(n9974), .ZN(n6069) );
  AOI21_X4 U4925 ( .B1(multOut[2]), .B2(net92392), .A(n5749), .ZN(net71394) );
  MUX2_X2 U4926 ( .A(multOut[6]), .B(n9662), .S(net73585), .Z(n9668) );
  OAI211_X4 U4927 ( .C1(n9673), .C2(net76646), .A(net70740), .B(n9672), .ZN(
        n9674) );
  INV_X2 U4928 ( .A(n9673), .ZN(dmem_addr_out[6]) );
  OAI21_X2 U4931 ( .B1(n6214), .B2(n6072), .A(n10048), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U4932 ( .B1(n10534), .B2(n6072), .A(n10050), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U4933 ( .B1(n10532), .B2(n6072), .A(n10049), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X1 U4935 ( .A1(n6100), .A2(\REGFILE/reg_out[13][1] ), .ZN(n10176) );
  INV_X16 U4936 ( .A(net77752), .ZN(net77746) );
  INV_X4 U4937 ( .A(net77436), .ZN(net77432) );
  INV_X8 U4938 ( .A(net77432), .ZN(net77414) );
  INV_X16 U4939 ( .A(net77432), .ZN(net77410) );
  INV_X8 U4940 ( .A(n4830), .ZN(n4897) );
  OAI21_X2 U4941 ( .B1(dmem_write_out[1]), .B2(net75427), .A(n10945), .ZN(
        net70921) );
  INV_X2 U4942 ( .A(net70921), .ZN(net36466) );
  INV_X8 U4943 ( .A(net80161), .ZN(n5576) );
  AND2_X4 U4944 ( .A1(net76270), .A2(n10521), .ZN(n4804) );
  AND2_X4 U4945 ( .A1(net76270), .A2(n10519), .ZN(n4805) );
  AND2_X4 U4946 ( .A1(n4874), .A2(n8673), .ZN(n4806) );
  INV_X32 U4947 ( .A(\PCLOGIC/imm26_32 [11]), .ZN(net87820) );
  XOR2_X1 U4948 ( .A(n9057), .B(n10463), .Z(n4807) );
  XOR2_X1 U4949 ( .A(n5762), .B(net77040), .Z(n4808) );
  AND2_X2 U4950 ( .A1(n5712), .A2(net70696), .ZN(n4809) );
  NAND2_X4 U4951 ( .A1(n10303), .A2(net70697), .ZN(net70710) );
  NAND2_X4 U4952 ( .A1(n8985), .A2(net70697), .ZN(n9606) );
  NAND2_X4 U4953 ( .A1(n8861), .A2(net70697), .ZN(n9854) );
  NAND2_X1 U4954 ( .A1(n6005), .A2(net71026), .ZN(n10544) );
  INV_X8 U4955 ( .A(n10544), .ZN(n6082) );
  NAND2_X1 U4956 ( .A1(net71026), .A2(n10099), .ZN(net70718) );
  XOR2_X1 U4957 ( .A(n5783), .B(net77038), .Z(n4810) );
  AND2_X2 U4958 ( .A1(n10465), .A2(net78051), .ZN(n4811) );
  AND4_X4 U4959 ( .A1(n9805), .A2(n8717), .A3(n8716), .A4(n8715), .ZN(n4812)
         );
  INV_X16 U4960 ( .A(n8679), .ZN(n6022) );
  NAND2_X4 U4961 ( .A1(net76270), .A2(n8668), .ZN(n8679) );
  XOR2_X1 U4962 ( .A(n10110), .B(n10404), .Z(n4813) );
  INV_X16 U4963 ( .A(n9325), .ZN(n6039) );
  NAND2_X4 U4964 ( .A1(net76270), .A2(n9320), .ZN(n9325) );
  INV_X16 U4965 ( .A(n8961), .ZN(n6028) );
  NAND2_X4 U4966 ( .A1(net76270), .A2(n8956), .ZN(n8961) );
  INV_X16 U4967 ( .A(n9579), .ZN(n6052) );
  NAND2_X4 U4968 ( .A1(net76270), .A2(n9573), .ZN(n9579) );
  XOR2_X1 U4969 ( .A(n4856), .B(net77038), .Z(n4814) );
  INV_X8 U4970 ( .A(dmem_write_out[19]), .ZN(n6529) );
  NAND2_X4 U4971 ( .A1(net76270), .A2(n9425), .ZN(n9426) );
  AND2_X2 U4972 ( .A1(multOut[2]), .A2(net92392), .ZN(n4815) );
  NAND2_X4 U4973 ( .A1(net76270), .A2(n9867), .ZN(n9868) );
  INV_X8 U4974 ( .A(net70541), .ZN(net76514) );
  NAND2_X4 U4975 ( .A1(net76270), .A2(n9113), .ZN(n4816) );
  INV_X8 U4976 ( .A(net77464), .ZN(net77452) );
  AOI22_X1 U4977 ( .A1(\REGFILE/reg_out[11][6] ), .A2(net77746), .B1(
        \REGFILE/reg_out[12][6] ), .B2(net83168), .ZN(n6769) );
  AOI22_X2 U4978 ( .A1(\REGFILE/reg_out[11][12] ), .A2(net77748), .B1(n4826), 
        .B2(net83168), .ZN(n6649) );
  AOI22_X4 U4979 ( .A1(\REGFILE/reg_out[9][10] ), .A2(net77698), .B1(
        \REGFILE/reg_out[8][10] ), .B2(net75454), .ZN(n6700) );
  NAND2_X1 U4980 ( .A1(\REGFILE/reg_out[3][10] ), .A2(net77414), .ZN(n7830) );
  INV_X4 U4981 ( .A(n5775), .ZN(n4817) );
  NAND4_X2 U4982 ( .A1(net75623), .A2(net75624), .A3(net75625), .A4(net75626), 
        .ZN(net75617) );
  AOI22_X2 U4983 ( .A1(\REGFILE/reg_out[19][26] ), .A2(net77814), .B1(
        \REGFILE/reg_out[1][26] ), .B2(net82631), .ZN(n6345) );
  INV_X32 U4984 ( .A(net77816), .ZN(net77814) );
  INV_X8 U4985 ( .A(net77640), .ZN(net77634) );
  AOI22_X4 U4986 ( .A1(\REGFILE/reg_out[29][16] ), .A2(net77652), .B1(n5787), 
        .B2(n6911), .ZN(n6579) );
  AOI22_X4 U4987 ( .A1(\REGFILE/reg_out[29][21] ), .A2(net77652), .B1(
        \REGFILE/reg_out[28][21] ), .B2(n6911), .ZN(n6475) );
  AOI22_X4 U4988 ( .A1(\REGFILE/reg_out[9][20] ), .A2(net77700), .B1(
        \REGFILE/reg_out[8][20] ), .B2(n4829), .ZN(n6494) );
  AOI22_X2 U4989 ( .A1(\REGFILE/reg_out[16][4] ), .A2(net77764), .B1(
        \REGFILE/reg_out[15][4] ), .B2(n5579), .ZN(n6814) );
  AOI22_X2 U4990 ( .A1(\REGFILE/reg_out[24][19] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][19] ), .B2(net75438), .ZN(n6520) );
  AOI22_X2 U4991 ( .A1(\REGFILE/reg_out[24][20] ), .A2(net75437), .B1(n4836), 
        .B2(net75438), .ZN(n6496) );
  INV_X8 U4992 ( .A(net75438), .ZN(net77616) );
  AOI22_X2 U4993 ( .A1(\REGFILE/reg_out[26][14] ), .A2(net75439), .B1(n5840), 
        .B2(net89184), .ZN(n6623) );
  AOI22_X2 U4994 ( .A1(\REGFILE/reg_out[16][18] ), .A2(net75467), .B1(
        \REGFILE/reg_out[15][18] ), .B2(net75468), .ZN(n6536) );
  AOI22_X2 U4995 ( .A1(\REGFILE/reg_out[16][16] ), .A2(net87506), .B1(n5666), 
        .B2(net75468), .ZN(n6568) );
  INV_X16 U4996 ( .A(net75465), .ZN(net77752) );
  INV_X8 U4997 ( .A(net76235), .ZN(net75465) );
  INV_X32 U4998 ( .A(net77752), .ZN(net77748) );
  INV_X4 U4999 ( .A(n5913), .ZN(n4818) );
  INV_X32 U5000 ( .A(net76201), .ZN(net75439) );
  NOR2_X4 U5001 ( .A1(n6420), .A2(n6419), .ZN(n6431) );
  INV_X4 U5002 ( .A(net81601), .ZN(net83408) );
  NOR2_X4 U5003 ( .A1(n6805), .A2(n6804), .ZN(n6806) );
  INV_X16 U5004 ( .A(\PCLOGIC/imm26_32 [12]), .ZN(net73533) );
  NAND4_X4 U5005 ( .A1(n6561), .A2(n6560), .A3(n6559), .A4(n6558), .ZN(
        net75847) );
  AOI22_X4 U5006 ( .A1(\REGFILE/reg_out[26][24] ), .A2(net77618), .B1(
        \REGFILE/reg_out[27][24] ), .B2(net77630), .ZN(n6402) );
  AOI22_X2 U5007 ( .A1(\REGFILE/reg_out[24][18] ), .A2(net75437), .B1(n5684), 
        .B2(net75438), .ZN(n6544) );
  NAND2_X1 U5008 ( .A1(\REGFILE/reg_out[13][15] ), .A2(net77454), .ZN(n7593)
         );
  NAND2_X1 U5009 ( .A1(n6100), .A2(\REGFILE/reg_out[13][12] ), .ZN(n9122) );
  NAND2_X1 U5010 ( .A1(\REGFILE/reg_out[13][12] ), .A2(net77452), .ZN(n7725)
         );
  BUF_X32 U5011 ( .A(n6505), .Z(n4819) );
  INV_X16 U5012 ( .A(net84760), .ZN(net84761) );
  NAND4_X2 U5013 ( .A1(n6959), .A2(n6958), .A3(n6957), .A4(n6956), .ZN(n6965)
         );
  NAND2_X4 U5014 ( .A1(\REGFILE/reg_out[1][29] ), .A2(net77516), .ZN(n6956) );
  INV_X32 U5015 ( .A(\PCLOGIC/imm26_32 [15]), .ZN(net82739) );
  AOI22_X4 U5016 ( .A1(\REGFILE/reg_out[0][17] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][17] ), .B2(net83203), .ZN(net75862) );
  BUF_X16 U5017 ( .A(n10916), .Z(n4864) );
  AOI22_X2 U5018 ( .A1(\REGFILE/reg_out[21][14] ), .A2(net77844), .B1(
        \REGFILE/reg_out[20][14] ), .B2(net77852), .ZN(n6611) );
  NAND2_X4 U5019 ( .A1(n6526), .A2(n6527), .ZN(dmem_write_out[19]) );
  NAND3_X4 U5020 ( .A1(n4842), .A2(\PCLOGIC/imm26_32 [15]), .A3(
        \PCLOGIC/imm26_32 [13]), .ZN(n4821) );
  NAND3_X2 U5021 ( .A1(n4842), .A2(\PCLOGIC/imm26_32 [15]), .A3(
        \PCLOGIC/imm26_32 [13]), .ZN(net76261) );
  NAND2_X4 U5022 ( .A1(n5642), .A2(net77272), .ZN(n4822) );
  INV_X32 U5023 ( .A(n4822), .ZN(n4963) );
  NAND2_X4 U5024 ( .A1(net73533), .A2(\PCLOGIC/imm26_32 [11]), .ZN(n4823) );
  INV_X8 U5025 ( .A(net77768), .ZN(net77764) );
  INV_X8 U5026 ( .A(net77768), .ZN(net77762) );
  INV_X2 U5027 ( .A(n4917), .ZN(n4824) );
  INV_X2 U5028 ( .A(n4825), .ZN(n4826) );
  AOI22_X2 U5029 ( .A1(\REGFILE/reg_out[26][10] ), .A2(net75439), .B1(
        \REGFILE/reg_out[27][10] ), .B2(net89184), .ZN(n6703) );
  NOR2_X4 U5030 ( .A1(n6525), .A2(n6524), .ZN(n6526) );
  NAND2_X1 U5031 ( .A1(\REGFILE/reg_out[28][18] ), .A2(net77384), .ZN(n7449)
         );
  INV_X2 U5032 ( .A(n5026), .ZN(n4827) );
  NAND4_X2 U5033 ( .A1(n6625), .A2(n6624), .A3(n6623), .A4(n6622), .ZN(n6626)
         );
  AOI22_X2 U5034 ( .A1(\REGFILE/reg_out[30][14] ), .A2(net77638), .B1(net82613), .B2(n4838), .ZN(n6624) );
  BUF_X32 U5035 ( .A(n10914), .Z(n4828) );
  INV_X16 U5037 ( .A(net76220), .ZN(n4829) );
  INV_X8 U5038 ( .A(net76220), .ZN(net75454) );
  NAND4_X4 U5039 ( .A1(n7041), .A2(n7040), .A3(n7039), .A4(n7038), .ZN(n8451)
         );
  NAND2_X2 U5040 ( .A1(n8451), .A2(net123282), .ZN(n5657) );
  INV_X32 U5041 ( .A(net77464), .ZN(net77456) );
  INV_X8 U5042 ( .A(net76251), .ZN(net76204) );
  NOR2_X4 U5044 ( .A1(n6515), .A2(n6514), .ZN(n6527) );
  AOI22_X2 U5045 ( .A1(n5921), .A2(net77406), .B1(n5968), .B2(n6014), .ZN(
        n6943) );
  AOI22_X4 U5046 ( .A1(\REGFILE/reg_out[26][7] ), .A2(net75439), .B1(
        \REGFILE/reg_out[27][7] ), .B2(net77626), .ZN(net75621) );
  NAND2_X4 U5047 ( .A1(\REGFILE/reg_out[31][29] ), .A2(net77498), .ZN(n6990)
         );
  AOI22_X4 U5048 ( .A1(\REGFILE/reg_out[0][15] ), .A2(net82342), .B1(n5853), 
        .B2(net83203), .ZN(n6588) );
  INV_X2 U5050 ( .A(n4831), .ZN(n4832) );
  INV_X1 U5051 ( .A(net73831), .ZN(n4833) );
  INV_X4 U5052 ( .A(n4833), .ZN(n4834) );
  NAND2_X1 U5053 ( .A1(n4884), .A2(\REGFILE/reg_out[18][16] ), .ZN(n9224) );
  INV_X4 U5054 ( .A(n5784), .ZN(n4835) );
  AOI22_X2 U5055 ( .A1(\REGFILE/reg_out[24][15] ), .A2(net75437), .B1(n4835), 
        .B2(net124970), .ZN(n6598) );
  NAND2_X2 U5056 ( .A1(n8411), .A2(net77272), .ZN(n6946) );
  INV_X16 U5057 ( .A(instruction[2]), .ZN(net74029) );
  INV_X16 U5058 ( .A(\PCLOGIC/imm26_32 [14]), .ZN(n4843) );
  AOI22_X2 U5059 ( .A1(\REGFILE/reg_out[30][17] ), .A2(net84761), .B1(
        \REGFILE/reg_out[2][17] ), .B2(net82613), .ZN(n5584) );
  AOI22_X2 U5061 ( .A1(\REGFILE/reg_out[30][15] ), .A2(net77638), .B1(n4837), 
        .B2(net82613), .ZN(n6600) );
  AOI22_X2 U5062 ( .A1(\REGFILE/reg_out[30][12] ), .A2(net84761), .B1(n5863), 
        .B2(net82613), .ZN(n6660) );
  AOI22_X2 U5063 ( .A1(\REGFILE/reg_out[30][9] ), .A2(net77634), .B1(
        \REGFILE/reg_out[2][9] ), .B2(net82613), .ZN(n6726) );
  AOI22_X2 U5064 ( .A1(\REGFILE/reg_out[30][7] ), .A2(net77634), .B1(
        \REGFILE/reg_out[2][7] ), .B2(net82613), .ZN(net75620) );
  AOI22_X2 U5065 ( .A1(\REGFILE/reg_out[30][8] ), .A2(net77634), .B1(n5912), 
        .B2(net75442), .ZN(n6748) );
  INV_X16 U5067 ( .A(net75418), .ZN(net77328) );
  INV_X16 U5068 ( .A(net74050), .ZN(net77512) );
  NOR2_X2 U5069 ( .A1(net87633), .A2(net77512), .ZN(net91561) );
  INV_X1 U5070 ( .A(net75464), .ZN(net77744) );
  AOI22_X2 U5071 ( .A1(\REGFILE/reg_out[0][20] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][20] ), .B2(net83203), .ZN(n6486) );
  INV_X4 U5072 ( .A(net77550), .ZN(net77576) );
  INV_X8 U5073 ( .A(net77576), .ZN(net77554) );
  INV_X4 U5074 ( .A(n5661), .ZN(n4836) );
  NAND2_X4 U5075 ( .A1(n6731), .A2(n6730), .ZN(dmem_write_out[9]) );
  INV_X4 U5076 ( .A(n5917), .ZN(n4837) );
  NAND2_X1 U5077 ( .A1(net77406), .A2(\REGFILE/reg_out[19][27] ), .ZN(n7059)
         );
  NAND2_X1 U5078 ( .A1(net77406), .A2(\REGFILE/reg_out[27][28] ), .ZN(n7005)
         );
  NAND2_X1 U5079 ( .A1(net77406), .A2(\REGFILE/reg_out[19][28] ), .ZN(n7015)
         );
  NAND2_X1 U5080 ( .A1(net77406), .A2(\REGFILE/reg_out[3][28] ), .ZN(n7035) );
  AOI22_X2 U5081 ( .A1(n4827), .A2(net77406), .B1(n5791), .B2(n6014), .ZN(
        n6922) );
  OAI21_X2 U5082 ( .B1(n7007), .B2(n7006), .A(n6011), .ZN(n7041) );
  INV_X4 U5084 ( .A(n5838), .ZN(n4838) );
  INV_X2 U5085 ( .A(n5683), .ZN(n4839) );
  INV_X16 U5086 ( .A(net77440), .ZN(net77436) );
  INV_X2 U5087 ( .A(net75437), .ZN(net77608) );
  AOI22_X4 U5088 ( .A1(\REGFILE/reg_out[11][14] ), .A2(net77748), .B1(n5846), 
        .B2(net83167), .ZN(n6613) );
  OAI21_X2 U5089 ( .B1(net76502), .B2(n10619), .A(n10618), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  AOI22_X4 U5090 ( .A1(\REGFILE/reg_out[16][22] ), .A2(net77764), .B1(
        \REGFILE/reg_out[15][22] ), .B2(n5579), .ZN(n6440) );
  NAND2_X1 U5091 ( .A1(\REGFILE/reg_out[30][13] ), .A2(net75441), .ZN(n5941)
         );
  AOI22_X1 U5092 ( .A1(\REGFILE/reg_out[19][28] ), .A2(net77814), .B1(
        \REGFILE/reg_out[1][28] ), .B2(net82631), .ZN(n6298) );
  AOI22_X1 U5093 ( .A1(\REGFILE/reg_out[19][27] ), .A2(net77814), .B1(
        \REGFILE/reg_out[1][27] ), .B2(net82631), .ZN(n6322) );
  AOI22_X2 U5095 ( .A1(\REGFILE/reg_out[16][14] ), .A2(net75467), .B1(n5884), 
        .B2(net75468), .ZN(n6614) );
  INV_X32 U5096 ( .A(net77624), .ZN(net77620) );
  INV_X16 U5097 ( .A(net75439), .ZN(net77624) );
  INV_X32 U5098 ( .A(\PCLOGIC/imm26_32 [14]), .ZN(n4840) );
  INV_X32 U5099 ( .A(\PCLOGIC/imm26_32 [14]), .ZN(n4841) );
  INV_X32 U5100 ( .A(\PCLOGIC/imm26_32 [14]), .ZN(n4842) );
  OAI21_X1 U5101 ( .B1(dmem_write_out[0]), .B2(net75427), .A(n10945), .ZN(
        net71027) );
  OAI21_X2 U5102 ( .B1(dmem_write_out[4]), .B2(net75427), .A(n10945), .ZN(
        n10400) );
  NAND2_X1 U5103 ( .A1(\REGFILE/reg_out[6][29] ), .A2(net77550), .ZN(n6963) );
  NAND2_X1 U5104 ( .A1(\REGFILE/reg_out[22][29] ), .A2(net77550), .ZN(n6981)
         );
  AOI22_X4 U5105 ( .A1(\REGFILE/reg_out[14][15] ), .A2(net77780), .B1(
        \REGFILE/reg_out[13][15] ), .B2(n5664), .ZN(n6591) );
  INV_X16 U5106 ( .A(n6074), .ZN(n6072) );
  INV_X16 U5107 ( .A(n6074), .ZN(n6073) );
  AOI22_X1 U5108 ( .A1(\REGFILE/reg_out[26][26] ), .A2(net77620), .B1(
        \REGFILE/reg_out[27][26] ), .B2(net89184), .ZN(n6359) );
  AOI22_X2 U5109 ( .A1(\REGFILE/reg_out[26][11] ), .A2(net75439), .B1(net89184), .B2(n5859), .ZN(n6681) );
  INV_X16 U5110 ( .A(net77776), .ZN(n5579) );
  NAND3_X2 U5111 ( .A1(\PCLOGIC/imm26_32 [15]), .A2(\PCLOGIC/imm26_32 [14]), 
        .A3(\PCLOGIC/imm26_32 [13]), .ZN(n4844) );
  INV_X8 U5112 ( .A(net75440), .ZN(net77632) );
  NAND3_X4 U5113 ( .A1(net87495), .A2(n4841), .A3(\PCLOGIC/imm26_32 [15]), 
        .ZN(net76252) );
  INV_X8 U5114 ( .A(net76252), .ZN(net76196) );
  AOI22_X2 U5115 ( .A1(\REGFILE/reg_out[24][5] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][5] ), .B2(net77610), .ZN(n6800) );
  AOI22_X2 U5116 ( .A1(\REGFILE/reg_out[24][29] ), .A2(net77602), .B1(
        \REGFILE/reg_out[25][29] ), .B2(net77610), .ZN(n6287) );
  AOI22_X2 U5117 ( .A1(n5935), .A2(net77478), .B1(n5974), .B2(net77550), .ZN(
        n6937) );
  OAI21_X4 U5118 ( .B1(n6964), .B2(n6965), .A(net73838), .ZN(n6997) );
  NAND4_X4 U5119 ( .A1(n6963), .A2(n6962), .A3(n6961), .A4(n6960), .ZN(n6964)
         );
  NAND2_X1 U5120 ( .A1(n4805), .A2(\REGFILE/reg_out[14][13] ), .ZN(n9437) );
  NAND2_X1 U5121 ( .A1(\REGFILE/reg_out[14][13] ), .A2(net77560), .ZN(n7684)
         );
  INV_X2 U5122 ( .A(n4845), .ZN(n4846) );
  NAND2_X1 U5123 ( .A1(n4875), .A2(\REGFILE/reg_out[24][13] ), .ZN(n9459) );
  NAND2_X1 U5124 ( .A1(\REGFILE/reg_out[24][13] ), .A2(net77308), .ZN(n7665)
         );
  INV_X1 U5125 ( .A(n4819), .ZN(dmem_write_out[20]) );
  OR2_X4 U5126 ( .A1(n10040), .A2(n10039), .ZN(dmem_addr_out[3]) );
  OAI22_X2 U5127 ( .A1(n10038), .A2(net70691), .B1(n10037), .B2(n5752), .ZN(
        n10039) );
  INV_X32 U5128 ( .A(instruction[1]), .ZN(net73496) );
  INV_X4 U5129 ( .A(net77550), .ZN(net77574) );
  INV_X8 U5130 ( .A(net77574), .ZN(net77564) );
  INV_X8 U5131 ( .A(net77574), .ZN(net77562) );
  INV_X8 U5132 ( .A(net77574), .ZN(net77560) );
  INV_X8 U5133 ( .A(net77574), .ZN(net77568) );
  INV_X8 U5134 ( .A(net77576), .ZN(net77566) );
  INV_X8 U5135 ( .A(net77576), .ZN(net77556) );
  INV_X8 U5136 ( .A(net77576), .ZN(net77558) );
  NAND4_X4 U5137 ( .A1(n6630), .A2(n6631), .A3(n6633), .A4(n6632), .ZN(
        net75759) );
  AOI22_X2 U5138 ( .A1(\REGFILE/reg_out[19][21] ), .A2(net77812), .B1(
        \REGFILE/reg_out[1][21] ), .B2(net75478), .ZN(n6459) );
  INV_X4 U5139 ( .A(n5680), .ZN(n4849) );
  AOI22_X2 U5140 ( .A1(\REGFILE/reg_out[3][30] ), .A2(net77406), .B1(n4849), 
        .B2(n6014), .ZN(n6939) );
  AND2_X2 U5141 ( .A1(n5654), .A2(n5655), .ZN(n6941) );
  INV_X2 U5142 ( .A(n4850), .ZN(n4851) );
  NAND2_X2 U5143 ( .A1(n10207), .A2(n10206), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  INV_X8 U5144 ( .A(n9835), .ZN(n10915) );
  INV_X16 U5145 ( .A(n5697), .ZN(net75456) );
  AOI22_X2 U5146 ( .A1(\REGFILE/reg_out[7][3] ), .A2(net75455), .B1(
        \REGFILE/reg_out[6][3] ), .B2(net75456), .ZN(n6843) );
  OAI21_X1 U5147 ( .B1(n6553), .B2(net78056), .A(n6552), .ZN(n4852) );
  INV_X8 U5148 ( .A(dmem_write_out[18]), .ZN(n6553) );
  AOI22_X2 U5149 ( .A1(\REGFILE/reg_out[24][14] ), .A2(net75437), .B1(n5880), 
        .B2(net124970), .ZN(n6622) );
  INV_X4 U5150 ( .A(n5843), .ZN(n4853) );
  AOI22_X4 U5151 ( .A1(\REGFILE/reg_out[11][13] ), .A2(net77748), .B1(n5608), 
        .B2(net83167), .ZN(net75763) );
  INV_X4 U5152 ( .A(n5915), .ZN(n5916) );
  NOR2_X2 U5153 ( .A1(n6501), .A2(n6500), .ZN(n6502) );
  INV_X4 U5154 ( .A(n5856), .ZN(n4854) );
  NAND2_X2 U5155 ( .A1(net77100), .A2(n4990), .ZN(n10171) );
  NAND2_X2 U5156 ( .A1(net77104), .A2(n4806), .ZN(n10207) );
  NAND2_X2 U5157 ( .A1(n10203), .A2(n10202), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U5158 ( .A1(n10197), .A2(n10196), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U5159 ( .A1(n10205), .A2(n10204), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U5160 ( .A1(n10191), .A2(n10190), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U5161 ( .A1(n10185), .A2(n10184), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U5162 ( .A1(n10169), .A2(n10168), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U5163 ( .A1(n10219), .A2(n10218), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U5164 ( .A1(n10221), .A2(n10220), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U5165 ( .A1(n10187), .A2(n10186), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U5166 ( .A1(n10171), .A2(n10170), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  INV_X8 U5167 ( .A(n5578), .ZN(net77454) );
  INV_X16 U5169 ( .A(net75467), .ZN(net77768) );
  INV_X16 U5170 ( .A(net77768), .ZN(net87506) );
  INV_X8 U5172 ( .A(net123382), .ZN(net76198) );
  NAND2_X1 U5173 ( .A1(n6175), .A2(\REGFILE/reg_out[28][15] ), .ZN(n10299) );
  NAND2_X1 U5174 ( .A1(net77382), .A2(\REGFILE/reg_out[28][15] ), .ZN(n7579)
         );
  NAND2_X2 U5176 ( .A1(net73851), .A2(n4963), .ZN(net75396) );
  OAI22_X4 U5177 ( .A1(net82515), .A2(n5648), .B1(net80208), .B2(net85371), 
        .ZN(net82513) );
  AOI22_X4 U5178 ( .A1(\REGFILE/reg_out[19][13] ), .A2(net77812), .B1(n4851), 
        .B2(net75478), .ZN(n6631) );
  AOI22_X2 U5179 ( .A1(\REGFILE/reg_out[16][17] ), .A2(net75467), .B1(
        \REGFILE/reg_out[15][17] ), .B2(net75468), .ZN(net75860) );
  NAND2_X4 U5180 ( .A1(net76238), .A2(n5607), .ZN(net76253) );
  AOI22_X2 U5181 ( .A1(\REGFILE/reg_out[0][10] ), .A2(net120684), .B1(n5876), 
        .B2(net83203), .ZN(n6692) );
  INV_X8 U5182 ( .A(net76194), .ZN(net75438) );
  INV_X8 U5183 ( .A(net77616), .ZN(net77610) );
  AOI22_X2 U5184 ( .A1(\REGFILE/reg_out[24][2] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][2] ), .B2(net77610), .ZN(n6866) );
  NOR2_X2 U5186 ( .A1(n6339), .A2(n6340), .ZN(n6341) );
  INV_X8 U5187 ( .A(n6000), .ZN(n6010) );
  INV_X16 U5188 ( .A(n6010), .ZN(n5664) );
  NAND4_X4 U5189 ( .A1(n6969), .A2(n6968), .A3(n6967), .A4(n6966), .ZN(n6975)
         );
  OAI21_X2 U5190 ( .B1(n6982), .B2(n6983), .A(net77588), .ZN(n6995) );
  AOI22_X2 U5191 ( .A1(\REGFILE/reg_out[16][5] ), .A2(net87506), .B1(
        \REGFILE/reg_out[15][5] ), .B2(net77774), .ZN(n6792) );
  NOR2_X2 U5192 ( .A1(n6795), .A2(n6794), .ZN(n6807) );
  INV_X4 U5193 ( .A(n5845), .ZN(n5846) );
  INV_X4 U5194 ( .A(n5996), .ZN(n5997) );
  INV_X2 U5195 ( .A(n9306), .ZN(n4856) );
  AOI22_X4 U5196 ( .A1(\REGFILE/reg_out[19][17] ), .A2(net77812), .B1(
        \REGFILE/reg_out[1][17] ), .B2(net75478), .ZN(n6555) );
  AOI22_X2 U5197 ( .A1(\REGFILE/reg_out[24][26] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][26] ), .B2(net77614), .ZN(n6358) );
  INV_X32 U5198 ( .A(\PCLOGIC/imm26_32 [14]), .ZN(net86793) );
  INV_X1 U5199 ( .A(n6994), .ZN(n4857) );
  INV_X4 U5200 ( .A(n4857), .ZN(n4858) );
  INV_X8 U5201 ( .A(n10288), .ZN(n5851) );
  INV_X2 U5202 ( .A(n4859), .ZN(n4860) );
  AOI22_X4 U5203 ( .A1(n5919), .A2(net77474), .B1(n5995), .B2(net77400), .ZN(
        n6948) );
  INV_X4 U5204 ( .A(n5994), .ZN(n5995) );
  INV_X4 U5205 ( .A(n8408), .ZN(n6952) );
  NAND2_X4 U5206 ( .A1(n5607), .A2(net122022), .ZN(net76235) );
  INV_X16 U5207 ( .A(n5689), .ZN(n5696) );
  NOR2_X4 U5208 ( .A1(n9963), .A2(n9962), .ZN(n9967) );
  OR2_X1 U5209 ( .A1(n5991), .A2(net75424), .ZN(n6971) );
  INV_X16 U5210 ( .A(net75424), .ZN(net77550) );
  OAI21_X2 U5211 ( .B1(n10532), .B2(net77114), .A(n10119), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  NOR2_X4 U5212 ( .A1(n6363), .A2(n6362), .ZN(n6364) );
  OAI21_X2 U5213 ( .B1(net70509), .B2(net77116), .A(n5690), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  INV_X8 U5214 ( .A(net86304), .ZN(net77506) );
  NAND2_X4 U5215 ( .A1(multOut[3]), .A2(n4861), .ZN(n4862) );
  NAND2_X4 U5216 ( .A1(n10032), .A2(net73585), .ZN(n4863) );
  NAND2_X4 U5217 ( .A1(n4862), .A2(n4863), .ZN(n10040) );
  INV_X4 U5218 ( .A(net73585), .ZN(n4861) );
  AOI22_X2 U5219 ( .A1(\REGFILE/reg_out[19][19] ), .A2(net77812), .B1(
        \REGFILE/reg_out[1][19] ), .B2(net75478), .ZN(n6507) );
  AOI22_X4 U5220 ( .A1(\REGFILE/reg_out[19][16] ), .A2(net77812), .B1(
        \REGFILE/reg_out[1][16] ), .B2(net75478), .ZN(n6563) );
  INV_X8 U5221 ( .A(net75478), .ZN(n5624) );
  AOI22_X1 U5222 ( .A1(\REGFILE/reg_out[16][0] ), .A2(net87506), .B1(
        \REGFILE/reg_out[15][0] ), .B2(net77774), .ZN(n6903) );
  AOI22_X1 U5223 ( .A1(\REGFILE/reg_out[16][2] ), .A2(net75467), .B1(
        \REGFILE/reg_out[15][2] ), .B2(net77774), .ZN(n6858) );
  AOI22_X1 U5224 ( .A1(\REGFILE/reg_out[16][27] ), .A2(net75467), .B1(
        \REGFILE/reg_out[15][27] ), .B2(net77774), .ZN(n6327) );
  AOI22_X1 U5225 ( .A1(\REGFILE/reg_out[16][29] ), .A2(net77762), .B1(
        \REGFILE/reg_out[15][29] ), .B2(net77774), .ZN(n6279) );
  AOI22_X1 U5226 ( .A1(\REGFILE/reg_out[16][26] ), .A2(net87506), .B1(
        \REGFILE/reg_out[15][26] ), .B2(n5579), .ZN(n6350) );
  AOI22_X1 U5227 ( .A1(\REGFILE/reg_out[16][3] ), .A2(net77764), .B1(
        \REGFILE/reg_out[15][3] ), .B2(n5579), .ZN(n6836) );
  INV_X4 U5228 ( .A(net88131), .ZN(net122022) );
  AOI22_X2 U5229 ( .A1(\REGFILE/reg_out[24][6] ), .A2(net75437), .B1(n5764), 
        .B2(net124970), .ZN(n6778) );
  AOI22_X4 U5230 ( .A1(\REGFILE/reg_out[19][24] ), .A2(net77814), .B1(
        \REGFILE/reg_out[1][24] ), .B2(net82631), .ZN(n5622) );
  NAND4_X4 U5231 ( .A1(net76031), .A2(net76032), .A3(n5622), .A4(net76034), 
        .ZN(net76025) );
  NOR2_X4 U5232 ( .A1(instruction[2]), .A2(instruction[4]), .ZN(n4865) );
  INV_X32 U5233 ( .A(net77392), .ZN(net77386) );
  NAND2_X2 U5234 ( .A1(\REGFILE/reg_out[5][29] ), .A2(net77444), .ZN(n6960) );
  INV_X16 U5235 ( .A(n5588), .ZN(net83203) );
  AOI22_X2 U5236 ( .A1(\REGFILE/reg_out[11][18] ), .A2(net77748), .B1(
        \REGFILE/reg_out[12][18] ), .B2(net83167), .ZN(n6535) );
  CLKBUF_X3 U5237 ( .A(net77272), .Z(n4866) );
  INV_X16 U5238 ( .A(net77464), .ZN(net77444) );
  INV_X16 U5239 ( .A(net77464), .ZN(net77458) );
  INV_X8 U5240 ( .A(net77272), .ZN(net77276) );
  NAND2_X1 U5241 ( .A1(\REGFILE/reg_out[25][26] ), .A2(net77514), .ZN(n7088)
         );
  NAND2_X1 U5242 ( .A1(\REGFILE/reg_out[17][26] ), .A2(net77514), .ZN(n7098)
         );
  NAND2_X1 U5243 ( .A1(\REGFILE/reg_out[9][26] ), .A2(net77514), .ZN(n7108) );
  NAND2_X1 U5244 ( .A1(\REGFILE/reg_out[1][26] ), .A2(net77514), .ZN(n7118) );
  NAND2_X1 U5245 ( .A1(net77514), .A2(\REGFILE/reg_out[17][27] ), .ZN(n7054)
         );
  NAND2_X1 U5246 ( .A1(net77514), .A2(\REGFILE/reg_out[25][28] ), .ZN(n7000)
         );
  NAND2_X1 U5247 ( .A1(net77514), .A2(\REGFILE/reg_out[17][28] ), .ZN(n7010)
         );
  AOI22_X2 U5248 ( .A1(n4824), .A2(net77514), .B1(n5779), .B2(net77298), .ZN(
        n6921) );
  INV_X4 U5249 ( .A(net77514), .ZN(net86238) );
  AOI22_X2 U5250 ( .A1(n5818), .A2(net77514), .B1(n5970), .B2(net77298), .ZN(
        n6942) );
  AOI22_X2 U5251 ( .A1(n5855), .A2(net77514), .B1(n5930), .B2(net77298), .ZN(
        n6934) );
  AOI22_X2 U5252 ( .A1(n5928), .A2(net77514), .B1(n5962), .B2(net77298), .ZN(
        n6950) );
  NAND2_X2 U5253 ( .A1(\REGFILE/reg_out[17][29] ), .A2(net77514), .ZN(n6976)
         );
  INV_X4 U5254 ( .A(net77320), .ZN(net77314) );
  INV_X4 U5255 ( .A(net77320), .ZN(net77316) );
  AOI22_X2 U5256 ( .A1(\REGFILE/reg_out[14][11] ), .A2(net77780), .B1(
        \REGFILE/reg_out[13][11] ), .B2(n5664), .ZN(n6673) );
  AOI22_X2 U5257 ( .A1(\REGFILE/reg_out[14][10] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][10] ), .B2(n5664), .ZN(n6695) );
  NAND2_X4 U5258 ( .A1(n9968), .A2(net76270), .ZN(n9974) );
  AOI22_X2 U5259 ( .A1(\REGFILE/reg_out[24][25] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][25] ), .B2(net77610), .ZN(n6382) );
  NAND2_X1 U5260 ( .A1(net77474), .A2(\REGFILE/reg_out[5][28] ), .ZN(n7028) );
  AOI22_X2 U5261 ( .A1(n5834), .A2(net77474), .B1(n5964), .B2(net77400), .ZN(
        n6944) );
  NOR2_X4 U5262 ( .A1(n10040), .A2(n10039), .ZN(n10045) );
  OAI21_X2 U5263 ( .B1(n6993), .B2(n6992), .A(n8411), .ZN(n6994) );
  NAND4_X4 U5264 ( .A1(n6987), .A2(n6986), .A3(n6985), .A4(n6984), .ZN(n6993)
         );
  NOR2_X2 U5265 ( .A1(n6491), .A2(n6490), .ZN(n6503) );
  AOI22_X2 U5266 ( .A1(\REGFILE/reg_out[24][10] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][10] ), .B2(net75438), .ZN(n6702) );
  AOI22_X2 U5267 ( .A1(\REGFILE/reg_out[24][9] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][9] ), .B2(net124970), .ZN(n6724) );
  INV_X16 U5268 ( .A(net76237), .ZN(net75467) );
  NAND4_X4 U5269 ( .A1(n6557), .A2(n6556), .A3(n6555), .A4(n6554), .ZN(
        net75857) );
  AOI22_X4 U5270 ( .A1(\REGFILE/reg_out[23][17] ), .A2(net77828), .B1(
        \REGFILE/reg_out[22][17] ), .B2(net77836), .ZN(n6556) );
  INV_X32 U5271 ( .A(net77816), .ZN(net77812) );
  INV_X32 U5272 ( .A(\PCLOGIC/imm26_32 [15]), .ZN(net73511) );
  NAND2_X4 U5273 ( .A1(multOut[0]), .A2(net105376), .ZN(net105318) );
  INV_X16 U5274 ( .A(n5588), .ZN(net75464) );
  NAND4_X4 U5275 ( .A1(net75849), .A2(n5584), .A3(n5586), .A4(n5585), .ZN(
        n5583) );
  NAND2_X1 U5276 ( .A1(net75844), .A2(\PCLOGIC/imm16_32 [30]), .ZN(n5639) );
  INV_X8 U5277 ( .A(n5645), .ZN(net77440) );
  OAI21_X2 U5278 ( .B1(n10367), .B2(n10366), .A(n10365), .ZN(n10370) );
  INV_X8 U5279 ( .A(n5646), .ZN(n5645) );
  INV_X16 U5280 ( .A(net77394), .ZN(net77384) );
  INV_X16 U5281 ( .A(net77394), .ZN(net77380) );
  INV_X4 U5282 ( .A(n10944), .ZN(n6505) );
  NAND3_X1 U5283 ( .A1(n8564), .A2(instruction[5]), .A3(net73496), .ZN(n8542)
         );
  INV_X16 U5284 ( .A(n6920), .ZN(n6014) );
  INV_X16 U5285 ( .A(net85371), .ZN(net77336) );
  NOR3_X1 U5286 ( .A1(n8438), .A2(n8437), .A3(n8436), .ZN(n8439) );
  NOR2_X1 U5287 ( .A1(net70868), .A2(net71273), .ZN(n8614) );
  OAI21_X2 U5288 ( .B1(n9033), .B2(n9032), .A(n9031), .ZN(n9053) );
  OAI21_X2 U5289 ( .B1(n9833), .B2(n9356), .A(n9355), .ZN(n10131) );
  AOI21_X2 U5290 ( .B1(net73638), .B2(net73646), .A(n8568), .ZN(n8569) );
  INV_X4 U5292 ( .A(n10385), .ZN(n10912) );
  NOR3_X2 U5293 ( .A1(n8559), .A2(instruction[2]), .A3(instruction[0]), .ZN(
        n8553) );
  INV_X4 U5294 ( .A(dmem_write_out[22]), .ZN(n6457) );
  OAI21_X2 U5295 ( .B1(n8270), .B2(n8269), .A(net77290), .ZN(n8271) );
  INV_X16 U5296 ( .A(net77360), .ZN(net77338) );
  OAI21_X1 U5297 ( .B1(n7214), .B2(n7213), .A(net77588), .ZN(n7215) );
  OAI21_X2 U5298 ( .B1(n7139), .B2(n7138), .A(n6011), .ZN(n7173) );
  OAI21_X1 U5299 ( .B1(n7259), .B2(n7258), .A(net77588), .ZN(n7260) );
  OAI21_X1 U5300 ( .B1(n7349), .B2(n7348), .A(net77588), .ZN(n7350) );
  INV_X8 U5301 ( .A(net75479), .ZN(net77832) );
  INV_X4 U5302 ( .A(net76257), .ZN(net75479) );
  INV_X8 U5303 ( .A(net75469), .ZN(net77784) );
  INV_X4 U5304 ( .A(net76241), .ZN(net75469) );
  OAI21_X1 U5305 ( .B1(net36488), .B2(net70535), .A(net70838), .ZN(net70837)
         );
  NOR2_X1 U5306 ( .A1(net70868), .A2(n10404), .ZN(n8611) );
  NOR2_X2 U5307 ( .A1(n8624), .A2(n8623), .ZN(n8625) );
  NOR2_X1 U5308 ( .A1(net70868), .A2(n9954), .ZN(n8623) );
  OAI21_X2 U5309 ( .B1(n8818), .B2(n10054), .A(n8817), .ZN(n9993) );
  NOR2_X1 U5310 ( .A1(net70868), .A2(n10109), .ZN(n8620) );
  OAI21_X2 U5311 ( .B1(n9511), .B2(n9510), .A(n9509), .ZN(n9611) );
  OAI21_X2 U5312 ( .B1(n9581), .B2(net71273), .A(n9580), .ZN(n10091) );
  OAI21_X2 U5313 ( .B1(net70535), .B2(n9581), .A(n9580), .ZN(net70727) );
  OAI21_X2 U5314 ( .B1(n7125), .B2(n7124), .A(net77290), .ZN(n7126) );
  OAI21_X2 U5315 ( .B1(n7428), .B2(n7427), .A(n6019), .ZN(n7440) );
  NOR3_X1 U5316 ( .A1(n8418), .A2(n8417), .A3(n8416), .ZN(n8429) );
  NOR3_X1 U5317 ( .A1(n8425), .A2(n8424), .A3(n8423), .ZN(n8426) );
  NOR2_X1 U5318 ( .A1(n8422), .A2(n8421), .ZN(n8427) );
  NOR2_X1 U5319 ( .A1(n8431), .A2(n8430), .ZN(n8442) );
  NOR2_X1 U5320 ( .A1(n8433), .A2(n8432), .ZN(n8441) );
  NOR2_X1 U5321 ( .A1(n8435), .A2(n8434), .ZN(n8440) );
  NOR2_X1 U5322 ( .A1(n10494), .A2(net73541), .ZN(n8580) );
  AOI222_X1 U5323 ( .A1(n6083), .A2(n8976), .B1(n8728), .B2(n10466), .C1(
        n10465), .C2(net71026), .ZN(n9801) );
  AOI222_X1 U5324 ( .A1(n6083), .A2(n8928), .B1(n8891), .B2(n8759), .C1(n8758), 
        .C2(net71026), .ZN(n9804) );
  NAND3_X2 U5325 ( .A1(n8853), .A2(n8852), .A3(n8851), .ZN(n9011) );
  INV_X4 U5326 ( .A(n5065), .ZN(net78003) );
  OAI21_X2 U5327 ( .B1(net70731), .B2(net70732), .A(n5627), .ZN(net70730) );
  OAI21_X2 U5328 ( .B1(instructionAddr_out[28]), .B2(instructionAddr_out[29]), 
        .A(n8337), .ZN(n8331) );
  OAI21_X1 U5329 ( .B1(n7452), .B2(n7451), .A(n6012), .ZN(n7486) );
  OAI21_X1 U5330 ( .B1(n7462), .B2(n7461), .A(net77588), .ZN(n7485) );
  OAI21_X1 U5331 ( .B1(n7482), .B2(n7481), .A(net77292), .ZN(n7483) );
  OAI21_X1 U5332 ( .B1(n7680), .B2(n7679), .A(net77588), .ZN(n7703) );
  OAI21_X1 U5333 ( .B1(n7670), .B2(n7669), .A(n6012), .ZN(n7704) );
  OAI21_X1 U5334 ( .B1(n7700), .B2(n7699), .A(net77292), .ZN(n7701) );
  AOI21_X2 U5335 ( .B1(n9531), .B2(net77030), .A(n9517), .ZN(n9518) );
  AOI21_X2 U5336 ( .B1(n9634), .B2(net77030), .A(n9633), .ZN(n9635) );
  AOI21_X1 U5337 ( .B1(n9671), .B2(net77030), .A(n9670), .ZN(n9672) );
  AOI21_X1 U5338 ( .B1(n9965), .B2(net77030), .A(n9964), .ZN(n9966) );
  AOI21_X1 U5339 ( .B1(n10043), .B2(net77030), .A(n10042), .ZN(n10044) );
  AOI21_X1 U5340 ( .B1(net71396), .B2(net77030), .A(n5693), .ZN(n5692) );
  AOI21_X1 U5341 ( .B1(n10139), .B2(net77030), .A(n10138), .ZN(n10140) );
  NAND3_X2 U5342 ( .A1(\SELECT_CORRECT_SEGMENTS/selHalf [16]), .A2(n4899), 
        .A3(net73170), .ZN(net70740) );
  NOR2_X2 U5343 ( .A1(n8592), .A2(net70691), .ZN(n8780) );
  OAI21_X2 U5344 ( .B1(n4909), .B2(n8379), .A(n5059), .ZN(n8297) );
  NOR2_X1 U5345 ( .A1(n10430), .A2(n10429), .ZN(n10440) );
  INV_X8 U5346 ( .A(net77336), .ZN(net77358) );
  INV_X4 U5347 ( .A(dmem_write_out[21]), .ZN(n6481) );
  NAND4_X2 U5348 ( .A1(n6950), .A2(n6949), .A3(n6948), .A4(n6947), .ZN(n8408)
         );
  NAND3_X2 U5349 ( .A1(n6930), .A2(net75401), .A3(n6931), .ZN(n5915) );
  NOR3_X2 U5350 ( .A1(n10308), .A2(n10307), .A3(n10394), .ZN(n10455) );
  NAND3_X1 U5351 ( .A1(n8564), .A2(net73496), .A3(net73503), .ZN(n8551) );
  NAND3_X2 U5352 ( .A1(n8553), .A2(net73498), .A3(net73503), .ZN(n8554) );
  NOR2_X2 U5353 ( .A1(\PCLOGIC/imm16_32 [31]), .A2(n8563), .ZN(n8552) );
  NAND3_X2 U5354 ( .A1(net73684), .A2(\PCLOGIC/imm16_32 [28]), .A3(n5605), 
        .ZN(net73695) );
  AOI21_X1 U5355 ( .B1(n8545), .B2(net73646), .A(n5252), .ZN(n8546) );
  NAND3_X1 U5356 ( .A1(n9066), .A2(n9093), .A3(n8850), .ZN(n9978) );
  OAI21_X2 U5357 ( .B1(n9683), .B2(n9614), .A(n9613), .ZN(n9663) );
  OAI21_X2 U5358 ( .B1(n7920), .B2(n7919), .A(net77290), .ZN(n7921) );
  OAI21_X2 U5359 ( .B1(n7962), .B2(n7961), .A(net77290), .ZN(n7963) );
  OAI21_X2 U5360 ( .B1(n8240), .B2(n8239), .A(n6011), .ZN(n8274) );
  OAI21_X2 U5361 ( .B1(n8260), .B2(n8259), .A(n6019), .ZN(n8272) );
  OAI21_X2 U5362 ( .B1(n8250), .B2(n8249), .A(net77588), .ZN(n8273) );
  OAI21_X2 U5363 ( .B1(n7876), .B2(n7875), .A(net77290), .ZN(n7877) );
  OAI21_X1 U5364 ( .B1(n7724), .B2(n7723), .A(net77588), .ZN(n7747) );
  OAI21_X1 U5365 ( .B1(n7714), .B2(n7713), .A(n6012), .ZN(n7748) );
  OAI21_X1 U5366 ( .B1(n7734), .B2(n7733), .A(n6019), .ZN(n7746) );
  OAI21_X1 U5367 ( .B1(n7184), .B2(n7183), .A(n6011), .ZN(n7218) );
  OAI21_X1 U5368 ( .B1(n7194), .B2(n7193), .A(net77290), .ZN(n7217) );
  OAI21_X1 U5369 ( .B1(n7204), .B2(n7203), .A(n6019), .ZN(n7216) );
  NAND4_X2 U5370 ( .A1(n6991), .A2(n6990), .A3(n6989), .A4(n6988), .ZN(n6992)
         );
  NAND4_X2 U5371 ( .A1(n6934), .A2(n6937), .A3(n6936), .A4(n6935), .ZN(
        net73831) );
  AOI22_X2 U5372 ( .A1(\REGFILE/reg_out[5][30] ), .A2(net77454), .B1(
        \REGFILE/reg_out[4][30] ), .B2(net77386), .ZN(n6940) );
  OAI21_X1 U5373 ( .B1(n7149), .B2(n7148), .A(net77290), .ZN(n7172) );
  OAI21_X1 U5374 ( .B1(n7159), .B2(n7158), .A(n6019), .ZN(n7171) );
  OAI21_X1 U5375 ( .B1(n7169), .B2(n7168), .A(net77588), .ZN(n7170) );
  NOR2_X2 U5376 ( .A1(net77999), .A2(n9373), .ZN(n8997) );
  NOR2_X2 U5377 ( .A1(net70811), .A2(n5597), .ZN(net72947) );
  AOI21_X1 U5378 ( .B1(n9000), .B2(net77030), .A(n8999), .ZN(n9001) );
  NOR2_X2 U5379 ( .A1(net76464), .A2(n8998), .ZN(n8999) );
  OAI21_X1 U5380 ( .B1(n7229), .B2(n7228), .A(n6012), .ZN(n7263) );
  OAI21_X1 U5381 ( .B1(n7239), .B2(n7238), .A(net77292), .ZN(n7262) );
  OAI21_X1 U5382 ( .B1(n7249), .B2(n7248), .A(n6019), .ZN(n7261) );
  OAI21_X1 U5383 ( .B1(n7822), .B2(n7821), .A(n6019), .ZN(n7834) );
  NOR2_X1 U5384 ( .A1(n8420), .A2(n8419), .ZN(n8428) );
  OAI21_X1 U5385 ( .B1(n7319), .B2(n7318), .A(n6012), .ZN(n7353) );
  OAI21_X1 U5386 ( .B1(n7329), .B2(n7328), .A(net77292), .ZN(n7352) );
  OAI21_X1 U5387 ( .B1(n7339), .B2(n7338), .A(n6019), .ZN(n7351) );
  OAI21_X2 U5388 ( .B1(n9393), .B2(n9062), .A(n9061), .ZN(n9353) );
  INV_X16 U5389 ( .A(net70718), .ZN(net77084) );
  NAND3_X2 U5390 ( .A1(n9584), .A2(n9583), .A3(n9582), .ZN(n9934) );
  AOI21_X2 U5391 ( .B1(n8728), .B2(n10013), .A(n5015), .ZN(n9582) );
  NOR2_X2 U5392 ( .A1(n10152), .A2(n9606), .ZN(n10105) );
  OAI21_X2 U5393 ( .B1(n8152), .B2(n8151), .A(n6011), .ZN(n8186) );
  OAI21_X2 U5394 ( .B1(n8162), .B2(n8161), .A(net77588), .ZN(n8185) );
  OAI21_X2 U5395 ( .B1(n8172), .B2(n8171), .A(n6019), .ZN(n8184) );
  OAI21_X2 U5396 ( .B1(n8064), .B2(n8063), .A(n6011), .ZN(n8098) );
  OAI21_X2 U5397 ( .B1(n8074), .B2(n8073), .A(net77588), .ZN(n8097) );
  OAI21_X2 U5398 ( .B1(n8084), .B2(n8083), .A(n6019), .ZN(n8096) );
  OAI21_X2 U5399 ( .B1(n8196), .B2(n8195), .A(n6011), .ZN(n8230) );
  OAI21_X2 U5400 ( .B1(n8216), .B2(n8215), .A(n6019), .ZN(n8228) );
  OAI21_X2 U5401 ( .B1(n8226), .B2(n8225), .A(net77290), .ZN(n8227) );
  OAI21_X2 U5402 ( .B1(n8108), .B2(n8107), .A(n6011), .ZN(n8142) );
  OAI21_X2 U5403 ( .B1(n8118), .B2(n8117), .A(net77588), .ZN(n8141) );
  OAI21_X1 U5404 ( .B1(n8128), .B2(n8127), .A(n6019), .ZN(n8140) );
  OAI21_X2 U5405 ( .B1(n8020), .B2(n8019), .A(n6011), .ZN(n8054) );
  OAI21_X1 U5406 ( .B1(n8030), .B2(n8029), .A(net77588), .ZN(n8053) );
  OAI21_X2 U5407 ( .B1(n8040), .B2(n8039), .A(n6019), .ZN(n8052) );
  OAI21_X2 U5408 ( .B1(n7976), .B2(n7975), .A(n6011), .ZN(n8010) );
  OAI21_X2 U5409 ( .B1(n7986), .B2(n7985), .A(net77588), .ZN(n8009) );
  OAI21_X2 U5410 ( .B1(n7996), .B2(n7995), .A(n6019), .ZN(n8008) );
  OAI21_X1 U5411 ( .B1(n7626), .B2(n7625), .A(n6012), .ZN(n7660) );
  OAI21_X1 U5412 ( .B1(n7636), .B2(n7635), .A(net77588), .ZN(n7659) );
  OAI21_X1 U5413 ( .B1(n7656), .B2(n7655), .A(net77292), .ZN(n7657) );
  OAI21_X1 U5414 ( .B1(n7582), .B2(n7581), .A(n6012), .ZN(n7616) );
  OAI21_X1 U5415 ( .B1(n7592), .B2(n7591), .A(net77588), .ZN(n7615) );
  OAI21_X1 U5416 ( .B1(n7612), .B2(n7611), .A(net77292), .ZN(n7613) );
  OAI21_X1 U5417 ( .B1(n7548), .B2(n7547), .A(net77588), .ZN(n7571) );
  OAI21_X1 U5418 ( .B1(n7558), .B2(n7557), .A(n6019), .ZN(n7570) );
  OAI21_X1 U5419 ( .B1(n7768), .B2(n7767), .A(net77588), .ZN(n7791) );
  OAI21_X1 U5420 ( .B1(n7758), .B2(n7757), .A(n6011), .ZN(n7792) );
  OAI21_X1 U5421 ( .B1(n7788), .B2(n7787), .A(net77290), .ZN(n7789) );
  NOR2_X2 U5422 ( .A1(n8661), .A2(n8660), .ZN(n8666) );
  OAI21_X2 U5423 ( .B1(n7095), .B2(n7094), .A(n6011), .ZN(n7129) );
  OAI21_X2 U5424 ( .B1(n7105), .B2(n7104), .A(net77588), .ZN(n7128) );
  OAI21_X2 U5425 ( .B1(n7115), .B2(n7114), .A(n6019), .ZN(n7127) );
  NAND4_X2 U5426 ( .A1(n7085), .A2(n7084), .A3(n7083), .A4(n7082), .ZN(n8450)
         );
  OAI21_X1 U5427 ( .B1(n7496), .B2(n7495), .A(n6012), .ZN(n7528) );
  OAI21_X1 U5428 ( .B1(n7506), .B2(n7505), .A(net77588), .ZN(n7527) );
  OAI21_X1 U5429 ( .B1(n7515), .B2(n7514), .A(n6019), .ZN(n7526) );
  NOR2_X2 U5430 ( .A1(n10000), .A2(n8949), .ZN(n8954) );
  OAI21_X2 U5431 ( .B1(n7274), .B2(n7273), .A(n6012), .ZN(n7308) );
  OAI21_X1 U5432 ( .B1(n7284), .B2(n7283), .A(net77292), .ZN(n7307) );
  OAI21_X1 U5433 ( .B1(n7294), .B2(n7293), .A(n6019), .ZN(n7306) );
  NOR2_X2 U5434 ( .A1(net77999), .A2(n5597), .ZN(net72876) );
  AOI21_X1 U5435 ( .B1(n9041), .B2(net77030), .A(n9040), .ZN(n9042) );
  NOR2_X2 U5436 ( .A1(net76464), .A2(n9039), .ZN(n9040) );
  AOI21_X2 U5437 ( .B1(\SELECT_CORRECT_SEGMENTS/selHalf [16]), .B2(n4911), .A(
        n10000), .ZN(n9204) );
  AOI222_X2 U5438 ( .A1(net76650), .A2(dmem_addr_out[16]), .B1(
        dmem_read_in[16]), .B2(net76468), .C1(n9203), .C2(net77030), .ZN(n9205) );
  OAI21_X2 U5439 ( .B1(n7408), .B2(n7407), .A(n6012), .ZN(n7442) );
  OAI21_X2 U5440 ( .B1(n7418), .B2(n7417), .A(net77588), .ZN(n7441) );
  OAI21_X2 U5441 ( .B1(n7438), .B2(n7437), .A(net77292), .ZN(n7439) );
  OAI21_X1 U5442 ( .B1(n7364), .B2(n7363), .A(n6012), .ZN(n7398) );
  OAI21_X1 U5443 ( .B1(n7374), .B2(n7373), .A(net77588), .ZN(n7397) );
  OAI21_X1 U5444 ( .B1(n7384), .B2(n7383), .A(n6019), .ZN(n7396) );
  NOR2_X2 U5445 ( .A1(n10000), .A2(n9313), .ZN(n9318) );
  AOI21_X2 U5446 ( .B1(n9375), .B2(net77030), .A(n9374), .ZN(n9376) );
  NOR2_X2 U5447 ( .A1(n10000), .A2(n9566), .ZN(n9571) );
  INV_X8 U5448 ( .A(n9800), .ZN(n6064) );
  NOR2_X2 U5449 ( .A1(n9788), .A2(net71906), .ZN(n9793) );
  INV_X16 U5450 ( .A(n10090), .ZN(n6077) );
  NOR2_X2 U5451 ( .A1(n10504), .A2(net76464), .ZN(n10293) );
  NAND3_X2 U5452 ( .A1(n4907), .A2(net73429), .A3(net73443), .ZN(n8677) );
  NAND4_X2 U5453 ( .A1(n6488), .A2(n6489), .A3(n6487), .A4(n6486), .ZN(n6490)
         );
  AOI22_X2 U5454 ( .A1(\REGFILE/reg_out[7][8] ), .A2(net77716), .B1(
        \REGFILE/reg_out[6][8] ), .B2(net75456), .ZN(n6745) );
  AOI22_X2 U5455 ( .A1(\REGFILE/reg_out[26][6] ), .A2(net77618), .B1(
        \REGFILE/reg_out[27][6] ), .B2(net77626), .ZN(n6779) );
  NOR3_X1 U5456 ( .A1(n8729), .A2(net71026), .A3(net78003), .ZN(n8730) );
  NOR2_X1 U5457 ( .A1(n4812), .A2(n9854), .ZN(n8718) );
  NOR3_X1 U5458 ( .A1(net78003), .A2(n10099), .A3(n10312), .ZN(n9806) );
  NOR2_X1 U5459 ( .A1(n10442), .A2(net78014), .ZN(n9811) );
  OAI21_X1 U5460 ( .B1(n9804), .B2(n10472), .A(n8764), .ZN(n8770) );
  NOR2_X1 U5461 ( .A1(n8601), .A2(net78014), .ZN(n8602) );
  NOR2_X1 U5462 ( .A1(n10336), .A2(net78014), .ZN(n9291) );
  NOR3_X1 U5463 ( .A1(n9306), .A2(n10334), .A3(net78003), .ZN(n9307) );
  NOR2_X1 U5464 ( .A1(n8921), .A2(net78014), .ZN(n8922) );
  NOR3_X1 U5465 ( .A1(n10338), .A2(n8967), .A3(net78003), .ZN(n8943) );
  NOR2_X1 U5466 ( .A1(n10343), .A2(net78014), .ZN(n9544) );
  NOR2_X1 U5467 ( .A1(n8833), .A2(net70710), .ZN(n8834) );
  AOI21_X2 U5468 ( .B1(n8863), .B2(n8862), .A(net72163), .ZN(n8864) );
  OAI21_X2 U5469 ( .B1(n8848), .B2(n9606), .A(n8847), .ZN(n8866) );
  OAI21_X2 U5470 ( .B1(n9414), .B2(n9854), .A(n9413), .ZN(n9415) );
  NOR2_X1 U5471 ( .A1(net70710), .A2(n9366), .ZN(n9367) );
  NOR2_X2 U5472 ( .A1(n9606), .A2(n9348), .ZN(n9350) );
  NOR2_X1 U5473 ( .A1(n10418), .A2(net78014), .ZN(n9349) );
  NOR2_X1 U5474 ( .A1(net70710), .A2(n9626), .ZN(n9627) );
  INV_X4 U5475 ( .A(net70691), .ZN(net71271) );
  NOR2_X2 U5476 ( .A1(n9606), .A2(n9605), .ZN(n9608) );
  NOR3_X1 U5477 ( .A1(net73630), .A2(n5605), .A3(net73532), .ZN(n5602) );
  NOR2_X1 U5478 ( .A1(n5604), .A2(net73629), .ZN(n5603) );
  NAND3_X2 U5479 ( .A1(net105361), .A2(n5637), .A3(n5636), .ZN(net105376) );
  AOI21_X2 U5480 ( .B1(n5710), .B2(net70701), .A(n4809), .ZN(net105361) );
  NOR2_X2 U5481 ( .A1(n10000), .A2(net73166), .ZN(n8875) );
  AOI21_X2 U5482 ( .B1(n8873), .B2(net77030), .A(n8872), .ZN(n8874) );
  NOR2_X2 U5483 ( .A1(n10000), .A2(n9999), .ZN(n10005) );
  AOI21_X1 U5484 ( .B1(n10003), .B2(net77030), .A(n10002), .ZN(n10004) );
  NOR2_X2 U5485 ( .A1(n5592), .A2(net70531), .ZN(net70529) );
  OAI21_X2 U5486 ( .B1(n8479), .B2(n8480), .A(n8395), .ZN(n8473) );
  OAI21_X2 U5487 ( .B1(n8493), .B2(n8494), .A(n8386), .ZN(n8487) );
  OAI21_X1 U5488 ( .B1(n4908), .B2(n8308), .A(n5060), .ZN(n8304) );
  OAI21_X2 U5489 ( .B1(n9107), .B2(n8372), .A(n8523), .ZN(n8373) );
  NOR2_X2 U5490 ( .A1(n8739), .A2(n8738), .ZN(n8740) );
  NOR2_X2 U5491 ( .A1(n8785), .A2(n8784), .ZN(n8790) );
  INV_X4 U5492 ( .A(n5002), .ZN(n6172) );
  OAI21_X2 U5493 ( .B1(n8502), .B2(n8503), .A(n8366), .ZN(n9388) );
  INV_X4 U5494 ( .A(n4992), .ZN(net76660) );
  INV_X4 U5495 ( .A(n4994), .ZN(n6158) );
  INV_X4 U5496 ( .A(n4999), .ZN(n6160) );
  INV_X4 U5497 ( .A(n5000), .ZN(n6162) );
  INV_X4 U5498 ( .A(n4997), .ZN(net76616) );
  INV_X4 U5499 ( .A(n4903), .ZN(n6208) );
  INV_X4 U5500 ( .A(n4904), .ZN(n6164) );
  INV_X4 U5501 ( .A(n4905), .ZN(n6166) );
  INV_X4 U5502 ( .A(n4906), .ZN(n6168) );
  INV_X4 U5503 ( .A(n4995), .ZN(n6170) );
  INV_X4 U5504 ( .A(n5003), .ZN(n6174) );
  INV_X4 U5505 ( .A(n5005), .ZN(net76550) );
  INV_X4 U5506 ( .A(n4996), .ZN(n6220) );
  INV_X4 U5507 ( .A(n5006), .ZN(n6183) );
  INV_X4 U5508 ( .A(n5007), .ZN(n6185) );
  INV_X4 U5509 ( .A(n4991), .ZN(n6187) );
  INV_X4 U5510 ( .A(n5008), .ZN(n6189) );
  INV_X4 U5511 ( .A(n4993), .ZN(n6199) );
  INV_X4 U5512 ( .A(n4998), .ZN(n6195) );
  INV_X4 U5513 ( .A(n5001), .ZN(n6204) );
  INV_X4 U5514 ( .A(n5004), .ZN(n6212) );
  INV_X4 U5515 ( .A(n5009), .ZN(net76320) );
  AOI21_X1 U5516 ( .B1(n9700), .B2(net77030), .A(n9699), .ZN(n9701) );
  NOR2_X2 U5517 ( .A1(n9819), .A2(n9818), .ZN(n9824) );
  INV_X4 U5518 ( .A(n4992), .ZN(net76658) );
  INV_X4 U5519 ( .A(n4990), .ZN(n6155) );
  INV_X4 U5520 ( .A(n4998), .ZN(n6194) );
  INV_X4 U5521 ( .A(n4993), .ZN(n6198) );
  INV_X4 U5522 ( .A(n4994), .ZN(n6157) );
  INV_X4 U5523 ( .A(n4999), .ZN(n6159) );
  INV_X4 U5524 ( .A(n5000), .ZN(n6161) );
  INV_X4 U5525 ( .A(n5001), .ZN(n6203) );
  INV_X4 U5526 ( .A(n4997), .ZN(net76614) );
  INV_X4 U5527 ( .A(n4903), .ZN(n6207) );
  INV_X4 U5528 ( .A(n4904), .ZN(n6163) );
  INV_X4 U5529 ( .A(n4905), .ZN(n6165) );
  INV_X4 U5530 ( .A(n4906), .ZN(n6167) );
  INV_X4 U5531 ( .A(n4995), .ZN(n6169) );
  INV_X4 U5532 ( .A(n5002), .ZN(n6171) );
  INV_X4 U5533 ( .A(n5003), .ZN(n6173) );
  INV_X4 U5534 ( .A(n5004), .ZN(n6211) );
  INV_X4 U5535 ( .A(n4806), .ZN(n6214) );
  INV_X4 U5536 ( .A(n5005), .ZN(net76548) );
  INV_X4 U5537 ( .A(n5009), .ZN(net76318) );
  INV_X4 U5538 ( .A(n4996), .ZN(n6219) );
  INV_X4 U5539 ( .A(n5006), .ZN(n6182) );
  INV_X4 U5540 ( .A(n5007), .ZN(n6184) );
  INV_X4 U5541 ( .A(n4991), .ZN(n6186) );
  INV_X4 U5542 ( .A(n5008), .ZN(n6188) );
  NAND2_X2 U5543 ( .A1(n6829), .A2(n6828), .ZN(dmem_write_out[4]) );
  NOR2_X1 U5544 ( .A1(n6005), .A2(n10312), .ZN(n10313) );
  NAND3_X2 U5545 ( .A1(net73509), .A2(\PCLOGIC/imm16_32 [26]), .A3(net73696), 
        .ZN(net73620) );
  INV_X4 U5546 ( .A(net77336), .ZN(net77360) );
  NAND3_X2 U5547 ( .A1(n10440), .A2(n10439), .A3(n10438), .ZN(n10451) );
  NAND3_X2 U5548 ( .A1(n8637), .A2(n9499), .A3(n8627), .ZN(n8892) );
  NOR2_X1 U5549 ( .A1(n8655), .A2(n8565), .ZN(n8566) );
  NAND3_X2 U5550 ( .A1(n8576), .A2(net73498), .A3(net73503), .ZN(n8535) );
  OAI21_X1 U5551 ( .B1(n7744), .B2(n7743), .A(net77292), .ZN(n7745) );
  NAND4_X2 U5552 ( .A1(n7011), .A2(n7010), .A3(n7009), .A4(n7008), .ZN(n7017)
         );
  NOR2_X1 U5553 ( .A1(instruction[2]), .A2(net73499), .ZN(net73504) );
  NAND4_X2 U5554 ( .A1(net75859), .A2(net75861), .A3(net75862), .A4(net75860), 
        .ZN(net75858) );
  OAI21_X1 U5555 ( .B1(net70868), .B2(n10247), .A(n9076), .ZN(n8708) );
  NOR2_X1 U5556 ( .A1(net70866), .A2(n9656), .ZN(n8709) );
  NAND3_X2 U5557 ( .A1(n9343), .A2(n8724), .A3(n8723), .ZN(n8978) );
  OAI21_X2 U5558 ( .B1(n6005), .B2(n8936), .A(n8935), .ZN(n9302) );
  NAND3_X1 U5559 ( .A1(n9070), .A2(n9069), .A3(n9068), .ZN(n9838) );
  NAND3_X1 U5560 ( .A1(n9341), .A2(n9340), .A3(n9339), .ZN(n9839) );
  OAI21_X2 U5561 ( .B1(n8576), .B2(net73637), .A(instruction[5]), .ZN(n8577)
         );
  OAI21_X2 U5562 ( .B1(net73638), .B2(net73616), .A(\PCLOGIC/imm16_32 [31]), 
        .ZN(n8578) );
  OAI21_X2 U5563 ( .B1(n9959), .B2(n9958), .A(n9957), .ZN(n10035) );
  NOR2_X1 U5564 ( .A1(n10093), .A2(n9606), .ZN(n10029) );
  NOR2_X2 U5565 ( .A1(n9941), .A2(n9940), .ZN(n9942) );
  OAI21_X2 U5566 ( .B1(n8182), .B2(n8181), .A(net77290), .ZN(n8183) );
  OAI21_X1 U5567 ( .B1(n8094), .B2(n8093), .A(net77290), .ZN(n8095) );
  OAI21_X2 U5568 ( .B1(n8206), .B2(n8205), .A(net77588), .ZN(n8229) );
  OAI21_X2 U5569 ( .B1(n8138), .B2(n8137), .A(net77290), .ZN(n8139) );
  OAI21_X2 U5570 ( .B1(n8050), .B2(n8049), .A(net77290), .ZN(n8051) );
  OAI21_X2 U5571 ( .B1(n8006), .B2(n8005), .A(net77290), .ZN(n8007) );
  OAI21_X1 U5572 ( .B1(n7646), .B2(n7645), .A(n6019), .ZN(n7658) );
  OAI21_X1 U5573 ( .B1(n7602), .B2(n7601), .A(n6019), .ZN(n7614) );
  OAI21_X1 U5574 ( .B1(n7568), .B2(n7567), .A(net77292), .ZN(n7569) );
  OAI21_X1 U5575 ( .B1(n7778), .B2(n7777), .A(n6019), .ZN(n7790) );
  NOR2_X2 U5576 ( .A1(net77999), .A2(n9516), .ZN(n8661) );
  NOR2_X2 U5577 ( .A1(net70811), .A2(n10540), .ZN(n8660) );
  AOI21_X2 U5578 ( .B1(n8664), .B2(net77030), .A(n8663), .ZN(n8665) );
  NOR2_X2 U5579 ( .A1(net76464), .A2(n8662), .ZN(n8663) );
  OAI21_X1 U5580 ( .B1(n7524), .B2(n7523), .A(net77292), .ZN(n7525) );
  OAI21_X1 U5581 ( .B1(n7472), .B2(n7471), .A(n6019), .ZN(n7484) );
  NOR2_X2 U5582 ( .A1(net77999), .A2(n9669), .ZN(n8949) );
  AOI21_X2 U5583 ( .B1(n8964), .B2(net77030), .A(n8952), .ZN(n8953) );
  NOR2_X2 U5584 ( .A1(net76464), .A2(n8951), .ZN(n8952) );
  OAI21_X1 U5585 ( .B1(n7304), .B2(n7303), .A(net77588), .ZN(n7305) );
  NOR2_X2 U5586 ( .A1(net76464), .A2(n9108), .ZN(n9109) );
  OAI21_X1 U5587 ( .B1(n7394), .B2(n7393), .A(net77292), .ZN(n7395) );
  NOR2_X2 U5588 ( .A1(net77999), .A2(n10505), .ZN(n9313) );
  AOI21_X1 U5589 ( .B1(n9316), .B2(net77030), .A(n9315), .ZN(n9317) );
  NOR2_X2 U5590 ( .A1(net76464), .A2(n9314), .ZN(n9315) );
  NOR2_X2 U5591 ( .A1(net76464), .A2(n9373), .ZN(n9374) );
  OAI21_X1 U5592 ( .B1(n7690), .B2(n7689), .A(n6019), .ZN(n7702) );
  AOI21_X2 U5593 ( .B1(n9422), .B2(net77030), .A(n9421), .ZN(n9423) );
  NOR2_X2 U5594 ( .A1(net76464), .A2(n9816), .ZN(n9421) );
  NOR2_X2 U5595 ( .A1(net76464), .A2(n9516), .ZN(n9517) );
  NOR2_X2 U5596 ( .A1(net77999), .A2(n9817), .ZN(n9566) );
  AOI21_X1 U5597 ( .B1(n9569), .B2(net77030), .A(n9568), .ZN(n9570) );
  NOR2_X2 U5598 ( .A1(net76464), .A2(n9567), .ZN(n9568) );
  NOR2_X2 U5599 ( .A1(net76464), .A2(n9817), .ZN(n9633) );
  NOR2_X2 U5600 ( .A1(net76464), .A2(n9669), .ZN(n9670) );
  NOR2_X2 U5601 ( .A1(net77999), .A2(n10137), .ZN(n9788) );
  NOR2_X2 U5602 ( .A1(net70811), .A2(n5694), .ZN(net71906) );
  AOI21_X1 U5603 ( .B1(n9791), .B2(net77030), .A(n9790), .ZN(n9792) );
  NOR2_X2 U5604 ( .A1(net76464), .A2(n9789), .ZN(n9790) );
  AOI21_X1 U5605 ( .B1(n9864), .B2(net77030), .A(n9863), .ZN(n9865) );
  NOR2_X2 U5606 ( .A1(net76464), .A2(n9862), .ZN(n9863) );
  NOR2_X2 U5607 ( .A1(net76464), .A2(n10083), .ZN(n9964) );
  NOR2_X2 U5608 ( .A1(net76464), .A2(n10041), .ZN(n10042) );
  NOR2_X2 U5609 ( .A1(net76464), .A2(n5694), .ZN(n5693) );
  NOR2_X2 U5610 ( .A1(net76464), .A2(n10137), .ZN(n10138) );
  NOR2_X1 U5611 ( .A1(n10484), .A2(net77040), .ZN(n10458) );
  AOI21_X2 U5612 ( .B1(n10495), .B2(n10494), .A(n10493), .ZN(n10496) );
  NOR2_X1 U5613 ( .A1(n10494), .A2(net77040), .ZN(n10492) );
  AOI21_X1 U5614 ( .B1(n10484), .B2(net77042), .A(n10494), .ZN(n10488) );
  NOR2_X2 U5615 ( .A1(n8575), .A2(n8581), .ZN(n8556) );
  NAND3_X2 U5616 ( .A1(n8619), .A2(n8618), .A3(n8617), .ZN(n9294) );
  NAND3_X2 U5617 ( .A1(n9981), .A2(n9980), .A3(n9979), .ZN(n10057) );
  NAND3_X2 U5618 ( .A1(n9551), .A2(n9550), .A3(n9549), .ZN(n10059) );
  AOI21_X1 U5619 ( .B1(net71085), .B2(n9182), .A(n9023), .ZN(n9024) );
  AOI21_X1 U5620 ( .B1(net71085), .B2(n10282), .A(n5058), .ZN(n10283) );
  AOI21_X2 U5621 ( .B1(net71085), .B2(n10248), .A(n5057), .ZN(n10249) );
  NAND3_X1 U5622 ( .A1(n9067), .A2(n9066), .A3(n10462), .ZN(n10239) );
  OAI21_X2 U5623 ( .B1(n9094), .B2(n10327), .A(n9017), .ZN(n10238) );
  OAI21_X2 U5624 ( .B1(n9094), .B2(net72312), .A(n9082), .ZN(n9395) );
  AOI21_X1 U5625 ( .B1(net71085), .B2(n10126), .A(n5056), .ZN(n10127) );
  AOI21_X2 U5626 ( .B1(net71085), .B2(n9685), .A(n5051), .ZN(n9503) );
  NAND3_X1 U5627 ( .A1(n9361), .A2(n9360), .A3(n9359), .ZN(n9945) );
  NAND3_X1 U5628 ( .A1(n9078), .A2(n9077), .A3(n9076), .ZN(n9500) );
  NAND3_X2 U5629 ( .A1(n9588), .A2(n9587), .A3(n9586), .ZN(n9655) );
  AOI21_X1 U5630 ( .B1(net77084), .B2(n9585), .A(n5015), .ZN(n9586) );
  AOI21_X1 U5631 ( .B1(net71085), .B2(n10016), .A(n5055), .ZN(n9950) );
  INV_X8 U5632 ( .A(net78003), .ZN(net71078) );
  NOR2_X1 U5633 ( .A1(net70709), .A2(n9606), .ZN(net71280) );
  AOI222_X1 U5634 ( .A1(n6083), .A2(n10103), .B1(n10102), .B2(n10541), .C1(
        net70713), .C2(net71026), .ZN(n10152) );
  OAI21_X1 U5635 ( .B1(net71299), .B2(net70718), .A(net71300), .ZN(n10151) );
  AOI21_X2 U5636 ( .B1(n5638), .B2(net70727), .A(net76452), .ZN(net70693) );
  OAI21_X1 U5637 ( .B1(net71027), .B2(net105349), .A(net72163), .ZN(n5712) );
  OAI21_X2 U5638 ( .B1(n7890), .B2(n7889), .A(n6011), .ZN(n7924) );
  OAI21_X1 U5639 ( .B1(n7900), .B2(n7899), .A(net77588), .ZN(n7923) );
  OAI21_X1 U5640 ( .B1(n7910), .B2(n7909), .A(n6019), .ZN(n7922) );
  NOR2_X2 U5641 ( .A1(net76464), .A2(n8871), .ZN(n8872) );
  NOR2_X2 U5642 ( .A1(net77999), .A2(n5694), .ZN(net73166) );
  NOR2_X2 U5643 ( .A1(net76464), .A2(n10001), .ZN(n10002) );
  NOR2_X2 U5644 ( .A1(net77999), .A2(n10041), .ZN(n9999) );
  OAI21_X2 U5645 ( .B1(n7934), .B2(n7933), .A(n6011), .ZN(n7966) );
  OAI21_X2 U5646 ( .B1(n7944), .B2(n7943), .A(net77588), .ZN(n7965) );
  OAI21_X2 U5647 ( .B1(n7954), .B2(n7953), .A(n6019), .ZN(n7964) );
  OAI21_X2 U5648 ( .B1(net76464), .B2(n5597), .A(net70740), .ZN(n5596) );
  AOI21_X1 U5649 ( .B1(net73878), .B2(n8295), .A(net73997), .ZN(n8385) );
  INV_X4 U5650 ( .A(net70531), .ZN(net73858) );
  OAI21_X2 U5651 ( .B1(n7846), .B2(n7845), .A(n6011), .ZN(n7880) );
  OAI21_X1 U5652 ( .B1(n7856), .B2(n7855), .A(net77588), .ZN(n7879) );
  OAI21_X1 U5653 ( .B1(n7866), .B2(n7865), .A(n6019), .ZN(n7878) );
  NAND4_X2 U5654 ( .A1(n6996), .A2(n6995), .A3(n6997), .A4(n6994), .ZN(n5936)
         );
  NOR2_X2 U5655 ( .A1(net76464), .A2(n8737), .ZN(n8738) );
  NOR2_X2 U5656 ( .A1(n5014), .A2(net70738), .ZN(n8739) );
  NOR2_X2 U5657 ( .A1(net77999), .A2(n9108), .ZN(n8785) );
  NOR2_X2 U5658 ( .A1(net70811), .A2(n10083), .ZN(n8784) );
  AOI21_X1 U5659 ( .B1(n8788), .B2(net77030), .A(n8787), .ZN(n8789) );
  NOR2_X2 U5660 ( .A1(net76464), .A2(n8786), .ZN(n8787) );
  AOI21_X1 U5661 ( .B1(n8908), .B2(net77030), .A(n8907), .ZN(n8909) );
  NOR2_X2 U5662 ( .A1(net76464), .A2(n8906), .ZN(n8907) );
  NOR2_X2 U5663 ( .A1(n8905), .A2(n8904), .ZN(n8910) );
  NOR2_X2 U5664 ( .A1(net70811), .A2(n10041), .ZN(n8904) );
  NOR2_X2 U5665 ( .A1(net77999), .A2(n9862), .ZN(n8905) );
  INV_X8 U5666 ( .A(n9009), .ZN(n6031) );
  NOR2_X2 U5667 ( .A1(n8997), .A2(net72947), .ZN(n9002) );
  OAI21_X2 U5668 ( .B1(n7802), .B2(n7801), .A(n6011), .ZN(n7836) );
  OAI21_X1 U5669 ( .B1(n7812), .B2(n7811), .A(net77588), .ZN(n7835) );
  OAI21_X2 U5670 ( .B1(n7832), .B2(n7831), .A(net77290), .ZN(n7833) );
  OAI21_X1 U5671 ( .B1(net73519), .B2(n8461), .A(net73780), .ZN(n8463) );
  NOR2_X2 U5672 ( .A1(n10505), .A2(net76464), .ZN(n9699) );
  NOR2_X2 U5673 ( .A1(net77999), .A2(n9816), .ZN(n9819) );
  NOR2_X2 U5674 ( .A1(net70811), .A2(n9817), .ZN(n9818) );
  NOR2_X2 U5675 ( .A1(n9822), .A2(n9821), .ZN(n9823) );
  NOR2_X1 U5676 ( .A1(instructionAddr_out[29]), .A2(net70738), .ZN(n9822) );
  NOR2_X2 U5677 ( .A1(net76464), .A2(n9820), .ZN(n9821) );
  OAI21_X1 U5678 ( .B1(net73496), .B2(net73780), .A(reset), .ZN(n10650) );
  NOR2_X2 U5679 ( .A1(net76646), .A2(n10503), .ZN(n10508) );
  NOR2_X2 U5680 ( .A1(net77999), .A2(n10504), .ZN(n10507) );
  NOR2_X2 U5681 ( .A1(net70811), .A2(n10505), .ZN(n10506) );
  NOR2_X1 U5682 ( .A1(net73503), .A2(net73499), .ZN(n8658) );
  NOR2_X1 U5683 ( .A1(net73498), .A2(net73499), .ZN(n8659) );
  NAND3_X1 U5684 ( .A1(n8655), .A2(net73170), .A3(n8654), .ZN(net70506) );
  NOR2_X2 U5685 ( .A1(instruction[1]), .A2(n8653), .ZN(n8654) );
  NAND4_X2 U5686 ( .A1(n6575), .A2(n6574), .A3(n6572), .A4(n6573), .ZN(n6581)
         );
  AOI22_X2 U5687 ( .A1(\REGFILE/reg_out[19][15] ), .A2(net77812), .B1(
        \REGFILE/reg_out[1][15] ), .B2(net75478), .ZN(n6585) );
  NAND3_X2 U5688 ( .A1(n10107), .A2(n5042), .A3(n10106), .ZN(n10108) );
  AOI21_X1 U5689 ( .B1(n10261), .B2(net77030), .A(n10260), .ZN(n10262) );
  NOR2_X2 U5690 ( .A1(net76464), .A2(n10259), .ZN(n10260) );
  NOR2_X2 U5691 ( .A1(n10000), .A2(net72876), .ZN(n9043) );
  INV_X4 U5692 ( .A(n4878), .ZN(n6132) );
  INV_X4 U5693 ( .A(n4867), .ZN(n6088) );
  INV_X4 U5694 ( .A(n4990), .ZN(n6156) );
  INV_X4 U5695 ( .A(n6093), .ZN(n6091) );
  INV_X4 U5696 ( .A(n6100), .ZN(n6097) );
  INV_X4 U5697 ( .A(n4804), .ZN(n6108) );
  INV_X4 U5698 ( .A(n4891), .ZN(n6112) );
  INV_X4 U5699 ( .A(n4892), .ZN(n6115) );
  INV_X4 U5700 ( .A(n4884), .ZN(n6118) );
  INV_X4 U5701 ( .A(n4877), .ZN(net76862) );
  INV_X4 U5702 ( .A(n4882), .ZN(n6121) );
  INV_X4 U5703 ( .A(n4888), .ZN(n6124) );
  INV_X4 U5704 ( .A(n4883), .ZN(n6127) );
  INV_X4 U5705 ( .A(n4875), .ZN(n6129) );
  INV_X4 U5706 ( .A(n4893), .ZN(n6136) );
  INV_X4 U5707 ( .A(n4879), .ZN(n6139) );
  INV_X4 U5708 ( .A(n4885), .ZN(n6144) );
  INV_X4 U5709 ( .A(n4889), .ZN(net76706) );
  INV_X4 U5710 ( .A(n4886), .ZN(net76692) );
  INV_X4 U5711 ( .A(n4890), .ZN(n6150) );
  INV_X4 U5712 ( .A(n4887), .ZN(n6153) );
  INV_X4 U5713 ( .A(n4876), .ZN(n6200) );
  INV_X4 U5714 ( .A(n4876), .ZN(n6202) );
  INV_X4 U5715 ( .A(n4867), .ZN(n6089) );
  INV_X4 U5716 ( .A(n6093), .ZN(n6092) );
  INV_X4 U5717 ( .A(n6100), .ZN(n6098) );
  INV_X4 U5718 ( .A(n4804), .ZN(n6109) );
  INV_X4 U5719 ( .A(n4891), .ZN(n6113) );
  INV_X4 U5720 ( .A(n4892), .ZN(n6116) );
  INV_X4 U5721 ( .A(n4884), .ZN(n6119) );
  INV_X4 U5722 ( .A(n4877), .ZN(net76864) );
  INV_X4 U5723 ( .A(n4882), .ZN(n6122) );
  INV_X4 U5724 ( .A(n4888), .ZN(n6125) );
  INV_X4 U5725 ( .A(n4883), .ZN(n6128) );
  INV_X4 U5726 ( .A(n4875), .ZN(n6130) );
  INV_X4 U5727 ( .A(n4878), .ZN(n6133) );
  INV_X4 U5728 ( .A(n4893), .ZN(n6137) );
  INV_X4 U5729 ( .A(n4879), .ZN(n6140) );
  INV_X4 U5730 ( .A(n4885), .ZN(n6145) );
  INV_X4 U5731 ( .A(n4889), .ZN(net76708) );
  INV_X4 U5732 ( .A(n4886), .ZN(net76694) );
  INV_X4 U5733 ( .A(n4890), .ZN(n6151) );
  INV_X4 U5734 ( .A(n4887), .ZN(n6154) );
  AOI21_X1 U5735 ( .B1(n10294), .B2(net77030), .A(n10293), .ZN(n10295) );
  INV_X4 U5736 ( .A(n4867), .ZN(n6090) );
  INV_X4 U5737 ( .A(n6100), .ZN(n6099) );
  INV_X4 U5738 ( .A(n6096), .ZN(n6094) );
  INV_X4 U5739 ( .A(n4804), .ZN(n6110) );
  INV_X4 U5740 ( .A(n6107), .ZN(n6105) );
  INV_X4 U5741 ( .A(n4876), .ZN(n6201) );
  INV_X4 U5742 ( .A(n4877), .ZN(net76866) );
  INV_X4 U5743 ( .A(n4875), .ZN(n6131) );
  INV_X4 U5744 ( .A(n4878), .ZN(n6134) );
  INV_X4 U5745 ( .A(n4879), .ZN(n6141) );
  INV_X4 U5746 ( .A(n6148), .ZN(n6146) );
  NOR2_X2 U5747 ( .A1(n6190), .A2(n10651), .ZN(n10652) );
  NOR2_X2 U5748 ( .A1(\PCLOGIC/imm16_32 [31]), .A2(n10650), .ZN(n10651) );
  NAND2_X2 U5749 ( .A1(n6408), .A2(n6407), .ZN(dmem_write_out[24]) );
  NAND2_X2 U5750 ( .A1(n6454), .A2(n6455), .ZN(dmem_write_out[22]) );
  NAND2_X2 U5751 ( .A1(n6479), .A2(n6478), .ZN(dmem_write_out[21]) );
  NAND2_X2 U5752 ( .A1(n6503), .A2(n6502), .ZN(n10944) );
  NAND2_X2 U5753 ( .A1(n6753), .A2(n6752), .ZN(dmem_write_out[8]) );
  NAND2_X2 U5754 ( .A1(n6850), .A2(n6851), .ZN(dmem_write_out[3]) );
  NAND2_X2 U5755 ( .A1(n6895), .A2(n6894), .ZN(dmem_write_out[1]) );
  NAND3_X2 U5756 ( .A1(n8734), .A2(n8733), .A3(n8732), .ZN(n8735) );
  NAND3_X2 U5757 ( .A1(n9815), .A2(n9814), .A3(n9813), .ZN(dmem_addr_out[29])
         );
  AOI21_X2 U5758 ( .B1(net71271), .B2(n9812), .A(n9811), .ZN(n9813) );
  OAI21_X2 U5759 ( .B1(n8770), .B2(n8769), .A(net70697), .ZN(n8782) );
  OAI21_X1 U5760 ( .B1(n8900), .B2(n8899), .A(net70697), .ZN(n8902) );
  AOI21_X2 U5761 ( .B1(net71271), .B2(n8889), .A(n8888), .ZN(n8903) );
  OAI21_X1 U5762 ( .B1(n9773), .B2(n9772), .A(net70697), .ZN(n9786) );
  AOI21_X2 U5763 ( .B1(n9784), .B2(n9783), .A(n9782), .ZN(n9785) );
  AOI21_X2 U5764 ( .B1(net71271), .B2(n8603), .A(n8602), .ZN(n8649) );
  AOI21_X2 U5765 ( .B1(net71271), .B2(n9292), .A(n9291), .ZN(n9312) );
  AOI21_X2 U5766 ( .B1(net71271), .B2(n8923), .A(n8922), .ZN(n8948) );
  AOI21_X2 U5767 ( .B1(net71271), .B2(n9545), .A(n9544), .ZN(n9565) );
  AOI21_X2 U5768 ( .B1(net71271), .B2(n8835), .A(n8834), .ZN(n8869) );
  AOI21_X1 U5769 ( .B1(n10064), .B2(n9182), .A(n9181), .ZN(n9200) );
  NOR2_X2 U5770 ( .A1(n9198), .A2(n9197), .ZN(n9199) );
  AOI21_X1 U5771 ( .B1(n10064), .B2(n10248), .A(n5050), .ZN(n9418) );
  AOI21_X1 U5772 ( .B1(n10064), .B2(n9403), .A(n5049), .ZN(n9104) );
  AOI21_X1 U5773 ( .B1(n10064), .B2(n9837), .A(n5054), .ZN(n9859) );
  AOI21_X1 U5774 ( .B1(net70697), .B2(n9338), .A(n9337), .ZN(n9372) );
  AOI21_X2 U5775 ( .B1(net71271), .B2(n9368), .A(n9367), .ZN(n9369) );
  AOI21_X1 U5776 ( .B1(n10064), .B2(n9685), .A(n5053), .ZN(n9696) );
  AOI21_X2 U5777 ( .B1(net71271), .B2(n9628), .A(n9627), .ZN(n9629) );
  AOI21_X1 U5778 ( .B1(n10649), .B2(n10642), .A(n6190), .ZN(n10646) );
  NOR2_X2 U5779 ( .A1(net73855), .A2(n8462), .ZN(n8468) );
  NOR2_X2 U5780 ( .A1(n8474), .A2(n8473), .ZN(n8478) );
  NOR2_X2 U5781 ( .A1(n8488), .A2(n8487), .ZN(n8492) );
  NOR2_X2 U5782 ( .A1(n8522), .A2(n8521), .ZN(n8526) );
  NAND3_X2 U5783 ( .A1(n8705), .A2(n8704), .A3(n8703), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  NAND3_X1 U5784 ( .A1(n10649), .A2(n8702), .A3(n8701), .ZN(n8704) );
  OAI21_X2 U5785 ( .B1(n6223), .B2(n6138), .A(n8753), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5786 ( .B1(n6223), .B2(n10534), .A(n8754), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5787 ( .B1(n6221), .B2(n10532), .A(n8793), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5788 ( .B1(n6221), .B2(n6142), .A(n8794), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5789 ( .B1(n6221), .B2(net70509), .A(n8795), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5790 ( .B1(n6213), .B2(n6023), .A(n8878), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5791 ( .B1(n6138), .B2(n6023), .A(n8879), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5792 ( .B1(n6142), .B2(n6023), .A(n8880), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5793 ( .B1(net76480), .B2(n6023), .A(n8881), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5794 ( .B1(n6213), .B2(n6025), .A(n8913), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5795 ( .B1(n6138), .B2(n6025), .A(n8914), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5796 ( .B1(n6142), .B2(n6025), .A(n8915), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5797 ( .B1(net76480), .B2(n6025), .A(n8916), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  NAND3_X2 U5798 ( .A1(n8973), .A2(n8972), .A3(n8971), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5799 ( .B1(n6213), .B2(n6032), .A(n9046), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5800 ( .B1(n6138), .B2(n6032), .A(n9047), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5801 ( .B1(n6142), .B2(n6032), .A(n9048), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5802 ( .B1(net76480), .B2(n6032), .A(n9049), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  NOR2_X1 U5803 ( .A1(n4968), .A2(n9271), .ZN(n9276) );
  NAND3_X2 U5804 ( .A1(n9288), .A2(n9287), .A3(n9286), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  NAND3_X2 U5805 ( .A1(n9541), .A2(n9540), .A3(n9539), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5806 ( .B1(n6056), .B2(n6138), .A(n9678), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5807 ( .B1(n6142), .B2(n4802), .A(n9679), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5808 ( .B1(net76480), .B2(n6057), .A(n9680), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5809 ( .B1(n6222), .B2(n10532), .A(n9829), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5810 ( .B1(n6222), .B2(n10534), .A(n9830), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5811 ( .B1(n6222), .B2(net70509), .A(n9831), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5812 ( .B1(n6214), .B2(n6068), .A(n9969), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5813 ( .B1(n10532), .B2(n4803), .A(n9970), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5814 ( .B1(n10534), .B2(n4803), .A(n9971), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5815 ( .B1(net70509), .B2(n6068), .A(n9972), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5816 ( .B1(n6214), .B2(n6070), .A(n10008), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5817 ( .B1(n10532), .B2(n6070), .A(n10009), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5818 ( .B1(n10534), .B2(n6070), .A(n10010), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5819 ( .B1(net70509), .B2(n6070), .A(n10011), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5820 ( .B1(n6214), .B2(n6085), .A(n10271), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5821 ( .B1(n10532), .B2(n6085), .A(n10272), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5822 ( .B1(n10534), .B2(n6085), .A(n10273), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5823 ( .B1(net70509), .B2(n6085), .A(n10274), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5824 ( .B1(n6214), .B2(n6087), .A(n10299), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5825 ( .B1(n10532), .B2(n6087), .A(n10300), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5826 ( .B1(n10534), .B2(n6087), .A(n10301), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5827 ( .B1(net70509), .B2(n6087), .A(n10302), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5828 ( .B1(n6214), .B2(n6191), .A(n10530), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5829 ( .B1(n6191), .B2(n6138), .A(n10531), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U5830 ( .B1(n6191), .B2(n6142), .A(n10533), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  NOR2_X2 U5831 ( .A1(net76278), .A2(net76658), .ZN(n10546) );
  NOR2_X2 U5832 ( .A1(net76278), .A2(n6155), .ZN(n10549) );
  NOR2_X2 U5833 ( .A1(n6194), .A2(net76274), .ZN(n10552) );
  NOR2_X2 U5834 ( .A1(n6198), .A2(net76274), .ZN(n10555) );
  NAND3_X2 U5835 ( .A1(n6096), .A2(reset), .A3(net76510), .ZN(n10559) );
  NAND3_X2 U5836 ( .A1(n6101), .A2(reset), .A3(net76510), .ZN(n10561) );
  NAND3_X2 U5837 ( .A1(n6107), .A2(reset), .A3(net76510), .ZN(n10563) );
  NOR2_X2 U5838 ( .A1(net76278), .A2(n6157), .ZN(n10564) );
  NOR2_X2 U5839 ( .A1(net76278), .A2(n6159), .ZN(n10567) );
  NOR2_X2 U5840 ( .A1(net76278), .A2(n6161), .ZN(n10570) );
  NOR2_X2 U5841 ( .A1(n6203), .A2(net76274), .ZN(n10573) );
  NOR2_X2 U5842 ( .A1(net76278), .A2(net76614), .ZN(n10576) );
  NOR2_X2 U5843 ( .A1(n6207), .A2(net76274), .ZN(n10579) );
  NOR2_X2 U5844 ( .A1(net76278), .A2(n6163), .ZN(n10582) );
  NOR2_X2 U5845 ( .A1(net76278), .A2(n6165), .ZN(n10585) );
  NOR2_X2 U5846 ( .A1(net76278), .A2(n6167), .ZN(n10588) );
  NOR2_X2 U5847 ( .A1(net76278), .A2(n6169), .ZN(n10591) );
  NOR2_X2 U5848 ( .A1(net76278), .A2(n6171), .ZN(n10594) );
  NOR2_X2 U5849 ( .A1(net76278), .A2(n6173), .ZN(n10597) );
  NOR2_X2 U5850 ( .A1(n6211), .A2(net76274), .ZN(n10600) );
  NOR2_X2 U5851 ( .A1(n6214), .A2(net76274), .ZN(n10603) );
  NAND3_X2 U5852 ( .A1(n10607), .A2(reset), .A3(net76510), .ZN(n10610) );
  NOR2_X2 U5853 ( .A1(net76278), .A2(net76548), .ZN(n10611) );
  NAND3_X2 U5854 ( .A1(n10614), .A2(reset), .A3(net76510), .ZN(n10617) );
  NAND3_X2 U5855 ( .A1(net70574), .A2(reset), .A3(net76510), .ZN(n10619) );
  NOR2_X2 U5856 ( .A1(net76318), .A2(net76274), .ZN(n10620) );
  NOR2_X2 U5857 ( .A1(n6219), .A2(net76274), .ZN(n10623) );
  NOR2_X2 U5858 ( .A1(net76278), .A2(n6182), .ZN(n10626) );
  NAND3_X2 U5859 ( .A1(n6148), .A2(reset), .A3(net76510), .ZN(n10630) );
  NOR2_X2 U5860 ( .A1(net76278), .A2(n6184), .ZN(n10631) );
  NOR2_X2 U5861 ( .A1(net76278), .A2(n6186), .ZN(n10634) );
  NOR2_X2 U5862 ( .A1(net76278), .A2(n6188), .ZN(n10637) );
  OAI21_X2 U5863 ( .B1(n6191), .B2(net76480), .A(n10656), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  AND2_X4 U5864 ( .A1(reset), .A2(net76660), .ZN(n4867) );
  AND2_X4 U5865 ( .A1(net76270), .A2(n6208), .ZN(n4868) );
  AND2_X4 U5866 ( .A1(net76270), .A2(n6195), .ZN(n4869) );
  AND2_X4 U5867 ( .A1(net76270), .A2(n6220), .ZN(n4870) );
  AND2_X4 U5868 ( .A1(net76270), .A2(net76320), .ZN(n4871) );
  AND2_X4 U5869 ( .A1(net76270), .A2(n6212), .ZN(n4872) );
  AND2_X4 U5870 ( .A1(net76270), .A2(n6199), .ZN(n4873) );
  AND2_X4 U5871 ( .A1(n8669), .A2(n8672), .ZN(n4874) );
  INV_X4 U5872 ( .A(n10604), .ZN(n6176) );
  INV_X16 U5873 ( .A(n9765), .ZN(n6061) );
  INV_X4 U5874 ( .A(n10012), .ZN(n6071) );
  INV_X16 U5875 ( .A(n6071), .ZN(n6070) );
  AND2_X4 U5876 ( .A1(net76270), .A2(n6170), .ZN(n4875) );
  AND2_X4 U5877 ( .A1(net76270), .A2(n6204), .ZN(n4876) );
  AND2_X4 U5878 ( .A1(net76270), .A2(net76616), .ZN(n4877) );
  AND2_X4 U5879 ( .A1(net76270), .A2(n6172), .ZN(n4878) );
  AND2_X4 U5880 ( .A1(net76270), .A2(net76550), .ZN(n4879) );
  AND2_X4 U5881 ( .A1(n6005), .A2(net78051), .ZN(n4880) );
  INV_X4 U5882 ( .A(n6101), .ZN(n6102) );
  INV_X4 U5883 ( .A(n6148), .ZN(n6147) );
  AND2_X4 U5884 ( .A1(net75791), .A2(net73697), .ZN(n4881) );
  INV_X8 U5885 ( .A(n5642), .ZN(n5644) );
  INV_X8 U5886 ( .A(n8402), .ZN(n6020) );
  INV_X4 U5887 ( .A(n10276), .ZN(n6086) );
  INV_X16 U5888 ( .A(n6086), .ZN(n6085) );
  INV_X4 U5889 ( .A(net76274), .ZN(net76270) );
  AND2_X4 U5890 ( .A1(net76270), .A2(n6164), .ZN(n4882) );
  AND2_X4 U5891 ( .A1(net76270), .A2(n6168), .ZN(n4883) );
  AND2_X4 U5892 ( .A1(net76270), .A2(n6162), .ZN(n4884) );
  AND2_X4 U5893 ( .A1(net76270), .A2(n6183), .ZN(n4885) );
  AND2_X4 U5894 ( .A1(net76270), .A2(n6185), .ZN(n4886) );
  AND2_X4 U5895 ( .A1(net76270), .A2(n6189), .ZN(n4887) );
  AND2_X4 U5896 ( .A1(net76270), .A2(n6166), .ZN(n4888) );
  AND2_X4 U5897 ( .A1(net76270), .A2(n10535), .ZN(n4889) );
  AND2_X4 U5898 ( .A1(net76270), .A2(n6187), .ZN(n4890) );
  AND2_X4 U5899 ( .A1(net76270), .A2(n6158), .ZN(n4891) );
  AND2_X4 U5900 ( .A1(net76270), .A2(n6160), .ZN(n4892) );
  AND2_X4 U5901 ( .A1(net76270), .A2(n6174), .ZN(n4893) );
  NAND4_X2 U5902 ( .A1(n6941), .A2(n6938), .A3(n6940), .A4(n6939), .ZN(
        net73837) );
  INV_X4 U5903 ( .A(net76650), .ZN(net76646) );
  INV_X4 U5904 ( .A(net73877), .ZN(net73997) );
  AND3_X4 U5905 ( .A1(n4900), .A2(net73429), .A3(net73443), .ZN(n4894) );
  NOR2_X2 U5906 ( .A1(n8677), .A2(net73434), .ZN(net70574) );
  NOR2_X2 U5907 ( .A1(n8677), .A2(net73439), .ZN(n10607) );
  NOR2_X2 U5908 ( .A1(n8677), .A2(net73436), .ZN(n10614) );
  AND3_X4 U5909 ( .A1(net73427), .A2(n4900), .A3(net73429), .ZN(n4895) );
  INV_X4 U5910 ( .A(n4872), .ZN(n6210) );
  INV_X4 U5911 ( .A(n4869), .ZN(n6193) );
  INV_X4 U5912 ( .A(n4868), .ZN(n6206) );
  INV_X4 U5913 ( .A(n4871), .ZN(n6216) );
  INV_X4 U5914 ( .A(n4870), .ZN(n6218) );
  INV_X4 U5915 ( .A(n4880), .ZN(n6084) );
  INV_X4 U5916 ( .A(n6084), .ZN(n6083) );
  AND2_X4 U5917 ( .A1(n8766), .A2(n8765), .ZN(n4896) );
  INV_X4 U5918 ( .A(n10544), .ZN(n6081) );
  INV_X4 U5920 ( .A(n8882), .ZN(n6024) );
  INV_X16 U5921 ( .A(n6024), .ZN(n6023) );
  INV_X4 U5922 ( .A(n9268), .ZN(n6037) );
  INV_X8 U5923 ( .A(n6037), .ZN(n6036) );
  INV_X8 U5924 ( .A(n6037), .ZN(n6035) );
  INV_X16 U5925 ( .A(n4816), .ZN(n6034) );
  INV_X16 U5926 ( .A(n4816), .ZN(n6033) );
  INV_X16 U5927 ( .A(n9426), .ZN(n6047) );
  INV_X16 U5928 ( .A(n9426), .ZN(n6046) );
  INV_X16 U5929 ( .A(n9868), .ZN(n6066) );
  INV_X16 U5930 ( .A(n9868), .ZN(n6065) );
  NAND2_X1 U5931 ( .A1(n4966), .A2(net73495), .ZN(net70738) );
  INV_X4 U5932 ( .A(net70738), .ZN(net77030) );
  INV_X4 U5933 ( .A(net80189), .ZN(net73608) );
  AND2_X4 U5934 ( .A1(net73494), .A2(net70507), .ZN(n4899) );
  AND2_X4 U5935 ( .A1(n5589), .A2(n5066), .ZN(n4900) );
  INV_X4 U5936 ( .A(net70718), .ZN(net105360) );
  AND2_X4 U5937 ( .A1(n5010), .A2(n4874), .ZN(n4903) );
  AND2_X4 U5938 ( .A1(n5010), .A2(net73416), .ZN(n4904) );
  AND2_X4 U5939 ( .A1(n5010), .A2(net73423), .ZN(n4905) );
  AND2_X4 U5940 ( .A1(n5010), .A2(net73421), .ZN(n4906) );
  NAND2_X2 U5941 ( .A1(n8464), .A2(n8463), .ZN(n9533) );
  INV_X4 U5942 ( .A(n9533), .ZN(n10649) );
  AND2_X4 U5943 ( .A1(n5066), .A2(net73468), .ZN(n4907) );
  AND2_X2 U5944 ( .A1(net70821), .A2(n8580), .ZN(n4910) );
  NAND2_X1 U5945 ( .A1(net78051), .A2(n10099), .ZN(n10094) );
  AND2_X4 U5946 ( .A1(dmem_dsize[1]), .A2(n4899), .ZN(n4911) );
  AND2_X2 U5947 ( .A1(n8728), .A2(n6041), .ZN(n4912) );
  AND2_X4 U5948 ( .A1(n5068), .A2(net73443), .ZN(n4913) );
  AND2_X4 U5949 ( .A1(n5067), .A2(net73443), .ZN(n4914) );
  NAND2_X2 U5950 ( .A1(net73500), .A2(net70738), .ZN(n4915) );
  INV_X4 U5951 ( .A(n8917), .ZN(n6026) );
  INV_X16 U5952 ( .A(n6026), .ZN(n6025) );
  AND2_X4 U5953 ( .A1(net73427), .A2(n5068), .ZN(n4916) );
  INV_X4 U5954 ( .A(reset), .ZN(net76274) );
  AND2_X4 U5955 ( .A1(n5067), .A2(net73427), .ZN(n4920) );
  AND2_X4 U5956 ( .A1(n8301), .A2(net73877), .ZN(n4921) );
  NAND2_X2 U5957 ( .A1(n4910), .A2(net73585), .ZN(net70691) );
  AND2_X4 U5958 ( .A1(n8768), .A2(n8767), .ZN(n4922) );
  NOR2_X2 U5959 ( .A1(net70574), .A2(net76274), .ZN(n5688) );
  NOR2_X2 U5960 ( .A1(n10607), .A2(net76274), .ZN(n10608) );
  NAND3_X2 U5961 ( .A1(reset), .A2(instruction[1]), .A3(n5591), .ZN(n4962) );
  INV_X4 U5962 ( .A(n10517), .ZN(n6100) );
  INV_X2 U5963 ( .A(net77276), .ZN(net123282) );
  INV_X16 U5964 ( .A(net77784), .ZN(net77780) );
  INV_X16 U5965 ( .A(net77832), .ZN(net77828) );
  INV_X16 U5966 ( .A(net75468), .ZN(net77776) );
  INV_X8 U5967 ( .A(n8411), .ZN(n6013) );
  INV_X16 U5968 ( .A(n6013), .ZN(n6012) );
  INV_X8 U5969 ( .A(net73838), .ZN(net77296) );
  INV_X16 U5970 ( .A(net77296), .ZN(net77292) );
  INV_X16 U5971 ( .A(net75443), .ZN(net77656) );
  AND2_X4 U5972 ( .A1(net76270), .A2(n9045), .ZN(n4964) );
  AND2_X4 U5973 ( .A1(reset), .A2(n10297), .ZN(n4965) );
  AND3_X4 U5974 ( .A1(instruction[4]), .A2(net74029), .A3(net73499), .ZN(n4966) );
  AND3_X4 U5975 ( .A1(net73684), .A2(\PCLOGIC/imm16_32 [29]), .A3(net73619), 
        .ZN(n4967) );
  XOR2_X2 U5976 ( .A(\PCLOGIC/imm16_32 [19]), .B(n10003), .Z(n4968) );
  AND4_X2 U5977 ( .A1(n5593), .A2(net71266), .A3(n5594), .A4(n5595), .ZN(n4970) );
  OR2_X2 U5978 ( .A1(\PCLOGIC/imm16_32 [28]), .A2(\PCLOGIC/imm16_32 [29]), 
        .ZN(n4971) );
  INV_X8 U5979 ( .A(n5628), .ZN(net77042) );
  INV_X4 U5980 ( .A(n5797), .ZN(n5955) );
  INV_X4 U5981 ( .A(net77504), .ZN(net77484) );
  INV_X8 U5982 ( .A(net77504), .ZN(net77482) );
  AND2_X4 U5983 ( .A1(net73423), .A2(n4913), .ZN(n4990) );
  AND2_X4 U5984 ( .A1(n4874), .A2(n4913), .ZN(n4991) );
  AND2_X4 U5985 ( .A1(n4916), .A2(n4874), .ZN(n4992) );
  AND2_X4 U5986 ( .A1(n4894), .A2(n4874), .ZN(n4993) );
  AND2_X4 U5987 ( .A1(n4920), .A2(n4874), .ZN(n4994) );
  AND2_X4 U5988 ( .A1(n4914), .A2(n4874), .ZN(n4995) );
  AND2_X4 U5989 ( .A1(n4895), .A2(n4874), .ZN(n4996) );
  AND2_X4 U5990 ( .A1(n4916), .A2(net73416), .ZN(n4997) );
  AND2_X4 U5991 ( .A1(n4913), .A2(net73421), .ZN(n4998) );
  AND2_X4 U5992 ( .A1(n4920), .A2(net73416), .ZN(n4999) );
  AND2_X4 U5993 ( .A1(n4920), .A2(net73423), .ZN(n5000) );
  AND2_X4 U5994 ( .A1(n4920), .A2(net73421), .ZN(n5001) );
  AND2_X4 U5995 ( .A1(n4914), .A2(net73416), .ZN(n5002) );
  AND2_X4 U5996 ( .A1(n4914), .A2(net73423), .ZN(n5003) );
  AND2_X4 U5997 ( .A1(n4914), .A2(net73421), .ZN(n5004) );
  AND2_X4 U5998 ( .A1(n4916), .A2(net73423), .ZN(n5005) );
  AND2_X4 U5999 ( .A1(n4895), .A2(net73416), .ZN(n5006) );
  AND2_X4 U6000 ( .A1(n4895), .A2(net73421), .ZN(n5007) );
  AND2_X4 U6001 ( .A1(n4913), .A2(net73416), .ZN(n5008) );
  AND2_X4 U6002 ( .A1(n4916), .A2(net73421), .ZN(n5009) );
  INV_X4 U6003 ( .A(n5577), .ZN(n5944) );
  AND3_X4 U6004 ( .A1(net73427), .A2(n4907), .A3(net73429), .ZN(n5010) );
  NAND3_X2 U6005 ( .A1(n8539), .A2(instruction[1]), .A3(net73170), .ZN(n8565)
         );
  AND2_X4 U6006 ( .A1(net76270), .A2(n8742), .ZN(n5011) );
  AND2_X4 U6007 ( .A1(net76270), .A2(n8792), .ZN(n5012) );
  AND2_X4 U6008 ( .A1(net76270), .A2(n9826), .ZN(n5013) );
  INV_X4 U6009 ( .A(n10400), .ZN(n10909) );
  AND2_X2 U6010 ( .A1(n4880), .A2(net70696), .ZN(n5015) );
  INV_X4 U6011 ( .A(net85047), .ZN(net84663) );
  AND2_X2 U6012 ( .A1(net70701), .A2(n10416), .ZN(n5039) );
  AND2_X2 U6013 ( .A1(net70701), .A2(n10415), .ZN(n5040) );
  AND2_X2 U6014 ( .A1(net70701), .A2(n10414), .ZN(n5041) );
  OR2_X4 U6015 ( .A1(n10093), .A2(net70710), .ZN(n5042) );
  NAND2_X2 U6016 ( .A1(n8464), .A2(n8463), .ZN(n6008) );
  AND2_X2 U6017 ( .A1(net70701), .A2(n10373), .ZN(n5049) );
  AND2_X2 U6018 ( .A1(net70701), .A2(n9402), .ZN(n5050) );
  AND2_X2 U6019 ( .A1(net70701), .A2(n10387), .ZN(n5051) );
  AND2_X2 U6020 ( .A1(net70701), .A2(n10394), .ZN(n5052) );
  AND2_X2 U6021 ( .A1(net70701), .A2(n10307), .ZN(n5053) );
  AND2_X2 U6022 ( .A1(net70701), .A2(n9836), .ZN(n5054) );
  AND2_X2 U6023 ( .A1(net70701), .A2(n10402), .ZN(n5055) );
  AND2_X2 U6024 ( .A1(net70701), .A2(n10380), .ZN(n5056) );
  AND2_X2 U6025 ( .A1(net70701), .A2(n10366), .ZN(n5057) );
  AND2_X2 U6026 ( .A1(net70701), .A2(n10281), .ZN(n5058) );
  AND3_X4 U6027 ( .A1(n8981), .A2(n8980), .A3(n8979), .ZN(n5061) );
  AND3_X4 U6028 ( .A1(n10542), .A2(net80189), .A3(net71094), .ZN(n5062) );
  AND2_X4 U6029 ( .A1(net70706), .A2(net73541), .ZN(n5065) );
  AND3_X4 U6030 ( .A1(n5590), .A2(net70506), .A3(net73519), .ZN(n5066) );
  AND2_X4 U6031 ( .A1(net73465), .A2(n4907), .ZN(n5067) );
  AND2_X4 U6032 ( .A1(net73465), .A2(n4900), .ZN(n5068) );
  AND2_X2 U6033 ( .A1(n8553), .A2(n8536), .ZN(n5252) );
  INV_X4 U6034 ( .A(n8527), .ZN(n6190) );
  INV_X4 U6035 ( .A(n4911), .ZN(net77999) );
  INV_X4 U6036 ( .A(n10608), .ZN(n6179) );
  INV_X4 U6037 ( .A(n6179), .ZN(n6178) );
  INV_X4 U6038 ( .A(n10615), .ZN(n6181) );
  NOR2_X2 U6039 ( .A1(n10614), .A2(net76274), .ZN(n10615) );
  INV_X4 U6040 ( .A(n6181), .ZN(n6180) );
  INV_X4 U6041 ( .A(n5688), .ZN(n5695) );
  INV_X4 U6042 ( .A(n5695), .ZN(net76488) );
  OR2_X4 U6043 ( .A1(n10152), .A2(net70710), .ZN(n5570) );
  INV_X1 U6044 ( .A(net148116), .ZN(net121580) );
  INV_X4 U6045 ( .A(n9330), .ZN(n6042) );
  INV_X8 U6046 ( .A(n6042), .ZN(n6040) );
  INV_X8 U6047 ( .A(n6042), .ZN(n6041) );
  AND2_X2 U6048 ( .A1(n10108), .A2(net73585), .ZN(n5571) );
  INV_X1 U6049 ( .A(n5867), .ZN(n5868) );
  INV_X4 U6050 ( .A(net70507), .ZN(net76468) );
  NAND3_X1 U6051 ( .A1(net73495), .A2(net73496), .A3(n8659), .ZN(net70507) );
  INV_X4 U6052 ( .A(net76468), .ZN(net76464) );
  INV_X4 U6053 ( .A(net70718), .ZN(net77086) );
  OR2_X4 U6054 ( .A1(net76464), .A2(n10540), .ZN(n5572) );
  INV_X4 U6055 ( .A(n10535), .ZN(n6148) );
  INV_X4 U6056 ( .A(n10519), .ZN(n6101) );
  OR2_X4 U6057 ( .A1(net76464), .A2(n10078), .ZN(n5573) );
  INV_X8 U6058 ( .A(net78050), .ZN(net78051) );
  INV_X1 U6059 ( .A(net78051), .ZN(net72962) );
  INV_X4 U6060 ( .A(n6176), .ZN(n6175) );
  INV_X4 U6061 ( .A(n6176), .ZN(n6177) );
  INV_X4 U6062 ( .A(n10607), .ZN(n6138) );
  INV_X4 U6063 ( .A(n10614), .ZN(n6142) );
  INV_X4 U6064 ( .A(net70574), .ZN(net76480) );
  INV_X4 U6065 ( .A(n10516), .ZN(n6096) );
  INV_X4 U6066 ( .A(n6096), .ZN(n6095) );
  INV_X4 U6067 ( .A(n10521), .ZN(n6107) );
  INV_X4 U6068 ( .A(n6107), .ZN(n6106) );
  INV_X4 U6069 ( .A(n4869), .ZN(n6192) );
  INV_X4 U6070 ( .A(n4873), .ZN(n6196) );
  INV_X4 U6071 ( .A(n4873), .ZN(n6197) );
  INV_X4 U6072 ( .A(n4868), .ZN(n6205) );
  INV_X4 U6073 ( .A(n4872), .ZN(n6209) );
  INV_X4 U6074 ( .A(n4871), .ZN(n6215) );
  INV_X4 U6075 ( .A(n4870), .ZN(n6217) );
  INV_X4 U6076 ( .A(n10512), .ZN(n6093) );
  INV_X4 U6077 ( .A(n4805), .ZN(n6103) );
  INV_X4 U6078 ( .A(n4805), .ZN(n6104) );
  INV_X4 U6079 ( .A(n4891), .ZN(n6111) );
  INV_X4 U6080 ( .A(n4892), .ZN(n6114) );
  INV_X4 U6081 ( .A(n4884), .ZN(n6117) );
  INV_X4 U6082 ( .A(n4882), .ZN(n6120) );
  INV_X4 U6083 ( .A(n4888), .ZN(n6123) );
  INV_X4 U6084 ( .A(n4883), .ZN(n6126) );
  INV_X4 U6085 ( .A(n4893), .ZN(n6135) );
  INV_X4 U6086 ( .A(n4885), .ZN(n6143) );
  INV_X4 U6087 ( .A(n4889), .ZN(net76716) );
  INV_X4 U6088 ( .A(n4886), .ZN(net76702) );
  INV_X4 U6089 ( .A(n4890), .ZN(n6149) );
  INV_X4 U6090 ( .A(n4887), .ZN(n6152) );
  INV_X4 U6091 ( .A(n4806), .ZN(n6213) );
  INV_X4 U6092 ( .A(n4915), .ZN(net76650) );
  INV_X4 U6093 ( .A(reset), .ZN(net76278) );
  INV_X16 U6094 ( .A(n10149), .ZN(n6080) );
  NAND2_X4 U6095 ( .A1(n10142), .A2(reset), .ZN(n10149) );
  OAI21_X2 U6096 ( .B1(n6078), .B2(net70509), .A(n10148), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6097 ( .B1(n6078), .B2(n6142), .A(n10147), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6098 ( .B1(n6078), .B2(n6214), .A(n10145), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6099 ( .B1(n6078), .B2(n6138), .A(n10146), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6100 ( .B1(net76480), .B2(n6043), .A(n9382), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6101 ( .B1(n6138), .B2(n6043), .A(n9380), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6102 ( .B1(n6213), .B2(n6043), .A(n9379), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6103 ( .B1(n6142), .B2(n6043), .A(n9381), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  INV_X16 U6104 ( .A(n6080), .ZN(n6079) );
  INV_X16 U6105 ( .A(n6080), .ZN(n6078) );
  INV_X16 U6106 ( .A(n6045), .ZN(n6043) );
  NAND2_X4 U6107 ( .A1(n9378), .A2(net76270), .ZN(n9383) );
  INV_X16 U6108 ( .A(n6045), .ZN(n6044) );
  MUX2_X2 U6109 ( .A(multOut[10]), .B(n10130), .S(net73585), .Z(n10136) );
  INV_X16 U6110 ( .A(n9383), .ZN(n6045) );
  OAI21_X2 U6112 ( .B1(net76480), .B2(n4801), .A(n9526), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6113 ( .B1(n6142), .B2(n4801), .A(n9525), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6114 ( .B1(n6138), .B2(n6048), .A(n9523), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6115 ( .B1(n6213), .B2(n6048), .A(n9522), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U6116 ( .A1(n5127), .A2(n6088), .B1(net76660), .B2(n6048), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X4 U6119 ( .A1(net76270), .A2(n9520), .ZN(n9528) );
  INV_X16 U6120 ( .A(n9704), .ZN(n9765) );
  NAND2_X4 U6121 ( .A1(net76270), .A2(n9703), .ZN(n9704) );
  OAI21_X2 U6122 ( .B1(n6213), .B2(n6056), .A(n9677), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  INV_X16 U6123 ( .A(n6058), .ZN(n6056) );
  NAND2_X4 U6124 ( .A1(n9674), .A2(net76270), .ZN(n9681) );
  INV_X16 U6125 ( .A(n6058), .ZN(n6057) );
  INV_X16 U6126 ( .A(n9681), .ZN(n6058) );
  OAI21_X2 U6127 ( .B1(n6053), .B2(net76480), .A(n9645), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6128 ( .B1(n6053), .B2(n6138), .A(n9643), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6129 ( .B1(n6053), .B2(n6213), .A(n9642), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6130 ( .B1(n6053), .B2(n6142), .A(n9644), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  INV_X16 U6131 ( .A(n6055), .ZN(n6054) );
  INV_X16 U6132 ( .A(n6055), .ZN(n6053) );
  NAND2_X1 U6133 ( .A1(n6178), .A2(\REGFILE/reg_out[29][3] ), .ZN(n10049) );
  INV_X16 U6134 ( .A(n9646), .ZN(n6055) );
  OAI21_X2 U6135 ( .B1(net76506), .B2(n10563), .A(n10562), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6136 ( .B1(net76506), .B2(n10596), .A(n10595), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6137 ( .B1(net76506), .B2(n10587), .A(n10586), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6138 ( .B1(net76506), .B2(n10584), .A(n10583), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6139 ( .B1(net76506), .B2(n10561), .A(n10560), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6140 ( .B1(net76506), .B2(n10559), .A(n10558), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6141 ( .B1(net76502), .B2(n10636), .A(n10635), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6142 ( .B1(net76502), .B2(n10630), .A(n10629), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6143 ( .B1(net76502), .B2(n10633), .A(n10632), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6144 ( .B1(net76502), .B2(n10639), .A(n10638), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6145 ( .B1(net76502), .B2(n10610), .A(n10609), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6146 ( .B1(net76506), .B2(n10617), .A(n10616), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6147 ( .B1(net76502), .B2(n10590), .A(n10589), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6148 ( .B1(net76506), .B2(n10578), .A(n10577), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6149 ( .B1(net76506), .B2(n10575), .A(n10574), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6150 ( .B1(net76502), .B2(n10628), .A(n10627), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  INV_X2 U6151 ( .A(n9519), .ZN(dmem_addr_out[8]) );
  OAI21_X2 U6152 ( .B1(net76506), .B2(n10572), .A(n10571), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6153 ( .B1(net76506), .B2(n10625), .A(n10624), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6154 ( .B1(net76506), .B2(n10566), .A(n10565), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6155 ( .B1(net76506), .B2(n10622), .A(n10621), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6156 ( .B1(net76506), .B2(n10557), .A(n10556), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6157 ( .B1(net76502), .B2(n10613), .A(n10612), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6158 ( .B1(net76506), .B2(n10554), .A(n10553), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6159 ( .B1(net76506), .B2(n10606), .A(n10605), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6160 ( .B1(net76506), .B2(n10602), .A(n10601), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6161 ( .B1(net76506), .B2(n10599), .A(n10598), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  OAI21_X2 U6162 ( .B1(net76506), .B2(n10551), .A(n10550), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X1 U6163 ( .A1(n4892), .A2(\REGFILE/reg_out[17][0] ), .ZN(n10568) );
  OAI21_X2 U6164 ( .B1(net76502), .B2(n10569), .A(n10568), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X1 U6165 ( .A1(n4867), .A2(\REGFILE/reg_out[0][0] ), .ZN(n10547) );
  OAI21_X2 U6166 ( .B1(net76502), .B2(n10548), .A(n10547), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X1 U6167 ( .A1(\REGFILE/reg_out[3][20] ), .A2(net77422), .ZN(n7392) );
  INV_X8 U6168 ( .A(net77632), .ZN(net77630) );
  AOI22_X2 U6169 ( .A1(\REGFILE/reg_out[26][19] ), .A2(net75439), .B1(
        \REGFILE/reg_out[27][19] ), .B2(net89184), .ZN(n6521) );
  INV_X8 U6170 ( .A(net75441), .ZN(net84760) );
  OAI21_X2 U6171 ( .B1(n6214), .B2(net77116), .A(n10118), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X1 U6172 ( .A1(n5009), .A2(n10947), .ZN(n10217) );
  INV_X16 U6173 ( .A(n5582), .ZN(net77106) );
  NAND2_X4 U6174 ( .A1(\PCLOGIC/imm26_32 [11]), .A2(\PCLOGIC/imm26_32 [12]), 
        .ZN(net80161) );
  AOI21_X4 U6175 ( .B1(net81874), .B2(n4970), .A(net76274), .ZN(n5582) );
  AOI22_X1 U6176 ( .A1(\REGFILE/reg_out[16][6] ), .A2(net77762), .B1(
        \REGFILE/reg_out[15][6] ), .B2(net75468), .ZN(n6770) );
  AOI22_X2 U6177 ( .A1(\REGFILE/reg_out[16][10] ), .A2(net75467), .B1(n5615), 
        .B2(net75468), .ZN(n6694) );
  AOI22_X2 U6178 ( .A1(n4846), .A2(net75467), .B1(net83261), .B2(net75468), 
        .ZN(n5606) );
  NAND2_X1 U6179 ( .A1(net92782), .A2(net81874), .ZN(dmem_addr_out[1]) );
  INV_X4 U6180 ( .A(net77300), .ZN(net93763) );
  NAND2_X1 U6181 ( .A1(\REGFILE/reg_out[2][10] ), .A2(net77342), .ZN(n7828) );
  BUF_X8 U6182 ( .A(n5943), .Z(n5577) );
  INV_X8 U6183 ( .A(net76194), .ZN(net124970) );
  AOI22_X4 U6184 ( .A1(\REGFILE/reg_out[23][15] ), .A2(net77828), .B1(
        \REGFILE/reg_out[22][15] ), .B2(net77836), .ZN(n6586) );
  INV_X4 U6185 ( .A(net77406), .ZN(n5648) );
  NAND3_X2 U6186 ( .A1(\PCLOGIC/imm26_32 [8]), .A2(net73989), .A3(
        \PCLOGIC/imm26_32 [10]), .ZN(n5578) );
  INV_X8 U6187 ( .A(net77776), .ZN(net77774) );
  INV_X8 U6188 ( .A(net72414), .ZN(net36470) );
  AOI22_X4 U6189 ( .A1(\REGFILE/reg_out[29][10] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][10] ), .B2(n5751), .ZN(n6705) );
  AOI22_X2 U6190 ( .A1(\REGFILE/reg_out[30][5] ), .A2(net77634), .B1(
        \REGFILE/reg_out[2][5] ), .B2(net75442), .ZN(n6802) );
  AOI22_X1 U6191 ( .A1(\REGFILE/reg_out[16][30] ), .A2(net77764), .B1(
        \REGFILE/reg_out[15][30] ), .B2(n5579), .ZN(n6257) );
  AOI22_X2 U6192 ( .A1(\REGFILE/reg_out[26][29] ), .A2(net77620), .B1(
        \REGFILE/reg_out[27][29] ), .B2(net77630), .ZN(n6288) );
  AOI22_X2 U6193 ( .A1(\REGFILE/reg_out[17][15] ), .A2(net77796), .B1(
        \REGFILE/reg_out[18][15] ), .B2(n5890), .ZN(n6584) );
  AOI22_X2 U6194 ( .A1(\REGFILE/reg_out[17][18] ), .A2(net77796), .B1(
        \REGFILE/reg_out[18][18] ), .B2(n6896), .ZN(n6530) );
  INV_X4 U6195 ( .A(n10943), .ZN(net75842) );
  AOI22_X4 U6196 ( .A1(\REGFILE/reg_out[7][13] ), .A2(net77714), .B1(
        \REGFILE/reg_out[6][13] ), .B2(net75456), .ZN(n6637) );
  AOI22_X4 U6197 ( .A1(\REGFILE/reg_out[17][10] ), .A2(net77794), .B1(
        \REGFILE/reg_out[18][10] ), .B2(n6896), .ZN(n6688) );
  AOI22_X2 U6198 ( .A1(\REGFILE/reg_out[19][29] ), .A2(net77814), .B1(
        \REGFILE/reg_out[1][29] ), .B2(net82631), .ZN(n6274) );
  NOR2_X2 U6199 ( .A1(n4806), .A2(net76274), .ZN(n10604) );
  INV_X16 U6200 ( .A(n5624), .ZN(net82631) );
  AOI22_X4 U6201 ( .A1(\REGFILE/reg_out[7][14] ), .A2(net77714), .B1(
        \REGFILE/reg_out[6][14] ), .B2(net75456), .ZN(n6621) );
  AOI22_X4 U6202 ( .A1(\REGFILE/reg_out[31][14] ), .A2(net77668), .B1(
        \REGFILE/reg_out[3][14] ), .B2(net77676), .ZN(n6618) );
  AOI22_X4 U6203 ( .A1(\REGFILE/reg_out[4][12] ), .A2(n5678), .B1(
        \REGFILE/reg_out[5][12] ), .B2(net75452), .ZN(n6655) );
  NAND2_X4 U6204 ( .A1(n5631), .A2(net77400), .ZN(net78105) );
  BUF_X32 U6205 ( .A(aluA[31]), .Z(net80189) );
  NAND2_X2 U6206 ( .A1(net71227), .A2(net71228), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U6207 ( .A1(n4877), .A2(\REGFILE/reg_out[1][1] ), .ZN(net71228) );
  NAND2_X1 U6208 ( .A1(net77420), .A2(\REGFILE/reg_out[27][18] ), .ZN(n7450)
         );
  INV_X32 U6209 ( .A(\PCLOGIC/imm26_32 [15]), .ZN(net82738) );
  INV_X8 U6210 ( .A(net77508), .ZN(net77502) );
  INV_X4 U6211 ( .A(net77508), .ZN(net77504) );
  OAI211_X1 U6212 ( .C1(n4865), .C2(net73170), .A(net73496), .B(n8658), .ZN(
        n8870) );
  NAND4_X1 U6213 ( .A1(n4865), .A2(net73503), .A3(n6607), .A4(net73496), .ZN(
        net75793) );
  NAND2_X2 U6214 ( .A1(n4898), .A2(n5581), .ZN(dmem_addr_out[2]) );
  INV_X1 U6215 ( .A(n10115), .ZN(n5581) );
  NAND2_X4 U6216 ( .A1(net75845), .A2(net75846), .ZN(n10943) );
  NOR2_X4 U6217 ( .A1(net75847), .A2(n5583), .ZN(net75846) );
  AOI22_X4 U6218 ( .A1(\REGFILE/reg_out[26][17] ), .A2(net75439), .B1(
        \REGFILE/reg_out[27][17] ), .B2(net75440), .ZN(n5585) );
  INV_X8 U6219 ( .A(net76199), .ZN(net75440) );
  AOI22_X4 U6220 ( .A1(\REGFILE/reg_out[24][17] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][17] ), .B2(net75438), .ZN(n5586) );
  INV_X32 U6221 ( .A(net76197), .ZN(net75437) );
  NAND2_X4 U6222 ( .A1(net84277), .A2(n5576), .ZN(net76197) );
  INV_X8 U6223 ( .A(net87982), .ZN(net84277) );
  AND2_X4 U6224 ( .A1(net91646), .A2(net76204), .ZN(net120684) );
  NAND2_X4 U6225 ( .A1(net84277), .A2(net76204), .ZN(net76233) );
  NAND3_X4 U6226 ( .A1(net92446), .A2(net86794), .A3(net87981), .ZN(net87982)
         );
  INV_X32 U6227 ( .A(\PCLOGIC/imm26_32 [13]), .ZN(net87981) );
  MUX2_X2 U6228 ( .A(net87981), .B(net73529), .S(net73509), .Z(net73527) );
  INV_X32 U6229 ( .A(\PCLOGIC/imm26_32 [14]), .ZN(net82933) );
  NAND3_X4 U6230 ( .A1(net73511), .A2(n4843), .A3(net82598), .ZN(net76239) );
  NAND3_X4 U6231 ( .A1(net73511), .A2(net82933), .A3(net82598), .ZN(net123382)
         );
  AOI21_X1 U6232 ( .B1(net73878), .B2(net86794), .A(net73997), .ZN(net73900)
         );
  INV_X32 U6233 ( .A(\PCLOGIC/imm26_32 [15]), .ZN(net92446) );
  NAND3_X4 U6234 ( .A1(net89734), .A2(net92446), .A3(\PCLOGIC/imm26_32 [14]), 
        .ZN(net90830) );
  NAND2_X4 U6235 ( .A1(net84754), .A2(n5576), .ZN(net76201) );
  INV_X16 U6236 ( .A(net76203), .ZN(net82613) );
  NOR2_X4 U6237 ( .A1(net75857), .A2(net75858), .ZN(net75845) );
  INV_X16 U6238 ( .A(net76236), .ZN(net75468) );
  NAND2_X4 U6239 ( .A1(net148494), .A2(net83408), .ZN(net76236) );
  NAND2_X2 U6240 ( .A1(net76206), .A2(net83408), .ZN(net76241) );
  NAND2_X2 U6241 ( .A1(net87806), .A2(n4797), .ZN(net76222) );
  NAND2_X4 U6242 ( .A1(net82618), .A2(\PCLOGIC/imm26_32 [12]), .ZN(net81601)
         );
  NAND2_X4 U6243 ( .A1(net87820), .A2(\PCLOGIC/imm26_32 [12]), .ZN(net88131)
         );
  INV_X8 U6244 ( .A(net76217), .ZN(net148494) );
  NAND2_X4 U6245 ( .A1(net148494), .A2(net76204), .ZN(net76224) );
  NAND2_X2 U6246 ( .A1(net91643), .A2(net148494), .ZN(net76257) );
  NAND2_X4 U6247 ( .A1(net91643), .A2(net76198), .ZN(net76237) );
  INV_X32 U6248 ( .A(\PCLOGIC/imm26_32 [13]), .ZN(net82598) );
  NAND3_X2 U6249 ( .A1(net82598), .A2(\PCLOGIC/imm26_32 [14]), .A3(
        \PCLOGIC/imm26_32 [15]), .ZN(net85731) );
  AOI21_X1 U6250 ( .B1(net73878), .B2(net73511), .A(net73997), .ZN(net73902)
         );
  INV_X16 U6251 ( .A(net76233), .ZN(net82342) );
  NAND2_X4 U6252 ( .A1(net88253), .A2(net82618), .ZN(net76251) );
  NAND2_X4 U6253 ( .A1(net88253), .A2(n4820), .ZN(net81164) );
  INV_X32 U6254 ( .A(\PCLOGIC/imm26_32 [12]), .ZN(net88253) );
  NAND2_X2 U6255 ( .A1(\REGFILE/reg_out[0][17] ), .A2(net77312), .ZN(net74799)
         );
  NAND2_X2 U6256 ( .A1(\REGFILE/reg_out[10][17] ), .A2(net77348), .ZN(net74808) );
  NAND2_X4 U6257 ( .A1(n5587), .A2(net76202), .ZN(n5588) );
  NAND2_X4 U6258 ( .A1(net76208), .A2(n5587), .ZN(net76234) );
  OAI21_X4 U6259 ( .B1(net75842), .B2(net73697), .A(net75843), .ZN(net36463)
         );
  BUF_X32 U6260 ( .A(net75842), .Z(net148116) );
  INV_X4 U6261 ( .A(net73439), .ZN(net73416) );
  NAND2_X2 U6262 ( .A1(n5591), .A2(net70738), .ZN(n5590) );
  INV_X4 U6263 ( .A(net73780), .ZN(n5591) );
  INV_X4 U6264 ( .A(net73468), .ZN(n5589) );
  NAND2_X2 U6265 ( .A1(net77104), .A2(n4997), .ZN(net71227) );
  INV_X4 U6266 ( .A(net73429), .ZN(net73465) );
  INV_X4 U6267 ( .A(net73443), .ZN(net73427) );
  INV_X16 U6268 ( .A(net77106), .ZN(net77102) );
  NAND2_X2 U6269 ( .A1(net71269), .A2(net76650), .ZN(n5595) );
  INV_X4 U6270 ( .A(net70502), .ZN(net71269) );
  NAND2_X2 U6271 ( .A1(n5592), .A2(net77030), .ZN(n5594) );
  INV_X4 U6272 ( .A(net73771), .ZN(n5592) );
  XNOR2_X2 U6273 ( .A(n5592), .B(net73858), .ZN(net73778) );
  INV_X4 U6274 ( .A(net70504), .ZN(net71266) );
  NOR2_X2 U6275 ( .A1(n5596), .A2(net71302), .ZN(n5593) );
  INV_X4 U6276 ( .A(net70503), .ZN(net71302) );
  INV_X4 U6277 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [17]), .ZN(n5597) );
  OAI211_X2 U6278 ( .C1(net73495), .C2(net73498), .A(net73496), .B(net73504), 
        .ZN(net73500) );
  INV_X4 U6279 ( .A(net73500), .ZN(net73494) );
  NOR2_X2 U6280 ( .A1(n5601), .A2(n5598), .ZN(net92782) );
  NAND2_X1 U6281 ( .A1(net70502), .A2(net70503), .ZN(n5598) );
  AND2_X2 U6282 ( .A1(net70504), .A2(net73585), .ZN(n5601) );
  NAND2_X4 U6283 ( .A1(multOut[1]), .A2(net81873), .ZN(net81874) );
  INV_X4 U6284 ( .A(net73585), .ZN(net81873) );
  NAND2_X2 U6285 ( .A1(net71271), .A2(n5599), .ZN(net70502) );
  XNOR2_X2 U6286 ( .A(net70731), .B(net70735), .ZN(n5599) );
  NAND3_X1 U6287 ( .A1(net71078), .A2(\WIRE_ALU_A/MUX2TO1_32BIT[1].MUX/N1 ), 
        .A3(net36466), .ZN(net70503) );
  INV_X4 U6288 ( .A(net71273), .ZN(\WIRE_ALU_A/MUX2TO1_32BIT[1].MUX/N1 ) );
  NAND3_X2 U6289 ( .A1(net71277), .A2(n5570), .A3(n5600), .ZN(net70504) );
  NOR2_X4 U6290 ( .A1(net71280), .A2(n5039), .ZN(n5600) );
  NAND2_X2 U6291 ( .A1(n5602), .A2(n5603), .ZN(net73585) );
  XNOR2_X2 U6292 ( .A(\PCLOGIC/imm16_32 [27]), .B(\PCLOGIC/imm16_32 [28]), 
        .ZN(n5604) );
  INV_X4 U6293 ( .A(\PCLOGIC/imm16_32 [29]), .ZN(n5605) );
  OAI22_X2 U6294 ( .A1(instructionAddr_out[29]), .A2(n5605), .B1(net73394), 
        .B2(net73938), .ZN(net73400) );
  INV_X16 U6295 ( .A(net73629), .ZN(net74011) );
  INV_X4 U6296 ( .A(net73630), .ZN(net73646) );
  OAI211_X4 U6297 ( .C1(net73532), .C2(net73622), .A(net75792), .B(net75793), 
        .ZN(net75791) );
  INV_X4 U6298 ( .A(net73532), .ZN(net73495) );
  NAND2_X4 U6299 ( .A1(net75748), .A2(net75747), .ZN(dmem_write_out[13]) );
  OAI21_X4 U6300 ( .B1(dmem_write_out[13]), .B2(net75427), .A(n10945), .ZN(
        net72414) );
  NOR2_X4 U6301 ( .A1(net75759), .A2(net75760), .ZN(net75747) );
  NAND4_X2 U6302 ( .A1(net75764), .A2(net75761), .A3(n5606), .A4(net75763), 
        .ZN(net75760) );
  INV_X8 U6303 ( .A(net76234), .ZN(net83167) );
  INV_X2 U6304 ( .A(net84518), .ZN(n5608) );
  INV_X8 U6305 ( .A(net77752), .ZN(net77750) );
  NAND2_X4 U6306 ( .A1(net122022), .A2(net91646), .ZN(net76220) );
  INV_X8 U6307 ( .A(net76254), .ZN(n5607) );
  NAND2_X4 U6308 ( .A1(net76195), .A2(n5607), .ZN(net76199) );
  NAND3_X4 U6309 ( .A1(net73528), .A2(\PCLOGIC/imm26_32 [14]), .A3(
        \PCLOGIC/imm26_32 [15]), .ZN(net76254) );
  INV_X32 U6310 ( .A(\PCLOGIC/imm26_32 [13]), .ZN(net73528) );
  NAND2_X1 U6311 ( .A1(net73878), .A2(net73528), .ZN(net73974) );
  INV_X4 U6312 ( .A(net76262), .ZN(net91643) );
  NAND2_X4 U6313 ( .A1(net91643), .A2(net121496), .ZN(net76258) );
  NAND2_X4 U6314 ( .A1(net73533), .A2(\PCLOGIC/imm26_32 [11]), .ZN(net76262)
         );
  INV_X8 U6315 ( .A(n4823), .ZN(net76238) );
  INV_X16 U6316 ( .A(net75791), .ZN(net75427) );
  INV_X2 U6317 ( .A(net83260), .ZN(net83261) );
  INV_X16 U6318 ( .A(net75481), .ZN(net77848) );
  INV_X8 U6319 ( .A(net77848), .ZN(net77846) );
  INV_X16 U6320 ( .A(n5704), .ZN(n5609) );
  NAND2_X1 U6321 ( .A1(n4888), .A2(\REGFILE/reg_out[22][16] ), .ZN(n9234) );
  AOI22_X4 U6322 ( .A1(\REGFILE/reg_out[17][16] ), .A2(net77796), .B1(
        \REGFILE/reg_out[18][16] ), .B2(n5890), .ZN(n6562) );
  AOI22_X4 U6323 ( .A1(\REGFILE/reg_out[4][16] ), .A2(n5678), .B1(n5756), .B2(
        net75452), .ZN(n6573) );
  INV_X2 U6324 ( .A(n5610), .ZN(n5611) );
  NAND2_X4 U6325 ( .A1(net77460), .A2(\REGFILE/reg_out[21][28] ), .ZN(n7008)
         );
  INV_X2 U6326 ( .A(n5612), .ZN(n5613) );
  OAI21_X2 U6327 ( .B1(n7027), .B2(n7026), .A(n6019), .ZN(n7039) );
  INV_X16 U6328 ( .A(\PCLOGIC/imm26_32 [9]), .ZN(net87097) );
  AOI22_X4 U6329 ( .A1(\REGFILE/reg_out[31][12] ), .A2(net77668), .B1(
        \REGFILE/reg_out[3][12] ), .B2(net77676), .ZN(n6654) );
  AOI22_X4 U6330 ( .A1(\REGFILE/reg_out[23][18] ), .A2(net77828), .B1(
        \REGFILE/reg_out[22][18] ), .B2(net77836), .ZN(n6532) );
  NAND2_X1 U6331 ( .A1(n4889), .A2(\REGFILE/reg_out[6][16] ), .ZN(n9262) );
  INV_X2 U6332 ( .A(n5614), .ZN(n5615) );
  AOI22_X4 U6333 ( .A1(\REGFILE/reg_out[31][10] ), .A2(net77666), .B1(
        \REGFILE/reg_out[3][10] ), .B2(n5609), .ZN(n6698) );
  AOI22_X2 U6334 ( .A1(\REGFILE/reg_out[24][8] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][8] ), .B2(net75438), .ZN(n6746) );
  AOI22_X1 U6335 ( .A1(\REGFILE/reg_out[24][4] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][4] ), .B2(net75438), .ZN(n6822) );
  AOI22_X2 U6336 ( .A1(\REGFILE/reg_out[19][10] ), .A2(net77810), .B1(
        \REGFILE/reg_out[1][10] ), .B2(net75478), .ZN(n6689) );
  AOI22_X2 U6337 ( .A1(\REGFILE/reg_out[24][22] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][22] ), .B2(net124970), .ZN(n6448) );
  AOI22_X2 U6338 ( .A1(\REGFILE/reg_out[0][9] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][9] ), .B2(net75464), .ZN(n6714) );
  INV_X16 U6339 ( .A(net77720), .ZN(net77716) );
  INV_X2 U6340 ( .A(n5617), .ZN(n5618) );
  NAND2_X1 U6341 ( .A1(\REGFILE/reg_out[20][0] ), .A2(net77386), .ZN(n8247) );
  NAND2_X1 U6342 ( .A1(\REGFILE/reg_out[20][1] ), .A2(net77386), .ZN(n8203) );
  NAND2_X1 U6343 ( .A1(\REGFILE/reg_out[28][19] ), .A2(net77386), .ZN(n7405)
         );
  NAND2_X1 U6344 ( .A1(\REGFILE/reg_out[28][20] ), .A2(net77386), .ZN(n7361)
         );
  NAND2_X1 U6345 ( .A1(\REGFILE/reg_out[20][20] ), .A2(net77386), .ZN(n7371)
         );
  NAND2_X1 U6346 ( .A1(\REGFILE/reg_out[12][20] ), .A2(net77386), .ZN(n7381)
         );
  NAND2_X1 U6347 ( .A1(\REGFILE/reg_out[4][20] ), .A2(net77386), .ZN(n7391) );
  NAND2_X1 U6348 ( .A1(\REGFILE/reg_out[28][21] ), .A2(net77386), .ZN(n7312)
         );
  NAND2_X1 U6349 ( .A1(\REGFILE/reg_out[4][21] ), .A2(net77386), .ZN(n7322) );
  NAND2_X1 U6350 ( .A1(\REGFILE/reg_out[12][21] ), .A2(net77386), .ZN(n7332)
         );
  NAND2_X1 U6351 ( .A1(\REGFILE/reg_out[20][21] ), .A2(net77386), .ZN(n7342)
         );
  NAND2_X1 U6352 ( .A1(\REGFILE/reg_out[4][22] ), .A2(net77386), .ZN(n7277) );
  NAND2_X1 U6353 ( .A1(\REGFILE/reg_out[12][22] ), .A2(net77386), .ZN(n7287)
         );
  NAND2_X1 U6354 ( .A1(\REGFILE/reg_out[20][22] ), .A2(net77386), .ZN(n7297)
         );
  NAND2_X1 U6355 ( .A1(net77386), .A2(\REGFILE/reg_out[28][27] ), .ZN(n7048)
         );
  NAND2_X1 U6356 ( .A1(net77386), .A2(\REGFILE/reg_out[12][27] ), .ZN(n7068)
         );
  NAND2_X1 U6357 ( .A1(net77386), .A2(\REGFILE/reg_out[4][27] ), .ZN(n7078) );
  NAND2_X1 U6358 ( .A1(net77386), .A2(\REGFILE/reg_out[12][28] ), .ZN(n7024)
         );
  INV_X16 U6359 ( .A(net77320), .ZN(net77318) );
  INV_X16 U6360 ( .A(n5703), .ZN(net77668) );
  INV_X16 U6361 ( .A(n5703), .ZN(net77666) );
  INV_X16 U6362 ( .A(n5703), .ZN(net77670) );
  NAND2_X1 U6363 ( .A1(\REGFILE/reg_out[5][18] ), .A2(net77456), .ZN(n7473) );
  AOI22_X2 U6364 ( .A1(\REGFILE/reg_out[4][18] ), .A2(net75451), .B1(
        \REGFILE/reg_out[5][18] ), .B2(net75452), .ZN(n6541) );
  AOI22_X4 U6365 ( .A1(\REGFILE/reg_out[9][16] ), .A2(net77700), .B1(n5668), 
        .B2(net75454), .ZN(n6574) );
  INV_X8 U6366 ( .A(net76239), .ZN(net91646) );
  AOI22_X2 U6367 ( .A1(\REGFILE/reg_out[9][13] ), .A2(net77700), .B1(n5716), 
        .B2(net75454), .ZN(n6636) );
  AOI22_X4 U6368 ( .A1(\REGFILE/reg_out[7][17] ), .A2(net77714), .B1(
        \REGFILE/reg_out[6][17] ), .B2(net75456), .ZN(n6561) );
  INV_X4 U6369 ( .A(net148735), .ZN(net148736) );
  NAND2_X1 U6370 ( .A1(n4891), .A2(\REGFILE/reg_out[16][13] ), .ZN(n9441) );
  NAND2_X1 U6371 ( .A1(net77308), .A2(\REGFILE/reg_out[16][13] ), .ZN(n7675)
         );
  BUF_X32 U6372 ( .A(net73851), .Z(n5619) );
  OAI22_X1 U6373 ( .A1(net78235), .A2(n6090), .B1(n6191), .B2(net76658), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X1 U6374 ( .A1(\REGFILE/reg_out[1][16] ), .A2(net77526), .ZN(n7561) );
  INV_X32 U6375 ( .A(net77800), .ZN(net77796) );
  INV_X16 U6376 ( .A(n6224), .ZN(n6896) );
  AOI22_X4 U6377 ( .A1(\REGFILE/reg_out[29][17] ), .A2(net77652), .B1(
        \REGFILE/reg_out[28][17] ), .B2(n5751), .ZN(net75849) );
  AOI22_X4 U6378 ( .A1(\REGFILE/reg_out[11][10] ), .A2(net77746), .B1(n4817), 
        .B2(net75466), .ZN(n6693) );
  NOR2_X4 U6379 ( .A1(n6453), .A2(n6452), .ZN(n6454) );
  NAND2_X1 U6381 ( .A1(\REGFILE/reg_out[28][12] ), .A2(n6177), .ZN(n9154) );
  NAND2_X1 U6382 ( .A1(\REGFILE/reg_out[28][12] ), .A2(net77380), .ZN(n7711)
         );
  NAND4_X2 U6383 ( .A1(n6924), .A2(n6923), .A3(n6921), .A4(n6922), .ZN(
        net73851) );
  NAND2_X1 U6384 ( .A1(\REGFILE/reg_out[18][16] ), .A2(net77346), .ZN(n7544)
         );
  INV_X8 U6385 ( .A(net77704), .ZN(net77702) );
  INV_X16 U6386 ( .A(net77704), .ZN(net77698) );
  INV_X16 U6387 ( .A(net75453), .ZN(net77704) );
  NAND2_X1 U6388 ( .A1(net77550), .A2(\REGFILE/reg_out[30][28] ), .ZN(n7001)
         );
  NAND2_X1 U6389 ( .A1(net77550), .A2(\REGFILE/reg_out[22][28] ), .ZN(n7011)
         );
  NAND2_X1 U6390 ( .A1(net77550), .A2(\REGFILE/reg_out[6][28] ), .ZN(n7031) );
  INV_X16 U6391 ( .A(net77848), .ZN(net77844) );
  INV_X16 U6392 ( .A(net77848), .ZN(net77842) );
  AOI22_X2 U6393 ( .A1(\REGFILE/reg_out[11][17] ), .A2(net77748), .B1(
        \REGFILE/reg_out[12][17] ), .B2(net75466), .ZN(net75861) );
  INV_X4 U6394 ( .A(n10378), .ZN(n10914) );
  NAND2_X4 U6395 ( .A1(n6551), .A2(n6550), .ZN(dmem_write_out[18]) );
  AOI22_X1 U6396 ( .A1(\REGFILE/reg_out[0][3] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][3] ), .B2(net75464), .ZN(n6834) );
  NAND2_X1 U6397 ( .A1(\REGFILE/reg_out[28][11] ), .A2(n6175), .ZN(n9909) );
  NAND2_X1 U6398 ( .A1(\REGFILE/reg_out[28][11] ), .A2(net77380), .ZN(n7755)
         );
  AOI22_X2 U6399 ( .A1(\REGFILE/reg_out[29][11] ), .A2(net77652), .B1(
        \REGFILE/reg_out[28][11] ), .B2(n5751), .ZN(n6683) );
  AOI22_X4 U6400 ( .A1(\REGFILE/reg_out[23][10] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][10] ), .B2(net77834), .ZN(n6690) );
  NAND2_X1 U6401 ( .A1(\REGFILE/reg_out[13][10] ), .A2(net77456), .ZN(n7813)
         );
  NAND2_X1 U6402 ( .A1(\REGFILE/reg_out[6][16] ), .A2(net77562), .ZN(n7562) );
  NAND2_X1 U6403 ( .A1(\REGFILE/reg_out[2][3] ), .A2(net77338), .ZN(n8134) );
  AOI22_X2 U6404 ( .A1(\REGFILE/reg_out[14][23] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][23] ), .B2(n6009), .ZN(n6418) );
  AOI22_X2 U6405 ( .A1(\REGFILE/reg_out[14][8] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][8] ), .B2(n6009), .ZN(n6739) );
  AOI22_X2 U6406 ( .A1(\REGFILE/reg_out[23][3] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][3] ), .B2(net77834), .ZN(n6832) );
  NAND2_X1 U6407 ( .A1(\REGFILE/reg_out[12][12] ), .A2(n4873), .ZN(n9120) );
  NAND2_X1 U6408 ( .A1(net77380), .A2(\REGFILE/reg_out[12][12] ), .ZN(n7731)
         );
  NAND3_X4 U6409 ( .A1(net92447), .A2(net82932), .A3(\PCLOGIC/imm26_32 [13]), 
        .ZN(net148091) );
  NAND2_X1 U6410 ( .A1(n4804), .A2(\REGFILE/reg_out[15][12] ), .ZN(n9126) );
  NAND2_X1 U6411 ( .A1(\REGFILE/reg_out[15][12] ), .A2(net77488), .ZN(n7726)
         );
  AOI22_X4 U6412 ( .A1(\REGFILE/reg_out[11][16] ), .A2(net77748), .B1(n5618), 
        .B2(net83168), .ZN(n6567) );
  INV_X16 U6413 ( .A(n5623), .ZN(net75478) );
  NAND2_X4 U6414 ( .A1(net76204), .A2(net87806), .ZN(n5623) );
  INV_X8 U6415 ( .A(net88102), .ZN(net87806) );
  NAND2_X4 U6416 ( .A1(net76238), .A2(net87806), .ZN(net76249) );
  NAND3_X4 U6417 ( .A1(net89734), .A2(n4840), .A3(\PCLOGIC/imm26_32 [15]), 
        .ZN(net88102) );
  INV_X32 U6418 ( .A(\PCLOGIC/imm26_32 [14]), .ZN(net82932) );
  INV_X16 U6419 ( .A(\PCLOGIC/imm26_32 [13]), .ZN(net89734) );
  INV_X16 U6420 ( .A(net75477), .ZN(net77816) );
  INV_X16 U6421 ( .A(net77816), .ZN(net77810) );
  INV_X8 U6422 ( .A(net76253), .ZN(net75477) );
  OR2_X2 U6423 ( .A1(n5578), .A2(net80211), .ZN(net78104) );
  AND2_X4 U6424 ( .A1(net78104), .A2(net78105), .ZN(net75415) );
  NAND3_X4 U6425 ( .A1(\PCLOGIC/imm26_32 [8]), .A2(net73989), .A3(
        \PCLOGIC/imm26_32 [10]), .ZN(net75423) );
  OAI22_X2 U6426 ( .A1(net78108), .A2(net77464), .B1(net78109), .B2(net75422), 
        .ZN(net78107) );
  INV_X16 U6427 ( .A(net75423), .ZN(net77474) );
  INV_X32 U6428 ( .A(\PCLOGIC/imm26_32 [9]), .ZN(net73989) );
  NAND2_X2 U6429 ( .A1(net105318), .A2(net70497), .ZN(dmem_addr_out[0]) );
  INV_X4 U6430 ( .A(net70689), .ZN(net70497) );
  NAND2_X2 U6431 ( .A1(net70685), .A2(net70497), .ZN(net70687) );
  OAI22_X2 U6432 ( .A1(net70690), .A2(net70691), .B1(net81873), .B2(net70692), 
        .ZN(net70689) );
  INV_X4 U6433 ( .A(net105376), .ZN(net70692) );
  AOI22_X2 U6434 ( .A1(net70692), .A2(net70684), .B1(net70685), .B2(n4915), 
        .ZN(net70541) );
  XNOR2_X2 U6435 ( .A(n5625), .B(n5626), .ZN(net70690) );
  INV_X4 U6436 ( .A(net70730), .ZN(n5626) );
  NAND2_X2 U6437 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[1].MUX/N1 ), .A2(net70734), 
        .ZN(n5627) );
  INV_X4 U6438 ( .A(net70735), .ZN(net70732) );
  XNOR2_X2 U6439 ( .A(net70729), .B(net71027), .ZN(n5625) );
  XNOR2_X2 U6440 ( .A(net77042), .B(net70535), .ZN(net70729) );
  NAND4_X2 U6441 ( .A1(net73611), .A2(net73612), .A3(net73613), .A4(n5629), 
        .ZN(n5628) );
  NOR3_X4 U6442 ( .A1(net73615), .A2(net73616), .A3(n5630), .ZN(n5629) );
  NOR3_X4 U6443 ( .A1(n4971), .A2(net73619), .A3(net73620), .ZN(n5630) );
  INV_X4 U6444 ( .A(\PCLOGIC/imm16_32 [30]), .ZN(net73619) );
  INV_X16 U6445 ( .A(net75422), .ZN(net77400) );
  INV_X2 U6446 ( .A(net80440), .ZN(n5631) );
  NAND3_X4 U6447 ( .A1(net73987), .A2(net87097), .A3(\PCLOGIC/imm26_32 [8]), 
        .ZN(net75422) );
  NAND2_X2 U6448 ( .A1(net73878), .A2(net87097), .ZN(net73988) );
  INV_X32 U6449 ( .A(\PCLOGIC/imm26_32 [10]), .ZN(net73987) );
  NOR2_X4 U6450 ( .A1(multOut[0]), .A2(net70687), .ZN(net70537) );
  NOR2_X4 U6451 ( .A1(n5634), .A2(n5635), .ZN(n5636) );
  INV_X4 U6452 ( .A(net70693), .ZN(n5635) );
  INV_X4 U6453 ( .A(net73585), .ZN(net76452) );
  NOR2_X4 U6454 ( .A1(n9854), .A2(net70718), .ZN(n5638) );
  NOR2_X4 U6455 ( .A1(net70709), .A2(net70710), .ZN(n5634) );
  INV_X4 U6456 ( .A(n5632), .ZN(n5637) );
  AOI21_X4 U6457 ( .B1(net105352), .B2(n5633), .A(n9606), .ZN(n5632) );
  NAND2_X2 U6458 ( .A1(net70713), .A2(net78051), .ZN(n5633) );
  INV_X4 U6459 ( .A(net36414), .ZN(net78050) );
  OAI21_X2 U6460 ( .B1(net76154), .B2(net78056), .A(n5639), .ZN(net36414) );
  INV_X8 U6461 ( .A(n5640), .ZN(net75844) );
  NAND2_X2 U6462 ( .A1(net77272), .A2(net78055), .ZN(n5640) );
  INV_X32 U6463 ( .A(net77280), .ZN(net77272) );
  INV_X16 U6464 ( .A(net73665), .ZN(net77280) );
  NOR2_X4 U6465 ( .A1(net77280), .A2(net73908), .ZN(net75792) );
  NAND2_X4 U6466 ( .A1(net76181), .A2(n5641), .ZN(net73665) );
  NOR3_X4 U6467 ( .A1(net74029), .A2(instruction[1]), .A3(instruction[0]), 
        .ZN(n5641) );
  NAND3_X4 U6468 ( .A1(net75397), .A2(net75395), .A3(net75396), .ZN(aluA[31])
         );
  AOI22_X4 U6469 ( .A1(net77276), .A2(\PCLOGIC/imm16_32 [30]), .B1(net73831), 
        .B2(n4963), .ZN(net75367) );
  NOR2_X4 U6470 ( .A1(n5643), .A2(net73503), .ZN(net76181) );
  NAND2_X4 U6471 ( .A1(instruction[3]), .A2(instruction[4]), .ZN(n5643) );
  INV_X32 U6472 ( .A(instruction[5]), .ZN(net73503) );
  INV_X32 U6473 ( .A(n5644), .ZN(net77588) );
  INV_X4 U6474 ( .A(net73836), .ZN(n5642) );
  AOI22_X4 U6475 ( .A1(net77276), .A2(\PCLOGIC/imm16_32 [31]), .B1(net73849), 
        .B2(n4897), .ZN(net75395) );
  NAND2_X4 U6476 ( .A1(net73837), .A2(n4897), .ZN(net75368) );
  INV_X32 U6477 ( .A(net77296), .ZN(net77290) );
  BUF_X32 U6478 ( .A(net73849), .Z(net80390) );
  INV_X4 U6479 ( .A(net78126), .ZN(net75414) );
  OAI22_X2 U6480 ( .A1(net78127), .A2(net77512), .B1(net78128), .B2(net75424), 
        .ZN(net78126) );
  INV_X32 U6481 ( .A(net77512), .ZN(net77508) );
  INV_X8 U6482 ( .A(net75425), .ZN(net74050) );
  INV_X4 U6483 ( .A(net82513), .ZN(net75416) );
  INV_X32 U6484 ( .A(n5647), .ZN(net77406) );
  INV_X8 U6485 ( .A(n5645), .ZN(n5647) );
  NAND3_X4 U6486 ( .A1(\PCLOGIC/imm26_32 [10]), .A2(net123931), .A3(
        \PCLOGIC/imm26_32 [9]), .ZN(n5646) );
  INV_X32 U6487 ( .A(\PCLOGIC/imm26_32 [8]), .ZN(net123931) );
  NAND3_X4 U6488 ( .A1(net123931), .A2(net73987), .A3(\PCLOGIC/imm26_32 [9]), 
        .ZN(net85371) );
  AOI22_X4 U6489 ( .A1(net82500), .A2(net77514), .B1(net80443), .B2(net77298), 
        .ZN(net75417) );
  INV_X16 U6490 ( .A(net77326), .ZN(net77298) );
  INV_X16 U6491 ( .A(net77328), .ZN(net77326) );
  INV_X16 U6492 ( .A(net77326), .ZN(net77300) );
  NAND2_X2 U6494 ( .A1(net76238), .A2(net84754), .ZN(n6224) );
  NAND2_X1 U6495 ( .A1(net77562), .A2(\REGFILE/reg_out[14][27] ), .ZN(n7065)
         );
  NAND2_X1 U6496 ( .A1(\REGFILE/reg_out[30][0] ), .A2(net77550), .ZN(n8234) );
  NAND2_X1 U6497 ( .A1(\REGFILE/reg_out[30][1] ), .A2(net77554), .ZN(n8190) );
  NAND2_X1 U6498 ( .A1(\REGFILE/reg_out[14][1] ), .A2(net77554), .ZN(n8210) );
  NAND2_X1 U6499 ( .A1(net77550), .A2(\REGFILE/reg_out[6][27] ), .ZN(n7075) );
  NAND2_X1 U6500 ( .A1(net77550), .A2(\REGFILE/reg_out[14][28] ), .ZN(n7021)
         );
  NAND2_X1 U6501 ( .A1(\REGFILE/reg_out[22][1] ), .A2(net77550), .ZN(n8200) );
  NAND2_X1 U6502 ( .A1(\REGFILE/reg_out[22][0] ), .A2(net77550), .ZN(n8244) );
  NAND2_X1 U6503 ( .A1(\REGFILE/reg_out[14][0] ), .A2(net77550), .ZN(n8254) );
  NAND2_X1 U6504 ( .A1(\REGFILE/reg_out[6][1] ), .A2(net77554), .ZN(n8220) );
  NAND2_X1 U6505 ( .A1(net77550), .A2(\REGFILE/reg_out[30][27] ), .ZN(n7045)
         );
  NAND4_X2 U6506 ( .A1(n6973), .A2(n6972), .A3(n6971), .A4(n6970), .ZN(n6974)
         );
  AOI22_X2 U6507 ( .A1(n5789), .A2(net77478), .B1(n5896), .B2(net77550), .ZN(
        n6927) );
  AOI22_X2 U6508 ( .A1(\REGFILE/reg_out[23][31] ), .A2(net77478), .B1(n5718), 
        .B2(net77550), .ZN(n6924) );
  AOI22_X2 U6509 ( .A1(n5795), .A2(net77478), .B1(n5926), .B2(net77550), .ZN(
        n6945) );
  INV_X16 U6510 ( .A(net77428), .ZN(net77422) );
  INV_X16 U6511 ( .A(net77400), .ZN(net77392) );
  INV_X16 U6512 ( .A(net77394), .ZN(net77382) );
  NOR2_X2 U6513 ( .A1(n5988), .A2(net77392), .ZN(n5754) );
  INV_X16 U6514 ( .A(\PCLOGIC/imm26_32 [13]), .ZN(net87495) );
  INV_X32 U6515 ( .A(net77720), .ZN(net77714) );
  NOR2_X2 U6516 ( .A1(n6751), .A2(n6750), .ZN(n6752) );
  INV_X16 U6517 ( .A(net77430), .ZN(net77424) );
  NAND2_X4 U6518 ( .A1(net88253), .A2(net87820), .ZN(n5706) );
  AOI22_X2 U6519 ( .A1(\REGFILE/reg_out[11][11] ), .A2(net77748), .B1(n5872), 
        .B2(net83168), .ZN(n6671) );
  NAND2_X4 U6520 ( .A1(net84754), .A2(net76238), .ZN(n5649) );
  AOI22_X1 U6521 ( .A1(\REGFILE/reg_out[0][4] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][4] ), .B2(net75464), .ZN(n6812) );
  NAND4_X2 U6522 ( .A1(n6393), .A2(n6394), .A3(n6395), .A4(n6392), .ZN(n6396)
         );
  INV_X4 U6523 ( .A(net77616), .ZN(net77614) );
  OAI21_X1 U6524 ( .B1(n6529), .B2(net78055), .A(n6528), .ZN(n5650) );
  OAI21_X1 U6525 ( .B1(dmem_write_out[27]), .B2(net78056), .A(n6343), .ZN(
        n5652) );
  OAI21_X2 U6526 ( .B1(n10355), .B2(n10354), .A(n10353), .ZN(n10358) );
  AOI22_X4 U6527 ( .A1(\REGFILE/reg_out[4][11] ), .A2(n5679), .B1(
        \REGFILE/reg_out[5][11] ), .B2(net84475), .ZN(n6677) );
  NAND2_X1 U6528 ( .A1(\REGFILE/reg_out[16][15] ), .A2(net77310), .ZN(n7587)
         );
  AOI22_X2 U6529 ( .A1(\REGFILE/reg_out[29][25] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][25] ), .B2(n6911), .ZN(n6385) );
  AOI22_X1 U6530 ( .A1(\REGFILE/reg_out[24][3] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][3] ), .B2(net75438), .ZN(n6844) );
  OAI211_X4 U6531 ( .C1(n10045), .C2(net76646), .A(net70740), .B(n10044), .ZN(
        n10046) );
  AOI22_X2 U6532 ( .A1(\REGFILE/reg_out[11][22] ), .A2(net77750), .B1(
        \REGFILE/reg_out[12][22] ), .B2(net75466), .ZN(n6439) );
  AOI22_X1 U6533 ( .A1(\REGFILE/reg_out[11][4] ), .A2(net77746), .B1(
        \REGFILE/reg_out[12][4] ), .B2(net75466), .ZN(n6813) );
  AOI22_X1 U6534 ( .A1(\REGFILE/reg_out[30][26] ), .A2(net77638), .B1(
        \REGFILE/reg_out[2][26] ), .B2(net75442), .ZN(n6360) );
  AOI22_X1 U6535 ( .A1(\REGFILE/reg_out[30][2] ), .A2(net77634), .B1(
        \REGFILE/reg_out[2][2] ), .B2(net75442), .ZN(n6868) );
  INV_X32 U6536 ( .A(\PCLOGIC/imm26_32 [8]), .ZN(net123932) );
  AOI22_X4 U6538 ( .A1(\REGFILE/reg_out[31][11] ), .A2(net77668), .B1(
        \REGFILE/reg_out[3][11] ), .B2(net77676), .ZN(n6676) );
  NAND2_X1 U6539 ( .A1(\REGFILE/reg_out[5][15] ), .A2(net77454), .ZN(n7603) );
  AOI22_X2 U6540 ( .A1(\REGFILE/reg_out[4][15] ), .A2(net75451), .B1(
        \REGFILE/reg_out[5][15] ), .B2(net84475), .ZN(n6595) );
  NAND2_X1 U6541 ( .A1(net73878), .A2(net90864), .ZN(n8380) );
  NAND2_X2 U6542 ( .A1(\REGFILE/reg_out[7][30] ), .A2(net77478), .ZN(n5654) );
  NAND2_X2 U6543 ( .A1(\REGFILE/reg_out[6][30] ), .A2(net77550), .ZN(n5655) );
  INV_X16 U6544 ( .A(net77506), .ZN(net77478) );
  NAND2_X1 U6545 ( .A1(net77298), .A2(\REGFILE/reg_out[24][28] ), .ZN(n7002)
         );
  NAND2_X1 U6548 ( .A1(\REGFILE/reg_out[27][17] ), .A2(net77420), .ZN(n7494)
         );
  INV_X8 U6549 ( .A(net76256), .ZN(net76206) );
  AOI22_X1 U6550 ( .A1(\REGFILE/reg_out[19][3] ), .A2(net77810), .B1(
        \REGFILE/reg_out[1][3] ), .B2(net75478), .ZN(n6831) );
  AOI22_X1 U6551 ( .A1(\REGFILE/reg_out[19][25] ), .A2(net77814), .B1(
        \REGFILE/reg_out[1][25] ), .B2(net75478), .ZN(n6369) );
  INV_X16 U6552 ( .A(net77832), .ZN(net77826) );
  NAND2_X1 U6553 ( .A1(\REGFILE/reg_out[29][0] ), .A2(net77444), .ZN(n8231) );
  NAND2_X1 U6554 ( .A1(\REGFILE/reg_out[21][0] ), .A2(net77444), .ZN(n8241) );
  NAND2_X1 U6555 ( .A1(\REGFILE/reg_out[13][0] ), .A2(net77444), .ZN(n8251) );
  NAND2_X1 U6556 ( .A1(\REGFILE/reg_out[29][1] ), .A2(net77444), .ZN(n8187) );
  NAND2_X1 U6557 ( .A1(\REGFILE/reg_out[21][1] ), .A2(net77444), .ZN(n8197) );
  NAND2_X1 U6558 ( .A1(\REGFILE/reg_out[13][1] ), .A2(net77444), .ZN(n8207) );
  NAND2_X1 U6559 ( .A1(\REGFILE/reg_out[5][1] ), .A2(net77444), .ZN(n8217) );
  NAND2_X1 U6560 ( .A1(net77444), .A2(\REGFILE/reg_out[29][27] ), .ZN(n7042)
         );
  NAND2_X1 U6561 ( .A1(net77444), .A2(\REGFILE/reg_out[13][27] ), .ZN(n7062)
         );
  NAND2_X1 U6562 ( .A1(net77444), .A2(\REGFILE/reg_out[5][27] ), .ZN(n7072) );
  NAND2_X1 U6563 ( .A1(net77444), .A2(\REGFILE/reg_out[13][28] ), .ZN(n7018)
         );
  BUF_X32 U6564 ( .A(n5851), .Z(n5931) );
  INV_X16 U6565 ( .A(net77800), .ZN(net77798) );
  AOI22_X4 U6566 ( .A1(\REGFILE/reg_out[9][15] ), .A2(net77700), .B1(
        \REGFILE/reg_out[8][15] ), .B2(n4829), .ZN(n6596) );
  INV_X32 U6567 ( .A(net77856), .ZN(net77852) );
  AOI22_X4 U6568 ( .A1(\REGFILE/reg_out[7][16] ), .A2(net77714), .B1(n4860), 
        .B2(net75456), .ZN(n6575) );
  NAND2_X1 U6569 ( .A1(net77382), .A2(\REGFILE/reg_out[12][16] ), .ZN(n7555)
         );
  AOI22_X1 U6570 ( .A1(\REGFILE/reg_out[7][4] ), .A2(net75455), .B1(
        \REGFILE/reg_out[6][4] ), .B2(net75456), .ZN(n6821) );
  AOI22_X1 U6571 ( .A1(\REGFILE/reg_out[7][5] ), .A2(net75455), .B1(
        \REGFILE/reg_out[6][5] ), .B2(net75456), .ZN(n6799) );
  INV_X1 U6572 ( .A(n4864), .ZN(n5805) );
  INV_X4 U6573 ( .A(dmem_write_out[24]), .ZN(n6410) );
  INV_X4 U6574 ( .A(net77324), .ZN(net77312) );
  INV_X4 U6575 ( .A(net77324), .ZN(net77310) );
  INV_X4 U6576 ( .A(net77324), .ZN(net77308) );
  AOI22_X2 U6577 ( .A1(\REGFILE/reg_out[17][24] ), .A2(net77798), .B1(
        \REGFILE/reg_out[18][24] ), .B2(n5890), .ZN(net76034) );
  AOI22_X4 U6578 ( .A1(\REGFILE/reg_out[29][18] ), .A2(net77652), .B1(
        \REGFILE/reg_out[28][18] ), .B2(n5751), .ZN(n6547) );
  NAND2_X2 U6579 ( .A1(\PCLOGIC/imm16_32 [28]), .A2(net77276), .ZN(n5658) );
  NAND2_X4 U6580 ( .A1(n5657), .A2(n5658), .ZN(aluA[28]) );
  INV_X8 U6581 ( .A(net77464), .ZN(net77460) );
  BUF_X8 U6582 ( .A(net36470), .Z(net85047) );
  INV_X4 U6583 ( .A(n10909), .ZN(n5659) );
  OAI22_X4 U6584 ( .A1(n5823), .A2(net86238), .B1(n5999), .B2(net93763), .ZN(
        n5822) );
  AOI22_X4 U6585 ( .A1(\REGFILE/reg_out[9][18] ), .A2(net77700), .B1(
        \REGFILE/reg_out[8][18] ), .B2(n4829), .ZN(n6542) );
  AOI22_X4 U6586 ( .A1(\REGFILE/reg_out[9][14] ), .A2(net77700), .B1(
        \REGFILE/reg_out[8][14] ), .B2(net75454), .ZN(n6620) );
  NAND2_X2 U6587 ( .A1(n6807), .A2(n6806), .ZN(dmem_write_out[5]) );
  AOI22_X2 U6588 ( .A1(\REGFILE/reg_out[11][5] ), .A2(net77746), .B1(
        \REGFILE/reg_out[12][5] ), .B2(net75466), .ZN(n6791) );
  NAND2_X1 U6589 ( .A1(n5902), .A2(net75464), .ZN(n5946) );
  AOI22_X2 U6590 ( .A1(\REGFILE/reg_out[0][14] ), .A2(net82342), .B1(n5829), 
        .B2(net83203), .ZN(n6612) );
  INV_X8 U6591 ( .A(net77324), .ZN(net77306) );
  INV_X8 U6592 ( .A(net77324), .ZN(net77304) );
  INV_X8 U6593 ( .A(net77324), .ZN(net77302) );
  AOI22_X4 U6594 ( .A1(\REGFILE/reg_out[9][17] ), .A2(net77700), .B1(
        \REGFILE/reg_out[8][17] ), .B2(net75454), .ZN(n6560) );
  AOI21_X1 U6595 ( .B1(n10418), .B2(n10384), .A(n10383), .ZN(n10388) );
  INV_X16 U6596 ( .A(n6010), .ZN(n5663) );
  INV_X8 U6597 ( .A(n6010), .ZN(n6009) );
  AOI22_X2 U6598 ( .A1(\REGFILE/reg_out[11][9] ), .A2(net77746), .B1(
        \REGFILE/reg_out[12][9] ), .B2(net75466), .ZN(n6715) );
  NAND2_X4 U6599 ( .A1(\REGFILE/reg_out[4][29] ), .A2(net77386), .ZN(n6961) );
  INV_X2 U6600 ( .A(n5665), .ZN(n5666) );
  INV_X2 U6601 ( .A(n5667), .ZN(n5668) );
  NAND2_X1 U6602 ( .A1(net73708), .A2(n6007), .ZN(n8694) );
  NAND2_X1 U6603 ( .A1(n10542), .A2(n6007), .ZN(n8766) );
  AOI22_X1 U6604 ( .A1(n9297), .A2(net72962), .B1(n4912), .B2(n6007), .ZN(
        n9769) );
  NAND2_X1 U6605 ( .A1(net70720), .A2(n6007), .ZN(n9081) );
  NAND2_X1 U6606 ( .A1(n9065), .A2(n6007), .ZN(n8837) );
  NAND2_X1 U6607 ( .A1(net70719), .A2(n6007), .ZN(n9943) );
  NAND2_X1 U6608 ( .A1(n6040), .A2(n6007), .ZN(n8711) );
  NAND2_X1 U6609 ( .A1(n6007), .A2(n10315), .ZN(n10316) );
  AOI21_X1 U6610 ( .B1(n8593), .B2(n6007), .A(n8592), .ZN(n8884) );
  XNOR2_X1 U6611 ( .A(n8591), .B(n6007), .ZN(n8773) );
  INV_X1 U6612 ( .A(n6007), .ZN(n8638) );
  NAND3_X2 U6613 ( .A1(n8694), .A2(n8693), .A3(n8692), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  NOR2_X2 U6614 ( .A1(n9769), .A2(n9770), .ZN(n8983) );
  OAI22_X1 U6615 ( .A1(n9771), .A2(n9770), .B1(n9769), .B2(n9802), .ZN(n9772)
         );
  NAND3_X2 U6616 ( .A1(n9081), .A2(n9080), .A3(n9079), .ZN(n9621) );
  NAND3_X2 U6617 ( .A1(n9944), .A2(n9943), .A3(n9942), .ZN(n10541) );
  OAI21_X2 U6618 ( .B1(n8884), .B2(n8883), .A(n8595), .ZN(n9776) );
  NOR2_X2 U6619 ( .A1(n6428), .A2(n6429), .ZN(n6430) );
  INV_X8 U6620 ( .A(net76259), .ZN(net121496) );
  INV_X4 U6621 ( .A(net148091), .ZN(net76208) );
  AOI22_X4 U6622 ( .A1(\REGFILE/reg_out[17][13] ), .A2(net77796), .B1(
        \REGFILE/reg_out[18][13] ), .B2(n6896), .ZN(n6630) );
  INV_X4 U6623 ( .A(n10392), .ZN(n10911) );
  NAND2_X2 U6624 ( .A1(\REGFILE/reg_out[15][6] ), .A2(net77484), .ZN(n7988) );
  AND2_X2 U6625 ( .A1(\REGFILE/reg_out[11][24] ), .A2(net77750), .ZN(n5669) );
  AND2_X2 U6626 ( .A1(\REGFILE/reg_out[12][24] ), .A2(net75466), .ZN(n5670) );
  NOR2_X2 U6627 ( .A1(n5669), .A2(n5670), .ZN(n6393) );
  INV_X2 U6628 ( .A(n5671), .ZN(n5672) );
  INV_X2 U6629 ( .A(n5673), .ZN(n5674) );
  AOI22_X2 U6630 ( .A1(\REGFILE/reg_out[24][13] ), .A2(net75437), .B1(n5940), 
        .B2(net124970), .ZN(n6638) );
  INV_X8 U6631 ( .A(net76255), .ZN(net77834) );
  AOI22_X1 U6632 ( .A1(\REGFILE/reg_out[9][28] ), .A2(net77702), .B1(
        \REGFILE/reg_out[8][28] ), .B2(n4829), .ZN(n6309) );
  AOI22_X2 U6633 ( .A1(\REGFILE/reg_out[16][15] ), .A2(net75467), .B1(n5782), 
        .B2(net75468), .ZN(n6590) );
  AOI22_X2 U6634 ( .A1(\REGFILE/reg_out[26][22] ), .A2(net75439), .B1(
        \REGFILE/reg_out[27][22] ), .B2(net89184), .ZN(n6449) );
  BUF_X16 U6635 ( .A(n10385), .Z(n5758) );
  NAND2_X2 U6636 ( .A1(\REGFILE/reg_out[6][7] ), .A2(net75456), .ZN(n5698) );
  OAI21_X1 U6637 ( .B1(n4819), .B2(net73697), .A(n6504), .ZN(n5675) );
  NAND2_X1 U6638 ( .A1(\REGFILE/reg_out[3][15] ), .A2(net77418), .ZN(n7610) );
  AOI22_X2 U6639 ( .A1(\REGFILE/reg_out[31][15] ), .A2(net77668), .B1(
        \REGFILE/reg_out[3][15] ), .B2(net77676), .ZN(n6594) );
  INV_X2 U6640 ( .A(n5676), .ZN(n5677) );
  AOI22_X2 U6641 ( .A1(\REGFILE/reg_out[7][24] ), .A2(net77716), .B1(
        \REGFILE/reg_out[6][24] ), .B2(net75456), .ZN(n6400) );
  NOR2_X2 U6642 ( .A1(n6827), .A2(n6826), .ZN(n6828) );
  NAND3_X1 U6643 ( .A1(net71078), .A2(n6007), .A3(n10926), .ZN(n8776) );
  XNOR2_X1 U6644 ( .A(n6007), .B(n10926), .ZN(n10441) );
  INV_X2 U6645 ( .A(n10926), .ZN(n10315) );
  NOR2_X4 U6646 ( .A1(n6539), .A2(n6538), .ZN(n6551) );
  NOR2_X4 U6647 ( .A1(n6549), .A2(n6548), .ZN(n6550) );
  AOI22_X1 U6648 ( .A1(\REGFILE/reg_out[4][26] ), .A2(n5678), .B1(
        \REGFILE/reg_out[5][26] ), .B2(net75452), .ZN(n6355) );
  AOI22_X2 U6649 ( .A1(\REGFILE/reg_out[4][14] ), .A2(n5678), .B1(
        \REGFILE/reg_out[5][14] ), .B2(net84475), .ZN(n6619) );
  NAND2_X4 U6650 ( .A1(net76206), .A2(net76195), .ZN(net76205) );
  AOI22_X2 U6651 ( .A1(\REGFILE/reg_out[29][19] ), .A2(net77652), .B1(
        \REGFILE/reg_out[28][19] ), .B2(n5751), .ZN(n6523) );
  INV_X8 U6652 ( .A(net76219), .ZN(n5678) );
  INV_X8 U6653 ( .A(net76219), .ZN(n5679) );
  INV_X8 U6654 ( .A(net76219), .ZN(net75451) );
  INV_X16 U6655 ( .A(n6239), .ZN(n6911) );
  NAND2_X1 U6656 ( .A1(net77346), .A2(\REGFILE/reg_out[2][15] ), .ZN(n7608) );
  NAND2_X1 U6657 ( .A1(n4804), .A2(\REGFILE/reg_out[15][16] ), .ZN(n9218) );
  OAI21_X4 U6658 ( .B1(n7037), .B2(n7036), .A(net77290), .ZN(n7038) );
  AOI22_X2 U6659 ( .A1(\REGFILE/reg_out[17][5] ), .A2(net77794), .B1(
        \REGFILE/reg_out[18][5] ), .B2(n5890), .ZN(n6786) );
  AOI22_X4 U6660 ( .A1(\REGFILE/reg_out[16][20] ), .A2(net77762), .B1(
        \REGFILE/reg_out[15][20] ), .B2(n5579), .ZN(n6488) );
  NAND2_X1 U6661 ( .A1(\REGFILE/reg_out[12][19] ), .A2(net77384), .ZN(n7425)
         );
  AOI22_X2 U6662 ( .A1(\REGFILE/reg_out[11][19] ), .A2(net77748), .B1(
        \REGFILE/reg_out[12][19] ), .B2(net83168), .ZN(n6511) );
  AOI22_X1 U6663 ( .A1(\REGFILE/reg_out[11][23] ), .A2(net77750), .B1(
        \REGFILE/reg_out[12][23] ), .B2(net83168), .ZN(n6416) );
  AOI22_X2 U6664 ( .A1(\REGFILE/reg_out[26][8] ), .A2(net75439), .B1(
        \REGFILE/reg_out[27][8] ), .B2(net89184), .ZN(n6747) );
  AOI22_X1 U6665 ( .A1(\REGFILE/reg_out[24][23] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][23] ), .B2(net124970), .ZN(n6425) );
  NAND2_X1 U6666 ( .A1(net77526), .A2(\REGFILE/reg_out[25][15] ), .ZN(n7575)
         );
  INV_X16 U6667 ( .A(n6006), .ZN(n6007) );
  AOI22_X1 U6668 ( .A1(\REGFILE/reg_out[30][4] ), .A2(net77634), .B1(
        \REGFILE/reg_out[2][4] ), .B2(net75442), .ZN(n6824) );
  INV_X2 U6669 ( .A(n5857), .ZN(n5684) );
  NAND2_X4 U6670 ( .A1(n10215), .A2(n10214), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  INV_X16 U6671 ( .A(net77784), .ZN(net77778) );
  AOI22_X4 U6672 ( .A1(\REGFILE/reg_out[11][15] ), .A2(net77748), .B1(n4854), 
        .B2(net83167), .ZN(n6589) );
  AOI22_X2 U6673 ( .A1(\REGFILE/reg_out[16][19] ), .A2(net77762), .B1(
        \REGFILE/reg_out[15][19] ), .B2(net75468), .ZN(n6512) );
  AOI22_X4 U6674 ( .A1(\REGFILE/reg_out[9][8] ), .A2(net77698), .B1(
        \REGFILE/reg_out[8][8] ), .B2(n4829), .ZN(n6744) );
  INV_X2 U6675 ( .A(n5686), .ZN(n5687) );
  AOI22_X2 U6676 ( .A1(\REGFILE/reg_out[0][25] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][25] ), .B2(net81764), .ZN(n6372) );
  INV_X16 U6677 ( .A(net77800), .ZN(net77794) );
  NOR2_X2 U6678 ( .A1(net91561), .A2(n5754), .ZN(n5753) );
  NAND2_X2 U6680 ( .A1(net76488), .A2(\REGFILE/reg_out[31][2] ), .ZN(n5690) );
  INV_X16 U6681 ( .A(n5696), .ZN(net77116) );
  INV_X16 U6682 ( .A(n5696), .ZN(net77114) );
  NAND2_X4 U6683 ( .A1(n5691), .A2(reset), .ZN(n5689) );
  OAI211_X4 U6684 ( .C1(net71394), .C2(net76646), .A(net70740), .B(n5692), 
        .ZN(n5691) );
  INV_X4 U6685 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [18]), .ZN(n5694) );
  AND2_X2 U6686 ( .A1(net80797), .A2(n5698), .ZN(net75623) );
  NAND2_X4 U6687 ( .A1(net76206), .A2(net83210), .ZN(n5697) );
  INV_X8 U6688 ( .A(net81164), .ZN(net83210) );
  NAND2_X4 U6689 ( .A1(net83210), .A2(net76202), .ZN(net76203) );
  NAND2_X4 U6690 ( .A1(net121496), .A2(net83210), .ZN(net76219) );
  NAND2_X4 U6691 ( .A1(net76238), .A2(net76206), .ZN(net76255) );
  NAND3_X4 U6692 ( .A1(net82738), .A2(\PCLOGIC/imm26_32 [14]), .A3(
        \PCLOGIC/imm26_32 [13]), .ZN(net76256) );
  MUX2_X2 U6693 ( .A(net82738), .B(net73512), .S(net73509), .Z(net73510) );
  NAND2_X1 U6694 ( .A1(\REGFILE/reg_out[7][7] ), .A2(net75455), .ZN(net80797)
         );
  INV_X8 U6695 ( .A(net76224), .ZN(net75455) );
  NAND2_X2 U6696 ( .A1(\REGFILE/reg_out[6][7] ), .A2(net77556), .ZN(net74359)
         );
  NAND2_X2 U6697 ( .A1(n4889), .A2(\REGFILE/reg_out[6][7] ), .ZN(net71936) );
  NAND2_X2 U6698 ( .A1(\REGFILE/reg_out[7][7] ), .A2(net77484), .ZN(net74361)
         );
  NAND2_X2 U6699 ( .A1(n4886), .A2(\REGFILE/reg_out[7][7] ), .ZN(net71934) );
  NAND2_X4 U6700 ( .A1(net75615), .A2(net75616), .ZN(dmem_write_out[7]) );
  OAI21_X4 U6701 ( .B1(dmem_write_out[7]), .B2(net75427), .A(n10945), .ZN(
        net72015) );
  NOR2_X4 U6702 ( .A1(net75617), .A2(net75618), .ZN(net75616) );
  NAND4_X2 U6703 ( .A1(net75619), .A2(net75620), .A3(net75621), .A4(n5699), 
        .ZN(net75618) );
  AOI22_X2 U6704 ( .A1(\REGFILE/reg_out[24][7] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][7] ), .B2(net124970), .ZN(n5699) );
  NAND2_X4 U6705 ( .A1(net76196), .A2(n5576), .ZN(net76194) );
  AOI22_X2 U6706 ( .A1(\REGFILE/reg_out[26][23] ), .A2(net77618), .B1(
        \REGFILE/reg_out[27][23] ), .B2(net77630), .ZN(net75995) );
  INV_X8 U6707 ( .A(net72015), .ZN(net36479) );
  AOI22_X2 U6708 ( .A1(\REGFILE/reg_out[31][7] ), .A2(net77666), .B1(
        \REGFILE/reg_out[3][7] ), .B2(n5609), .ZN(net75626) );
  INV_X32 U6709 ( .A(n5704), .ZN(net77676) );
  INV_X8 U6710 ( .A(n5705), .ZN(n5704) );
  NOR2_X4 U6711 ( .A1(net85731), .A2(n5706), .ZN(n5705) );
  INV_X8 U6712 ( .A(n5700), .ZN(n5703) );
  NOR2_X4 U6713 ( .A1(n4844), .A2(net87489), .ZN(n5700) );
  AOI22_X2 U6714 ( .A1(\REGFILE/reg_out[4][7] ), .A2(n5678), .B1(
        \REGFILE/reg_out[5][7] ), .B2(net84475), .ZN(net75625) );
  INV_X16 U6715 ( .A(n5702), .ZN(net84475) );
  NAND2_X4 U6716 ( .A1(net76204), .A2(n5701), .ZN(n5702) );
  INV_X8 U6717 ( .A(n4821), .ZN(n5701) );
  NAND2_X2 U6718 ( .A1(net76204), .A2(n5701), .ZN(net91311) );
  NAND2_X2 U6719 ( .A1(n5701), .A2(net76195), .ZN(net76209) );
  NAND2_X2 U6720 ( .A1(net76238), .A2(n5701), .ZN(net76260) );
  INV_X4 U6721 ( .A(net70868), .ZN(net70720) );
  INV_X4 U6722 ( .A(net72163), .ZN(net70697) );
  INV_X4 U6723 ( .A(net71027), .ZN(net36488) );
  INV_X4 U6724 ( .A(net71300), .ZN(net70696) );
  NAND2_X2 U6725 ( .A1(n5707), .A2(net73543), .ZN(net78014) );
  INV_X4 U6726 ( .A(aluA[16]), .ZN(n5708) );
  INV_X4 U6727 ( .A(net70706), .ZN(net105349) );
  AOI21_X4 U6728 ( .B1(n5709), .B2(net105360), .A(net70714), .ZN(net105352) );
  INV_X4 U6729 ( .A(net70845), .ZN(n5707) );
  INV_X4 U6730 ( .A(net70703), .ZN(n5710) );
  INV_X4 U6731 ( .A(net78014), .ZN(net70701) );
  NAND2_X2 U6732 ( .A1(net70719), .A2(net36391), .ZN(n5711) );
  OAI211_X2 U6733 ( .C1(net70868), .C2(n5708), .A(n5711), .B(net70717), .ZN(
        n5709) );
  NAND2_X1 U6734 ( .A1(\REGFILE/reg_out[12][15] ), .A2(net77382), .ZN(n7599)
         );
  NAND2_X1 U6735 ( .A1(\REGFILE/reg_out[26][13] ), .A2(net77344), .ZN(n7666)
         );
  NAND2_X1 U6736 ( .A1(n4893), .A2(\REGFILE/reg_out[26][13] ), .ZN(n9463) );
  AOI22_X2 U6737 ( .A1(\REGFILE/reg_out[26][13] ), .A2(net75439), .B1(n5938), 
        .B2(net75440), .ZN(n6639) );
  INV_X1 U6738 ( .A(n4828), .ZN(n5713) );
  NAND2_X4 U6739 ( .A1(n9637), .A2(net76270), .ZN(n9646) );
  OAI211_X4 U6740 ( .C1(n9636), .C2(net76646), .A(net70740), .B(n9635), .ZN(
        n9637) );
  INV_X2 U6741 ( .A(n5715), .ZN(n5716) );
  AOI22_X1 U6742 ( .A1(\REGFILE/reg_out[9][1] ), .A2(net77698), .B1(
        \REGFILE/reg_out[8][1] ), .B2(n4829), .ZN(n6886) );
  AOI22_X1 U6743 ( .A1(\REGFILE/reg_out[9][3] ), .A2(net77698), .B1(
        \REGFILE/reg_out[8][3] ), .B2(n4829), .ZN(n6842) );
  AOI22_X1 U6744 ( .A1(\REGFILE/reg_out[9][0] ), .A2(net77698), .B1(
        \REGFILE/reg_out[8][0] ), .B2(n4829), .ZN(n6909) );
  AOI22_X1 U6745 ( .A1(\REGFILE/reg_out[9][2] ), .A2(net77698), .B1(
        \REGFILE/reg_out[8][2] ), .B2(n4829), .ZN(n6864) );
  AOI22_X1 U6746 ( .A1(\REGFILE/reg_out[9][26] ), .A2(net77702), .B1(
        \REGFILE/reg_out[8][26] ), .B2(n4829), .ZN(n6356) );
  AOI22_X1 U6747 ( .A1(\REGFILE/reg_out[9][29] ), .A2(net77702), .B1(
        \REGFILE/reg_out[8][29] ), .B2(n4829), .ZN(n6285) );
  AOI22_X1 U6748 ( .A1(\REGFILE/reg_out[9][25] ), .A2(net77702), .B1(
        \REGFILE/reg_out[8][25] ), .B2(n4829), .ZN(n6380) );
  AOI22_X2 U6749 ( .A1(\REGFILE/reg_out[0][24] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][24] ), .B2(net75464), .ZN(n6392) );
  INV_X2 U6750 ( .A(n8810), .ZN(n8599) );
  NAND2_X1 U6751 ( .A1(net36391), .A2(n10331), .ZN(n10332) );
  NOR3_X1 U6752 ( .A1(n10331), .A2(net72312), .A3(net78003), .ZN(n8644) );
  XNOR2_X1 U6753 ( .A(net36391), .B(n8599), .ZN(n8808) );
  NOR3_X2 U6754 ( .A1(n8646), .A2(n8645), .A3(n8644), .ZN(n8647) );
  INV_X1 U6755 ( .A(n10430), .ZN(n8601) );
  NAND2_X2 U6757 ( .A1(net77422), .A2(\REGFILE/reg_out[27][20] ), .ZN(n7362)
         );
  AOI22_X2 U6758 ( .A1(\REGFILE/reg_out[31][13] ), .A2(net77668), .B1(n5802), 
        .B2(net77676), .ZN(n6634) );
  OAI21_X4 U6759 ( .B1(n6553), .B2(net78056), .A(n6552), .ZN(n5759) );
  INV_X2 U6760 ( .A(n5717), .ZN(n5718) );
  INV_X8 U6761 ( .A(net90830), .ZN(net84754) );
  AOI22_X4 U6762 ( .A1(\REGFILE/reg_out[17][17] ), .A2(net77796), .B1(
        \REGFILE/reg_out[18][17] ), .B2(n6896), .ZN(n6554) );
  AOI22_X1 U6763 ( .A1(\REGFILE/reg_out[29][31] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][31] ), .B2(n6911), .ZN(n6243) );
  AOI22_X1 U6764 ( .A1(\REGFILE/reg_out[29][0] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][0] ), .B2(n6911), .ZN(n6915) );
  AOI22_X1 U6765 ( .A1(\REGFILE/reg_out[29][30] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][30] ), .B2(n6911), .ZN(n6268) );
  AOI22_X1 U6766 ( .A1(\REGFILE/reg_out[29][28] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][28] ), .B2(n6911), .ZN(n6314) );
  AOI22_X1 U6767 ( .A1(\REGFILE/reg_out[29][26] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][26] ), .B2(n6911), .ZN(n6361) );
  AOI22_X1 U6768 ( .A1(\REGFILE/reg_out[29][27] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][27] ), .B2(n6911), .ZN(n6338) );
  AOI22_X1 U6769 ( .A1(\REGFILE/reg_out[29][3] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][3] ), .B2(n6911), .ZN(n6847) );
  INV_X2 U6770 ( .A(n5719), .ZN(n5720) );
  NAND2_X1 U6771 ( .A1(\REGFILE/reg_out[10][19] ), .A2(net77348), .ZN(n7424)
         );
  AOI22_X2 U6772 ( .A1(\REGFILE/reg_out[19][2] ), .A2(net77810), .B1(
        \REGFILE/reg_out[1][2] ), .B2(net82631), .ZN(n6853) );
  AOI22_X2 U6773 ( .A1(\REGFILE/reg_out[16][11] ), .A2(net75467), .B1(n5909), 
        .B2(net75468), .ZN(n6672) );
  NAND2_X1 U6774 ( .A1(\REGFILE/reg_out[18][15] ), .A2(net77346), .ZN(n7588)
         );
  NAND2_X1 U6775 ( .A1(\REGFILE/reg_out[22][15] ), .A2(net77562), .ZN(n7586)
         );
  OAI21_X2 U6776 ( .B1(n10403), .B2(n10402), .A(n10401), .ZN(n10406) );
  NAND2_X4 U6777 ( .A1(\REGFILE/reg_out[27][29] ), .A2(net77426), .ZN(n6986)
         );
  AOI21_X2 U6778 ( .B1(n10391), .B2(n10390), .A(n10389), .ZN(n10395) );
  OAI21_X1 U6779 ( .B1(n9692), .B2(n9854), .A(n9691), .ZN(n9693) );
  NOR2_X2 U6780 ( .A1(n9694), .A2(n9693), .ZN(n9695) );
  AOI22_X2 U6781 ( .A1(\REGFILE/reg_out[4][4] ), .A2(net75451), .B1(
        \REGFILE/reg_out[5][4] ), .B2(net75452), .ZN(n6819) );
  AOI22_X2 U6782 ( .A1(\REGFILE/reg_out[16][25] ), .A2(net75467), .B1(
        \REGFILE/reg_out[15][25] ), .B2(net77774), .ZN(n6374) );
  AOI22_X1 U6783 ( .A1(\REGFILE/reg_out[11][25] ), .A2(net77750), .B1(
        \REGFILE/reg_out[12][25] ), .B2(net75466), .ZN(n6373) );
  AOI22_X2 U6784 ( .A1(\REGFILE/reg_out[11][8] ), .A2(net77746), .B1(n5951), 
        .B2(net75466), .ZN(n6737) );
  NAND2_X1 U6785 ( .A1(\REGFILE/reg_out[6][13] ), .A2(net77560), .ZN(n7694) );
  NAND2_X1 U6786 ( .A1(net77308), .A2(\REGFILE/reg_out[8][13] ), .ZN(n7685) );
  NAND2_X4 U6787 ( .A1(net77100), .A2(n10607), .ZN(n10209) );
  NAND2_X4 U6788 ( .A1(net77102), .A2(n10614), .ZN(n10213) );
  INV_X16 U6789 ( .A(n10052), .ZN(n6074) );
  NAND4_X1 U6790 ( .A1(n6996), .A2(n4858), .A3(n6997), .A4(n6995), .ZN(n5748)
         );
  OR2_X4 U6791 ( .A1(n10115), .A2(n5571), .ZN(n5749) );
  OAI22_X2 U6792 ( .A1(n10114), .A2(net70691), .B1(n10113), .B2(n10408), .ZN(
        n10115) );
  NAND2_X4 U6793 ( .A1(net77104), .A2(net70574), .ZN(n10215) );
  NAND2_X4 U6794 ( .A1(n10213), .A2(n10212), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X4 U6795 ( .A1(n10209), .A2(n10208), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  INV_X16 U6796 ( .A(n6069), .ZN(n6067) );
  INV_X16 U6797 ( .A(n6069), .ZN(n6068) );
  INV_X1 U6798 ( .A(n9967), .ZN(dmem_addr_out[4]) );
  INV_X32 U6799 ( .A(\PCLOGIC/imm26_32 [15]), .ZN(net92447) );
  INV_X16 U6800 ( .A(net77392), .ZN(net77388) );
  NAND2_X2 U6801 ( .A1(net77478), .A2(\REGFILE/reg_out[7][28] ), .ZN(n7029) );
  INV_X4 U6802 ( .A(net73585), .ZN(net92392) );
  INV_X8 U6803 ( .A(n6239), .ZN(n5751) );
  OAI21_X1 U6804 ( .B1(dmem_write_out[3]), .B2(net75427), .A(n10945), .ZN(
        n5752) );
  INV_X2 U6805 ( .A(n5755), .ZN(n5756) );
  NAND2_X1 U6806 ( .A1(\REGFILE/reg_out[3][16] ), .A2(n4871), .ZN(n9256) );
  AOI22_X2 U6807 ( .A1(\REGFILE/reg_out[23][5] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][5] ), .B2(net77834), .ZN(n6788) );
  AOI22_X4 U6808 ( .A1(n5812), .A2(net77452), .B1(n5894), .B2(net77388), .ZN(
        n6926) );
  INV_X8 U6809 ( .A(net91311), .ZN(net75452) );
  BUF_X4 U6810 ( .A(n10392), .Z(n5757) );
  AOI22_X4 U6811 ( .A1(\REGFILE/reg_out[31][16] ), .A2(net77668), .B1(n5677), 
        .B2(net77676), .ZN(n6572) );
  AOI22_X1 U6812 ( .A1(\REGFILE/reg_out[23][4] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][4] ), .B2(net77834), .ZN(n6810) );
  AOI22_X2 U6813 ( .A1(\REGFILE/reg_out[23][0] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][0] ), .B2(net77834), .ZN(n6899) );
  AOI22_X2 U6814 ( .A1(\REGFILE/reg_out[23][6] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][6] ), .B2(net77834), .ZN(n6766) );
  AOI22_X2 U6815 ( .A1(\REGFILE/reg_out[7][6] ), .A2(net77714), .B1(
        \REGFILE/reg_out[6][6] ), .B2(net75456), .ZN(n6777) );
  AOI22_X2 U6816 ( .A1(\REGFILE/reg_out[7][21] ), .A2(net77714), .B1(
        \REGFILE/reg_out[6][21] ), .B2(net75456), .ZN(n6471) );
  AOI22_X1 U6817 ( .A1(\REGFILE/reg_out[7][1] ), .A2(net75455), .B1(
        \REGFILE/reg_out[6][1] ), .B2(net75456), .ZN(n6887) );
  AOI22_X4 U6818 ( .A1(n5960), .A2(net77406), .B1(n5997), .B2(n6014), .ZN(
        n6947) );
  AOI22_X1 U6819 ( .A1(\REGFILE/reg_out[11][2] ), .A2(net77746), .B1(
        \REGFILE/reg_out[12][2] ), .B2(net83168), .ZN(n6857) );
  NAND4_X2 U6820 ( .A1(n6673), .A2(n6671), .A3(n6670), .A4(n6672), .ZN(n6674)
         );
  AOI22_X2 U6821 ( .A1(\REGFILE/reg_out[4][20] ), .A2(n5679), .B1(
        \REGFILE/reg_out[5][20] ), .B2(net84475), .ZN(n6493) );
  AOI22_X2 U6822 ( .A1(\REGFILE/reg_out[4][8] ), .A2(net75451), .B1(n5687), 
        .B2(net84475), .ZN(n6743) );
  AOI22_X4 U6823 ( .A1(\REGFILE/reg_out[29][9] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][9] ), .B2(n5751), .ZN(n6727) );
  NAND2_X4 U6824 ( .A1(\PCLOGIC/imm26_32 [11]), .A2(\PCLOGIC/imm26_32 [12]), 
        .ZN(net87489) );
  INV_X8 U6825 ( .A(aluA[27]), .ZN(n5760) );
  INV_X16 U6826 ( .A(n5760), .ZN(n5761) );
  OAI21_X4 U6827 ( .B1(n6974), .B2(n6975), .A(n6019), .ZN(n6996) );
  INV_X16 U6828 ( .A(net74051), .ZN(net77548) );
  INV_X16 U6829 ( .A(net77542), .ZN(net77516) );
  INV_X32 U6830 ( .A(\PCLOGIC/imm26_32 [8]), .ZN(net90864) );
  AOI22_X4 U6831 ( .A1(\REGFILE/reg_out[4][17] ), .A2(net75451), .B1(
        \REGFILE/reg_out[5][17] ), .B2(net75452), .ZN(n6559) );
  AOI22_X4 U6832 ( .A1(n5796), .A2(net77406), .B1(n5972), .B2(n6014), .ZN(
        n6935) );
  NOR2_X2 U6835 ( .A1(n6260), .A2(n6259), .ZN(n6272) );
  INV_X2 U6836 ( .A(n5765), .ZN(n5766) );
  AOI22_X2 U6837 ( .A1(\REGFILE/reg_out[24][16] ), .A2(net75437), .B1(n5613), 
        .B2(net124970), .ZN(n6576) );
  INV_X1 U6838 ( .A(n10420), .ZN(n9836) );
  NAND4_X2 U6839 ( .A1(n6591), .A2(n6589), .A3(n6588), .A4(n6590), .ZN(n6592)
         );
  AOI22_X2 U6840 ( .A1(\REGFILE/reg_out[19][14] ), .A2(net77812), .B1(
        \REGFILE/reg_out[1][14] ), .B2(net75478), .ZN(n6609) );
  AOI22_X2 U6841 ( .A1(\REGFILE/reg_out[19][11] ), .A2(net77812), .B1(
        \REGFILE/reg_out[1][11] ), .B2(net75478), .ZN(n6667) );
  INV_X2 U6842 ( .A(n5767), .ZN(n5768) );
  NAND2_X1 U6843 ( .A1(\REGFILE/reg_out[1][13] ), .A2(net77524), .ZN(n7693) );
  NAND2_X1 U6844 ( .A1(n4877), .A2(\REGFILE/reg_out[1][13] ), .ZN(n9449) );
  OAI21_X2 U6845 ( .B1(n9100), .B2(n9854), .A(n9099), .ZN(n9101) );
  INV_X2 U6846 ( .A(n5847), .ZN(n5769) );
  NOR2_X2 U6847 ( .A1(n10447), .A2(net78014), .ZN(n9181) );
  INV_X2 U6848 ( .A(n9054), .ZN(n9055) );
  XNOR2_X1 U6849 ( .A(n9054), .B(aluA[16]), .ZN(n9178) );
  OAI21_X2 U6850 ( .B1(n9196), .B2(n9854), .A(n9195), .ZN(n9197) );
  XNOR2_X1 U6851 ( .A(n10930), .B(n8989), .ZN(n10435) );
  XNOR2_X1 U6852 ( .A(n10930), .B(n4808), .ZN(n8988) );
  NOR3_X2 U6853 ( .A1(n10437), .A2(n10436), .A3(n10435), .ZN(n10438) );
  NAND2_X1 U6854 ( .A1(net70701), .A2(n10435), .ZN(n8991) );
  AOI21_X2 U6855 ( .B1(net71271), .B2(n8993), .A(n8992), .ZN(n8995) );
  NAND2_X1 U6856 ( .A1(n8816), .A2(aluA[20]), .ZN(n8817) );
  NOR3_X2 U6857 ( .A1(n10451), .A2(n10450), .A3(n10449), .ZN(n10452) );
  AOI21_X2 U6858 ( .B1(net71271), .B2(n10056), .A(n10055), .ZN(n10077) );
  NOR3_X2 U6859 ( .A1(n10074), .A2(n10073), .A3(n10072), .ZN(n10075) );
  AOI22_X2 U6860 ( .A1(\REGFILE/reg_out[26][30] ), .A2(net77620), .B1(
        \REGFILE/reg_out[27][30] ), .B2(net77630), .ZN(n6266) );
  INV_X8 U6861 ( .A(net76199), .ZN(net89184) );
  INV_X1 U6862 ( .A(n10922), .ZN(n9306) );
  AOI22_X4 U6863 ( .A1(\REGFILE/reg_out[21][13] ), .A2(net77844), .B1(n5720), 
        .B2(net77852), .ZN(n6633) );
  NAND2_X4 U6864 ( .A1(instruction[5]), .A2(net73170), .ZN(net73532) );
  NAND2_X1 U6865 ( .A1(n4966), .A2(net73170), .ZN(net73780) );
  INV_X32 U6866 ( .A(instruction[3]), .ZN(net73170) );
  INV_X4 U6867 ( .A(n8410), .ZN(n5815) );
  INV_X8 U6868 ( .A(n10036), .ZN(n10908) );
  AOI22_X2 U6869 ( .A1(\REGFILE/reg_out[11][3] ), .A2(net77746), .B1(
        \REGFILE/reg_out[12][3] ), .B2(net83167), .ZN(n6835) );
  AOI22_X1 U6870 ( .A1(\REGFILE/reg_out[30][25] ), .A2(net77638), .B1(
        \REGFILE/reg_out[2][25] ), .B2(net75442), .ZN(n6384) );
  NAND2_X1 U6871 ( .A1(\REGFILE/reg_out[0][14] ), .A2(net77310), .ZN(n7651) );
  NAND2_X1 U6872 ( .A1(\REGFILE/reg_out[12][16] ), .A2(n4873), .ZN(n9212) );
  INV_X2 U6873 ( .A(n5771), .ZN(n5772) );
  AOI22_X2 U6874 ( .A1(\REGFILE/reg_out[26][15] ), .A2(net75439), .B1(n4839), 
        .B2(net75440), .ZN(n6599) );
  NAND4_X2 U6875 ( .A1(n6945), .A2(n6942), .A3(n6944), .A4(n6943), .ZN(n8410)
         );
  AOI22_X1 U6876 ( .A1(\REGFILE/reg_out[23][31] ), .A2(net77828), .B1(
        \REGFILE/reg_out[22][31] ), .B2(net77836), .ZN(n6227) );
  AOI22_X2 U6877 ( .A1(n5825), .A2(net77406), .B1(n5828), .B2(n6014), .ZN(
        n6925) );
  INV_X32 U6878 ( .A(\PCLOGIC/imm26_32 [14]), .ZN(net86794) );
  NOR2_X4 U6879 ( .A1(n6763), .A2(n6762), .ZN(net75615) );
  NAND2_X4 U6880 ( .A1(\REGFILE/reg_out[25][29] ), .A2(net77514), .ZN(n6984)
         );
  INV_X2 U6881 ( .A(n5776), .ZN(n5777) );
  INV_X2 U6882 ( .A(n5778), .ZN(n5779) );
  INV_X2 U6883 ( .A(n5780), .ZN(n5781) );
  NAND4_X2 U6884 ( .A1(n6547), .A2(n6546), .A3(n6544), .A4(n6545), .ZN(n6548)
         );
  NOR2_X4 U6885 ( .A1(n6580), .A2(n6581), .ZN(n6582) );
  OAI22_X1 U6886 ( .A1(n9961), .A2(net70691), .B1(n9960), .B2(n5659), .ZN(
        n9962) );
  XNOR2_X1 U6887 ( .A(n5659), .B(net77040), .ZN(n10033) );
  NAND2_X1 U6888 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[4].MUX/N1 ), .A2(n5659), .ZN(
        n10401) );
  XNOR2_X1 U6889 ( .A(n5659), .B(n9954), .ZN(n10306) );
  INV_X8 U6890 ( .A(net76203), .ZN(net75442) );
  AOI22_X2 U6891 ( .A1(\REGFILE/reg_out[26][2] ), .A2(net77620), .B1(
        \REGFILE/reg_out[27][2] ), .B2(net77630), .ZN(n6867) );
  AOI22_X2 U6892 ( .A1(\REGFILE/reg_out[17][19] ), .A2(net77796), .B1(
        \REGFILE/reg_out[18][19] ), .B2(n6896), .ZN(n6506) );
  NAND2_X1 U6893 ( .A1(net77298), .A2(\REGFILE/reg_out[16][27] ), .ZN(n7056)
         );
  AOI22_X2 U6894 ( .A1(n5793), .A2(net77514), .B1(n5892), .B2(net77298), .ZN(
        n6928) );
  NOR2_X4 U6896 ( .A1(n6729), .A2(n6728), .ZN(n6730) );
  AOI22_X2 U6897 ( .A1(\REGFILE/reg_out[16][21] ), .A2(net87506), .B1(
        \REGFILE/reg_out[15][21] ), .B2(n5579), .ZN(n6464) );
  AOI22_X1 U6898 ( .A1(\REGFILE/reg_out[16][28] ), .A2(net87506), .B1(
        \REGFILE/reg_out[15][28] ), .B2(n5579), .ZN(n6303) );
  AOI22_X2 U6899 ( .A1(\REGFILE/reg_out[0][16] ), .A2(net82342), .B1(n5772), 
        .B2(net83203), .ZN(n6566) );
  NAND2_X2 U6900 ( .A1(n6431), .A2(n6430), .ZN(dmem_write_out[23]) );
  AOI22_X2 U6901 ( .A1(\REGFILE/reg_out[26][3] ), .A2(net77620), .B1(
        \REGFILE/reg_out[27][3] ), .B2(net77630), .ZN(n6845) );
  INV_X2 U6902 ( .A(n5866), .ZN(n5782) );
  OAI21_X1 U6903 ( .B1(n6481), .B2(net78056), .A(n6480), .ZN(n5783) );
  NAND2_X1 U6904 ( .A1(\REGFILE/reg_out[18][13] ), .A2(net77344), .ZN(n7676)
         );
  NAND2_X1 U6905 ( .A1(\REGFILE/reg_out[10][22] ), .A2(n6015), .ZN(n7286) );
  INV_X1 U6906 ( .A(n10923), .ZN(n10331) );
  INV_X4 U6907 ( .A(net77624), .ZN(net77618) );
  INV_X8 U6908 ( .A(n5931), .ZN(n5870) );
  OAI21_X2 U6909 ( .B1(n7538), .B2(n7537), .A(n6012), .ZN(n7572) );
  INV_X2 U6910 ( .A(n5786), .ZN(n5787) );
  OAI22_X2 U6911 ( .A1(n5948), .A2(net77506), .B1(n5949), .B2(net75424), .ZN(
        n5947) );
  NAND2_X4 U6912 ( .A1(n5916), .A2(n6929), .ZN(n8403) );
  INV_X4 U6913 ( .A(net77608), .ZN(net77602) );
  AOI22_X2 U6914 ( .A1(\REGFILE/reg_out[26][21] ), .A2(net75439), .B1(
        \REGFILE/reg_out[27][21] ), .B2(net89184), .ZN(n6473) );
  INV_X2 U6915 ( .A(n5788), .ZN(n5789) );
  INV_X2 U6916 ( .A(n5790), .ZN(n5791) );
  NOR2_X1 U6917 ( .A1(net73850), .A2(net73836), .ZN(n8406) );
  INV_X2 U6918 ( .A(n5792), .ZN(n5793) );
  INV_X1 U6919 ( .A(n5672), .ZN(n10936) );
  INV_X2 U6920 ( .A(n5794), .ZN(n5795) );
  OAI21_X2 U6921 ( .B1(n6223), .B2(net76480), .A(n8755), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U6922 ( .A(n5898), .ZN(n5796) );
  AND2_X2 U6923 ( .A1(n5899), .A2(n5900), .ZN(n5797) );
  NAND2_X2 U6924 ( .A1(\PCLOGIC/imm16_32 [29]), .A2(net77276), .ZN(n5900) );
  AOI22_X2 U6925 ( .A1(\REGFILE/reg_out[17][11] ), .A2(net77796), .B1(
        \REGFILE/reg_out[18][11] ), .B2(n6896), .ZN(n6666) );
  AOI22_X1 U6926 ( .A1(\REGFILE/reg_out[7][25] ), .A2(net77714), .B1(
        \REGFILE/reg_out[6][25] ), .B2(net75456), .ZN(n6381) );
  NOR2_X2 U6927 ( .A1(n6467), .A2(n6466), .ZN(n6479) );
  AOI22_X2 U6928 ( .A1(\REGFILE/reg_out[0][22] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][22] ), .B2(net83203), .ZN(n6438) );
  AOI22_X2 U6929 ( .A1(\REGFILE/reg_out[30][21] ), .A2(net84761), .B1(
        \REGFILE/reg_out[2][21] ), .B2(net75442), .ZN(n6474) );
  INV_X2 U6930 ( .A(\REGFILE/reg_out[15][31] ), .ZN(n10522) );
  NAND4_X2 U6931 ( .A1(n6641), .A2(n6640), .A3(n6638), .A4(n6639), .ZN(n6642)
         );
  AOI22_X2 U6932 ( .A1(\REGFILE/reg_out[23][11] ), .A2(net77828), .B1(
        \REGFILE/reg_out[22][11] ), .B2(net77836), .ZN(n6668) );
  AOI22_X1 U6933 ( .A1(\REGFILE/reg_out[0][27] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][27] ), .B2(net75464), .ZN(n6325) );
  AOI22_X2 U6934 ( .A1(\REGFILE/reg_out[19][12] ), .A2(net77812), .B1(
        \REGFILE/reg_out[1][12] ), .B2(net75478), .ZN(n6645) );
  BUF_X32 U6935 ( .A(aluA[30]), .Z(n5798) );
  INV_X32 U6936 ( .A(\PCLOGIC/imm26_32 [9]), .ZN(net87098) );
  OAI22_X2 U6937 ( .A1(n6002), .A2(net77440), .B1(n6003), .B2(net85371), .ZN(
        n6001) );
  NAND4_X2 U6938 ( .A1(n6451), .A2(n6450), .A3(n6449), .A4(n6448), .ZN(n6452)
         );
  INV_X8 U6939 ( .A(net75425), .ZN(net86304) );
  INV_X4 U6940 ( .A(n5947), .ZN(n6931) );
  INV_X1 U6941 ( .A(\REGFILE/reg_out[20][31] ), .ZN(n10525) );
  AOI22_X1 U6942 ( .A1(\REGFILE/reg_out[21][31] ), .A2(net77846), .B1(
        \REGFILE/reg_out[20][31] ), .B2(net77854), .ZN(n6228) );
  INV_X2 U6943 ( .A(n5799), .ZN(n5800) );
  INV_X2 U6944 ( .A(n5801), .ZN(n5802) );
  INV_X2 U6945 ( .A(n5803), .ZN(n5804) );
  AOI22_X2 U6946 ( .A1(\REGFILE/reg_out[0][13] ), .A2(net82342), .B1(n5814), 
        .B2(net75464), .ZN(net75764) );
  NOR2_X2 U6948 ( .A1(n6477), .A2(n6476), .ZN(n6478) );
  NOR2_X1 U6949 ( .A1(n4856), .A2(n10334), .ZN(n10335) );
  AOI22_X1 U6950 ( .A1(\REGFILE/reg_out[11][27] ), .A2(net77750), .B1(
        \REGFILE/reg_out[12][27] ), .B2(net75466), .ZN(n6326) );
  INV_X4 U6951 ( .A(dmem_write_out[23]), .ZN(n6433) );
  INV_X2 U6952 ( .A(n10323), .ZN(n5806) );
  NAND2_X1 U6953 ( .A1(\REGFILE/reg_out[25][21] ), .A2(net77530), .ZN(n7316)
         );
  AOI22_X2 U6954 ( .A1(\REGFILE/reg_out[24][21] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][21] ), .B2(net75438), .ZN(n6472) );
  INV_X2 U6955 ( .A(\REGFILE/reg_out[18][31] ), .ZN(n10524) );
  INV_X2 U6956 ( .A(n5808), .ZN(n5809) );
  INV_X2 U6957 ( .A(n5811), .ZN(n5812) );
  INV_X2 U6958 ( .A(n5813), .ZN(n5814) );
  AOI22_X2 U6959 ( .A1(\REGFILE/reg_out[30][11] ), .A2(net84761), .B1(n5874), 
        .B2(net82613), .ZN(n6682) );
  INV_X2 U6960 ( .A(n5816), .ZN(n5817) );
  INV_X4 U6961 ( .A(n5924), .ZN(n5818) );
  NOR2_X2 U6963 ( .A1(n6443), .A2(n6442), .ZN(n6455) );
  INV_X8 U6964 ( .A(net77632), .ZN(net77626) );
  NAND2_X1 U6965 ( .A1(\REGFILE/reg_out[27][19] ), .A2(net77422), .ZN(n7406)
         );
  OAI21_X2 U6966 ( .B1(n10388), .B2(n10387), .A(n10386), .ZN(n10390) );
  AND2_X2 U6967 ( .A1(n5916), .A2(n6929), .ZN(n5820) );
  INV_X8 U6968 ( .A(n5822), .ZN(n6929) );
  AOI22_X2 U6969 ( .A1(\REGFILE/reg_out[21][8] ), .A2(net77842), .B1(
        \REGFILE/reg_out[20][8] ), .B2(net77850), .ZN(n6735) );
  NOR2_X4 U6970 ( .A1(n6719), .A2(n6718), .ZN(n6731) );
  NAND2_X1 U6971 ( .A1(net77346), .A2(\REGFILE/reg_out[2][14] ), .ZN(n7652) );
  INV_X1 U6972 ( .A(\REGFILE/reg_out[13][31] ), .ZN(n10518) );
  INV_X2 U6973 ( .A(n5824), .ZN(n5825) );
  INV_X1 U6974 ( .A(\REGFILE/reg_out[9][31] ), .ZN(n10537) );
  AOI22_X1 U6975 ( .A1(\REGFILE/reg_out[9][31] ), .A2(net77702), .B1(
        \REGFILE/reg_out[8][31] ), .B2(n4829), .ZN(n6237) );
  INV_X4 U6976 ( .A(n6946), .ZN(n6932) );
  AOI22_X2 U6977 ( .A1(\REGFILE/reg_out[24][12] ), .A2(net75437), .B1(n5865), 
        .B2(net124970), .ZN(n6658) );
  AOI22_X2 U6978 ( .A1(\REGFILE/reg_out[24][11] ), .A2(net75437), .B1(n5882), 
        .B2(net124970), .ZN(n6680) );
  INV_X1 U6979 ( .A(n10913), .ZN(n5826) );
  NAND2_X1 U6980 ( .A1(\REGFILE/reg_out[3][8] ), .A2(net77414), .ZN(n7918) );
  NAND2_X2 U6981 ( .A1(\REGFILE/reg_out[25][20] ), .A2(net77530), .ZN(n7357)
         );
  NAND4_X2 U6982 ( .A1(n6495), .A2(n6494), .A3(n6493), .A4(n6492), .ZN(n6501)
         );
  AOI22_X2 U6983 ( .A1(\REGFILE/reg_out[7][19] ), .A2(net77714), .B1(
        \REGFILE/reg_out[6][19] ), .B2(net75456), .ZN(n6519) );
  NOR3_X1 U6985 ( .A1(n10352), .A2(n8849), .A3(net78003), .ZN(n8865) );
  AOI22_X1 U6986 ( .A1(\REGFILE/reg_out[7][30] ), .A2(net77714), .B1(
        \REGFILE/reg_out[6][30] ), .B2(net75456), .ZN(n6264) );
  AOI22_X1 U6987 ( .A1(\REGFILE/reg_out[7][28] ), .A2(net77716), .B1(
        \REGFILE/reg_out[6][28] ), .B2(net75456), .ZN(n6310) );
  AOI22_X1 U6988 ( .A1(\REGFILE/reg_out[7][27] ), .A2(net77716), .B1(
        \REGFILE/reg_out[6][27] ), .B2(net75456), .ZN(n6334) );
  AOI22_X2 U6989 ( .A1(\REGFILE/reg_out[26][20] ), .A2(net75439), .B1(
        \REGFILE/reg_out[27][20] ), .B2(net89184), .ZN(n6497) );
  AOI22_X1 U6990 ( .A1(\REGFILE/reg_out[24][30] ), .A2(net77602), .B1(
        \REGFILE/reg_out[25][30] ), .B2(net77610), .ZN(n6265) );
  NAND2_X1 U6991 ( .A1(\REGFILE/reg_out[27][21] ), .A2(net77422), .ZN(n7313)
         );
  AOI22_X2 U6992 ( .A1(\REGFILE/reg_out[17][12] ), .A2(net77796), .B1(
        \REGFILE/reg_out[18][12] ), .B2(n6896), .ZN(n6644) );
  NOR2_X2 U6993 ( .A1(n6377), .A2(n6376), .ZN(n6389) );
  NAND2_X4 U6994 ( .A1(n5990), .A2(net77462), .ZN(n6988) );
  XNOR2_X1 U6995 ( .A(n5806), .B(aluA[26]), .ZN(n10444) );
  INV_X1 U6996 ( .A(n10925), .ZN(n10323) );
  XNOR2_X1 U6997 ( .A(n5806), .B(net77040), .ZN(n8596) );
  AOI22_X1 U6998 ( .A1(\REGFILE/reg_out[0][5] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][5] ), .B2(net75464), .ZN(n6790) );
  AOI22_X2 U6999 ( .A1(\REGFILE/reg_out[26][25] ), .A2(net77620), .B1(
        \REGFILE/reg_out[27][25] ), .B2(net77626), .ZN(n6383) );
  NAND4_X2 U7000 ( .A1(n6499), .A2(n6497), .A3(n6498), .A4(n6496), .ZN(n6500)
         );
  NAND2_X1 U7001 ( .A1(\REGFILE/reg_out[8][14] ), .A2(net77310), .ZN(n7641) );
  NAND2_X1 U7002 ( .A1(n5781), .A2(net77382), .ZN(n7633) );
  NAND2_X1 U7003 ( .A1(\REGFILE/reg_out[28][14] ), .A2(n6175), .ZN(n10271) );
  NAND2_X1 U7004 ( .A1(\REGFILE/reg_out[28][14] ), .A2(net77382), .ZN(n7623)
         );
  OAI21_X4 U7005 ( .B1(n6296), .B2(net73697), .A(n6295), .ZN(n10927) );
  INV_X16 U7006 ( .A(n10927), .ZN(n6004) );
  NAND2_X1 U7007 ( .A1(net76488), .A2(\REGFILE/reg_out[31][30] ), .ZN(n8755)
         );
  AOI22_X1 U7008 ( .A1(\REGFILE/reg_out[31][30] ), .A2(net77670), .B1(
        \REGFILE/reg_out[3][30] ), .B2(n5609), .ZN(n6261) );
  NAND2_X1 U7009 ( .A1(\REGFILE/reg_out[1][15] ), .A2(net77526), .ZN(n7605) );
  AOI22_X2 U7010 ( .A1(\REGFILE/reg_out[0][7] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][7] ), .B2(net75464), .ZN(n6758) );
  INV_X2 U7011 ( .A(n5827), .ZN(n5828) );
  INV_X8 U7012 ( .A(net77506), .ZN(net77480) );
  INV_X4 U7013 ( .A(n5844), .ZN(n5829) );
  NAND4_X2 U7014 ( .A1(n6637), .A2(n6636), .A3(n6635), .A4(n6634), .ZN(n6643)
         );
  NAND2_X1 U7015 ( .A1(n10926), .A2(n5652), .ZN(n9094) );
  NAND2_X1 U7016 ( .A1(n5652), .A2(n10315), .ZN(n9581) );
  XNOR2_X1 U7017 ( .A(n5761), .B(n5652), .ZN(n10436) );
  XNOR2_X1 U7018 ( .A(net77040), .B(n5652), .ZN(n8594) );
  INV_X4 U7019 ( .A(n5918), .ZN(n5830) );
  NAND2_X1 U7020 ( .A1(\REGFILE/reg_out[3][14] ), .A2(net77418), .ZN(n7654) );
  INV_X4 U7021 ( .A(n5831), .ZN(n5832) );
  INV_X2 U7022 ( .A(n5833), .ZN(n5834) );
  AOI22_X2 U7023 ( .A1(\REGFILE/reg_out[26][4] ), .A2(net77620), .B1(
        \REGFILE/reg_out[27][4] ), .B2(net77626), .ZN(n6823) );
  NAND2_X1 U7024 ( .A1(n4890), .A2(\REGFILE/reg_out[8][13] ), .ZN(n9487) );
  INV_X2 U7025 ( .A(n5835), .ZN(n5836) );
  AOI22_X2 U7026 ( .A1(\REGFILE/reg_out[0][11] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][11] ), .B2(net75464), .ZN(n6670) );
  AOI22_X2 U7027 ( .A1(\REGFILE/reg_out[0][19] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][19] ), .B2(net83203), .ZN(n6510) );
  INV_X16 U7028 ( .A(net77500), .ZN(net77496) );
  INV_X16 U7029 ( .A(net77500), .ZN(net77494) );
  AOI22_X4 U7030 ( .A1(\REGFILE/reg_out[23][13] ), .A2(net77828), .B1(n5800), 
        .B2(net77836), .ZN(n6632) );
  NAND3_X1 U7031 ( .A1(n10929), .A2(n5761), .A3(net71078), .ZN(n8886) );
  NAND2_X1 U7032 ( .A1(n10929), .A2(net70696), .ZN(n9093) );
  NAND2_X1 U7033 ( .A1(n10929), .A2(n10926), .ZN(net70866) );
  NAND2_X1 U7034 ( .A1(n10929), .A2(n10315), .ZN(net70868) );
  NOR2_X1 U7035 ( .A1(n10929), .A2(n10319), .ZN(n10320) );
  NAND2_X1 U7036 ( .A1(net73708), .A2(aluA[26]), .ZN(n8683) );
  NAND3_X1 U7037 ( .A1(net71078), .A2(aluA[26]), .A3(n5806), .ZN(n9780) );
  NOR2_X1 U7038 ( .A1(n8449), .A2(n8448), .ZN(n8453) );
  NAND2_X1 U7039 ( .A1(n8937), .A2(aluA[26]), .ZN(n8938) );
  NAND2_X1 U7040 ( .A1(n9065), .A2(aluA[26]), .ZN(n8843) );
  NAND2_X1 U7041 ( .A1(net70720), .A2(aluA[26]), .ZN(n9359) );
  NAND2_X1 U7042 ( .A1(net70719), .A2(aluA[26]), .ZN(n10097) );
  NAND2_X1 U7043 ( .A1(n6040), .A2(aluA[26]), .ZN(n8714) );
  INV_X2 U7044 ( .A(aluA[26]), .ZN(n8597) );
  XNOR2_X1 U7045 ( .A(n8596), .B(aluA[26]), .ZN(n9777) );
  NAND2_X1 U7046 ( .A1(\REGFILE/reg_out[28][13] ), .A2(n6177), .ZN(n9467) );
  NAND2_X1 U7047 ( .A1(\REGFILE/reg_out[28][13] ), .A2(net77380), .ZN(n7667)
         );
  NAND2_X1 U7048 ( .A1(\REGFILE/reg_out[2][20] ), .A2(n6015), .ZN(n7390) );
  AOI22_X4 U7049 ( .A1(\REGFILE/reg_out[29][14] ), .A2(net77652), .B1(n4832), 
        .B2(n6911), .ZN(n6625) );
  INV_X2 U7050 ( .A(n5839), .ZN(n5840) );
  AOI22_X4 U7051 ( .A1(\REGFILE/reg_out[23][14] ), .A2(net77828), .B1(
        \REGFILE/reg_out[22][14] ), .B2(net77836), .ZN(n6610) );
  AOI22_X2 U7052 ( .A1(\REGFILE/reg_out[30][24] ), .A2(net77638), .B1(
        \REGFILE/reg_out[2][24] ), .B2(net75442), .ZN(n6403) );
  AOI22_X2 U7053 ( .A1(\REGFILE/reg_out[30][19] ), .A2(net84761), .B1(
        \REGFILE/reg_out[2][19] ), .B2(net75442), .ZN(n6522) );
  XNOR2_X1 U7054 ( .A(n10923), .B(net77038), .ZN(n8810) );
  XNOR2_X1 U7055 ( .A(n10408), .B(net77040), .ZN(n10165) );
  NAND2_X1 U7056 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[2].MUX/N1 ), .A2(n10408), 
        .ZN(n10409) );
  XNOR2_X1 U7057 ( .A(n10408), .B(n10109), .ZN(n10104) );
  AOI22_X4 U7058 ( .A1(\REGFILE/reg_out[17][14] ), .A2(net77796), .B1(n10953), 
        .B2(n5890), .ZN(n6608) );
  XNOR2_X1 U7059 ( .A(n5752), .B(net77040), .ZN(n10110) );
  XNOR2_X1 U7060 ( .A(n5752), .B(n10404), .ZN(n10407) );
  INV_X8 U7061 ( .A(net76205), .ZN(net75441) );
  NAND4_X2 U7062 ( .A1(n6661), .A2(n6659), .A3(n6660), .A4(n6658), .ZN(n6662)
         );
  INV_X8 U7063 ( .A(net76248), .ZN(net76202) );
  INV_X1 U7064 ( .A(n10917), .ZN(n5847) );
  NAND2_X1 U7065 ( .A1(net77550), .A2(\REGFILE/reg_out[22][27] ), .ZN(n7055)
         );
  NAND2_X1 U7066 ( .A1(net77348), .A2(\REGFILE/reg_out[2][17] ), .ZN(n7520) );
  NAND2_X1 U7067 ( .A1(\REGFILE/reg_out[25][17] ), .A2(net77528), .ZN(n7489)
         );
  AOI22_X1 U7068 ( .A1(\REGFILE/reg_out[11][0] ), .A2(net77746), .B1(
        \REGFILE/reg_out[12][0] ), .B2(net75466), .ZN(n6902) );
  AOI22_X2 U7069 ( .A1(\REGFILE/reg_out[26][27] ), .A2(net77620), .B1(
        \REGFILE/reg_out[27][27] ), .B2(net77630), .ZN(n6336) );
  AOI22_X2 U7070 ( .A1(\REGFILE/reg_out[17][21] ), .A2(net77796), .B1(
        \REGFILE/reg_out[18][21] ), .B2(n6896), .ZN(n6458) );
  AOI22_X2 U7071 ( .A1(\REGFILE/reg_out[4][9] ), .A2(n5678), .B1(
        \REGFILE/reg_out[5][9] ), .B2(net84475), .ZN(n6721) );
  NOR2_X2 U7072 ( .A1(n6387), .A2(n6386), .ZN(n6388) );
  NAND2_X1 U7073 ( .A1(net73878), .A2(net88253), .ZN(n8306) );
  AOI22_X2 U7074 ( .A1(\REGFILE/reg_out[17][20] ), .A2(net77796), .B1(
        \REGFILE/reg_out[18][20] ), .B2(n6896), .ZN(n6482) );
  AOI22_X2 U7075 ( .A1(\REGFILE/reg_out[30][18] ), .A2(net84761), .B1(
        \REGFILE/reg_out[2][18] ), .B2(net82613), .ZN(n6546) );
  AOI22_X1 U7076 ( .A1(\REGFILE/reg_out[7][31] ), .A2(net77716), .B1(
        \REGFILE/reg_out[6][31] ), .B2(net75456), .ZN(n6238) );
  AOI22_X1 U7077 ( .A1(\REGFILE/reg_out[7][29] ), .A2(net77714), .B1(
        \REGFILE/reg_out[6][29] ), .B2(net75456), .ZN(n6286) );
  AOI22_X1 U7078 ( .A1(\REGFILE/reg_out[7][26] ), .A2(net77714), .B1(
        \REGFILE/reg_out[6][26] ), .B2(net75456), .ZN(n6357) );
  AOI22_X1 U7079 ( .A1(\REGFILE/reg_out[7][23] ), .A2(net77714), .B1(
        \REGFILE/reg_out[6][23] ), .B2(net75456), .ZN(n6424) );
  INV_X8 U7080 ( .A(net76234), .ZN(net75466) );
  INV_X2 U7081 ( .A(n10352), .ZN(n5848) );
  NAND4_X2 U7082 ( .A1(n6441), .A2(n6440), .A3(n6439), .A4(n6438), .ZN(n6442)
         );
  AOI22_X4 U7083 ( .A1(\REGFILE/reg_out[14][14] ), .A2(net77780), .B1(n4853), 
        .B2(n5664), .ZN(n6615) );
  AOI22_X2 U7084 ( .A1(\REGFILE/reg_out[26][5] ), .A2(net77620), .B1(
        \REGFILE/reg_out[27][5] ), .B2(net77626), .ZN(n6801) );
  AOI22_X1 U7085 ( .A1(\REGFILE/reg_out[4][5] ), .A2(net75451), .B1(
        \REGFILE/reg_out[5][5] ), .B2(net75452), .ZN(n6797) );
  NAND2_X1 U7086 ( .A1(net77344), .A2(\REGFILE/reg_out[2][13] ), .ZN(n7696) );
  INV_X2 U7087 ( .A(n5849), .ZN(n5850) );
  INV_X16 U7088 ( .A(net75475), .ZN(net77800) );
  AOI22_X1 U7089 ( .A1(\REGFILE/reg_out[11][1] ), .A2(net77746), .B1(
        \REGFILE/reg_out[12][1] ), .B2(net75466), .ZN(n6879) );
  AOI22_X2 U7090 ( .A1(\REGFILE/reg_out[11][7] ), .A2(net77746), .B1(
        \REGFILE/reg_out[12][7] ), .B2(net75466), .ZN(n6759) );
  AOI22_X2 U7091 ( .A1(\REGFILE/reg_out[11][20] ), .A2(net77748), .B1(
        \REGFILE/reg_out[12][20] ), .B2(net83168), .ZN(n6487) );
  INV_X8 U7092 ( .A(net75441), .ZN(net77640) );
  INV_X2 U7093 ( .A(n5852), .ZN(n5853) );
  INV_X2 U7094 ( .A(n5854), .ZN(n5855) );
  AOI22_X4 U7095 ( .A1(\REGFILE/reg_out[29][15] ), .A2(net77652), .B1(n10951), 
        .B2(n6911), .ZN(n6601) );
  AOI22_X2 U7096 ( .A1(\REGFILE/reg_out[30][10] ), .A2(net77634), .B1(
        \REGFILE/reg_out[2][10] ), .B2(net82613), .ZN(n6704) );
  AOI22_X4 U7097 ( .A1(\REGFILE/reg_out[29][13] ), .A2(net77652), .B1(n5768), 
        .B2(n5751), .ZN(n6641) );
  NAND2_X1 U7098 ( .A1(\REGFILE/reg_out[27][8] ), .A2(net77414), .ZN(n7888) );
  INV_X1 U7099 ( .A(\REGFILE/reg_out[27][14] ), .ZN(n10270) );
  AOI22_X1 U7100 ( .A1(\REGFILE/reg_out[26][31] ), .A2(net77620), .B1(
        \REGFILE/reg_out[27][31] ), .B2(net89184), .ZN(n6241) );
  AOI22_X2 U7101 ( .A1(\REGFILE/reg_out[0][21] ), .A2(net120684), .B1(n5809), 
        .B2(net75464), .ZN(n6462) );
  AOI22_X2 U7102 ( .A1(\REGFILE/reg_out[11][21] ), .A2(net77748), .B1(
        \REGFILE/reg_out[12][21] ), .B2(net83168), .ZN(n6463) );
  INV_X1 U7103 ( .A(\REGFILE/reg_out[16][31] ), .ZN(n10523) );
  AOI22_X1 U7104 ( .A1(\REGFILE/reg_out[16][31] ), .A2(net75467), .B1(
        \REGFILE/reg_out[15][31] ), .B2(net77774), .ZN(n6231) );
  NAND2_X1 U7105 ( .A1(\REGFILE/reg_out[2][18] ), .A2(net77348), .ZN(n7478) );
  AOI22_X1 U7106 ( .A1(\REGFILE/reg_out[30][23] ), .A2(net77638), .B1(
        \REGFILE/reg_out[2][23] ), .B2(net75442), .ZN(n6426) );
  INV_X2 U7107 ( .A(n5858), .ZN(n5859) );
  INV_X2 U7108 ( .A(n5860), .ZN(n5861) );
  INV_X2 U7109 ( .A(n5862), .ZN(n5863) );
  INV_X2 U7110 ( .A(n5864), .ZN(n5865) );
  INV_X2 U7111 ( .A(\REGFILE/reg_out[10][15] ), .ZN(n10298) );
  INV_X2 U7112 ( .A(n9057), .ZN(n9058) );
  INV_X1 U7113 ( .A(n10424), .ZN(n10281) );
  AOI22_X1 U7114 ( .A1(\REGFILE/reg_out[17][27] ), .A2(net77798), .B1(
        \REGFILE/reg_out[18][27] ), .B2(n5890), .ZN(n6321) );
  AOI22_X1 U7115 ( .A1(\REGFILE/reg_out[17][23] ), .A2(net77798), .B1(
        \REGFILE/reg_out[18][23] ), .B2(n5890), .ZN(n6411) );
  AOI22_X2 U7116 ( .A1(\REGFILE/reg_out[16][7] ), .A2(net77762), .B1(
        \REGFILE/reg_out[15][7] ), .B2(net75468), .ZN(n6760) );
  INV_X32 U7117 ( .A(net77500), .ZN(net77498) );
  INV_X16 U7118 ( .A(net77856), .ZN(net77850) );
  INV_X1 U7119 ( .A(n10915), .ZN(n5867) );
  INV_X8 U7120 ( .A(net76258), .ZN(net75482) );
  AOI22_X2 U7121 ( .A1(\REGFILE/reg_out[9][7] ), .A2(net77698), .B1(
        \REGFILE/reg_out[8][7] ), .B2(n4829), .ZN(net75624) );
  NAND2_X1 U7122 ( .A1(\REGFILE/reg_out[27][11] ), .A2(n4872), .ZN(n9907) );
  NAND2_X1 U7123 ( .A1(\REGFILE/reg_out[27][11] ), .A2(net77416), .ZN(n7756)
         );
  INV_X1 U7124 ( .A(\REGFILE/reg_out[15][10] ), .ZN(n10144) );
  NAND2_X1 U7125 ( .A1(\REGFILE/reg_out[15][10] ), .A2(net77484), .ZN(n7814)
         );
  NAND2_X1 U7126 ( .A1(n6100), .A2(\REGFILE/reg_out[13][11] ), .ZN(n9877) );
  NAND2_X1 U7127 ( .A1(\REGFILE/reg_out[13][11] ), .A2(net77452), .ZN(n7769)
         );
  NAND2_X2 U7128 ( .A1(\REGFILE/reg_out[25][8] ), .A2(net77522), .ZN(n7883) );
  OAI22_X1 U7129 ( .A1(n8729), .A2(n8823), .B1(n6005), .B2(n8714), .ZN(n9297)
         );
  AOI22_X1 U7130 ( .A1(\REGFILE/reg_out[26][28] ), .A2(net77620), .B1(
        \REGFILE/reg_out[27][28] ), .B2(net89184), .ZN(n6312) );
  AOI22_X1 U7131 ( .A1(\REGFILE/reg_out[26][0] ), .A2(net77620), .B1(
        \REGFILE/reg_out[27][0] ), .B2(net89184), .ZN(n6913) );
  AOI22_X1 U7132 ( .A1(\REGFILE/reg_out[26][1] ), .A2(net77620), .B1(
        \REGFILE/reg_out[27][1] ), .B2(net77630), .ZN(n6889) );
  NAND4_X2 U7133 ( .A1(n6523), .A2(n6522), .A3(n6521), .A4(n6520), .ZN(n6524)
         );
  NAND2_X2 U7134 ( .A1(\REGFILE/reg_out[10][14] ), .A2(net77346), .ZN(n7642)
         );
  AOI22_X2 U7136 ( .A1(\REGFILE/reg_out[16][9] ), .A2(net87506), .B1(
        \REGFILE/reg_out[15][9] ), .B2(net75468), .ZN(n6716) );
  INV_X16 U7137 ( .A(net77640), .ZN(net77638) );
  INV_X8 U7138 ( .A(net76234), .ZN(net83168) );
  INV_X2 U7139 ( .A(n5871), .ZN(n5872) );
  INV_X2 U7140 ( .A(n5873), .ZN(n5874) );
  AOI22_X1 U7141 ( .A1(\REGFILE/reg_out[0][23] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][23] ), .B2(net75464), .ZN(n6415) );
  NAND2_X1 U7142 ( .A1(net77376), .A2(\REGFILE/reg_out[12][10] ), .ZN(n7819)
         );
  OAI21_X1 U7143 ( .B1(n9855), .B2(n9854), .A(n9853), .ZN(n9856) );
  OAI21_X2 U7144 ( .B1(n10381), .B2(n10380), .A(n10379), .ZN(n10384) );
  INV_X2 U7145 ( .A(n9029), .ZN(n9030) );
  XNOR2_X1 U7146 ( .A(n9029), .B(aluA[18]), .ZN(n9028) );
  NAND2_X1 U7147 ( .A1(aluA[18]), .A2(n10352), .ZN(n10353) );
  NOR2_X1 U7148 ( .A1(n5931), .A2(n10463), .ZN(n10362) );
  AOI21_X2 U7149 ( .B1(n10424), .B2(n10363), .A(n10362), .ZN(n10367) );
  INV_X2 U7150 ( .A(n5875), .ZN(n5876) );
  NAND2_X1 U7151 ( .A1(net73878), .A2(net73987), .ZN(n8301) );
  INV_X8 U7152 ( .A(n10371), .ZN(n5943) );
  NAND2_X4 U7153 ( .A1(net121496), .A2(net76195), .ZN(n6239) );
  NAND2_X1 U7154 ( .A1(\REGFILE/reg_out[25][10] ), .A2(net77522), .ZN(n7795)
         );
  NAND2_X1 U7155 ( .A1(\REGFILE/reg_out[12][11] ), .A2(net77380), .ZN(n7775)
         );
  NAND2_X1 U7156 ( .A1(\REGFILE/reg_out[12][11] ), .A2(n4873), .ZN(n9875) );
  INV_X2 U7157 ( .A(n5879), .ZN(n5880) );
  INV_X2 U7158 ( .A(n5881), .ZN(n5882) );
  NAND2_X1 U7159 ( .A1(n4878), .A2(\REGFILE/reg_out[25][16] ), .ZN(n9240) );
  NAND2_X1 U7160 ( .A1(net77528), .A2(\REGFILE/reg_out[25][16] ), .ZN(n7531)
         );
  INV_X2 U7161 ( .A(n5883), .ZN(n5884) );
  NOR2_X2 U7162 ( .A1(n9857), .A2(n9856), .ZN(n9858) );
  INV_X1 U7163 ( .A(n10422), .ZN(n9402) );
  AOI21_X2 U7164 ( .B1(n10422), .B2(n10370), .A(n10369), .ZN(n10374) );
  NAND3_X1 U7165 ( .A1(net71078), .A2(\WIRE_ALU_A/MUX2TO1_32BIT[13].MUX/N1 ), 
        .A3(net85047), .ZN(n9413) );
  NOR2_X1 U7166 ( .A1(net85047), .A2(n10368), .ZN(n10369) );
  AOI22_X4 U7167 ( .A1(\REGFILE/reg_out[31][18] ), .A2(net77668), .B1(
        \REGFILE/reg_out[3][18] ), .B2(net77676), .ZN(n6540) );
  AOI22_X2 U7168 ( .A1(\REGFILE/reg_out[7][10] ), .A2(net75455), .B1(
        \REGFILE/reg_out[6][10] ), .B2(net75456), .ZN(n6701) );
  AOI22_X1 U7169 ( .A1(\REGFILE/reg_out[24][0] ), .A2(net77602), .B1(
        \REGFILE/reg_out[25][0] ), .B2(net77614), .ZN(n6912) );
  AOI22_X1 U7170 ( .A1(\REGFILE/reg_out[24][1] ), .A2(net77602), .B1(
        \REGFILE/reg_out[25][1] ), .B2(net77610), .ZN(n6888) );
  AOI22_X1 U7171 ( .A1(\REGFILE/reg_out[24][28] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][28] ), .B2(net77610), .ZN(n6311) );
  NAND4_X2 U7172 ( .A1(n6427), .A2(n6426), .A3(net75995), .A4(n6425), .ZN(
        n6428) );
  OAI21_X1 U7173 ( .B1(net148116), .B2(net73697), .A(net75843), .ZN(n5885) );
  NAND2_X1 U7174 ( .A1(\REGFILE/reg_out[25][9] ), .A2(net77522), .ZN(n7839) );
  NAND2_X1 U7175 ( .A1(\REGFILE/reg_out[2][9] ), .A2(net77342), .ZN(n7872) );
  NAND2_X1 U7176 ( .A1(\REGFILE/reg_out[12][18] ), .A2(net77384), .ZN(n7469)
         );
  AOI22_X1 U7177 ( .A1(\REGFILE/reg_out[29][1] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][1] ), .B2(n6911), .ZN(n6891) );
  NAND4_X2 U7178 ( .A1(n6891), .A2(n6890), .A3(n6889), .A4(n6888), .ZN(n6892)
         );
  INV_X16 U7179 ( .A(n5649), .ZN(n5890) );
  NOR2_X2 U7180 ( .A1(net76261), .A2(net88131), .ZN(n6000) );
  AOI22_X2 U7181 ( .A1(\REGFILE/reg_out[26][12] ), .A2(net75439), .B1(n5861), 
        .B2(net75440), .ZN(n6659) );
  AOI22_X2 U7182 ( .A1(\REGFILE/reg_out[26][16] ), .A2(net75439), .B1(
        \REGFILE/reg_out[27][16] ), .B2(net89184), .ZN(n6577) );
  INV_X8 U7183 ( .A(n8885), .ZN(n10929) );
  INV_X2 U7184 ( .A(n5891), .ZN(n5892) );
  AOI22_X2 U7185 ( .A1(\REGFILE/reg_out[17][22] ), .A2(net77798), .B1(
        \REGFILE/reg_out[18][22] ), .B2(n5890), .ZN(n6434) );
  INV_X2 U7186 ( .A(n5893), .ZN(n5894) );
  INV_X2 U7187 ( .A(n5895), .ZN(n5896) );
  INV_X2 U7188 ( .A(net82499), .ZN(net82500) );
  INV_X16 U7189 ( .A(net77106), .ZN(net77100) );
  NAND4_X2 U7190 ( .A1(n6465), .A2(n6464), .A3(n6462), .A4(n6463), .ZN(n6466)
         );
  NAND2_X4 U7191 ( .A1(n6342), .A2(n6341), .ZN(dmem_write_out[27]) );
  INV_X1 U7192 ( .A(n5762), .ZN(n8989) );
  NOR2_X1 U7193 ( .A1(n5762), .A2(n10327), .ZN(n10328) );
  NAND3_X1 U7194 ( .A1(n10930), .A2(n5762), .A3(net71078), .ZN(n8990) );
  OAI21_X1 U7195 ( .B1(n6457), .B2(net78055), .A(n6456), .ZN(n5897) );
  NOR2_X2 U7196 ( .A1(n6406), .A2(n6405), .ZN(n6407) );
  INV_X8 U7197 ( .A(net76222), .ZN(net75453) );
  INV_X8 U7198 ( .A(net76209), .ZN(net75443) );
  NAND2_X4 U7199 ( .A1(n6583), .A2(n6582), .ZN(dmem_write_out[16]) );
  AOI22_X1 U7200 ( .A1(\REGFILE/reg_out[17][25] ), .A2(net77798), .B1(
        \REGFILE/reg_out[18][25] ), .B2(n5890), .ZN(n6368) );
  AOI22_X2 U7201 ( .A1(\REGFILE/reg_out[17][8] ), .A2(net77794), .B1(
        \REGFILE/reg_out[18][8] ), .B2(n6896), .ZN(n6732) );
  INV_X8 U7202 ( .A(aluA[28]), .ZN(n6006) );
  AOI22_X4 U7203 ( .A1(\REGFILE/reg_out[4][13] ), .A2(n5679), .B1(n5817), .B2(
        net84475), .ZN(n6635) );
  XNOR2_X1 U7204 ( .A(n5870), .B(net77038), .ZN(n9057) );
  XNOR2_X1 U7205 ( .A(n5870), .B(n10463), .ZN(n10424) );
  INV_X16 U7206 ( .A(net76255), .ZN(net77836) );
  XNOR2_X1 U7207 ( .A(n9615), .B(n9656), .ZN(n9664) );
  OAI21_X2 U7208 ( .B1(n10395), .B2(n10394), .A(n10393), .ZN(n10398) );
  NAND2_X4 U7209 ( .A1(n5936), .A2(net123282), .ZN(n5899) );
  NAND2_X4 U7210 ( .A1(n5899), .A2(n5900), .ZN(aluA[29]) );
  NAND3_X2 U7211 ( .A1(n6980), .A2(n6981), .A3(n5753), .ZN(n6982) );
  NAND2_X1 U7212 ( .A1(\REGFILE/reg_out[21][29] ), .A2(net77462), .ZN(n6980)
         );
  NAND2_X1 U7214 ( .A1(\REGFILE/reg_out[12][13] ), .A2(n4873), .ZN(n9433) );
  NAND2_X1 U7215 ( .A1(\REGFILE/reg_out[12][13] ), .A2(net77380), .ZN(n7687)
         );
  AOI22_X1 U7216 ( .A1(\REGFILE/reg_out[4][29] ), .A2(n5678), .B1(
        \REGFILE/reg_out[5][29] ), .B2(net84475), .ZN(n6284) );
  NAND2_X1 U7217 ( .A1(n6093), .A2(\REGFILE/reg_out[10][13] ), .ZN(n9429) );
  NAND2_X1 U7218 ( .A1(\REGFILE/reg_out[10][13] ), .A2(net77344), .ZN(n7686)
         );
  INV_X4 U7219 ( .A(n5903), .ZN(n5904) );
  INV_X1 U7220 ( .A(n10910), .ZN(n5905) );
  NAND2_X1 U7221 ( .A1(n5904), .A2(n4872), .ZN(n9244) );
  NAND2_X1 U7222 ( .A1(\REGFILE/reg_out[5][5] ), .A2(net77456), .ZN(n8041) );
  NAND2_X1 U7223 ( .A1(\REGFILE/reg_out[27][16] ), .A2(net77420), .ZN(n7536)
         );
  NAND2_X1 U7224 ( .A1(aluA[16]), .A2(n5847), .ZN(n10359) );
  NAND2_X1 U7225 ( .A1(\REGFILE/reg_out[10][5] ), .A2(net77338), .ZN(n8036) );
  NAND2_X1 U7226 ( .A1(\REGFILE/reg_out[2][5] ), .A2(net77338), .ZN(n8046) );
  INV_X2 U7227 ( .A(n9050), .ZN(n9051) );
  XNOR2_X1 U7228 ( .A(n9050), .B(aluA[17]), .ZN(n9052) );
  AOI21_X2 U7229 ( .B1(n10448), .B2(n10358), .A(n10357), .ZN(n10361) );
  NOR2_X2 U7230 ( .A1(n10448), .A2(net78014), .ZN(n9023) );
  NAND2_X1 U7231 ( .A1(n6180), .A2(n5850), .ZN(n9473) );
  NAND2_X1 U7232 ( .A1(n5850), .A2(net77560), .ZN(n7664) );
  INV_X4 U7233 ( .A(n5906), .ZN(n5907) );
  INV_X2 U7234 ( .A(n5908), .ZN(n5909) );
  INV_X1 U7235 ( .A(n5897), .ZN(n10338) );
  AOI22_X1 U7236 ( .A1(\REGFILE/reg_out[11][30] ), .A2(net77750), .B1(
        \REGFILE/reg_out[12][30] ), .B2(net83168), .ZN(n6256) );
  AOI22_X1 U7237 ( .A1(\REGFILE/reg_out[11][28] ), .A2(net77750), .B1(
        \REGFILE/reg_out[12][28] ), .B2(net83168), .ZN(n6302) );
  AOI22_X1 U7238 ( .A1(\REGFILE/reg_out[11][29] ), .A2(net77750), .B1(
        \REGFILE/reg_out[12][29] ), .B2(net83168), .ZN(n6278) );
  AOI22_X1 U7239 ( .A1(\REGFILE/reg_out[11][26] ), .A2(net77750), .B1(
        \REGFILE/reg_out[12][26] ), .B2(net83168), .ZN(n6349) );
  XNOR2_X1 U7240 ( .A(n5905), .B(n10396), .ZN(n10399) );
  XNOR2_X1 U7241 ( .A(n5905), .B(net77038), .ZN(n9956) );
  NOR3_X1 U7242 ( .A1(net78003), .A2(n5905), .A3(n10396), .ZN(n9591) );
  NOR2_X1 U7243 ( .A1(n10910), .A2(n10396), .ZN(n10397) );
  AOI21_X2 U7244 ( .B1(n10399), .B2(n10398), .A(n10397), .ZN(n10403) );
  NOR2_X1 U7245 ( .A1(n10399), .A2(net78014), .ZN(n9607) );
  NAND2_X1 U7246 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[5].MUX/N1 ), .A2(n9956), .ZN(
        n9957) );
  AOI21_X2 U7247 ( .B1(n9592), .B2(net70697), .A(n9591), .ZN(n9632) );
  AOI22_X4 U7248 ( .A1(\REGFILE/reg_out[31][8] ), .A2(net77666), .B1(
        \REGFILE/reg_out[3][8] ), .B2(n5609), .ZN(n6742) );
  INV_X2 U7249 ( .A(n5911), .ZN(n5912) );
  XNOR2_X1 U7250 ( .A(n10933), .B(n9559), .ZN(n10431) );
  NOR2_X2 U7251 ( .A1(n10432), .A2(n10431), .ZN(n10439) );
  INV_X2 U7252 ( .A(\REGFILE/reg_out[2][8] ), .ZN(n9524) );
  NAND2_X1 U7253 ( .A1(\REGFILE/reg_out[2][8] ), .A2(net77342), .ZN(n7916) );
  INV_X4 U7254 ( .A(net36479), .ZN(net81810) );
  AOI21_X2 U7255 ( .B1(n10344), .B2(n10343), .A(n10342), .ZN(n10348) );
  NOR3_X1 U7256 ( .A1(n9559), .A2(n10341), .A3(net78003), .ZN(n9560) );
  XNOR2_X1 U7257 ( .A(n10933), .B(n4810), .ZN(n9543) );
  OAI21_X2 U7258 ( .B1(n10348), .B2(n10347), .A(n10346), .ZN(n10351) );
  NOR3_X2 U7259 ( .A1(n9562), .A2(n9561), .A3(n9560), .ZN(n9563) );
  INV_X1 U7260 ( .A(n5783), .ZN(n9559) );
  AOI22_X1 U7261 ( .A1(\REGFILE/reg_out[30][0] ), .A2(net77634), .B1(
        \REGFILE/reg_out[2][0] ), .B2(net75442), .ZN(n6914) );
  AOI22_X1 U7262 ( .A1(\REGFILE/reg_out[30][29] ), .A2(net77638), .B1(
        \REGFILE/reg_out[2][29] ), .B2(net75442), .ZN(n6289) );
  AOI22_X1 U7263 ( .A1(\REGFILE/reg_out[30][28] ), .A2(net77638), .B1(
        \REGFILE/reg_out[2][28] ), .B2(net75442), .ZN(n6313) );
  XNOR2_X1 U7264 ( .A(n5897), .B(net77038), .ZN(n8813) );
  AOI22_X1 U7265 ( .A1(\REGFILE/reg_out[7][0] ), .A2(net77716), .B1(
        \REGFILE/reg_out[6][0] ), .B2(net75456), .ZN(n6910) );
  AOI22_X2 U7266 ( .A1(\REGFILE/reg_out[7][15] ), .A2(net77714), .B1(
        \REGFILE/reg_out[6][15] ), .B2(net75456), .ZN(n6597) );
  AOI22_X2 U7267 ( .A1(\REGFILE/reg_out[17][9] ), .A2(net77794), .B1(
        \REGFILE/reg_out[18][9] ), .B2(n6896), .ZN(n6710) );
  AOI22_X2 U7268 ( .A1(\REGFILE/reg_out[19][9] ), .A2(net77810), .B1(
        \REGFILE/reg_out[1][9] ), .B2(net75478), .ZN(n6711) );
  AOI22_X1 U7269 ( .A1(\REGFILE/reg_out[0][2] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][2] ), .B2(net75464), .ZN(n6856) );
  AOI22_X1 U7270 ( .A1(\REGFILE/reg_out[17][31] ), .A2(net77798), .B1(
        \REGFILE/reg_out[18][31] ), .B2(n5890), .ZN(n6225) );
  AOI22_X1 U7271 ( .A1(\REGFILE/reg_out[17][30] ), .A2(net77798), .B1(
        \REGFILE/reg_out[18][30] ), .B2(n5890), .ZN(n6251) );
  AOI22_X1 U7272 ( .A1(\REGFILE/reg_out[17][29] ), .A2(net77798), .B1(
        \REGFILE/reg_out[18][29] ), .B2(n5890), .ZN(n6273) );
  AOI22_X1 U7273 ( .A1(\REGFILE/reg_out[17][28] ), .A2(net77798), .B1(
        \REGFILE/reg_out[18][28] ), .B2(n5890), .ZN(n6297) );
  AOI22_X1 U7274 ( .A1(\REGFILE/reg_out[17][26] ), .A2(net77798), .B1(
        \REGFILE/reg_out[18][26] ), .B2(n5890), .ZN(n6344) );
  INV_X1 U7275 ( .A(n4852), .ZN(n10352) );
  NAND2_X4 U7276 ( .A1(n10046), .A2(net76270), .ZN(n10052) );
  NAND2_X1 U7277 ( .A1(n6093), .A2(\REGFILE/reg_out[10][7] ), .ZN(n9707) );
  NAND2_X1 U7278 ( .A1(\REGFILE/reg_out[10][7] ), .A2(net77338), .ZN(n7950) );
  INV_X2 U7279 ( .A(n5846), .ZN(n10266) );
  NAND2_X1 U7280 ( .A1(n5846), .A2(net77382), .ZN(n7643) );
  NAND2_X1 U7281 ( .A1(\REGFILE/reg_out[27][14] ), .A2(net77418), .ZN(n7624)
         );
  NAND2_X1 U7282 ( .A1(n4879), .A2(\REGFILE/reg_out[2][7] ), .ZN(n9749) );
  NAND2_X1 U7283 ( .A1(\REGFILE/reg_out[2][7] ), .A2(net77338), .ZN(n7958) );
  NAND2_X1 U7284 ( .A1(\REGFILE/reg_out[27][7] ), .A2(n4872), .ZN(n9743) );
  OR2_X2 U7285 ( .A1(n5914), .A2(net77506), .ZN(n6970) );
  INV_X2 U7286 ( .A(\REGFILE/reg_out[25][14] ), .ZN(n10269) );
  NAND2_X1 U7287 ( .A1(\REGFILE/reg_out[25][14] ), .A2(net77526), .ZN(n7619)
         );
  INV_X2 U7288 ( .A(\REGFILE/reg_out[14][31] ), .ZN(n10520) );
  AOI22_X1 U7289 ( .A1(\REGFILE/reg_out[14][31] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][31] ), .B2(n6009), .ZN(n6232) );
  INV_X1 U7290 ( .A(n5619), .ZN(net73850) );
  INV_X2 U7291 ( .A(\REGFILE/reg_out[12][31] ), .ZN(n10515) );
  AOI22_X1 U7292 ( .A1(\REGFILE/reg_out[11][31] ), .A2(net77750), .B1(
        \REGFILE/reg_out[12][31] ), .B2(net83167), .ZN(n6230) );
  NAND2_X2 U7293 ( .A1(\REGFILE/reg_out[8][29] ), .A2(net77318), .ZN(n6973) );
  AOI21_X2 U7294 ( .B1(n10446), .B2(n10351), .A(n10350), .ZN(n10355) );
  NAND4_X1 U7295 ( .A1(n10448), .A2(n10447), .A3(n10446), .A4(n10445), .ZN(
        n10449) );
  NOR2_X2 U7296 ( .A1(n10446), .A2(net78014), .ZN(n9985) );
  INV_X2 U7297 ( .A(n8819), .ZN(n8820) );
  XNOR2_X1 U7298 ( .A(n8819), .B(aluA[19]), .ZN(n9992) );
  AOI22_X2 U7299 ( .A1(\REGFILE/reg_out[17][7] ), .A2(net77794), .B1(
        \REGFILE/reg_out[18][7] ), .B2(n5890), .ZN(n6754) );
  INV_X1 U7300 ( .A(n5650), .ZN(n9995) );
  NOR2_X1 U7301 ( .A1(n5783), .A2(n10341), .ZN(n10342) );
  INV_X2 U7302 ( .A(n8815), .ZN(n8816) );
  XNOR2_X1 U7303 ( .A(n8815), .B(aluA[20]), .ZN(n10053) );
  NAND4_X1 U7304 ( .A1(n10444), .A2(n10443), .A3(n10442), .A4(n10441), .ZN(
        n10450) );
  NOR2_X2 U7305 ( .A1(n10443), .A2(net78014), .ZN(n10055) );
  NAND2_X1 U7306 ( .A1(aluA[20]), .A2(n10345), .ZN(n10346) );
  NOR3_X2 U7307 ( .A1(n10345), .A2(n10071), .A3(net78003), .ZN(n10072) );
  AOI22_X1 U7308 ( .A1(\REGFILE/reg_out[17][0] ), .A2(net77794), .B1(
        \REGFILE/reg_out[18][0] ), .B2(n5890), .ZN(n6897) );
  AOI22_X1 U7309 ( .A1(\REGFILE/reg_out[17][1] ), .A2(net77794), .B1(
        \REGFILE/reg_out[18][1] ), .B2(n5890), .ZN(n6874) );
  AOI22_X1 U7310 ( .A1(\REGFILE/reg_out[17][2] ), .A2(net77794), .B1(
        \REGFILE/reg_out[18][2] ), .B2(n5890), .ZN(n6852) );
  AOI22_X1 U7311 ( .A1(\REGFILE/reg_out[17][4] ), .A2(net77794), .B1(
        \REGFILE/reg_out[18][4] ), .B2(n5890), .ZN(n6808) );
  AOI22_X1 U7312 ( .A1(\REGFILE/reg_out[17][3] ), .A2(net77794), .B1(
        \REGFILE/reg_out[18][3] ), .B2(n5890), .ZN(n6830) );
  XNOR2_X1 U7313 ( .A(n5675), .B(net77038), .ZN(n8815) );
  XNOR2_X1 U7314 ( .A(n5675), .B(aluA[20]), .ZN(n10443) );
  INV_X1 U7315 ( .A(n5675), .ZN(n10345) );
  XNOR2_X1 U7316 ( .A(n5848), .B(aluA[18]), .ZN(n10445) );
  XNOR2_X1 U7317 ( .A(n5848), .B(net77038), .ZN(n9029) );
  NOR2_X1 U7318 ( .A1(n5650), .A2(n10349), .ZN(n10350) );
  XNOR2_X1 U7319 ( .A(n5650), .B(aluA[19]), .ZN(n10446) );
  XNOR2_X1 U7320 ( .A(n5650), .B(net77038), .ZN(n8819) );
  NAND2_X1 U7321 ( .A1(\REGFILE/reg_out[27][7] ), .A2(net77410), .ZN(n7932) );
  NAND2_X1 U7322 ( .A1(net77418), .A2(\REGFILE/reg_out[27][15] ), .ZN(n7580)
         );
  NAND2_X2 U7323 ( .A1(\REGFILE/reg_out[0][6] ), .A2(net120684), .ZN(n5945) );
  NOR2_X2 U7324 ( .A1(n6839), .A2(n6838), .ZN(n6851) );
  AOI22_X1 U7325 ( .A1(\REGFILE/reg_out[30][3] ), .A2(net77634), .B1(
        \REGFILE/reg_out[2][3] ), .B2(net82613), .ZN(n6846) );
  NOR2_X1 U7326 ( .A1(net36479), .A2(n10464), .ZN(n10389) );
  NAND3_X1 U7327 ( .A1(net71078), .A2(\WIRE_ALU_A/MUX2TO1_32BIT[7].MUX/N1 ), 
        .A3(net36479), .ZN(n9691) );
  AOI22_X2 U7328 ( .A1(\REGFILE/reg_out[4][6] ), .A2(n5678), .B1(
        \REGFILE/reg_out[5][6] ), .B2(net84475), .ZN(n6775) );
  NAND2_X1 U7329 ( .A1(n4878), .A2(\REGFILE/reg_out[25][7] ), .ZN(n9739) );
  NAND2_X1 U7330 ( .A1(\REGFILE/reg_out[25][7] ), .A2(net77520), .ZN(n7927) );
  AOI22_X1 U7331 ( .A1(net73838), .A2(n10949), .B1(n6019), .B2(n5998), .ZN(
        n8413) );
  INV_X4 U7332 ( .A(n5958), .ZN(n5919) );
  INV_X2 U7333 ( .A(n5920), .ZN(n5921) );
  INV_X2 U7334 ( .A(n5922), .ZN(n5923) );
  INV_X2 U7335 ( .A(n5925), .ZN(n5926) );
  INV_X2 U7336 ( .A(n5927), .ZN(n5928) );
  INV_X2 U7337 ( .A(n5929), .ZN(n5930) );
  NAND2_X1 U7338 ( .A1(n10423), .A2(n10422), .ZN(n10427) );
  AOI22_X4 U7339 ( .A1(\REGFILE/reg_out[4][10] ), .A2(net75451), .B1(n4798), 
        .B2(net84475), .ZN(n6699) );
  XNOR2_X1 U7340 ( .A(n5885), .B(net77038), .ZN(n9050) );
  XNOR2_X1 U7341 ( .A(n5885), .B(aluA[17]), .ZN(n10448) );
  NOR2_X1 U7342 ( .A1(n5885), .A2(n10356), .ZN(n10357) );
  INV_X1 U7343 ( .A(n5885), .ZN(n9035) );
  NAND3_X4 U7344 ( .A1(net75368), .A2(n6955), .A3(net75367), .ZN(aluA[30]) );
  AOI22_X1 U7345 ( .A1(\REGFILE/reg_out[4][1] ), .A2(n5678), .B1(
        \REGFILE/reg_out[5][1] ), .B2(net84475), .ZN(n6885) );
  AOI22_X1 U7346 ( .A1(\REGFILE/reg_out[4][2] ), .A2(n5679), .B1(
        \REGFILE/reg_out[5][2] ), .B2(net75452), .ZN(n6863) );
  AOI22_X1 U7347 ( .A1(\REGFILE/reg_out[4][3] ), .A2(net75451), .B1(
        \REGFILE/reg_out[5][3] ), .B2(net75452), .ZN(n6841) );
  NOR2_X4 U7348 ( .A1(n6571), .A2(n6570), .ZN(n6583) );
  OAI22_X1 U7349 ( .A1(n10290), .A2(net70691), .B1(n10289), .B2(n5870), .ZN(
        n10291) );
  INV_X4 U7350 ( .A(net77386), .ZN(net77396) );
  INV_X4 U7351 ( .A(net77386), .ZN(net77394) );
  AOI22_X1 U7352 ( .A1(\REGFILE/reg_out[16][1] ), .A2(net87506), .B1(
        \REGFILE/reg_out[15][1] ), .B2(n5579), .ZN(n6880) );
  XNOR2_X1 U7353 ( .A(net81810), .B(net77040), .ZN(n9612) );
  XNOR2_X1 U7354 ( .A(net81810), .B(n10464), .ZN(n10391) );
  AOI22_X1 U7355 ( .A1(\REGFILE/reg_out[14][0] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][0] ), .B2(n6009), .ZN(n6904) );
  AOI22_X1 U7356 ( .A1(\REGFILE/reg_out[14][1] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][1] ), .B2(n5663), .ZN(n6881) );
  AOI22_X1 U7357 ( .A1(\REGFILE/reg_out[14][2] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][2] ), .B2(n5663), .ZN(n6859) );
  AOI22_X1 U7358 ( .A1(\REGFILE/reg_out[14][3] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][3] ), .B2(n5664), .ZN(n6837) );
  AOI22_X1 U7359 ( .A1(\REGFILE/reg_out[14][4] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][4] ), .B2(n6009), .ZN(n6815) );
  AOI22_X4 U7360 ( .A1(\REGFILE/reg_out[31][17] ), .A2(net77668), .B1(
        \REGFILE/reg_out[3][17] ), .B2(net77676), .ZN(n6558) );
  XNOR2_X1 U7361 ( .A(n5805), .B(net77038), .ZN(n9059) );
  XNOR2_X1 U7362 ( .A(n5805), .B(n10247), .ZN(n10425) );
  AND3_X4 U7364 ( .A1(\PCLOGIC/imm16_32 [16]), .A2(net77272), .A3(net78056), 
        .ZN(n5933) );
  AOI22_X1 U7365 ( .A1(\REGFILE/reg_out[19][30] ), .A2(net77814), .B1(
        \REGFILE/reg_out[1][30] ), .B2(net82631), .ZN(n6252) );
  INV_X2 U7366 ( .A(n5934), .ZN(n5935) );
  XNOR2_X1 U7367 ( .A(n5867), .B(n10375), .ZN(n10420) );
  XNOR2_X1 U7368 ( .A(n5867), .B(net77040), .ZN(n9354) );
  NAND4_X1 U7369 ( .A1(n10421), .A2(n10420), .A3(n10419), .A4(n10418), .ZN(
        n10428) );
  AOI21_X2 U7370 ( .B1(n10420), .B2(n10377), .A(n10376), .ZN(n10381) );
  NAND2_X1 U7371 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[11].MUX/N1 ), .A2(n9354), 
        .ZN(n9355) );
  INV_X2 U7372 ( .A(\REGFILE/reg_out[9][30] ), .ZN(n8757) );
  INV_X2 U7373 ( .A(\REGFILE/reg_out[1][31] ), .ZN(net70780) );
  AOI22_X1 U7374 ( .A1(\REGFILE/reg_out[19][31] ), .A2(net77814), .B1(
        \REGFILE/reg_out[1][31] ), .B2(net82631), .ZN(n6226) );
  NAND2_X1 U7375 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[14].MUX/N1 ), .A2(n5805), 
        .ZN(n10365) );
  AOI22_X4 U7376 ( .A1(\REGFILE/reg_out[31][9] ), .A2(net77666), .B1(
        \REGFILE/reg_out[3][9] ), .B2(net77676), .ZN(n6720) );
  INV_X8 U7377 ( .A(n9616), .ZN(n10910) );
  AOI22_X1 U7378 ( .A1(\REGFILE/reg_out[7][2] ), .A2(net75455), .B1(
        \REGFILE/reg_out[6][2] ), .B2(net75456), .ZN(n6865) );
  NOR2_X1 U7379 ( .A1(n10375), .A2(n10915), .ZN(n10376) );
  NAND3_X1 U7380 ( .A1(net71078), .A2(\WIRE_ALU_A/MUX2TO1_32BIT[11].MUX/N1 ), 
        .A3(n5868), .ZN(n9853) );
  XNOR2_X1 U7381 ( .A(net84663), .B(net77040), .ZN(n9060) );
  XNOR2_X1 U7382 ( .A(net84663), .B(n10368), .ZN(n10422) );
  NAND2_X1 U7383 ( .A1(n4879), .A2(\REGFILE/reg_out[2][13] ), .ZN(n9471) );
  INV_X2 U7384 ( .A(n5937), .ZN(n5938) );
  INV_X2 U7385 ( .A(n5939), .ZN(n5940) );
  AND2_X2 U7386 ( .A1(n5942), .A2(n5941), .ZN(n6640) );
  NAND3_X1 U7387 ( .A1(net71078), .A2(aluA[16]), .A3(n5769), .ZN(n9195) );
  XNOR2_X1 U7388 ( .A(n5769), .B(net77038), .ZN(n9054) );
  XNOR2_X1 U7389 ( .A(n5769), .B(aluA[16]), .ZN(n10447) );
  NAND2_X4 U7390 ( .A1(n6604), .A2(n6605), .ZN(dmem_write_out[15]) );
  AOI22_X1 U7391 ( .A1(\REGFILE/reg_out[31][1] ), .A2(net77666), .B1(
        \REGFILE/reg_out[3][1] ), .B2(n5609), .ZN(n6884) );
  AOI22_X1 U7392 ( .A1(\REGFILE/reg_out[31][3] ), .A2(net77666), .B1(
        \REGFILE/reg_out[3][3] ), .B2(n5609), .ZN(n6840) );
  NAND2_X4 U7393 ( .A1(n6628), .A2(n6629), .ZN(dmem_write_out[14]) );
  NAND2_X1 U7394 ( .A1(n10615), .A2(\REGFILE/reg_out[30][30] ), .ZN(n8754) );
  AOI22_X1 U7395 ( .A1(\REGFILE/reg_out[30][30] ), .A2(net77638), .B1(
        \REGFILE/reg_out[2][30] ), .B2(net75442), .ZN(n6267) );
  AND2_X2 U7396 ( .A1(n5946), .A2(n5945), .ZN(n6768) );
  AOI22_X2 U7397 ( .A1(\REGFILE/reg_out[30][6] ), .A2(net77634), .B1(
        \REGFILE/reg_out[2][6] ), .B2(net75442), .ZN(n6780) );
  INV_X16 U7398 ( .A(n10946), .ZN(net77104) );
  NAND3_X1 U7399 ( .A1(net71078), .A2(\WIRE_ALU_A/MUX2TO1_32BIT[12].MUX/N1 ), 
        .A3(n5577), .ZN(n9099) );
  AOI22_X1 U7400 ( .A1(\REGFILE/reg_out[0][30] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][30] ), .B2(net81764), .ZN(n6255) );
  AOI22_X1 U7401 ( .A1(\REGFILE/reg_out[0][28] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][28] ), .B2(net75464), .ZN(n6301) );
  AOI22_X1 U7402 ( .A1(\REGFILE/reg_out[0][29] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][29] ), .B2(net75464), .ZN(n6277) );
  AOI22_X1 U7403 ( .A1(\REGFILE/reg_out[0][26] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][26] ), .B2(net75464), .ZN(n6348) );
  AOI22_X1 U7404 ( .A1(\REGFILE/reg_out[0][0] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][0] ), .B2(net81764), .ZN(n6901) );
  OAI22_X1 U7405 ( .A1(n10256), .A2(net70691), .B1(n10255), .B2(n5805), .ZN(
        n10257) );
  INV_X8 U7406 ( .A(n10364), .ZN(n10916) );
  INV_X2 U7407 ( .A(\REGFILE/reg_out[10][31] ), .ZN(n10513) );
  AOI22_X1 U7408 ( .A1(\REGFILE/reg_out[0][31] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][31] ), .B2(net81764), .ZN(n6229) );
  AOI22_X2 U7409 ( .A1(\REGFILE/reg_out[16][8] ), .A2(net87506), .B1(
        \REGFILE/reg_out[15][8] ), .B2(net75468), .ZN(n6738) );
  INV_X2 U7410 ( .A(n5950), .ZN(n5951) );
  XNOR2_X1 U7411 ( .A(n5826), .B(net77040), .ZN(n9508) );
  XNOR2_X1 U7412 ( .A(n5826), .B(n10382), .ZN(n10418) );
  NOR3_X1 U7413 ( .A1(net78003), .A2(n5826), .A3(n10382), .ZN(n9337) );
  NOR2_X1 U7414 ( .A1(n10913), .A2(n10382), .ZN(n10383) );
  AOI22_X2 U7415 ( .A1(\REGFILE/reg_out[0][8] ), .A2(net120684), .B1(
        \REGFILE/reg_out[10][8] ), .B2(net75464), .ZN(n6736) );
  NOR2_X2 U7416 ( .A1(n6849), .A2(n6848), .ZN(n6850) );
  AOI22_X1 U7417 ( .A1(\REGFILE/reg_out[30][1] ), .A2(net77634), .B1(
        \REGFILE/reg_out[2][1] ), .B2(net75442), .ZN(n6890) );
  AOI22_X1 U7418 ( .A1(\REGFILE/reg_out[0][1] ), .A2(net82342), .B1(
        \REGFILE/reg_out[10][1] ), .B2(net81764), .ZN(n6878) );
  XNOR2_X1 U7419 ( .A(n5944), .B(net77038), .ZN(n9351) );
  NAND2_X1 U7420 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[12].MUX/N1 ), .A2(n5944), 
        .ZN(n10372) );
  XNOR2_X1 U7421 ( .A(n5944), .B(n9075), .ZN(n10423) );
  OAI22_X1 U7422 ( .A1(n10134), .A2(net70691), .B1(n10133), .B2(n5713), .ZN(
        n10135) );
  XNOR2_X1 U7423 ( .A(n5713), .B(net77040), .ZN(n9357) );
  NAND2_X1 U7424 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[10].MUX/N1 ), .A2(n5713), 
        .ZN(n10379) );
  XNOR2_X1 U7425 ( .A(n5713), .B(n10125), .ZN(n10421) );
  INV_X1 U7426 ( .A(n5815), .ZN(n5952) );
  INV_X4 U7427 ( .A(net78235), .ZN(net80443) );
  AOI22_X2 U7429 ( .A1(\REGFILE/reg_out[19][5] ), .A2(net77810), .B1(
        \REGFILE/reg_out[1][5] ), .B2(net82631), .ZN(n6787) );
  AOI22_X2 U7430 ( .A1(\REGFILE/reg_out[31][5] ), .A2(net77666), .B1(
        \REGFILE/reg_out[3][5] ), .B2(n5609), .ZN(n6796) );
  INV_X2 U7431 ( .A(n5956), .ZN(n5957) );
  INV_X1 U7432 ( .A(\REGFILE/reg_out[16][30] ), .ZN(n8745) );
  XNOR2_X1 U7433 ( .A(n8587), .B(n5955), .ZN(n9809) );
  NAND2_X1 U7434 ( .A1(net73708), .A2(n5955), .ZN(n8696) );
  NAND2_X1 U7435 ( .A1(n6040), .A2(n5955), .ZN(n8726) );
  NAND2_X1 U7436 ( .A1(n10542), .A2(n5955), .ZN(n8768) );
  NAND2_X1 U7437 ( .A1(n9065), .A2(n5955), .ZN(n8822) );
  AOI22_X1 U7438 ( .A1(n8974), .A2(net72962), .B1(n4912), .B2(n5955), .ZN(
        n9771) );
  NAND2_X1 U7439 ( .A1(net70720), .A2(n5955), .ZN(n9070) );
  NAND2_X1 U7440 ( .A1(net70719), .A2(n5955), .ZN(n9599) );
  INV_X1 U7441 ( .A(n5955), .ZN(n10312) );
  XNOR2_X1 U7442 ( .A(n5955), .B(n6005), .ZN(n10442) );
  NAND2_X1 U7443 ( .A1(n8588), .A2(n5955), .ZN(n8589) );
  AOI22_X2 U7444 ( .A1(\REGFILE/reg_out[19][1] ), .A2(net77810), .B1(
        \REGFILE/reg_out[1][1] ), .B2(net82631), .ZN(n6875) );
  INV_X16 U7445 ( .A(net75455), .ZN(net77720) );
  INV_X8 U7446 ( .A(n10408), .ZN(n10907) );
  AOI21_X2 U7447 ( .B1(n10407), .B2(n10406), .A(n10405), .ZN(n10410) );
  OAI21_X2 U7448 ( .B1(n10410), .B2(n10414), .A(n10409), .ZN(n10411) );
  AOI22_X2 U7449 ( .A1(\REGFILE/reg_out[21][2] ), .A2(net77842), .B1(
        \REGFILE/reg_out[20][2] ), .B2(net77850), .ZN(n6855) );
  NOR2_X1 U7450 ( .A1(n10908), .A2(n10404), .ZN(n10405) );
  NAND4_X2 U7451 ( .A1(n6868), .A2(n6869), .A3(n6867), .A4(n6866), .ZN(n6870)
         );
  NAND2_X4 U7452 ( .A1(n8539), .A2(net73496), .ZN(net73622) );
  INV_X8 U7453 ( .A(net76249), .ZN(net75475) );
  NOR2_X4 U7454 ( .A1(n6883), .A2(n6882), .ZN(n6895) );
  NAND2_X4 U7455 ( .A1(n6665), .A2(n6664), .ZN(dmem_write_out[12]) );
  NAND2_X4 U7456 ( .A1(n6687), .A2(n6686), .ZN(dmem_write_out[11]) );
  NAND2_X4 U7457 ( .A1(n6708), .A2(n6709), .ZN(dmem_write_out[10]) );
  INV_X2 U7458 ( .A(n5959), .ZN(n5960) );
  OAI22_X1 U7459 ( .A1(net73608), .A2(n8823), .B1(n10319), .B2(n8634), .ZN(
        n8974) );
  AOI21_X1 U7460 ( .B1(n10305), .B2(n10304), .A(net73608), .ZN(n10461) );
  INV_X2 U7461 ( .A(n5961), .ZN(n5962) );
  AOI21_X1 U7462 ( .B1(n6019), .B2(n8401), .A(n8400), .ZN(n8415) );
  NOR2_X4 U7463 ( .A1(n6952), .A2(n6951), .ZN(n6953) );
  INV_X2 U7464 ( .A(n5963), .ZN(n5964) );
  INV_X2 U7465 ( .A(n5965), .ZN(n5966) );
  INV_X2 U7466 ( .A(n5967), .ZN(n5968) );
  INV_X2 U7467 ( .A(n5969), .ZN(n5970) );
  XNOR2_X1 U7468 ( .A(n5758), .B(n9535), .ZN(n10419) );
  XNOR2_X1 U7469 ( .A(n5758), .B(net77040), .ZN(n9609) );
  OAI22_X1 U7470 ( .A1(n9513), .A2(net70691), .B1(n9512), .B2(n5758), .ZN(
        n9514) );
  NAND2_X1 U7471 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[8].MUX/N1 ), .A2(n5758), .ZN(
        n10386) );
  XNOR2_X1 U7472 ( .A(n9609), .B(n9535), .ZN(n9610) );
  INV_X2 U7473 ( .A(n5971), .ZN(n5972) );
  NOR2_X1 U7474 ( .A1(net73842), .A2(net73848), .ZN(n8405) );
  NOR3_X2 U7475 ( .A1(n8406), .A2(n8405), .A3(n8404), .ZN(n8414) );
  INV_X2 U7476 ( .A(n5973), .ZN(n5974) );
  AOI22_X4 U7477 ( .A1(n5923), .A2(net77444), .B1(n5966), .B2(net77400), .ZN(
        n6936) );
  INV_X1 U7478 ( .A(net80390), .ZN(net73848) );
  AOI22_X1 U7479 ( .A1(\REGFILE/reg_out[4][0] ), .A2(n5678), .B1(
        \REGFILE/reg_out[5][0] ), .B2(net84475), .ZN(n6908) );
  AOI22_X4 U7480 ( .A1(\REGFILE/reg_out[29][8] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][8] ), .B2(n6911), .ZN(n6749) );
  OAI22_X1 U7481 ( .A1(n9666), .A2(net70691), .B1(n9665), .B2(n5757), .ZN(
        n9667) );
  XNOR2_X1 U7482 ( .A(n5757), .B(net77040), .ZN(n9615) );
  NAND2_X1 U7483 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[6].MUX/N1 ), .A2(n5757), .ZN(
        n10393) );
  XNOR2_X1 U7484 ( .A(n5757), .B(n9656), .ZN(n9657) );
  NAND2_X2 U7485 ( .A1(\REGFILE/reg_out[19][4] ), .A2(net77810), .ZN(n5975) );
  NAND2_X1 U7486 ( .A1(\REGFILE/reg_out[1][4] ), .A2(net75478), .ZN(n5976) );
  AND2_X2 U7487 ( .A1(n5975), .A2(n5976), .ZN(n6809) );
  NOR2_X4 U7488 ( .A1(n5815), .A2(n6946), .ZN(n6954) );
  INV_X2 U7489 ( .A(\REGFILE/reg_out[8][30] ), .ZN(n8756) );
  AOI22_X1 U7490 ( .A1(\REGFILE/reg_out[9][30] ), .A2(net77702), .B1(
        \REGFILE/reg_out[8][30] ), .B2(n4829), .ZN(n6263) );
  NAND2_X1 U7491 ( .A1(\REGFILE/reg_out[3][3] ), .A2(net77410), .ZN(n8136) );
  NAND2_X1 U7493 ( .A1(\REGFILE/reg_out[1][4] ), .A2(net77518), .ZN(n8087) );
  INV_X2 U7496 ( .A(n5985), .ZN(n5986) );
  OR2_X2 U7497 ( .A1(n5987), .A2(net77542), .ZN(n6972) );
  INV_X16 U7498 ( .A(net74051), .ZN(net77542) );
  NAND2_X1 U7499 ( .A1(net76488), .A2(\REGFILE/reg_out[31][29] ), .ZN(n9831)
         );
  AOI22_X1 U7500 ( .A1(\REGFILE/reg_out[31][29] ), .A2(net77670), .B1(
        \REGFILE/reg_out[3][29] ), .B2(n5609), .ZN(n6283) );
  INV_X1 U7501 ( .A(\REGFILE/reg_out[23][29] ), .ZN(net71824) );
  AOI22_X1 U7502 ( .A1(\REGFILE/reg_out[23][29] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][29] ), .B2(net77834), .ZN(n6275) );
  INV_X2 U7503 ( .A(n5989), .ZN(n5990) );
  INV_X1 U7504 ( .A(\REGFILE/reg_out[15][29] ), .ZN(n9828) );
  AOI22_X1 U7505 ( .A1(\REGFILE/reg_out[21][29] ), .A2(net77846), .B1(
        \REGFILE/reg_out[20][29] ), .B2(net77854), .ZN(n6276) );
  INV_X1 U7506 ( .A(\REGFILE/reg_out[28][29] ), .ZN(n10934) );
  AOI22_X1 U7507 ( .A1(\REGFILE/reg_out[29][29] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][29] ), .B2(n6911), .ZN(n6290) );
  AOI22_X1 U7508 ( .A1(\REGFILE/reg_out[19][0] ), .A2(net77810), .B1(
        \REGFILE/reg_out[1][0] ), .B2(net82631), .ZN(n6898) );
  AOI22_X1 U7509 ( .A1(\REGFILE/reg_out[31][0] ), .A2(net77666), .B1(
        \REGFILE/reg_out[3][0] ), .B2(n5609), .ZN(n6907) );
  AOI22_X1 U7510 ( .A1(\REGFILE/reg_out[31][2] ), .A2(net77666), .B1(
        \REGFILE/reg_out[3][2] ), .B2(n5609), .ZN(n6862) );
  AOI22_X1 U7511 ( .A1(\REGFILE/reg_out[31][4] ), .A2(net77666), .B1(n5982), 
        .B2(n5609), .ZN(n6818) );
  INV_X8 U7512 ( .A(n9358), .ZN(n10913) );
  AOI22_X2 U7513 ( .A1(\REGFILE/reg_out[31][6] ), .A2(net77666), .B1(
        \REGFILE/reg_out[3][6] ), .B2(n5609), .ZN(n6774) );
  AOI22_X2 U7514 ( .A1(\REGFILE/reg_out[17][6] ), .A2(net77794), .B1(
        \REGFILE/reg_out[18][6] ), .B2(n5890), .ZN(n6764) );
  NOR2_X4 U7515 ( .A1(n6817), .A2(n6816), .ZN(n6829) );
  NAND2_X4 U7516 ( .A1(n6248), .A2(n4865), .ZN(net73629) );
  INV_X32 U7517 ( .A(instruction[4]), .ZN(net73498) );
  INV_X8 U7518 ( .A(net76211), .ZN(net76195) );
  NAND2_X4 U7519 ( .A1(\REGFILE/reg_out[24][29] ), .A2(net77318), .ZN(n6985)
         );
  NAND2_X4 U7520 ( .A1(n6785), .A2(n6784), .ZN(dmem_write_out[6]) );
  NAND2_X4 U7521 ( .A1(n6873), .A2(n6872), .ZN(dmem_write_out[2]) );
  NOR3_X1 U7522 ( .A1(n8451), .A2(n5748), .A3(n8450), .ZN(n8452) );
  AOI22_X1 U7523 ( .A1(\REGFILE/reg_out[24][31] ), .A2(net77602), .B1(
        \REGFILE/reg_out[25][31] ), .B2(net77610), .ZN(n6240) );
  XNOR2_X1 U7524 ( .A(n8584), .B(net80189), .ZN(n8583) );
  INV_X4 U7525 ( .A(net78107), .ZN(net75401) );
  INV_X2 U7526 ( .A(n5992), .ZN(n5993) );
  AOI22_X1 U7527 ( .A1(net77588), .A2(n4834), .B1(n8411), .B2(n5952), .ZN(
        n8412) );
  AOI22_X4 U7528 ( .A1(n5830), .A2(net77478), .B1(n5993), .B2(net77550), .ZN(
        n6949) );
  INV_X1 U7529 ( .A(n6952), .ZN(n5998) );
  NAND2_X1 U7530 ( .A1(net73708), .A2(net80189), .ZN(n10655) );
  NAND3_X2 U7531 ( .A1(n10470), .A2(net80189), .A3(n10542), .ZN(n10471) );
  NAND2_X1 U7532 ( .A1(n9065), .A2(net80189), .ZN(n8827) );
  NAND2_X1 U7533 ( .A1(n4912), .A2(net80189), .ZN(n8767) );
  INV_X4 U7534 ( .A(n6001), .ZN(n6930) );
  INV_X2 U7535 ( .A(\REGFILE/reg_out[4][31] ), .ZN(net70757) );
  AOI22_X1 U7536 ( .A1(\REGFILE/reg_out[4][31] ), .A2(net75451), .B1(
        \REGFILE/reg_out[5][31] ), .B2(net75452), .ZN(n6236) );
  INV_X1 U7537 ( .A(\REGFILE/reg_out[2][31] ), .ZN(net70761) );
  AOI22_X1 U7538 ( .A1(\REGFILE/reg_out[30][31] ), .A2(net84761), .B1(
        \REGFILE/reg_out[2][31] ), .B2(net75442), .ZN(n6242) );
  INV_X16 U7539 ( .A(net70537), .ZN(net76508) );
  INV_X16 U7540 ( .A(net75419), .ZN(net74051) );
  NAND2_X4 U7541 ( .A1(n5574), .A2(\PCLOGIC/imm26_32 [12]), .ZN(net76242) );
  NOR2_X4 U7542 ( .A1(n6893), .A2(n6892), .ZN(n6894) );
  NOR2_X2 U7543 ( .A1(n8409), .A2(n5820), .ZN(n8404) );
  NAND4_X2 U7544 ( .A1(n6881), .A2(n6880), .A3(n6879), .A4(n6878), .ZN(n6882)
         );
  NAND2_X4 U7545 ( .A1(\PCLOGIC/imm26_32 [11]), .A2(\PCLOGIC/imm26_32 [12]), 
        .ZN(net76211) );
  XNOR2_X1 U7546 ( .A(net70921), .B(net77040), .ZN(net70734) );
  NAND2_X1 U7547 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[1].MUX/N1 ), .A2(net70921), 
        .ZN(n10412) );
  XNOR2_X1 U7548 ( .A(net70921), .B(net71273), .ZN(n10164) );
  NAND2_X1 U7549 ( .A1(n5798), .A2(net71026), .ZN(n10309) );
  NAND2_X1 U7550 ( .A1(net70719), .A2(n5798), .ZN(n9619) );
  NAND2_X1 U7551 ( .A1(net70720), .A2(n5798), .ZN(n9078) );
  NAND2_X1 U7552 ( .A1(n9065), .A2(n5798), .ZN(n8841) );
  NAND2_X1 U7553 ( .A1(n4912), .A2(n5798), .ZN(n8765) );
  INV_X1 U7554 ( .A(n5798), .ZN(n8729) );
  NAND2_X1 U7555 ( .A1(net73708), .A2(n5798), .ZN(n8703) );
  XNOR2_X1 U7556 ( .A(n8585), .B(n5798), .ZN(n8706) );
  AOI22_X4 U7557 ( .A1(n8401), .A2(n6933), .B1(n8403), .B2(n6932), .ZN(
        net75397) );
  NAND3_X4 U7558 ( .A1(net74011), .A2(net73503), .A3(net73170), .ZN(net78055)
         );
  NAND3_X4 U7559 ( .A1(net74011), .A2(net73503), .A3(net73170), .ZN(net78056)
         );
  INV_X32 U7560 ( .A(n6004), .ZN(n6005) );
  INV_X16 U7561 ( .A(n10327), .ZN(n10930) );
  NAND2_X4 U7562 ( .A1(net74009), .A2(\PCLOGIC/imm16_32 [16]), .ZN(net73878)
         );
  NAND4_X4 U7563 ( .A1(n8572), .A2(n8571), .A3(n8570), .A4(n8569), .ZN(n10494)
         );
  INV_X16 U7564 ( .A(n6005), .ZN(n10099) );
  INV_X16 U7565 ( .A(net78051), .ZN(net71026) );
  INV_X8 U7566 ( .A(n9803), .ZN(n10058) );
  INV_X16 U7567 ( .A(n9094), .ZN(n9065) );
  INV_X8 U7568 ( .A(net70866), .ZN(net70719) );
  NAND2_X4 U7569 ( .A1(n10494), .A2(n10470), .ZN(n10472) );
  INV_X8 U7570 ( .A(net70710), .ZN(n10064) );
  INV_X8 U7571 ( .A(n9606), .ZN(n10066) );
  INV_X8 U7572 ( .A(net70710), .ZN(net71094) );
  INV_X8 U7573 ( .A(n9854), .ZN(net71092) );
  INV_X8 U7574 ( .A(n9012), .ZN(n10280) );
  INV_X32 U7575 ( .A(net75482), .ZN(net77856) );
  INV_X32 U7576 ( .A(net77704), .ZN(net77700) );
  INV_X32 U7577 ( .A(net77656), .ZN(net77650) );
  INV_X32 U7578 ( .A(net77656), .ZN(net77652) );
  INV_X32 U7579 ( .A(n6013), .ZN(n6011) );
  INV_X32 U7580 ( .A(net77548), .ZN(net77544) );
  INV_X32 U7581 ( .A(net77542), .ZN(net77514) );
  INV_X32 U7582 ( .A(net77540), .ZN(net77518) );
  INV_X32 U7583 ( .A(net77540), .ZN(net77520) );
  INV_X32 U7584 ( .A(net77540), .ZN(net77522) );
  INV_X32 U7585 ( .A(net77538), .ZN(net77524) );
  INV_X32 U7586 ( .A(net77538), .ZN(net77526) );
  INV_X32 U7587 ( .A(net77538), .ZN(net77528) );
  INV_X32 U7588 ( .A(net77538), .ZN(net77530) );
  INV_X32 U7589 ( .A(net77548), .ZN(net77532) );
  INV_X32 U7590 ( .A(net77544), .ZN(net77538) );
  INV_X32 U7591 ( .A(net77544), .ZN(net77540) );
  INV_X32 U7592 ( .A(net77502), .ZN(net77488) );
  INV_X32 U7593 ( .A(net77502), .ZN(net77490) );
  INV_X32 U7594 ( .A(net77502), .ZN(net77492) );
  INV_X32 U7595 ( .A(net77508), .ZN(net77500) );
  INV_X32 U7596 ( .A(net77464), .ZN(net77462) );
  INV_X32 U7597 ( .A(net77474), .ZN(net77464) );
  INV_X32 U7598 ( .A(net77428), .ZN(net77426) );
  INV_X32 U7599 ( .A(net77396), .ZN(net77376) );
  INV_X32 U7600 ( .A(net77360), .ZN(net77342) );
  INV_X32 U7601 ( .A(net77358), .ZN(net77344) );
  INV_X32 U7602 ( .A(net77358), .ZN(net77346) );
  INV_X32 U7603 ( .A(net77358), .ZN(net77348) );
  INV_X32 U7604 ( .A(n6018), .ZN(n6015) );
  INV_X32 U7605 ( .A(n6018), .ZN(n6016) );
  INV_X32 U7606 ( .A(n6018), .ZN(n6017) );
  INV_X32 U7607 ( .A(n6014), .ZN(n6018) );
  INV_X32 U7608 ( .A(n6020), .ZN(n6019) );
  INV_X32 U7609 ( .A(n6022), .ZN(n6021) );
  INV_X32 U7610 ( .A(n6028), .ZN(n6027) );
  INV_X32 U7611 ( .A(n6031), .ZN(n6029) );
  INV_X32 U7612 ( .A(n6031), .ZN(n6030) );
  INV_X32 U7613 ( .A(n4964), .ZN(n6032) );
  INV_X32 U7614 ( .A(n6039), .ZN(n6038) );
  INV_X32 U7615 ( .A(n6052), .ZN(n6051) );
  INV_X32 U7616 ( .A(n6061), .ZN(n6059) );
  INV_X32 U7617 ( .A(n6061), .ZN(n6060) );
  INV_X32 U7618 ( .A(n6064), .ZN(n6062) );
  INV_X32 U7619 ( .A(n6064), .ZN(n6063) );
  INV_X32 U7620 ( .A(n6077), .ZN(n6075) );
  INV_X32 U7621 ( .A(n6077), .ZN(n6076) );
  INV_X32 U7622 ( .A(n4965), .ZN(n6087) );
  INV_X32 U7623 ( .A(net77042), .ZN(net77038) );
  INV_X32 U7624 ( .A(net77042), .ZN(net77040) );
  INV_X32 U7625 ( .A(net76514), .ZN(net76510) );
  INV_X32 U7627 ( .A(net76508), .ZN(net76506) );
  INV_X32 U7628 ( .A(n10511), .ZN(n6191) );
  INV_X32 U7629 ( .A(n5012), .ZN(n6221) );
  INV_X32 U7630 ( .A(n5013), .ZN(n6222) );
  INV_X32 U7631 ( .A(n5011), .ZN(n6223) );
  NAND3_X4 U7632 ( .A1(net92447), .A2(net86793), .A3(\PCLOGIC/imm26_32 [13]), 
        .ZN(net76259) );
  NAND3_X4 U7633 ( .A1(\PCLOGIC/imm26_32 [15]), .A2(\PCLOGIC/imm26_32 [14]), 
        .A3(\PCLOGIC/imm26_32 [13]), .ZN(net76217) );
  NAND3_X4 U7634 ( .A1(net87495), .A2(net82739), .A3(\PCLOGIC/imm26_32 [14]), 
        .ZN(net76248) );
  NAND4_X2 U7635 ( .A1(n6228), .A2(n6227), .A3(n6226), .A4(n6225), .ZN(n6234)
         );
  NAND4_X2 U7636 ( .A1(n6232), .A2(n6231), .A3(n6230), .A4(n6229), .ZN(n6233)
         );
  NOR2_X4 U7637 ( .A1(n6234), .A2(n6233), .ZN(n6247) );
  AOI22_X2 U7638 ( .A1(\REGFILE/reg_out[31][31] ), .A2(net77670), .B1(
        \REGFILE/reg_out[3][31] ), .B2(n5609), .ZN(n6235) );
  NAND4_X2 U7639 ( .A1(n6238), .A2(n6237), .A3(n6236), .A4(n6235), .ZN(n6245)
         );
  NAND4_X2 U7640 ( .A1(n6243), .A2(n6242), .A3(n6241), .A4(n6240), .ZN(n6244)
         );
  NOR2_X4 U7641 ( .A1(n6245), .A2(n6244), .ZN(n6246) );
  NAND2_X2 U7642 ( .A1(n6247), .A2(n6246), .ZN(dmem_write_out[31]) );
  INV_X4 U7643 ( .A(dmem_write_out[31]), .ZN(n6250) );
  NOR2_X4 U7644 ( .A1(instruction[1]), .A2(instruction[0]), .ZN(n6248) );
  NAND3_X4 U7645 ( .A1(net74011), .A2(net73503), .A3(net73170), .ZN(net73697)
         );
  NAND2_X2 U7646 ( .A1(\PCLOGIC/imm16_32 [31]), .A2(net75844), .ZN(n6249) );
  OAI21_X4 U7647 ( .B1(n6250), .B2(net78055), .A(n6249), .ZN(n10928) );
  AOI22_X2 U7648 ( .A1(\REGFILE/reg_out[21][30] ), .A2(net77846), .B1(
        \REGFILE/reg_out[20][30] ), .B2(net77854), .ZN(n6254) );
  AOI22_X2 U7649 ( .A1(\REGFILE/reg_out[23][30] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][30] ), .B2(net77836), .ZN(n6253) );
  NAND4_X2 U7650 ( .A1(n6254), .A2(n6253), .A3(n6252), .A4(n6251), .ZN(n6260)
         );
  AOI22_X2 U7651 ( .A1(\REGFILE/reg_out[14][30] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][30] ), .B2(n6009), .ZN(n6258) );
  NAND4_X2 U7652 ( .A1(n6255), .A2(n6257), .A3(n6256), .A4(n6258), .ZN(n6259)
         );
  AOI22_X2 U7653 ( .A1(n5672), .A2(n5679), .B1(\REGFILE/reg_out[5][30] ), .B2(
        net84475), .ZN(n6262) );
  NAND4_X2 U7654 ( .A1(n6264), .A2(n6263), .A3(n6262), .A4(n6261), .ZN(n6270)
         );
  NAND4_X2 U7655 ( .A1(n6265), .A2(n6267), .A3(n6266), .A4(n6268), .ZN(n6269)
         );
  NOR2_X4 U7656 ( .A1(n6270), .A2(n6269), .ZN(n6271) );
  NAND2_X2 U7657 ( .A1(n6272), .A2(n6271), .ZN(dmem_write_out[30]) );
  INV_X4 U7658 ( .A(dmem_write_out[30]), .ZN(net76154) );
  NAND4_X2 U7659 ( .A1(n6276), .A2(n6275), .A3(n6274), .A4(n6273), .ZN(n6282)
         );
  AOI22_X2 U7660 ( .A1(\REGFILE/reg_out[14][29] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][29] ), .B2(n5663), .ZN(n6280) );
  NAND4_X2 U7661 ( .A1(n6280), .A2(n6279), .A3(n6278), .A4(n6277), .ZN(n6281)
         );
  NOR2_X4 U7662 ( .A1(n6282), .A2(n6281), .ZN(n6294) );
  NAND4_X2 U7663 ( .A1(n6286), .A2(n6285), .A3(n6284), .A4(n6283), .ZN(n6292)
         );
  NAND4_X2 U7664 ( .A1(n6288), .A2(n6289), .A3(n6290), .A4(n6287), .ZN(n6291)
         );
  NOR2_X4 U7665 ( .A1(n6292), .A2(n6291), .ZN(n6293) );
  NAND2_X2 U7666 ( .A1(n6294), .A2(n6293), .ZN(dmem_write_out[29]) );
  INV_X4 U7667 ( .A(dmem_write_out[29]), .ZN(n6296) );
  NAND2_X2 U7668 ( .A1(net75844), .A2(\PCLOGIC/imm16_32 [29]), .ZN(n6295) );
  AOI22_X2 U7669 ( .A1(\REGFILE/reg_out[21][28] ), .A2(net77846), .B1(
        \REGFILE/reg_out[20][28] ), .B2(net77854), .ZN(n6300) );
  AOI22_X2 U7670 ( .A1(\REGFILE/reg_out[23][28] ), .A2(net77828), .B1(
        \REGFILE/reg_out[22][28] ), .B2(net77834), .ZN(n6299) );
  NAND4_X2 U7671 ( .A1(n6300), .A2(n6299), .A3(n6298), .A4(n6297), .ZN(n6306)
         );
  NAND4_X2 U7672 ( .A1(n6304), .A2(n6303), .A3(n6302), .A4(n6301), .ZN(n6305)
         );
  NOR2_X4 U7673 ( .A1(n6306), .A2(n6305), .ZN(n6318) );
  AOI22_X2 U7674 ( .A1(\REGFILE/reg_out[4][28] ), .A2(net75451), .B1(
        \REGFILE/reg_out[5][28] ), .B2(net84475), .ZN(n6308) );
  AOI22_X2 U7675 ( .A1(\REGFILE/reg_out[31][28] ), .A2(net77670), .B1(
        \REGFILE/reg_out[3][28] ), .B2(n5609), .ZN(n6307) );
  NAND4_X2 U7676 ( .A1(n6310), .A2(n6309), .A3(n6308), .A4(n6307), .ZN(n6316)
         );
  NAND4_X2 U7677 ( .A1(n6312), .A2(n6311), .A3(n6314), .A4(n6313), .ZN(n6315)
         );
  NOR2_X4 U7678 ( .A1(n6316), .A2(n6315), .ZN(n6317) );
  NAND2_X2 U7679 ( .A1(n6318), .A2(n6317), .ZN(dmem_write_out[28]) );
  INV_X4 U7680 ( .A(dmem_write_out[28]), .ZN(n6320) );
  NAND2_X2 U7681 ( .A1(net75844), .A2(\PCLOGIC/imm16_32 [28]), .ZN(n6319) );
  OAI21_X4 U7682 ( .B1(n6320), .B2(net78055), .A(n6319), .ZN(n10926) );
  AOI22_X2 U7683 ( .A1(\REGFILE/reg_out[21][27] ), .A2(net77846), .B1(
        \REGFILE/reg_out[20][27] ), .B2(net77854), .ZN(n6324) );
  AOI22_X2 U7684 ( .A1(\REGFILE/reg_out[23][27] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][27] ), .B2(net77836), .ZN(n6323) );
  NAND4_X2 U7685 ( .A1(n6324), .A2(n6323), .A3(n6322), .A4(n6321), .ZN(n6330)
         );
  AOI22_X2 U7686 ( .A1(\REGFILE/reg_out[14][27] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][27] ), .B2(n5663), .ZN(n6328) );
  NAND4_X2 U7687 ( .A1(n6328), .A2(n6327), .A3(n6326), .A4(n6325), .ZN(n6329)
         );
  NOR2_X4 U7688 ( .A1(n6330), .A2(n6329), .ZN(n6342) );
  AOI22_X2 U7689 ( .A1(\REGFILE/reg_out[9][27] ), .A2(net77702), .B1(
        \REGFILE/reg_out[8][27] ), .B2(n4829), .ZN(n6333) );
  AOI22_X2 U7690 ( .A1(\REGFILE/reg_out[4][27] ), .A2(n5679), .B1(
        \REGFILE/reg_out[5][27] ), .B2(net84475), .ZN(n6332) );
  AOI22_X2 U7691 ( .A1(\REGFILE/reg_out[31][27] ), .A2(net77670), .B1(
        \REGFILE/reg_out[3][27] ), .B2(n5609), .ZN(n6331) );
  NAND4_X2 U7692 ( .A1(n6334), .A2(n6333), .A3(n6332), .A4(n6331), .ZN(n6340)
         );
  AOI22_X2 U7693 ( .A1(\REGFILE/reg_out[24][27] ), .A2(net77602), .B1(
        \REGFILE/reg_out[25][27] ), .B2(net77614), .ZN(n6335) );
  NAND4_X2 U7694 ( .A1(n6335), .A2(n6337), .A3(n6336), .A4(n6338), .ZN(n6339)
         );
  INV_X4 U7695 ( .A(\PCLOGIC/imm16_32 [27]), .ZN(net73696) );
  NAND2_X2 U7696 ( .A1(net75844), .A2(net73696), .ZN(n6343) );
  OAI21_X4 U7697 ( .B1(dmem_write_out[27]), .B2(net78056), .A(n6343), .ZN(
        n8885) );
  AOI22_X2 U7698 ( .A1(\REGFILE/reg_out[21][26] ), .A2(net77846), .B1(
        \REGFILE/reg_out[20][26] ), .B2(net77854), .ZN(n6347) );
  AOI22_X2 U7699 ( .A1(\REGFILE/reg_out[23][26] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][26] ), .B2(net77834), .ZN(n6346) );
  NAND4_X2 U7700 ( .A1(n6347), .A2(n6346), .A3(n6345), .A4(n6344), .ZN(n6353)
         );
  AOI22_X2 U7701 ( .A1(\REGFILE/reg_out[14][26] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][26] ), .B2(n5663), .ZN(n6351) );
  NAND4_X2 U7702 ( .A1(n6351), .A2(n6350), .A3(n6349), .A4(n6348), .ZN(n6352)
         );
  NOR2_X4 U7703 ( .A1(n6353), .A2(n6352), .ZN(n6365) );
  AOI22_X2 U7704 ( .A1(\REGFILE/reg_out[31][26] ), .A2(net77670), .B1(
        \REGFILE/reg_out[3][26] ), .B2(n5609), .ZN(n6354) );
  NAND4_X2 U7705 ( .A1(n6357), .A2(n6356), .A3(n6355), .A4(n6354), .ZN(n6363)
         );
  NAND4_X2 U7706 ( .A1(n6361), .A2(n6360), .A3(n6359), .A4(n6358), .ZN(n6362)
         );
  NAND2_X2 U7707 ( .A1(n6365), .A2(n6364), .ZN(dmem_write_out[26]) );
  INV_X4 U7708 ( .A(dmem_write_out[26]), .ZN(n6367) );
  NAND2_X2 U7709 ( .A1(net75844), .A2(\PCLOGIC/imm16_32 [26]), .ZN(n6366) );
  OAI21_X4 U7710 ( .B1(n6367), .B2(net73697), .A(n6366), .ZN(n10925) );
  AOI22_X2 U7711 ( .A1(\REGFILE/reg_out[21][25] ), .A2(net77846), .B1(
        \REGFILE/reg_out[20][25] ), .B2(net77854), .ZN(n6371) );
  AOI22_X2 U7712 ( .A1(\REGFILE/reg_out[23][25] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][25] ), .B2(net77836), .ZN(n6370) );
  NAND4_X2 U7713 ( .A1(n6371), .A2(n6370), .A3(n6369), .A4(n6368), .ZN(n6377)
         );
  AOI22_X2 U7714 ( .A1(\REGFILE/reg_out[14][25] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][25] ), .B2(n5663), .ZN(n6375) );
  NAND4_X2 U7715 ( .A1(n6372), .A2(n6373), .A3(n6375), .A4(n6374), .ZN(n6376)
         );
  AOI22_X2 U7716 ( .A1(\REGFILE/reg_out[4][25] ), .A2(n5679), .B1(
        \REGFILE/reg_out[5][25] ), .B2(net84475), .ZN(n6379) );
  AOI22_X2 U7717 ( .A1(\REGFILE/reg_out[31][25] ), .A2(net77670), .B1(
        \REGFILE/reg_out[3][25] ), .B2(n5609), .ZN(n6378) );
  NAND4_X2 U7718 ( .A1(n6380), .A2(n6381), .A3(n6379), .A4(n6378), .ZN(n6387)
         );
  NAND4_X2 U7719 ( .A1(n6384), .A2(n6385), .A3(n6383), .A4(n6382), .ZN(n6386)
         );
  NAND2_X2 U7720 ( .A1(n6389), .A2(n6388), .ZN(dmem_write_out[25]) );
  INV_X4 U7721 ( .A(dmem_write_out[25]), .ZN(n6391) );
  NAND2_X2 U7722 ( .A1(\PCLOGIC/imm16_32 [25]), .A2(net75844), .ZN(n6390) );
  OAI21_X4 U7723 ( .B1(n6391), .B2(net78055), .A(n6390), .ZN(n10924) );
  AOI22_X2 U7724 ( .A1(\REGFILE/reg_out[21][24] ), .A2(net77846), .B1(
        \REGFILE/reg_out[20][24] ), .B2(net77854), .ZN(net76031) );
  AOI22_X2 U7725 ( .A1(\REGFILE/reg_out[23][24] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][24] ), .B2(net77836), .ZN(net76032) );
  AOI22_X2 U7726 ( .A1(\REGFILE/reg_out[14][24] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][24] ), .B2(n5663), .ZN(n6395) );
  AOI22_X2 U7727 ( .A1(\REGFILE/reg_out[16][24] ), .A2(net77764), .B1(
        \REGFILE/reg_out[15][24] ), .B2(n5579), .ZN(n6394) );
  NOR2_X4 U7728 ( .A1(net76025), .A2(n6396), .ZN(n6408) );
  AOI22_X2 U7729 ( .A1(\REGFILE/reg_out[9][24] ), .A2(net77702), .B1(
        \REGFILE/reg_out[8][24] ), .B2(n4829), .ZN(n6399) );
  AOI22_X2 U7730 ( .A1(\REGFILE/reg_out[4][24] ), .A2(n5678), .B1(
        \REGFILE/reg_out[5][24] ), .B2(net84475), .ZN(n6398) );
  AOI22_X2 U7731 ( .A1(\REGFILE/reg_out[31][24] ), .A2(net77670), .B1(
        \REGFILE/reg_out[3][24] ), .B2(n5609), .ZN(n6397) );
  NAND4_X2 U7732 ( .A1(n6400), .A2(n6399), .A3(n6398), .A4(n6397), .ZN(n6406)
         );
  AOI22_X2 U7733 ( .A1(\REGFILE/reg_out[29][24] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][24] ), .B2(n6911), .ZN(n6404) );
  AOI22_X2 U7734 ( .A1(\REGFILE/reg_out[24][24] ), .A2(net75437), .B1(
        \REGFILE/reg_out[25][24] ), .B2(net75438), .ZN(n6401) );
  NAND4_X2 U7735 ( .A1(n6404), .A2(n6403), .A3(n6402), .A4(n6401), .ZN(n6405)
         );
  NAND2_X2 U7736 ( .A1(\PCLOGIC/imm16_32 [24]), .A2(net75844), .ZN(n6409) );
  OAI21_X4 U7737 ( .B1(n6410), .B2(net78056), .A(n6409), .ZN(n10923) );
  AOI22_X2 U7738 ( .A1(\REGFILE/reg_out[21][23] ), .A2(net77846), .B1(
        \REGFILE/reg_out[20][23] ), .B2(net77854), .ZN(n6414) );
  AOI22_X2 U7739 ( .A1(\REGFILE/reg_out[23][23] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][23] ), .B2(net77836), .ZN(n6413) );
  AOI22_X2 U7740 ( .A1(\REGFILE/reg_out[19][23] ), .A2(net77814), .B1(
        \REGFILE/reg_out[1][23] ), .B2(net82631), .ZN(n6412) );
  NAND4_X2 U7741 ( .A1(n6414), .A2(n6413), .A3(n6412), .A4(n6411), .ZN(n6420)
         );
  AOI22_X2 U7742 ( .A1(\REGFILE/reg_out[16][23] ), .A2(net87506), .B1(
        \REGFILE/reg_out[15][23] ), .B2(n5579), .ZN(n6417) );
  NAND4_X2 U7743 ( .A1(n6415), .A2(n6417), .A3(n6416), .A4(n6418), .ZN(n6419)
         );
  AOI22_X2 U7744 ( .A1(\REGFILE/reg_out[9][23] ), .A2(net77702), .B1(
        \REGFILE/reg_out[8][23] ), .B2(n4829), .ZN(n6423) );
  AOI22_X2 U7745 ( .A1(\REGFILE/reg_out[4][23] ), .A2(n5679), .B1(
        \REGFILE/reg_out[5][23] ), .B2(net84475), .ZN(n6422) );
  AOI22_X2 U7746 ( .A1(\REGFILE/reg_out[31][23] ), .A2(net77670), .B1(
        \REGFILE/reg_out[3][23] ), .B2(n5609), .ZN(n6421) );
  NAND4_X2 U7747 ( .A1(n6424), .A2(n6423), .A3(n6422), .A4(n6421), .ZN(n6429)
         );
  AOI22_X2 U7748 ( .A1(\REGFILE/reg_out[29][23] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][23] ), .B2(n6911), .ZN(n6427) );
  NAND2_X2 U7749 ( .A1(\PCLOGIC/imm16_32 [23]), .A2(net75844), .ZN(n6432) );
  OAI21_X4 U7750 ( .B1(n6433), .B2(net73697), .A(n6432), .ZN(n10922) );
  AOI22_X2 U7751 ( .A1(\REGFILE/reg_out[21][22] ), .A2(net77846), .B1(
        \REGFILE/reg_out[20][22] ), .B2(net77854), .ZN(n6437) );
  AOI22_X2 U7752 ( .A1(\REGFILE/reg_out[23][22] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][22] ), .B2(net77836), .ZN(n6436) );
  AOI22_X2 U7753 ( .A1(\REGFILE/reg_out[19][22] ), .A2(net77814), .B1(
        \REGFILE/reg_out[1][22] ), .B2(net75478), .ZN(n6435) );
  NAND4_X2 U7754 ( .A1(n6437), .A2(n6436), .A3(n6435), .A4(n6434), .ZN(n6443)
         );
  AOI22_X2 U7755 ( .A1(\REGFILE/reg_out[14][22] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][22] ), .B2(n5663), .ZN(n6441) );
  AOI22_X2 U7756 ( .A1(\REGFILE/reg_out[7][22] ), .A2(net77716), .B1(
        \REGFILE/reg_out[6][22] ), .B2(net75456), .ZN(n6447) );
  AOI22_X2 U7757 ( .A1(\REGFILE/reg_out[9][22] ), .A2(net77702), .B1(
        \REGFILE/reg_out[8][22] ), .B2(n4829), .ZN(n6446) );
  AOI22_X2 U7758 ( .A1(\REGFILE/reg_out[4][22] ), .A2(n5679), .B1(
        \REGFILE/reg_out[5][22] ), .B2(net84475), .ZN(n6445) );
  AOI22_X2 U7759 ( .A1(\REGFILE/reg_out[31][22] ), .A2(net77670), .B1(
        \REGFILE/reg_out[3][22] ), .B2(n5609), .ZN(n6444) );
  NAND4_X2 U7760 ( .A1(n6447), .A2(n6446), .A3(n6444), .A4(n6445), .ZN(n6453)
         );
  AOI22_X2 U7761 ( .A1(\REGFILE/reg_out[29][22] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][22] ), .B2(n6911), .ZN(n6451) );
  AOI22_X2 U7762 ( .A1(\REGFILE/reg_out[30][22] ), .A2(net77638), .B1(
        \REGFILE/reg_out[2][22] ), .B2(net82613), .ZN(n6450) );
  NAND2_X2 U7763 ( .A1(\PCLOGIC/imm16_32 [22]), .A2(net75844), .ZN(n6456) );
  OAI21_X4 U7764 ( .B1(n6457), .B2(net78055), .A(n6456), .ZN(n10921) );
  AOI22_X2 U7765 ( .A1(\REGFILE/reg_out[21][21] ), .A2(net77844), .B1(
        \REGFILE/reg_out[20][21] ), .B2(net77852), .ZN(n6461) );
  AOI22_X2 U7766 ( .A1(\REGFILE/reg_out[23][21] ), .A2(net77828), .B1(
        \REGFILE/reg_out[22][21] ), .B2(net77836), .ZN(n6460) );
  NAND4_X2 U7767 ( .A1(n6461), .A2(n6460), .A3(n6459), .A4(n6458), .ZN(n6467)
         );
  AOI22_X2 U7768 ( .A1(\REGFILE/reg_out[14][21] ), .A2(net77780), .B1(
        \REGFILE/reg_out[13][21] ), .B2(n5663), .ZN(n6465) );
  AOI22_X2 U7769 ( .A1(\REGFILE/reg_out[9][21] ), .A2(net77700), .B1(
        \REGFILE/reg_out[8][21] ), .B2(n4829), .ZN(n6470) );
  AOI22_X2 U7770 ( .A1(\REGFILE/reg_out[4][21] ), .A2(n5679), .B1(
        \REGFILE/reg_out[5][21] ), .B2(net84475), .ZN(n6469) );
  AOI22_X2 U7771 ( .A1(\REGFILE/reg_out[31][21] ), .A2(net77668), .B1(
        \REGFILE/reg_out[3][21] ), .B2(n5609), .ZN(n6468) );
  NAND4_X2 U7772 ( .A1(n6471), .A2(n6470), .A3(n6469), .A4(n6468), .ZN(n6477)
         );
  NAND4_X2 U7773 ( .A1(n6474), .A2(n6473), .A3(n6475), .A4(n6472), .ZN(n6476)
         );
  NAND2_X2 U7774 ( .A1(\PCLOGIC/imm16_32 [21]), .A2(net75844), .ZN(n6480) );
  OAI21_X4 U7775 ( .B1(n6481), .B2(net78056), .A(n6480), .ZN(n10920) );
  AOI22_X2 U7776 ( .A1(\REGFILE/reg_out[21][20] ), .A2(net77844), .B1(
        \REGFILE/reg_out[20][20] ), .B2(net77852), .ZN(n6485) );
  AOI22_X2 U7777 ( .A1(\REGFILE/reg_out[23][20] ), .A2(net77828), .B1(
        \REGFILE/reg_out[22][20] ), .B2(net77836), .ZN(n6484) );
  AOI22_X2 U7778 ( .A1(\REGFILE/reg_out[19][20] ), .A2(net77812), .B1(
        \REGFILE/reg_out[1][20] ), .B2(net75478), .ZN(n6483) );
  NAND4_X2 U7779 ( .A1(n6485), .A2(n6484), .A3(n6483), .A4(n6482), .ZN(n6491)
         );
  AOI22_X2 U7780 ( .A1(\REGFILE/reg_out[14][20] ), .A2(net77780), .B1(
        \REGFILE/reg_out[13][20] ), .B2(n5664), .ZN(n6489) );
  AOI22_X2 U7781 ( .A1(\REGFILE/reg_out[7][20] ), .A2(net77716), .B1(
        \REGFILE/reg_out[6][20] ), .B2(net75456), .ZN(n6495) );
  AOI22_X2 U7782 ( .A1(\REGFILE/reg_out[31][20] ), .A2(net77668), .B1(
        \REGFILE/reg_out[3][20] ), .B2(net77676), .ZN(n6492) );
  AOI22_X2 U7783 ( .A1(\REGFILE/reg_out[29][20] ), .A2(net77652), .B1(
        \REGFILE/reg_out[28][20] ), .B2(n5751), .ZN(n6499) );
  NAND2_X2 U7784 ( .A1(net75844), .A2(\PCLOGIC/imm16_32 [20]), .ZN(n6504) );
  OAI21_X4 U7785 ( .B1(n6505), .B2(net73697), .A(n6504), .ZN(n10919) );
  AOI22_X2 U7786 ( .A1(\REGFILE/reg_out[21][19] ), .A2(net77844), .B1(
        \REGFILE/reg_out[20][19] ), .B2(net77852), .ZN(n6509) );
  AOI22_X2 U7787 ( .A1(\REGFILE/reg_out[23][19] ), .A2(net77828), .B1(
        \REGFILE/reg_out[22][19] ), .B2(net77836), .ZN(n6508) );
  NAND4_X2 U7788 ( .A1(n6509), .A2(n6508), .A3(n6506), .A4(n6507), .ZN(n6515)
         );
  AOI22_X2 U7789 ( .A1(\REGFILE/reg_out[14][19] ), .A2(net77780), .B1(
        \REGFILE/reg_out[13][19] ), .B2(n5663), .ZN(n6513) );
  NAND4_X2 U7790 ( .A1(n6513), .A2(n6512), .A3(n6511), .A4(n6510), .ZN(n6514)
         );
  AOI22_X2 U7791 ( .A1(\REGFILE/reg_out[9][19] ), .A2(net77700), .B1(
        \REGFILE/reg_out[8][19] ), .B2(net75454), .ZN(n6518) );
  AOI22_X2 U7792 ( .A1(\REGFILE/reg_out[4][19] ), .A2(n5679), .B1(
        \REGFILE/reg_out[5][19] ), .B2(net84475), .ZN(n6517) );
  AOI22_X2 U7793 ( .A1(\REGFILE/reg_out[31][19] ), .A2(net77668), .B1(
        \REGFILE/reg_out[3][19] ), .B2(net77676), .ZN(n6516) );
  NAND4_X2 U7794 ( .A1(n6519), .A2(n6518), .A3(n6517), .A4(n6516), .ZN(n6525)
         );
  NAND2_X2 U7795 ( .A1(net75844), .A2(\PCLOGIC/imm16_32 [19]), .ZN(n6528) );
  OAI21_X4 U7796 ( .B1(n6529), .B2(net78055), .A(n6528), .ZN(n10918) );
  AOI22_X2 U7797 ( .A1(\REGFILE/reg_out[21][18] ), .A2(net77844), .B1(
        \REGFILE/reg_out[20][18] ), .B2(net77852), .ZN(n6533) );
  AOI22_X2 U7798 ( .A1(\REGFILE/reg_out[19][18] ), .A2(net77812), .B1(
        \REGFILE/reg_out[1][18] ), .B2(net75478), .ZN(n6531) );
  NAND4_X2 U7799 ( .A1(n6533), .A2(n6532), .A3(n6531), .A4(n6530), .ZN(n6539)
         );
  NAND4_X2 U7800 ( .A1(n6537), .A2(n6535), .A3(n6536), .A4(n6534), .ZN(n6538)
         );
  AOI22_X2 U7801 ( .A1(\REGFILE/reg_out[7][18] ), .A2(net77714), .B1(
        \REGFILE/reg_out[6][18] ), .B2(net75456), .ZN(n6543) );
  NAND2_X2 U7802 ( .A1(net75844), .A2(\PCLOGIC/imm16_32 [18]), .ZN(n6552) );
  AOI22_X2 U7803 ( .A1(\REGFILE/reg_out[21][17] ), .A2(net77844), .B1(
        \REGFILE/reg_out[20][17] ), .B2(net77852), .ZN(n6557) );
  NAND2_X2 U7804 ( .A1(net75844), .A2(\PCLOGIC/imm16_32 [17]), .ZN(net75843)
         );
  AOI22_X2 U7805 ( .A1(\REGFILE/reg_out[21][16] ), .A2(net77844), .B1(
        \REGFILE/reg_out[20][16] ), .B2(net77852), .ZN(n6565) );
  AOI22_X2 U7806 ( .A1(\REGFILE/reg_out[23][16] ), .A2(net77828), .B1(
        \REGFILE/reg_out[22][16] ), .B2(net77836), .ZN(n6564) );
  NAND4_X2 U7807 ( .A1(n6565), .A2(n6564), .A3(n6563), .A4(n6562), .ZN(n6571)
         );
  NAND4_X2 U7808 ( .A1(n6568), .A2(n6567), .A3(n6569), .A4(n6566), .ZN(n6570)
         );
  AOI22_X2 U7809 ( .A1(\REGFILE/reg_out[30][16] ), .A2(net77638), .B1(
        \REGFILE/reg_out[2][16] ), .B2(net82613), .ZN(n6578) );
  NAND4_X2 U7810 ( .A1(n6578), .A2(n6579), .A3(n6577), .A4(n6576), .ZN(n6580)
         );
  AOI22_X2 U7811 ( .A1(\REGFILE/reg_out[21][15] ), .A2(net77844), .B1(
        \REGFILE/reg_out[20][15] ), .B2(net77852), .ZN(n6587) );
  NAND4_X2 U7812 ( .A1(n6587), .A2(n6585), .A3(n6586), .A4(n6584), .ZN(n6593)
         );
  NOR2_X4 U7813 ( .A1(n6593), .A2(n6592), .ZN(n6605) );
  NAND4_X2 U7814 ( .A1(n6597), .A2(n6596), .A3(n6595), .A4(n6594), .ZN(n6603)
         );
  NAND4_X2 U7815 ( .A1(n6601), .A2(n6600), .A3(n6598), .A4(n6599), .ZN(n6602)
         );
  NOR2_X4 U7816 ( .A1(n6603), .A2(n6602), .ZN(n6604) );
  INV_X4 U7817 ( .A(instruction[0]), .ZN(net73499) );
  NAND2_X2 U7818 ( .A1(instruction[2]), .A2(net73499), .ZN(n6606) );
  INV_X4 U7819 ( .A(n6606), .ZN(n8539) );
  NOR2_X4 U7820 ( .A1(instruction[3]), .A2(instruction[0]), .ZN(n6607) );
  OAI21_X4 U7821 ( .B1(dmem_write_out[15]), .B2(net75427), .A(net78042), .ZN(
        n10288) );
  NAND4_X2 U7822 ( .A1(n6609), .A2(n6610), .A3(n6611), .A4(n6608), .ZN(n6617)
         );
  NAND4_X2 U7823 ( .A1(n6612), .A2(n6615), .A3(n6613), .A4(n6614), .ZN(n6616)
         );
  NOR2_X4 U7824 ( .A1(n6617), .A2(n6616), .ZN(n6629) );
  NAND4_X2 U7825 ( .A1(n6621), .A2(n6620), .A3(n6618), .A4(n6619), .ZN(n6627)
         );
  NOR2_X4 U7826 ( .A1(n6627), .A2(n6626), .ZN(n6628) );
  OAI21_X4 U7827 ( .B1(dmem_write_out[14]), .B2(net75427), .A(net78042), .ZN(
        n10364) );
  NOR2_X4 U7828 ( .A1(n6643), .A2(n6642), .ZN(net75748) );
  AOI22_X2 U7829 ( .A1(\REGFILE/reg_out[21][12] ), .A2(net77844), .B1(
        \REGFILE/reg_out[20][12] ), .B2(net77852), .ZN(n6647) );
  AOI22_X2 U7830 ( .A1(\REGFILE/reg_out[23][12] ), .A2(net77828), .B1(
        \REGFILE/reg_out[22][12] ), .B2(net77836), .ZN(n6646) );
  NAND4_X2 U7831 ( .A1(n6647), .A2(n6646), .A3(n6645), .A4(n6644), .ZN(n6653)
         );
  AOI22_X2 U7832 ( .A1(\REGFILE/reg_out[14][12] ), .A2(net77780), .B1(
        \REGFILE/reg_out[13][12] ), .B2(n5664), .ZN(n6651) );
  AOI22_X2 U7833 ( .A1(\REGFILE/reg_out[0][12] ), .A2(net82342), .B1(n5674), 
        .B2(net83203), .ZN(n6648) );
  NAND4_X2 U7834 ( .A1(n6651), .A2(n6650), .A3(n6649), .A4(n6648), .ZN(n6652)
         );
  NOR2_X4 U7835 ( .A1(n6653), .A2(n6652), .ZN(n6665) );
  AOI22_X2 U7836 ( .A1(\REGFILE/reg_out[7][12] ), .A2(net77714), .B1(
        \REGFILE/reg_out[6][12] ), .B2(net75456), .ZN(n6657) );
  AOI22_X2 U7837 ( .A1(\REGFILE/reg_out[9][12] ), .A2(net77700), .B1(
        \REGFILE/reg_out[8][12] ), .B2(net75454), .ZN(n6656) );
  NAND4_X2 U7838 ( .A1(n6657), .A2(n6656), .A3(n6655), .A4(n6654), .ZN(n6663)
         );
  AOI22_X2 U7839 ( .A1(\REGFILE/reg_out[29][12] ), .A2(net77652), .B1(
        \REGFILE/reg_out[28][12] ), .B2(n6911), .ZN(n6661) );
  NOR2_X4 U7840 ( .A1(n6663), .A2(n6662), .ZN(n6664) );
  OAI21_X4 U7841 ( .B1(dmem_write_out[12]), .B2(net75427), .A(net78042), .ZN(
        n10371) );
  AOI22_X2 U7842 ( .A1(\REGFILE/reg_out[21][11] ), .A2(net77844), .B1(
        \REGFILE/reg_out[20][11] ), .B2(net77852), .ZN(n6669) );
  NAND4_X2 U7843 ( .A1(n6669), .A2(n6666), .A3(n6667), .A4(n6668), .ZN(n6675)
         );
  NOR2_X4 U7844 ( .A1(n6675), .A2(n6674), .ZN(n6687) );
  AOI22_X2 U7845 ( .A1(\REGFILE/reg_out[7][11] ), .A2(net77716), .B1(
        \REGFILE/reg_out[6][11] ), .B2(net75456), .ZN(n6679) );
  AOI22_X2 U7846 ( .A1(\REGFILE/reg_out[9][11] ), .A2(net77700), .B1(
        \REGFILE/reg_out[8][11] ), .B2(net75454), .ZN(n6678) );
  NAND4_X2 U7847 ( .A1(n6679), .A2(n6678), .A3(n6677), .A4(n6676), .ZN(n6685)
         );
  NAND4_X2 U7848 ( .A1(n6683), .A2(n6682), .A3(n6681), .A4(n6680), .ZN(n6684)
         );
  NOR2_X4 U7849 ( .A1(n6685), .A2(n6684), .ZN(n6686) );
  OAI21_X4 U7850 ( .B1(dmem_write_out[11]), .B2(net75427), .A(net78042), .ZN(
        n9835) );
  AOI22_X2 U7851 ( .A1(\REGFILE/reg_out[21][10] ), .A2(net77842), .B1(
        \REGFILE/reg_out[20][10] ), .B2(net77850), .ZN(n6691) );
  NAND4_X2 U7852 ( .A1(n6691), .A2(n6690), .A3(n6689), .A4(n6688), .ZN(n6697)
         );
  NAND4_X2 U7853 ( .A1(n6695), .A2(n6694), .A3(n6693), .A4(n6692), .ZN(n6696)
         );
  NOR2_X4 U7854 ( .A1(n6697), .A2(n6696), .ZN(n6709) );
  NAND4_X2 U7855 ( .A1(n6701), .A2(n6700), .A3(n6699), .A4(n6698), .ZN(n6707)
         );
  NAND4_X2 U7856 ( .A1(n6705), .A2(n6702), .A3(n6704), .A4(n6703), .ZN(n6706)
         );
  NOR2_X4 U7857 ( .A1(n6706), .A2(n6707), .ZN(n6708) );
  OAI21_X4 U7858 ( .B1(dmem_write_out[10]), .B2(net75427), .A(net78042), .ZN(
        n10378) );
  AOI22_X2 U7859 ( .A1(\REGFILE/reg_out[21][9] ), .A2(net77842), .B1(
        \REGFILE/reg_out[20][9] ), .B2(net77850), .ZN(n6713) );
  AOI22_X2 U7860 ( .A1(\REGFILE/reg_out[23][9] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][9] ), .B2(net77834), .ZN(n6712) );
  NAND4_X2 U7861 ( .A1(n6713), .A2(n6712), .A3(n6711), .A4(n6710), .ZN(n6719)
         );
  AOI22_X2 U7862 ( .A1(\REGFILE/reg_out[14][9] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][9] ), .B2(n5664), .ZN(n6717) );
  NAND4_X2 U7863 ( .A1(n6717), .A2(n6716), .A3(n6715), .A4(n6714), .ZN(n6718)
         );
  AOI22_X2 U7864 ( .A1(\REGFILE/reg_out[7][9] ), .A2(net75455), .B1(
        \REGFILE/reg_out[6][9] ), .B2(net75456), .ZN(n6723) );
  AOI22_X2 U7865 ( .A1(\REGFILE/reg_out[9][9] ), .A2(net77698), .B1(
        \REGFILE/reg_out[8][9] ), .B2(n4829), .ZN(n6722) );
  NAND4_X2 U7866 ( .A1(n6723), .A2(n6722), .A3(n6721), .A4(n6720), .ZN(n6729)
         );
  AOI22_X2 U7867 ( .A1(\REGFILE/reg_out[26][9] ), .A2(net75439), .B1(
        \REGFILE/reg_out[27][9] ), .B2(net89184), .ZN(n6725) );
  NAND4_X2 U7868 ( .A1(n6727), .A2(n6725), .A3(n6726), .A4(n6724), .ZN(n6728)
         );
  OAI21_X4 U7869 ( .B1(dmem_write_out[9]), .B2(net75427), .A(n10945), .ZN(
        n9358) );
  AOI22_X2 U7870 ( .A1(\REGFILE/reg_out[23][8] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][8] ), .B2(net77834), .ZN(n6734) );
  NAND4_X2 U7871 ( .A1(n6733), .A2(n6734), .A3(n6735), .A4(n6732), .ZN(n6741)
         );
  NAND4_X2 U7872 ( .A1(n6739), .A2(n6738), .A3(n6737), .A4(n6736), .ZN(n6740)
         );
  NOR2_X4 U7873 ( .A1(n6741), .A2(n6740), .ZN(n6753) );
  NAND4_X2 U7874 ( .A1(n6745), .A2(n6744), .A3(n6743), .A4(n6742), .ZN(n6751)
         );
  NAND4_X2 U7875 ( .A1(n6749), .A2(n6748), .A3(n6746), .A4(n6747), .ZN(n6750)
         );
  OAI21_X4 U7876 ( .B1(dmem_write_out[8]), .B2(net75427), .A(net78042), .ZN(
        n10385) );
  AOI22_X2 U7877 ( .A1(\REGFILE/reg_out[21][7] ), .A2(net77842), .B1(
        \REGFILE/reg_out[20][7] ), .B2(net77850), .ZN(n6757) );
  AOI22_X2 U7878 ( .A1(\REGFILE/reg_out[23][7] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][7] ), .B2(net77834), .ZN(n6756) );
  AOI22_X2 U7879 ( .A1(\REGFILE/reg_out[19][7] ), .A2(net77810), .B1(
        \REGFILE/reg_out[1][7] ), .B2(net75478), .ZN(n6755) );
  NAND4_X2 U7880 ( .A1(n6757), .A2(n6756), .A3(n6755), .A4(n6754), .ZN(n6763)
         );
  AOI22_X2 U7881 ( .A1(\REGFILE/reg_out[14][7] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][7] ), .B2(n5664), .ZN(n6761) );
  NAND4_X2 U7882 ( .A1(n6759), .A2(n6760), .A3(n6761), .A4(n6758), .ZN(n6762)
         );
  AOI22_X2 U7883 ( .A1(\REGFILE/reg_out[29][7] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][7] ), .B2(n5751), .ZN(net75619) );
  AOI22_X2 U7884 ( .A1(\REGFILE/reg_out[21][6] ), .A2(net77842), .B1(
        \REGFILE/reg_out[20][6] ), .B2(net77850), .ZN(n6767) );
  AOI22_X2 U7885 ( .A1(\REGFILE/reg_out[19][6] ), .A2(net77810), .B1(
        \REGFILE/reg_out[1][6] ), .B2(net75478), .ZN(n6765) );
  NAND4_X2 U7886 ( .A1(n6767), .A2(n6766), .A3(n6765), .A4(n6764), .ZN(n6773)
         );
  AOI22_X2 U7887 ( .A1(\REGFILE/reg_out[14][6] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][6] ), .B2(n6009), .ZN(n6771) );
  NAND4_X2 U7888 ( .A1(n6770), .A2(n6771), .A3(n6769), .A4(n6768), .ZN(n6772)
         );
  NOR2_X4 U7889 ( .A1(n6772), .A2(n6773), .ZN(n6785) );
  AOI22_X2 U7890 ( .A1(\REGFILE/reg_out[9][6] ), .A2(net77698), .B1(
        \REGFILE/reg_out[8][6] ), .B2(n4829), .ZN(n6776) );
  NAND4_X2 U7891 ( .A1(n6777), .A2(n6776), .A3(n6775), .A4(n6774), .ZN(n6783)
         );
  AOI22_X2 U7892 ( .A1(\REGFILE/reg_out[29][6] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][6] ), .B2(n6911), .ZN(n6781) );
  NAND4_X2 U7893 ( .A1(n6780), .A2(n6781), .A3(n6779), .A4(n6778), .ZN(n6782)
         );
  NOR2_X4 U7894 ( .A1(n6783), .A2(n6782), .ZN(n6784) );
  OAI21_X4 U7895 ( .B1(dmem_write_out[6]), .B2(net75427), .A(n10945), .ZN(
        n10392) );
  AOI22_X2 U7896 ( .A1(\REGFILE/reg_out[21][5] ), .A2(net77842), .B1(
        \REGFILE/reg_out[20][5] ), .B2(net77850), .ZN(n6789) );
  NAND4_X2 U7897 ( .A1(n6789), .A2(n6788), .A3(n6787), .A4(n6786), .ZN(n6795)
         );
  AOI22_X2 U7898 ( .A1(\REGFILE/reg_out[14][5] ), .A2(net77778), .B1(
        \REGFILE/reg_out[13][5] ), .B2(n6009), .ZN(n6793) );
  NAND4_X2 U7899 ( .A1(n6790), .A2(n6792), .A3(n6791), .A4(n6793), .ZN(n6794)
         );
  AOI22_X2 U7900 ( .A1(\REGFILE/reg_out[9][5] ), .A2(net77698), .B1(
        \REGFILE/reg_out[8][5] ), .B2(n4829), .ZN(n6798) );
  NAND4_X2 U7901 ( .A1(n6799), .A2(n6798), .A3(n6797), .A4(n6796), .ZN(n6805)
         );
  AOI22_X2 U7902 ( .A1(\REGFILE/reg_out[29][5] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][5] ), .B2(n6911), .ZN(n6803) );
  NAND4_X2 U7903 ( .A1(n6803), .A2(n6802), .A3(n6801), .A4(n6800), .ZN(n6804)
         );
  OAI21_X4 U7904 ( .B1(dmem_write_out[5]), .B2(net75427), .A(n10945), .ZN(
        n9616) );
  AOI22_X2 U7905 ( .A1(\REGFILE/reg_out[21][4] ), .A2(net77842), .B1(
        \REGFILE/reg_out[20][4] ), .B2(net77850), .ZN(n6811) );
  NAND4_X2 U7906 ( .A1(n6811), .A2(n6810), .A3(n6809), .A4(n6808), .ZN(n6817)
         );
  NAND4_X2 U7907 ( .A1(n6815), .A2(n6812), .A3(n6813), .A4(n6814), .ZN(n6816)
         );
  AOI22_X2 U7908 ( .A1(\REGFILE/reg_out[9][4] ), .A2(net77698), .B1(
        \REGFILE/reg_out[8][4] ), .B2(n4829), .ZN(n6820) );
  NAND4_X2 U7909 ( .A1(n6821), .A2(n6820), .A3(n6819), .A4(n6818), .ZN(n6827)
         );
  AOI22_X2 U7910 ( .A1(\REGFILE/reg_out[29][4] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][4] ), .B2(n6911), .ZN(n6825) );
  NAND4_X2 U7911 ( .A1(n6824), .A2(n6825), .A3(n6823), .A4(n6822), .ZN(n6826)
         );
  AOI22_X2 U7912 ( .A1(\REGFILE/reg_out[21][3] ), .A2(net77842), .B1(
        \REGFILE/reg_out[20][3] ), .B2(net77850), .ZN(n6833) );
  NAND4_X2 U7913 ( .A1(n6833), .A2(n6832), .A3(n6830), .A4(n6831), .ZN(n6839)
         );
  NAND4_X2 U7914 ( .A1(n6836), .A2(n6834), .A3(n6835), .A4(n6837), .ZN(n6838)
         );
  NAND4_X2 U7915 ( .A1(n6840), .A2(n6842), .A3(n6841), .A4(n6843), .ZN(n6849)
         );
  NAND4_X2 U7916 ( .A1(n6847), .A2(n6846), .A3(n6845), .A4(n6844), .ZN(n6848)
         );
  OAI21_X4 U7917 ( .B1(dmem_write_out[3]), .B2(net75427), .A(n10945), .ZN(
        n10036) );
  AOI22_X2 U7918 ( .A1(\REGFILE/reg_out[23][2] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][2] ), .B2(net77834), .ZN(n6854) );
  NAND4_X2 U7919 ( .A1(n6853), .A2(n6854), .A3(n6855), .A4(n6852), .ZN(n6861)
         );
  NAND4_X2 U7920 ( .A1(n6859), .A2(n6858), .A3(n6857), .A4(n6856), .ZN(n6860)
         );
  NOR2_X4 U7921 ( .A1(n6861), .A2(n6860), .ZN(n6873) );
  NAND4_X2 U7922 ( .A1(n6862), .A2(n6864), .A3(n6863), .A4(n6865), .ZN(n6871)
         );
  AOI22_X2 U7923 ( .A1(\REGFILE/reg_out[29][2] ), .A2(net77650), .B1(
        \REGFILE/reg_out[28][2] ), .B2(n6911), .ZN(n6869) );
  NOR2_X4 U7924 ( .A1(n6871), .A2(n6870), .ZN(n6872) );
  OAI21_X4 U7925 ( .B1(dmem_write_out[2]), .B2(net75427), .A(n10945), .ZN(
        n10408) );
  AOI22_X2 U7926 ( .A1(\REGFILE/reg_out[21][1] ), .A2(net77842), .B1(
        \REGFILE/reg_out[20][1] ), .B2(net77850), .ZN(n6877) );
  AOI22_X2 U7927 ( .A1(\REGFILE/reg_out[23][1] ), .A2(net77826), .B1(
        \REGFILE/reg_out[22][1] ), .B2(net77834), .ZN(n6876) );
  NAND4_X2 U7928 ( .A1(n6877), .A2(n6876), .A3(n6875), .A4(n6874), .ZN(n6883)
         );
  NAND4_X2 U7929 ( .A1(n6884), .A2(n6886), .A3(n6885), .A4(n6887), .ZN(n6893)
         );
  AOI22_X2 U7930 ( .A1(\REGFILE/reg_out[21][0] ), .A2(net77842), .B1(
        \REGFILE/reg_out[20][0] ), .B2(net77850), .ZN(n6900) );
  NAND4_X2 U7931 ( .A1(n6900), .A2(n6899), .A3(n6898), .A4(n6897), .ZN(n6906)
         );
  NAND4_X2 U7932 ( .A1(n6901), .A2(n6903), .A3(n6902), .A4(n6904), .ZN(n6905)
         );
  NOR2_X4 U7933 ( .A1(n6906), .A2(n6905), .ZN(n6919) );
  NAND4_X2 U7934 ( .A1(n6910), .A2(n6909), .A3(n6908), .A4(n6907), .ZN(n6917)
         );
  NAND4_X2 U7935 ( .A1(n6915), .A2(n6914), .A3(n6913), .A4(n6912), .ZN(n6916)
         );
  NOR2_X4 U7936 ( .A1(n6917), .A2(n6916), .ZN(n6918) );
  NAND2_X2 U7937 ( .A1(n6919), .A2(n6918), .ZN(dmem_write_out[0]) );
  INV_X4 U7938 ( .A(\PCLOGIC/imm26_32 [7]), .ZN(n8295) );
  INV_X4 U7939 ( .A(\PCLOGIC/imm26_32 [6]), .ZN(n8287) );
  NAND2_X2 U7940 ( .A1(n8295), .A2(n8287), .ZN(net73842) );
  NAND3_X4 U7941 ( .A1(\PCLOGIC/imm26_32 [10]), .A2(\PCLOGIC/imm26_32 [8]), 
        .A3(\PCLOGIC/imm26_32 [9]), .ZN(net75425) );
  NAND3_X4 U7942 ( .A1(\PCLOGIC/imm26_32 [8]), .A2(net73987), .A3(
        \PCLOGIC/imm26_32 [9]), .ZN(net75424) );
  NAND3_X4 U7943 ( .A1(net90864), .A2(net73987), .A3(\PCLOGIC/imm26_32 [9]), 
        .ZN(n6920) );
  NAND3_X4 U7944 ( .A1(net123932), .A2(net87098), .A3(\PCLOGIC/imm26_32 [10]), 
        .ZN(net75419) );
  NAND3_X4 U7945 ( .A1(net73987), .A2(net87098), .A3(net73879), .ZN(net75418)
         );
  NAND2_X2 U7946 ( .A1(\PCLOGIC/imm26_32 [6]), .A2(n8295), .ZN(net73836) );
  NAND2_X2 U7947 ( .A1(\PCLOGIC/imm26_32 [7]), .A2(n8287), .ZN(n8407) );
  INV_X4 U7948 ( .A(n8407), .ZN(n8402) );
  NAND2_X2 U7949 ( .A1(n8402), .A2(net77272), .ZN(n6951) );
  INV_X4 U7950 ( .A(n6951), .ZN(n6933) );
  NAND2_X2 U7951 ( .A1(\PCLOGIC/imm26_32 [7]), .A2(\PCLOGIC/imm26_32 [6]), 
        .ZN(n8409) );
  NOR2_X4 U7952 ( .A1(n6954), .A2(n6953), .ZN(n6955) );
  NAND2_X2 U7953 ( .A1(\REGFILE/reg_out[2][29] ), .A2(net77336), .ZN(n6959) );
  NAND2_X2 U7954 ( .A1(\REGFILE/reg_out[3][29] ), .A2(net77406), .ZN(n6958) );
  NAND2_X2 U7955 ( .A1(\REGFILE/reg_out[0][29] ), .A2(net77300), .ZN(n6957) );
  NAND2_X2 U7956 ( .A1(\REGFILE/reg_out[7][29] ), .A2(net77480), .ZN(n6962) );
  NAND2_X2 U7957 ( .A1(\REGFILE/reg_out[12][29] ), .A2(net77388), .ZN(n6969)
         );
  NAND2_X2 U7958 ( .A1(\REGFILE/reg_out[13][29] ), .A2(net77462), .ZN(n6968)
         );
  NAND2_X2 U7959 ( .A1(\REGFILE/reg_out[10][29] ), .A2(n6017), .ZN(n6967) );
  NAND2_X2 U7960 ( .A1(\REGFILE/reg_out[11][29] ), .A2(net77426), .ZN(n6966)
         );
  NAND2_X2 U7961 ( .A1(\REGFILE/reg_out[18][29] ), .A2(n6017), .ZN(n6979) );
  NAND2_X2 U7962 ( .A1(\REGFILE/reg_out[19][29] ), .A2(net77426), .ZN(n6978)
         );
  NAND2_X2 U7963 ( .A1(\REGFILE/reg_out[16][29] ), .A2(net77318), .ZN(n6977)
         );
  NAND4_X2 U7964 ( .A1(n6979), .A2(n6978), .A3(n6977), .A4(n6976), .ZN(n6983)
         );
  NAND2_X2 U7965 ( .A1(\REGFILE/reg_out[26][29] ), .A2(n6017), .ZN(n6987) );
  NAND2_X2 U7966 ( .A1(\REGFILE/reg_out[30][29] ), .A2(net77550), .ZN(n6991)
         );
  NAND2_X2 U7967 ( .A1(n5986), .A2(net77400), .ZN(n6989) );
  NAND2_X2 U7968 ( .A1(net77478), .A2(\REGFILE/reg_out[31][28] ), .ZN(n6999)
         );
  NAND2_X2 U7969 ( .A1(net77456), .A2(\REGFILE/reg_out[29][28] ), .ZN(n6998)
         );
  NAND4_X2 U7970 ( .A1(n7001), .A2(n7000), .A3(n6999), .A4(n6998), .ZN(n7007)
         );
  NAND2_X2 U7971 ( .A1(net77388), .A2(\REGFILE/reg_out[28][28] ), .ZN(n7004)
         );
  NAND2_X2 U7972 ( .A1(n6014), .A2(\REGFILE/reg_out[26][28] ), .ZN(n7003) );
  NAND4_X2 U7973 ( .A1(n7005), .A2(n7004), .A3(n7003), .A4(n7002), .ZN(n7006)
         );
  NAND2_X2 U7974 ( .A1(net77478), .A2(\REGFILE/reg_out[23][28] ), .ZN(n7009)
         );
  NAND2_X2 U7975 ( .A1(net77388), .A2(\REGFILE/reg_out[20][28] ), .ZN(n7014)
         );
  NAND2_X2 U7976 ( .A1(n6014), .A2(\REGFILE/reg_out[18][28] ), .ZN(n7013) );
  NAND4_X2 U7977 ( .A1(n7015), .A2(n7014), .A3(n7013), .A4(n7012), .ZN(n7016)
         );
  OAI21_X4 U7978 ( .B1(n7017), .B2(n7016), .A(net77588), .ZN(n7040) );
  NAND2_X2 U7979 ( .A1(net77516), .A2(\REGFILE/reg_out[9][28] ), .ZN(n7020) );
  NAND2_X2 U7980 ( .A1(net77480), .A2(\REGFILE/reg_out[15][28] ), .ZN(n7019)
         );
  NAND4_X2 U7981 ( .A1(n7021), .A2(n7020), .A3(n7019), .A4(n7018), .ZN(n7027)
         );
  NAND2_X2 U7982 ( .A1(net77422), .A2(\REGFILE/reg_out[11][28] ), .ZN(n7025)
         );
  NAND2_X2 U7983 ( .A1(net77336), .A2(\REGFILE/reg_out[10][28] ), .ZN(n7023)
         );
  NAND2_X2 U7984 ( .A1(net77300), .A2(\REGFILE/reg_out[8][28] ), .ZN(n7022) );
  NAND4_X2 U7985 ( .A1(n7025), .A2(n7024), .A3(n7023), .A4(n7022), .ZN(n7026)
         );
  NAND2_X2 U7986 ( .A1(net77514), .A2(\REGFILE/reg_out[1][28] ), .ZN(n7030) );
  NAND4_X2 U7987 ( .A1(n7031), .A2(n7030), .A3(n7029), .A4(n7028), .ZN(n7037)
         );
  NAND2_X2 U7988 ( .A1(net77388), .A2(\REGFILE/reg_out[4][28] ), .ZN(n7034) );
  NAND2_X2 U7989 ( .A1(n6014), .A2(\REGFILE/reg_out[2][28] ), .ZN(n7033) );
  NAND4_X2 U7990 ( .A1(n7035), .A2(n7034), .A3(n7033), .A4(n7032), .ZN(n7036)
         );
  NAND2_X2 U7991 ( .A1(net77516), .A2(\REGFILE/reg_out[25][27] ), .ZN(n7044)
         );
  NAND2_X2 U7992 ( .A1(net77480), .A2(\REGFILE/reg_out[31][27] ), .ZN(n7043)
         );
  NAND4_X2 U7993 ( .A1(n7045), .A2(n7044), .A3(n7043), .A4(n7042), .ZN(n7051)
         );
  NAND2_X2 U7994 ( .A1(net77414), .A2(\REGFILE/reg_out[27][27] ), .ZN(n7049)
         );
  NAND2_X2 U7995 ( .A1(net77336), .A2(\REGFILE/reg_out[26][27] ), .ZN(n7047)
         );
  NAND2_X2 U7996 ( .A1(net77300), .A2(\REGFILE/reg_out[24][27] ), .ZN(n7046)
         );
  NAND4_X2 U7997 ( .A1(n7049), .A2(n7048), .A3(n7047), .A4(n7046), .ZN(n7050)
         );
  OAI21_X4 U7998 ( .B1(n7051), .B2(n7050), .A(n6012), .ZN(n7085) );
  NAND2_X2 U7999 ( .A1(net77478), .A2(\REGFILE/reg_out[23][27] ), .ZN(n7053)
         );
  NAND2_X2 U8000 ( .A1(net77456), .A2(\REGFILE/reg_out[21][27] ), .ZN(n7052)
         );
  NAND4_X2 U8001 ( .A1(n7055), .A2(n7054), .A3(n7053), .A4(n7052), .ZN(n7061)
         );
  NAND2_X2 U8003 ( .A1(n6014), .A2(\REGFILE/reg_out[18][27] ), .ZN(n7057) );
  NAND4_X2 U8004 ( .A1(n7059), .A2(n7058), .A3(n7057), .A4(n7056), .ZN(n7060)
         );
  OAI21_X4 U8005 ( .B1(n7061), .B2(n7060), .A(net77588), .ZN(n7084) );
  NAND2_X2 U8006 ( .A1(net77516), .A2(\REGFILE/reg_out[9][27] ), .ZN(n7064) );
  NAND2_X2 U8007 ( .A1(net77480), .A2(\REGFILE/reg_out[15][27] ), .ZN(n7063)
         );
  NAND4_X2 U8008 ( .A1(n7065), .A2(n7064), .A3(n7063), .A4(n7062), .ZN(n7071)
         );
  NAND2_X2 U8009 ( .A1(net77420), .A2(\REGFILE/reg_out[11][27] ), .ZN(n7069)
         );
  NAND2_X2 U8010 ( .A1(net77336), .A2(\REGFILE/reg_out[10][27] ), .ZN(n7067)
         );
  NAND2_X2 U8011 ( .A1(net77300), .A2(\REGFILE/reg_out[8][27] ), .ZN(n7066) );
  NAND4_X2 U8012 ( .A1(n7069), .A2(n7068), .A3(n7067), .A4(n7066), .ZN(n7070)
         );
  OAI21_X4 U8013 ( .B1(n7071), .B2(n7070), .A(n6019), .ZN(n7083) );
  NAND2_X2 U8014 ( .A1(net77516), .A2(\REGFILE/reg_out[1][27] ), .ZN(n7074) );
  NAND2_X2 U8015 ( .A1(net77480), .A2(\REGFILE/reg_out[7][27] ), .ZN(n7073) );
  NAND4_X2 U8016 ( .A1(n7075), .A2(n7074), .A3(n7073), .A4(n7072), .ZN(n7081)
         );
  NAND2_X2 U8017 ( .A1(net77418), .A2(\REGFILE/reg_out[3][27] ), .ZN(n7079) );
  NAND2_X2 U8018 ( .A1(net77336), .A2(\REGFILE/reg_out[2][27] ), .ZN(n7077) );
  NAND4_X2 U8020 ( .A1(n7079), .A2(n7078), .A3(n7077), .A4(n7076), .ZN(n7080)
         );
  OAI21_X4 U8021 ( .B1(n7081), .B2(n7080), .A(net77292), .ZN(n7082) );
  MUX2_X2 U8022 ( .A(n8450), .B(\PCLOGIC/imm16_32 [27]), .S(net77276), .Z(
        aluA[27]) );
  NAND2_X2 U8023 ( .A1(\REGFILE/reg_out[30][26] ), .A2(net77564), .ZN(n7089)
         );
  NAND2_X2 U8024 ( .A1(\REGFILE/reg_out[31][26] ), .A2(net77498), .ZN(n7087)
         );
  NAND2_X2 U8025 ( .A1(\REGFILE/reg_out[29][26] ), .A2(net77462), .ZN(n7086)
         );
  NAND4_X2 U8026 ( .A1(n7089), .A2(n7088), .A3(n7087), .A4(n7086), .ZN(n7095)
         );
  NAND2_X2 U8027 ( .A1(\REGFILE/reg_out[27][26] ), .A2(net77426), .ZN(n7093)
         );
  NAND2_X2 U8028 ( .A1(\REGFILE/reg_out[28][26] ), .A2(net77376), .ZN(n7092)
         );
  NAND2_X2 U8029 ( .A1(\REGFILE/reg_out[26][26] ), .A2(n6017), .ZN(n7091) );
  NAND2_X2 U8030 ( .A1(\REGFILE/reg_out[24][26] ), .A2(net77318), .ZN(n7090)
         );
  NAND4_X2 U8031 ( .A1(n7093), .A2(n7092), .A3(n7091), .A4(n7090), .ZN(n7094)
         );
  NAND2_X2 U8032 ( .A1(\REGFILE/reg_out[22][26] ), .A2(net77566), .ZN(n7099)
         );
  NAND2_X2 U8033 ( .A1(\REGFILE/reg_out[23][26] ), .A2(net77498), .ZN(n7097)
         );
  NAND2_X2 U8034 ( .A1(\REGFILE/reg_out[21][26] ), .A2(net77462), .ZN(n7096)
         );
  NAND4_X2 U8035 ( .A1(n7099), .A2(n7098), .A3(n7097), .A4(n7096), .ZN(n7105)
         );
  NAND2_X2 U8036 ( .A1(\REGFILE/reg_out[19][26] ), .A2(net77426), .ZN(n7103)
         );
  NAND2_X2 U8037 ( .A1(\REGFILE/reg_out[20][26] ), .A2(net77384), .ZN(n7102)
         );
  NAND2_X2 U8038 ( .A1(\REGFILE/reg_out[18][26] ), .A2(n6017), .ZN(n7101) );
  NAND2_X2 U8039 ( .A1(\REGFILE/reg_out[16][26] ), .A2(net77318), .ZN(n7100)
         );
  NAND4_X2 U8040 ( .A1(n7103), .A2(n7102), .A3(n7101), .A4(n7100), .ZN(n7104)
         );
  NAND2_X2 U8041 ( .A1(\REGFILE/reg_out[14][26] ), .A2(net77568), .ZN(n7109)
         );
  NAND2_X2 U8042 ( .A1(\REGFILE/reg_out[15][26] ), .A2(net77498), .ZN(n7107)
         );
  NAND2_X2 U8043 ( .A1(\REGFILE/reg_out[13][26] ), .A2(net77462), .ZN(n7106)
         );
  NAND4_X2 U8044 ( .A1(n7109), .A2(n7108), .A3(n7107), .A4(n7106), .ZN(n7115)
         );
  NAND2_X2 U8045 ( .A1(\REGFILE/reg_out[11][26] ), .A2(net77426), .ZN(n7113)
         );
  NAND2_X2 U8046 ( .A1(\REGFILE/reg_out[12][26] ), .A2(net77380), .ZN(n7112)
         );
  NAND2_X2 U8047 ( .A1(\REGFILE/reg_out[10][26] ), .A2(n6017), .ZN(n7111) );
  NAND2_X2 U8048 ( .A1(\REGFILE/reg_out[8][26] ), .A2(net77318), .ZN(n7110) );
  NAND4_X2 U8049 ( .A1(n7113), .A2(n7112), .A3(n7111), .A4(n7110), .ZN(n7114)
         );
  NAND2_X2 U8050 ( .A1(\REGFILE/reg_out[6][26] ), .A2(net77560), .ZN(n7119) );
  NAND2_X2 U8051 ( .A1(\REGFILE/reg_out[7][26] ), .A2(net77498), .ZN(n7117) );
  NAND2_X2 U8052 ( .A1(\REGFILE/reg_out[5][26] ), .A2(net77462), .ZN(n7116) );
  NAND4_X2 U8053 ( .A1(n7119), .A2(n7118), .A3(n7117), .A4(n7116), .ZN(n7125)
         );
  NAND2_X2 U8054 ( .A1(\REGFILE/reg_out[3][26] ), .A2(net77426), .ZN(n7123) );
  NAND2_X2 U8055 ( .A1(\REGFILE/reg_out[4][26] ), .A2(net77382), .ZN(n7122) );
  NAND2_X2 U8056 ( .A1(\REGFILE/reg_out[2][26] ), .A2(n6017), .ZN(n7121) );
  NAND2_X2 U8057 ( .A1(\REGFILE/reg_out[0][26] ), .A2(net77318), .ZN(n7120) );
  NAND4_X2 U8058 ( .A1(n7123), .A2(n7122), .A3(n7121), .A4(n7120), .ZN(n7124)
         );
  NAND4_X2 U8059 ( .A1(n7129), .A2(n7128), .A3(n7127), .A4(n7126), .ZN(n8448)
         );
  MUX2_X2 U8060 ( .A(n8448), .B(\PCLOGIC/imm16_32 [26]), .S(net77276), .Z(
        aluA[26]) );
  NAND2_X2 U8061 ( .A1(\REGFILE/reg_out[27][25] ), .A2(net77426), .ZN(n7133)
         );
  NAND2_X2 U8062 ( .A1(\REGFILE/reg_out[28][25] ), .A2(net77376), .ZN(n7132)
         );
  NAND2_X2 U8063 ( .A1(\REGFILE/reg_out[26][25] ), .A2(n6017), .ZN(n7131) );
  NAND2_X2 U8064 ( .A1(\REGFILE/reg_out[24][25] ), .A2(net77318), .ZN(n7130)
         );
  NAND4_X2 U8065 ( .A1(n7133), .A2(n7132), .A3(n7131), .A4(n7130), .ZN(n7139)
         );
  NAND2_X2 U8066 ( .A1(\REGFILE/reg_out[30][25] ), .A2(net77558), .ZN(n7137)
         );
  NAND2_X2 U8067 ( .A1(\REGFILE/reg_out[25][25] ), .A2(net77544), .ZN(n7136)
         );
  NAND2_X2 U8068 ( .A1(\REGFILE/reg_out[31][25] ), .A2(net77498), .ZN(n7135)
         );
  NAND2_X2 U8069 ( .A1(\REGFILE/reg_out[29][25] ), .A2(net77462), .ZN(n7134)
         );
  NAND4_X2 U8070 ( .A1(n7137), .A2(n7136), .A3(n7135), .A4(n7134), .ZN(n7138)
         );
  NAND2_X2 U8071 ( .A1(\REGFILE/reg_out[3][25] ), .A2(net77424), .ZN(n7143) );
  NAND2_X2 U8073 ( .A1(\REGFILE/reg_out[2][25] ), .A2(n6016), .ZN(n7141) );
  NAND2_X2 U8074 ( .A1(\REGFILE/reg_out[0][25] ), .A2(net77316), .ZN(n7140) );
  NAND4_X2 U8075 ( .A1(n7143), .A2(n7142), .A3(n7141), .A4(n7140), .ZN(n7149)
         );
  NAND2_X2 U8076 ( .A1(\REGFILE/reg_out[6][25] ), .A2(net77568), .ZN(n7147) );
  NAND2_X2 U8077 ( .A1(\REGFILE/reg_out[1][25] ), .A2(net77532), .ZN(n7146) );
  NAND2_X2 U8078 ( .A1(\REGFILE/reg_out[7][25] ), .A2(net77496), .ZN(n7145) );
  NAND2_X2 U8079 ( .A1(\REGFILE/reg_out[5][25] ), .A2(net77460), .ZN(n7144) );
  NAND4_X2 U8080 ( .A1(n7147), .A2(n7146), .A3(n7145), .A4(n7144), .ZN(n7148)
         );
  NAND2_X2 U8081 ( .A1(\REGFILE/reg_out[11][25] ), .A2(net77424), .ZN(n7153)
         );
  NAND2_X2 U8083 ( .A1(\REGFILE/reg_out[10][25] ), .A2(n6016), .ZN(n7151) );
  NAND2_X2 U8084 ( .A1(\REGFILE/reg_out[8][25] ), .A2(net77316), .ZN(n7150) );
  NAND4_X2 U8085 ( .A1(n7153), .A2(n7152), .A3(n7151), .A4(n7150), .ZN(n7159)
         );
  NAND2_X2 U8086 ( .A1(\REGFILE/reg_out[14][25] ), .A2(net77568), .ZN(n7157)
         );
  NAND2_X2 U8087 ( .A1(\REGFILE/reg_out[9][25] ), .A2(net77532), .ZN(n7156) );
  NAND2_X2 U8088 ( .A1(\REGFILE/reg_out[15][25] ), .A2(net77496), .ZN(n7155)
         );
  NAND2_X2 U8089 ( .A1(\REGFILE/reg_out[13][25] ), .A2(net77460), .ZN(n7154)
         );
  NAND4_X2 U8090 ( .A1(n7157), .A2(n7156), .A3(n7155), .A4(n7154), .ZN(n7158)
         );
  NAND2_X2 U8091 ( .A1(\REGFILE/reg_out[19][25] ), .A2(net77424), .ZN(n7163)
         );
  NAND2_X2 U8093 ( .A1(\REGFILE/reg_out[18][25] ), .A2(n6016), .ZN(n7161) );
  NAND2_X2 U8094 ( .A1(\REGFILE/reg_out[16][25] ), .A2(net77316), .ZN(n7160)
         );
  NAND4_X2 U8095 ( .A1(n7163), .A2(n7162), .A3(n7161), .A4(n7160), .ZN(n7169)
         );
  NAND2_X2 U8096 ( .A1(\REGFILE/reg_out[22][25] ), .A2(net77568), .ZN(n7167)
         );
  NAND2_X2 U8097 ( .A1(\REGFILE/reg_out[17][25] ), .A2(net77532), .ZN(n7166)
         );
  NAND2_X2 U8098 ( .A1(\REGFILE/reg_out[23][25] ), .A2(net77496), .ZN(n7165)
         );
  NAND2_X2 U8099 ( .A1(\REGFILE/reg_out[21][25] ), .A2(net77460), .ZN(n7164)
         );
  NAND4_X2 U8100 ( .A1(n7167), .A2(n7166), .A3(n7165), .A4(n7164), .ZN(n7168)
         );
  NAND4_X2 U8101 ( .A1(n7173), .A2(n7172), .A3(n7171), .A4(n7170), .ZN(n8419)
         );
  INV_X4 U8102 ( .A(n8419), .ZN(n7174) );
  INV_X4 U8103 ( .A(\PCLOGIC/imm16_32 [25]), .ZN(n8329) );
  MUX2_X2 U8104 ( .A(n7174), .B(n8329), .S(net77276), .Z(n10327) );
  NAND2_X2 U8105 ( .A1(\REGFILE/reg_out[27][24] ), .A2(net77424), .ZN(n7178)
         );
  NAND2_X2 U8107 ( .A1(\REGFILE/reg_out[26][24] ), .A2(n6016), .ZN(n7176) );
  NAND2_X2 U8108 ( .A1(\REGFILE/reg_out[24][24] ), .A2(net77316), .ZN(n7175)
         );
  NAND4_X2 U8109 ( .A1(n7178), .A2(n7177), .A3(n7176), .A4(n7175), .ZN(n7184)
         );
  NAND2_X2 U8110 ( .A1(\REGFILE/reg_out[30][24] ), .A2(net77568), .ZN(n7182)
         );
  NAND2_X2 U8111 ( .A1(\REGFILE/reg_out[25][24] ), .A2(net77532), .ZN(n7181)
         );
  NAND2_X2 U8112 ( .A1(\REGFILE/reg_out[31][24] ), .A2(net77496), .ZN(n7180)
         );
  NAND2_X2 U8113 ( .A1(\REGFILE/reg_out[29][24] ), .A2(net77460), .ZN(n7179)
         );
  NAND4_X2 U8114 ( .A1(n7182), .A2(n7181), .A3(n7180), .A4(n7179), .ZN(n7183)
         );
  NAND2_X2 U8115 ( .A1(\REGFILE/reg_out[3][24] ), .A2(net77424), .ZN(n7188) );
  NAND2_X2 U8117 ( .A1(\REGFILE/reg_out[2][24] ), .A2(n6016), .ZN(n7186) );
  NAND2_X2 U8118 ( .A1(\REGFILE/reg_out[0][24] ), .A2(net77316), .ZN(n7185) );
  NAND4_X2 U8119 ( .A1(n7188), .A2(n7187), .A3(n7186), .A4(n7185), .ZN(n7194)
         );
  NAND2_X2 U8120 ( .A1(\REGFILE/reg_out[6][24] ), .A2(net77568), .ZN(n7192) );
  NAND2_X2 U8121 ( .A1(\REGFILE/reg_out[1][24] ), .A2(net77532), .ZN(n7191) );
  NAND2_X2 U8122 ( .A1(\REGFILE/reg_out[7][24] ), .A2(net77496), .ZN(n7190) );
  NAND2_X2 U8123 ( .A1(\REGFILE/reg_out[5][24] ), .A2(net77460), .ZN(n7189) );
  NAND4_X2 U8124 ( .A1(n7192), .A2(n7191), .A3(n7190), .A4(n7189), .ZN(n7193)
         );
  NAND2_X2 U8125 ( .A1(\REGFILE/reg_out[11][24] ), .A2(net77424), .ZN(n7198)
         );
  NAND2_X2 U8127 ( .A1(\REGFILE/reg_out[10][24] ), .A2(n6016), .ZN(n7196) );
  NAND2_X2 U8128 ( .A1(\REGFILE/reg_out[8][24] ), .A2(net77316), .ZN(n7195) );
  NAND4_X2 U8129 ( .A1(n7198), .A2(n7197), .A3(n7196), .A4(n7195), .ZN(n7204)
         );
  NAND2_X2 U8130 ( .A1(\REGFILE/reg_out[14][24] ), .A2(net77568), .ZN(n7202)
         );
  NAND2_X2 U8131 ( .A1(\REGFILE/reg_out[9][24] ), .A2(net77532), .ZN(n7201) );
  NAND2_X2 U8132 ( .A1(\REGFILE/reg_out[15][24] ), .A2(net77496), .ZN(n7200)
         );
  NAND2_X2 U8133 ( .A1(\REGFILE/reg_out[13][24] ), .A2(net77460), .ZN(n7199)
         );
  NAND4_X2 U8134 ( .A1(n7202), .A2(n7201), .A3(n7200), .A4(n7199), .ZN(n7203)
         );
  NAND2_X2 U8135 ( .A1(\REGFILE/reg_out[19][24] ), .A2(net77424), .ZN(n7208)
         );
  NAND2_X2 U8137 ( .A1(\REGFILE/reg_out[18][24] ), .A2(n6016), .ZN(n7206) );
  NAND2_X2 U8138 ( .A1(\REGFILE/reg_out[16][24] ), .A2(net77316), .ZN(n7205)
         );
  NAND4_X2 U8139 ( .A1(n7208), .A2(n7207), .A3(n7206), .A4(n7205), .ZN(n7214)
         );
  NAND2_X2 U8140 ( .A1(\REGFILE/reg_out[22][24] ), .A2(net77568), .ZN(n7212)
         );
  NAND2_X2 U8141 ( .A1(\REGFILE/reg_out[17][24] ), .A2(net77532), .ZN(n7211)
         );
  NAND2_X2 U8142 ( .A1(\REGFILE/reg_out[23][24] ), .A2(net77496), .ZN(n7210)
         );
  NAND2_X2 U8143 ( .A1(\REGFILE/reg_out[21][24] ), .A2(net77460), .ZN(n7209)
         );
  NAND4_X2 U8144 ( .A1(n7212), .A2(n7211), .A3(n7210), .A4(n7209), .ZN(n7213)
         );
  NAND4_X2 U8145 ( .A1(n7218), .A2(n7217), .A3(n7216), .A4(n7215), .ZN(n8420)
         );
  INV_X4 U8146 ( .A(n8420), .ZN(n7219) );
  INV_X4 U8147 ( .A(\PCLOGIC/imm16_32 [24]), .ZN(n8351) );
  MUX2_X2 U8148 ( .A(n7219), .B(n8351), .S(net77276), .Z(net72312) );
  INV_X4 U8149 ( .A(net72312), .ZN(net36391) );
  NAND2_X2 U8150 ( .A1(\REGFILE/reg_out[27][23] ), .A2(net77424), .ZN(n7223)
         );
  NAND2_X2 U8152 ( .A1(\REGFILE/reg_out[26][23] ), .A2(n6016), .ZN(n7221) );
  NAND2_X2 U8153 ( .A1(\REGFILE/reg_out[24][23] ), .A2(net77316), .ZN(n7220)
         );
  NAND4_X2 U8154 ( .A1(n7223), .A2(n7222), .A3(n7221), .A4(n7220), .ZN(n7229)
         );
  NAND2_X2 U8155 ( .A1(\REGFILE/reg_out[30][23] ), .A2(net77568), .ZN(n7227)
         );
  NAND2_X2 U8156 ( .A1(\REGFILE/reg_out[25][23] ), .A2(net77532), .ZN(n7226)
         );
  NAND2_X2 U8157 ( .A1(\REGFILE/reg_out[31][23] ), .A2(net77496), .ZN(n7225)
         );
  NAND2_X2 U8158 ( .A1(\REGFILE/reg_out[29][23] ), .A2(net77460), .ZN(n7224)
         );
  NAND4_X2 U8159 ( .A1(n7227), .A2(n7226), .A3(n7225), .A4(n7224), .ZN(n7228)
         );
  NAND2_X2 U8160 ( .A1(\REGFILE/reg_out[3][23] ), .A2(net77424), .ZN(n7233) );
  NAND2_X2 U8162 ( .A1(\REGFILE/reg_out[2][23] ), .A2(n6016), .ZN(n7231) );
  NAND2_X2 U8163 ( .A1(\REGFILE/reg_out[0][23] ), .A2(net77316), .ZN(n7230) );
  NAND4_X2 U8164 ( .A1(n7233), .A2(n7232), .A3(n7231), .A4(n7230), .ZN(n7239)
         );
  NAND2_X2 U8165 ( .A1(\REGFILE/reg_out[6][23] ), .A2(net77568), .ZN(n7237) );
  NAND2_X2 U8166 ( .A1(\REGFILE/reg_out[1][23] ), .A2(net77532), .ZN(n7236) );
  NAND2_X2 U8167 ( .A1(\REGFILE/reg_out[7][23] ), .A2(net77496), .ZN(n7235) );
  NAND2_X2 U8168 ( .A1(\REGFILE/reg_out[5][23] ), .A2(net77460), .ZN(n7234) );
  NAND4_X2 U8169 ( .A1(n7237), .A2(n7236), .A3(n7235), .A4(n7234), .ZN(n7238)
         );
  NAND2_X2 U8170 ( .A1(\REGFILE/reg_out[11][23] ), .A2(net77424), .ZN(n7243)
         );
  NAND2_X2 U8172 ( .A1(\REGFILE/reg_out[10][23] ), .A2(n6016), .ZN(n7241) );
  NAND2_X2 U8173 ( .A1(\REGFILE/reg_out[8][23] ), .A2(net77316), .ZN(n7240) );
  NAND4_X2 U8174 ( .A1(n7243), .A2(n7242), .A3(n7241), .A4(n7240), .ZN(n7249)
         );
  NAND2_X2 U8175 ( .A1(\REGFILE/reg_out[14][23] ), .A2(net77568), .ZN(n7247)
         );
  NAND2_X2 U8176 ( .A1(\REGFILE/reg_out[9][23] ), .A2(net77532), .ZN(n7246) );
  NAND2_X2 U8177 ( .A1(\REGFILE/reg_out[15][23] ), .A2(net77496), .ZN(n7245)
         );
  NAND2_X2 U8178 ( .A1(\REGFILE/reg_out[13][23] ), .A2(net77460), .ZN(n7244)
         );
  NAND4_X2 U8179 ( .A1(n7247), .A2(n7246), .A3(n7245), .A4(n7244), .ZN(n7248)
         );
  NAND2_X2 U8180 ( .A1(\REGFILE/reg_out[19][23] ), .A2(net77424), .ZN(n7253)
         );
  NAND2_X2 U8182 ( .A1(\REGFILE/reg_out[18][23] ), .A2(n6016), .ZN(n7251) );
  NAND2_X2 U8183 ( .A1(\REGFILE/reg_out[16][23] ), .A2(net77316), .ZN(n7250)
         );
  NAND4_X2 U8184 ( .A1(n7253), .A2(n7252), .A3(n7251), .A4(n7250), .ZN(n7259)
         );
  NAND2_X2 U8185 ( .A1(\REGFILE/reg_out[22][23] ), .A2(net77568), .ZN(n7257)
         );
  NAND2_X2 U8186 ( .A1(\REGFILE/reg_out[17][23] ), .A2(net77532), .ZN(n7256)
         );
  NAND2_X2 U8187 ( .A1(\REGFILE/reg_out[23][23] ), .A2(net77496), .ZN(n7255)
         );
  NAND2_X2 U8188 ( .A1(\REGFILE/reg_out[21][23] ), .A2(net77460), .ZN(n7254)
         );
  NAND4_X2 U8189 ( .A1(n7257), .A2(n7256), .A3(n7255), .A4(n7254), .ZN(n7258)
         );
  NAND4_X2 U8190 ( .A1(n7263), .A2(n7262), .A3(n7261), .A4(n7260), .ZN(n8418)
         );
  INV_X4 U8191 ( .A(n8418), .ZN(n7264) );
  INV_X4 U8192 ( .A(\PCLOGIC/imm16_32 [23]), .ZN(n8324) );
  MUX2_X2 U8193 ( .A(n7264), .B(n8324), .S(net77276), .Z(n10334) );
  INV_X4 U8194 ( .A(n10334), .ZN(n10931) );
  NAND2_X2 U8195 ( .A1(\REGFILE/reg_out[27][22] ), .A2(net77424), .ZN(n7268)
         );
  NAND2_X2 U8197 ( .A1(\REGFILE/reg_out[26][22] ), .A2(n6016), .ZN(n7266) );
  NAND2_X2 U8198 ( .A1(\REGFILE/reg_out[24][22] ), .A2(net77316), .ZN(n7265)
         );
  NAND4_X2 U8199 ( .A1(n7268), .A2(n7267), .A3(n7266), .A4(n7265), .ZN(n7274)
         );
  NAND2_X2 U8200 ( .A1(\REGFILE/reg_out[30][22] ), .A2(net77568), .ZN(n7272)
         );
  NAND2_X2 U8201 ( .A1(\REGFILE/reg_out[25][22] ), .A2(net77532), .ZN(n7271)
         );
  NAND2_X2 U8202 ( .A1(\REGFILE/reg_out[31][22] ), .A2(net77496), .ZN(n7270)
         );
  NAND2_X2 U8203 ( .A1(\REGFILE/reg_out[29][22] ), .A2(net77460), .ZN(n7269)
         );
  NAND4_X2 U8204 ( .A1(n7272), .A2(n7271), .A3(n7270), .A4(n7269), .ZN(n7273)
         );
  NAND2_X2 U8205 ( .A1(\REGFILE/reg_out[3][22] ), .A2(net77422), .ZN(n7278) );
  NAND2_X2 U8206 ( .A1(\REGFILE/reg_out[2][22] ), .A2(n6015), .ZN(n7276) );
  NAND2_X2 U8207 ( .A1(\REGFILE/reg_out[0][22] ), .A2(net77314), .ZN(n7275) );
  NAND4_X2 U8208 ( .A1(n7278), .A2(n7277), .A3(n7276), .A4(n7275), .ZN(n7284)
         );
  NAND2_X2 U8209 ( .A1(\REGFILE/reg_out[6][22] ), .A2(net77566), .ZN(n7282) );
  NAND2_X2 U8210 ( .A1(\REGFILE/reg_out[1][22] ), .A2(net77530), .ZN(n7281) );
  NAND2_X2 U8211 ( .A1(\REGFILE/reg_out[7][22] ), .A2(net77494), .ZN(n7280) );
  NAND2_X2 U8212 ( .A1(\REGFILE/reg_out[5][22] ), .A2(net77458), .ZN(n7279) );
  NAND4_X2 U8213 ( .A1(n7282), .A2(n7281), .A3(n7280), .A4(n7279), .ZN(n7283)
         );
  NAND2_X2 U8214 ( .A1(\REGFILE/reg_out[11][22] ), .A2(net77422), .ZN(n7288)
         );
  NAND2_X2 U8215 ( .A1(\REGFILE/reg_out[8][22] ), .A2(net77314), .ZN(n7285) );
  NAND4_X2 U8216 ( .A1(n7288), .A2(n7287), .A3(n7286), .A4(n7285), .ZN(n7294)
         );
  NAND2_X2 U8217 ( .A1(\REGFILE/reg_out[14][22] ), .A2(net77566), .ZN(n7292)
         );
  NAND2_X2 U8218 ( .A1(\REGFILE/reg_out[9][22] ), .A2(net77530), .ZN(n7291) );
  NAND2_X2 U8219 ( .A1(\REGFILE/reg_out[15][22] ), .A2(net77494), .ZN(n7290)
         );
  NAND2_X2 U8220 ( .A1(\REGFILE/reg_out[13][22] ), .A2(net77458), .ZN(n7289)
         );
  NAND4_X2 U8221 ( .A1(n7292), .A2(n7291), .A3(n7290), .A4(n7289), .ZN(n7293)
         );
  NAND2_X2 U8222 ( .A1(\REGFILE/reg_out[19][22] ), .A2(net77422), .ZN(n7298)
         );
  NAND2_X2 U8223 ( .A1(\REGFILE/reg_out[18][22] ), .A2(n6015), .ZN(n7296) );
  NAND2_X2 U8224 ( .A1(\REGFILE/reg_out[16][22] ), .A2(net77314), .ZN(n7295)
         );
  NAND4_X2 U8225 ( .A1(n7298), .A2(n7297), .A3(n7296), .A4(n7295), .ZN(n7304)
         );
  NAND2_X2 U8226 ( .A1(\REGFILE/reg_out[22][22] ), .A2(net77566), .ZN(n7302)
         );
  NAND2_X2 U8227 ( .A1(\REGFILE/reg_out[17][22] ), .A2(net77530), .ZN(n7301)
         );
  NAND2_X2 U8228 ( .A1(\REGFILE/reg_out[23][22] ), .A2(net77494), .ZN(n7300)
         );
  NAND2_X2 U8229 ( .A1(\REGFILE/reg_out[21][22] ), .A2(net77458), .ZN(n7299)
         );
  NAND4_X2 U8230 ( .A1(n7302), .A2(n7301), .A3(n7300), .A4(n7299), .ZN(n7303)
         );
  NAND4_X2 U8231 ( .A1(n7308), .A2(n7307), .A3(n7306), .A4(n7305), .ZN(n8400)
         );
  INV_X4 U8232 ( .A(n8400), .ZN(n7309) );
  INV_X4 U8233 ( .A(\PCLOGIC/imm16_32 [22]), .ZN(n8355) );
  MUX2_X2 U8234 ( .A(n7309), .B(n8355), .S(net77276), .Z(n8967) );
  INV_X4 U8235 ( .A(n8967), .ZN(n10932) );
  NAND2_X2 U8236 ( .A1(\REGFILE/reg_out[26][21] ), .A2(n6015), .ZN(n7311) );
  NAND2_X2 U8237 ( .A1(\REGFILE/reg_out[24][21] ), .A2(net77314), .ZN(n7310)
         );
  NAND4_X2 U8238 ( .A1(n7313), .A2(n7312), .A3(n7311), .A4(n7310), .ZN(n7319)
         );
  NAND2_X2 U8239 ( .A1(\REGFILE/reg_out[30][21] ), .A2(net77566), .ZN(n7317)
         );
  NAND2_X2 U8240 ( .A1(\REGFILE/reg_out[31][21] ), .A2(net77494), .ZN(n7315)
         );
  NAND2_X2 U8241 ( .A1(\REGFILE/reg_out[29][21] ), .A2(net77458), .ZN(n7314)
         );
  NAND4_X2 U8242 ( .A1(n7317), .A2(n7316), .A3(n7315), .A4(n7314), .ZN(n7318)
         );
  NAND2_X2 U8243 ( .A1(\REGFILE/reg_out[3][21] ), .A2(net77422), .ZN(n7323) );
  NAND2_X2 U8244 ( .A1(\REGFILE/reg_out[2][21] ), .A2(n6015), .ZN(n7321) );
  NAND2_X2 U8245 ( .A1(\REGFILE/reg_out[0][21] ), .A2(net77314), .ZN(n7320) );
  NAND4_X2 U8246 ( .A1(n7323), .A2(n7322), .A3(n7321), .A4(n7320), .ZN(n7329)
         );
  NAND2_X2 U8247 ( .A1(\REGFILE/reg_out[6][21] ), .A2(net77566), .ZN(n7327) );
  NAND2_X2 U8248 ( .A1(\REGFILE/reg_out[1][21] ), .A2(net77530), .ZN(n7326) );
  NAND2_X2 U8249 ( .A1(\REGFILE/reg_out[7][21] ), .A2(net77494), .ZN(n7325) );
  NAND2_X2 U8250 ( .A1(\REGFILE/reg_out[5][21] ), .A2(net77458), .ZN(n7324) );
  NAND4_X2 U8251 ( .A1(n7327), .A2(n7326), .A3(n7325), .A4(n7324), .ZN(n7328)
         );
  NAND2_X2 U8252 ( .A1(\REGFILE/reg_out[11][21] ), .A2(net77422), .ZN(n7333)
         );
  NAND2_X2 U8253 ( .A1(\REGFILE/reg_out[10][21] ), .A2(n6015), .ZN(n7331) );
  NAND2_X2 U8254 ( .A1(\REGFILE/reg_out[8][21] ), .A2(net77314), .ZN(n7330) );
  NAND4_X2 U8255 ( .A1(n7333), .A2(n7332), .A3(n7331), .A4(n7330), .ZN(n7339)
         );
  NAND2_X2 U8256 ( .A1(\REGFILE/reg_out[14][21] ), .A2(net77566), .ZN(n7337)
         );
  NAND2_X2 U8257 ( .A1(\REGFILE/reg_out[9][21] ), .A2(net77530), .ZN(n7336) );
  NAND2_X2 U8258 ( .A1(\REGFILE/reg_out[15][21] ), .A2(net77494), .ZN(n7335)
         );
  NAND2_X2 U8259 ( .A1(\REGFILE/reg_out[13][21] ), .A2(net77458), .ZN(n7334)
         );
  NAND4_X2 U8260 ( .A1(n7337), .A2(n7336), .A3(n7335), .A4(n7334), .ZN(n7338)
         );
  NAND2_X2 U8261 ( .A1(\REGFILE/reg_out[19][21] ), .A2(net77422), .ZN(n7343)
         );
  NAND2_X2 U8262 ( .A1(\REGFILE/reg_out[18][21] ), .A2(n6015), .ZN(n7341) );
  NAND2_X2 U8263 ( .A1(\REGFILE/reg_out[16][21] ), .A2(net77314), .ZN(n7340)
         );
  NAND4_X2 U8264 ( .A1(n7343), .A2(n7342), .A3(n7341), .A4(n7340), .ZN(n7349)
         );
  NAND2_X2 U8265 ( .A1(\REGFILE/reg_out[22][21] ), .A2(net77566), .ZN(n7347)
         );
  NAND2_X2 U8266 ( .A1(\REGFILE/reg_out[17][21] ), .A2(net77530), .ZN(n7346)
         );
  NAND2_X2 U8267 ( .A1(\REGFILE/reg_out[23][21] ), .A2(net77494), .ZN(n7345)
         );
  NAND2_X2 U8268 ( .A1(\REGFILE/reg_out[21][21] ), .A2(net77458), .ZN(n7344)
         );
  NAND4_X2 U8269 ( .A1(n7347), .A2(n7346), .A3(n7345), .A4(n7344), .ZN(n7348)
         );
  NAND4_X2 U8270 ( .A1(n7353), .A2(n7352), .A3(n7351), .A4(n7350), .ZN(n8417)
         );
  INV_X4 U8271 ( .A(n8417), .ZN(n7354) );
  INV_X4 U8272 ( .A(\PCLOGIC/imm16_32 [21]), .ZN(n8319) );
  MUX2_X2 U8273 ( .A(n7354), .B(n8319), .S(net77276), .Z(n10341) );
  INV_X4 U8274 ( .A(n10341), .ZN(n10933) );
  NAND2_X2 U8275 ( .A1(\REGFILE/reg_out[30][20] ), .A2(net77566), .ZN(n7358)
         );
  NAND2_X2 U8276 ( .A1(\REGFILE/reg_out[31][20] ), .A2(net77494), .ZN(n7356)
         );
  NAND2_X2 U8277 ( .A1(\REGFILE/reg_out[29][20] ), .A2(net77458), .ZN(n7355)
         );
  NAND4_X2 U8278 ( .A1(n7358), .A2(n7357), .A3(n7356), .A4(n7355), .ZN(n7364)
         );
  NAND2_X2 U8279 ( .A1(\REGFILE/reg_out[26][20] ), .A2(n6015), .ZN(n7360) );
  NAND2_X2 U8280 ( .A1(\REGFILE/reg_out[24][20] ), .A2(net77314), .ZN(n7359)
         );
  NAND4_X2 U8281 ( .A1(n7362), .A2(n7361), .A3(n7360), .A4(n7359), .ZN(n7363)
         );
  NAND2_X2 U8282 ( .A1(\REGFILE/reg_out[22][20] ), .A2(net77566), .ZN(n7368)
         );
  NAND2_X2 U8283 ( .A1(\REGFILE/reg_out[17][20] ), .A2(net77530), .ZN(n7367)
         );
  NAND2_X2 U8284 ( .A1(\REGFILE/reg_out[23][20] ), .A2(net77494), .ZN(n7366)
         );
  NAND2_X2 U8285 ( .A1(\REGFILE/reg_out[21][20] ), .A2(net77458), .ZN(n7365)
         );
  NAND4_X2 U8286 ( .A1(n7368), .A2(n7367), .A3(n7366), .A4(n7365), .ZN(n7374)
         );
  NAND2_X2 U8287 ( .A1(\REGFILE/reg_out[19][20] ), .A2(net77422), .ZN(n7372)
         );
  NAND2_X2 U8288 ( .A1(\REGFILE/reg_out[18][20] ), .A2(n6015), .ZN(n7370) );
  NAND2_X2 U8289 ( .A1(\REGFILE/reg_out[16][20] ), .A2(net77314), .ZN(n7369)
         );
  NAND4_X2 U8290 ( .A1(n7372), .A2(n7371), .A3(n7370), .A4(n7369), .ZN(n7373)
         );
  NAND2_X2 U8291 ( .A1(\REGFILE/reg_out[14][20] ), .A2(net77566), .ZN(n7378)
         );
  NAND2_X2 U8292 ( .A1(\REGFILE/reg_out[9][20] ), .A2(net77530), .ZN(n7377) );
  NAND2_X2 U8293 ( .A1(\REGFILE/reg_out[15][20] ), .A2(net77494), .ZN(n7376)
         );
  NAND2_X2 U8294 ( .A1(\REGFILE/reg_out[13][20] ), .A2(net77458), .ZN(n7375)
         );
  NAND4_X2 U8295 ( .A1(n7378), .A2(n7377), .A3(n7376), .A4(n7375), .ZN(n7384)
         );
  NAND2_X2 U8296 ( .A1(\REGFILE/reg_out[11][20] ), .A2(net77422), .ZN(n7382)
         );
  NAND2_X2 U8297 ( .A1(\REGFILE/reg_out[10][20] ), .A2(n6015), .ZN(n7380) );
  NAND2_X2 U8298 ( .A1(\REGFILE/reg_out[8][20] ), .A2(net77314), .ZN(n7379) );
  NAND4_X2 U8299 ( .A1(n7382), .A2(n7381), .A3(n7380), .A4(n7379), .ZN(n7383)
         );
  NAND2_X2 U8300 ( .A1(\REGFILE/reg_out[6][20] ), .A2(net77566), .ZN(n7388) );
  NAND2_X2 U8301 ( .A1(\REGFILE/reg_out[1][20] ), .A2(net77530), .ZN(n7387) );
  NAND2_X2 U8302 ( .A1(\REGFILE/reg_out[7][20] ), .A2(net77494), .ZN(n7386) );
  NAND2_X2 U8303 ( .A1(\REGFILE/reg_out[5][20] ), .A2(net77458), .ZN(n7385) );
  NAND4_X2 U8304 ( .A1(n7388), .A2(n7387), .A3(n7386), .A4(n7385), .ZN(n7394)
         );
  NAND2_X2 U8305 ( .A1(\REGFILE/reg_out[0][20] ), .A2(net77314), .ZN(n7389) );
  NAND4_X2 U8306 ( .A1(n7392), .A2(n7391), .A3(n7390), .A4(n7389), .ZN(n7393)
         );
  NAND4_X2 U8307 ( .A1(n7398), .A2(n7397), .A3(n7396), .A4(n7395), .ZN(n8449)
         );
  MUX2_X2 U8308 ( .A(n8449), .B(\PCLOGIC/imm16_32 [20]), .S(net77276), .Z(
        aluA[20]) );
  NAND2_X2 U8309 ( .A1(\REGFILE/reg_out[30][19] ), .A2(net77566), .ZN(n7402)
         );
  NAND2_X2 U8310 ( .A1(\REGFILE/reg_out[25][19] ), .A2(net77530), .ZN(n7401)
         );
  NAND2_X2 U8311 ( .A1(\REGFILE/reg_out[31][19] ), .A2(net77494), .ZN(n7400)
         );
  NAND2_X2 U8312 ( .A1(\REGFILE/reg_out[29][19] ), .A2(net77458), .ZN(n7399)
         );
  NAND4_X2 U8313 ( .A1(n7402), .A2(n7401), .A3(n7400), .A4(n7399), .ZN(n7408)
         );
  NAND2_X2 U8314 ( .A1(\REGFILE/reg_out[26][19] ), .A2(n6015), .ZN(n7404) );
  NAND2_X2 U8315 ( .A1(\REGFILE/reg_out[24][19] ), .A2(net77314), .ZN(n7403)
         );
  NAND4_X2 U8316 ( .A1(n7406), .A2(n7405), .A3(n7404), .A4(n7403), .ZN(n7407)
         );
  NAND2_X2 U8317 ( .A1(\REGFILE/reg_out[22][19] ), .A2(net77564), .ZN(n7412)
         );
  NAND2_X2 U8318 ( .A1(\REGFILE/reg_out[17][19] ), .A2(net77528), .ZN(n7411)
         );
  NAND2_X2 U8319 ( .A1(\REGFILE/reg_out[23][19] ), .A2(net77492), .ZN(n7410)
         );
  NAND2_X2 U8320 ( .A1(\REGFILE/reg_out[21][19] ), .A2(net77456), .ZN(n7409)
         );
  NAND4_X2 U8321 ( .A1(n7412), .A2(n7411), .A3(n7410), .A4(n7409), .ZN(n7418)
         );
  NAND2_X2 U8322 ( .A1(\REGFILE/reg_out[19][19] ), .A2(net77420), .ZN(n7416)
         );
  NAND2_X2 U8323 ( .A1(\REGFILE/reg_out[20][19] ), .A2(net77384), .ZN(n7415)
         );
  NAND2_X2 U8324 ( .A1(\REGFILE/reg_out[18][19] ), .A2(net77348), .ZN(n7414)
         );
  NAND2_X2 U8325 ( .A1(\REGFILE/reg_out[16][19] ), .A2(net77312), .ZN(n7413)
         );
  NAND4_X2 U8326 ( .A1(n7416), .A2(n7415), .A3(n7414), .A4(n7413), .ZN(n7417)
         );
  NAND2_X2 U8327 ( .A1(\REGFILE/reg_out[14][19] ), .A2(net77564), .ZN(n7422)
         );
  NAND2_X2 U8328 ( .A1(\REGFILE/reg_out[9][19] ), .A2(net77528), .ZN(n7421) );
  NAND2_X2 U8329 ( .A1(\REGFILE/reg_out[15][19] ), .A2(net77492), .ZN(n7420)
         );
  NAND2_X2 U8330 ( .A1(\REGFILE/reg_out[13][19] ), .A2(net77456), .ZN(n7419)
         );
  NAND4_X2 U8331 ( .A1(n7422), .A2(n7421), .A3(n7420), .A4(n7419), .ZN(n7428)
         );
  NAND2_X2 U8332 ( .A1(\REGFILE/reg_out[11][19] ), .A2(net77420), .ZN(n7426)
         );
  NAND2_X2 U8333 ( .A1(\REGFILE/reg_out[8][19] ), .A2(net77312), .ZN(n7423) );
  NAND4_X2 U8334 ( .A1(n7426), .A2(n7425), .A3(n7424), .A4(n7423), .ZN(n7427)
         );
  NAND2_X2 U8335 ( .A1(\REGFILE/reg_out[6][19] ), .A2(net77564), .ZN(n7432) );
  NAND2_X2 U8336 ( .A1(\REGFILE/reg_out[1][19] ), .A2(net77528), .ZN(n7431) );
  NAND2_X2 U8337 ( .A1(\REGFILE/reg_out[7][19] ), .A2(net77492), .ZN(n7430) );
  NAND2_X2 U8338 ( .A1(\REGFILE/reg_out[5][19] ), .A2(net77456), .ZN(n7429) );
  NAND4_X2 U8339 ( .A1(n7432), .A2(n7431), .A3(n7430), .A4(n7429), .ZN(n7438)
         );
  NAND2_X2 U8340 ( .A1(\REGFILE/reg_out[3][19] ), .A2(net77420), .ZN(n7436) );
  NAND2_X2 U8341 ( .A1(\REGFILE/reg_out[4][19] ), .A2(net77384), .ZN(n7435) );
  NAND2_X2 U8342 ( .A1(\REGFILE/reg_out[2][19] ), .A2(net77348), .ZN(n7434) );
  NAND2_X2 U8343 ( .A1(\REGFILE/reg_out[0][19] ), .A2(net77312), .ZN(n7433) );
  NAND4_X2 U8344 ( .A1(n7436), .A2(n7435), .A3(n7434), .A4(n7433), .ZN(n7437)
         );
  NAND4_X2 U8345 ( .A1(n7442), .A2(n7441), .A3(n7440), .A4(n7439), .ZN(n8444)
         );
  MUX2_X2 U8346 ( .A(n8444), .B(\PCLOGIC/imm16_32 [19]), .S(net77276), .Z(
        aluA[19]) );
  NAND2_X2 U8347 ( .A1(\REGFILE/reg_out[30][18] ), .A2(net77564), .ZN(n7446)
         );
  NAND2_X2 U8348 ( .A1(net77528), .A2(\REGFILE/reg_out[25][18] ), .ZN(n7445)
         );
  NAND2_X2 U8349 ( .A1(\REGFILE/reg_out[31][18] ), .A2(net77492), .ZN(n7444)
         );
  NAND2_X2 U8350 ( .A1(\REGFILE/reg_out[29][18] ), .A2(net77456), .ZN(n7443)
         );
  NAND4_X2 U8351 ( .A1(n7446), .A2(n7445), .A3(n7444), .A4(n7443), .ZN(n7452)
         );
  NAND2_X2 U8352 ( .A1(\REGFILE/reg_out[26][18] ), .A2(net77348), .ZN(n7448)
         );
  NAND2_X2 U8353 ( .A1(\REGFILE/reg_out[24][18] ), .A2(net77312), .ZN(n7447)
         );
  NAND4_X2 U8354 ( .A1(n7450), .A2(n7449), .A3(n7448), .A4(n7447), .ZN(n7451)
         );
  NAND2_X2 U8355 ( .A1(\REGFILE/reg_out[22][18] ), .A2(net77564), .ZN(n7456)
         );
  NAND2_X2 U8356 ( .A1(\REGFILE/reg_out[17][18] ), .A2(net77528), .ZN(n7455)
         );
  NAND2_X2 U8357 ( .A1(\REGFILE/reg_out[23][18] ), .A2(net77492), .ZN(n7454)
         );
  NAND2_X2 U8358 ( .A1(\REGFILE/reg_out[21][18] ), .A2(net77456), .ZN(n7453)
         );
  NAND4_X2 U8359 ( .A1(n7456), .A2(n7455), .A3(n7454), .A4(n7453), .ZN(n7462)
         );
  NAND2_X2 U8360 ( .A1(\REGFILE/reg_out[19][18] ), .A2(net77420), .ZN(n7460)
         );
  NAND2_X2 U8361 ( .A1(\REGFILE/reg_out[20][18] ), .A2(net77384), .ZN(n7459)
         );
  NAND2_X2 U8362 ( .A1(\REGFILE/reg_out[18][18] ), .A2(net77348), .ZN(n7458)
         );
  NAND2_X2 U8363 ( .A1(\REGFILE/reg_out[16][18] ), .A2(net77312), .ZN(n7457)
         );
  NAND4_X2 U8364 ( .A1(n7460), .A2(n7459), .A3(n7458), .A4(n7457), .ZN(n7461)
         );
  NAND2_X2 U8365 ( .A1(\REGFILE/reg_out[14][18] ), .A2(net77564), .ZN(n7466)
         );
  NAND2_X2 U8366 ( .A1(\REGFILE/reg_out[9][18] ), .A2(net77528), .ZN(n7465) );
  NAND2_X2 U8367 ( .A1(\REGFILE/reg_out[15][18] ), .A2(net77492), .ZN(n7464)
         );
  NAND2_X2 U8368 ( .A1(\REGFILE/reg_out[13][18] ), .A2(net77456), .ZN(n7463)
         );
  NAND4_X2 U8369 ( .A1(n7466), .A2(n7465), .A3(n7464), .A4(n7463), .ZN(n7472)
         );
  NAND2_X2 U8370 ( .A1(\REGFILE/reg_out[11][18] ), .A2(net77420), .ZN(n7470)
         );
  NAND2_X2 U8371 ( .A1(\REGFILE/reg_out[10][18] ), .A2(net77348), .ZN(n7468)
         );
  NAND2_X2 U8372 ( .A1(\REGFILE/reg_out[8][18] ), .A2(net77312), .ZN(n7467) );
  NAND4_X2 U8373 ( .A1(n7470), .A2(n7469), .A3(n7468), .A4(n7467), .ZN(n7471)
         );
  NAND2_X2 U8374 ( .A1(\REGFILE/reg_out[6][18] ), .A2(net77564), .ZN(n7476) );
  NAND2_X2 U8375 ( .A1(\REGFILE/reg_out[1][18] ), .A2(net77528), .ZN(n7475) );
  NAND2_X2 U8376 ( .A1(\REGFILE/reg_out[7][18] ), .A2(net77492), .ZN(n7474) );
  NAND4_X2 U8377 ( .A1(n7476), .A2(n7475), .A3(n7474), .A4(n7473), .ZN(n7482)
         );
  NAND2_X2 U8378 ( .A1(\REGFILE/reg_out[3][18] ), .A2(net77420), .ZN(n7480) );
  NAND2_X2 U8379 ( .A1(\REGFILE/reg_out[4][18] ), .A2(net77384), .ZN(n7479) );
  NAND2_X2 U8380 ( .A1(\REGFILE/reg_out[0][18] ), .A2(net77312), .ZN(n7477) );
  NAND4_X2 U8381 ( .A1(n7480), .A2(n7479), .A3(n7478), .A4(n7477), .ZN(n7481)
         );
  NAND4_X2 U8382 ( .A1(n7486), .A2(n7485), .A3(n7484), .A4(n7483), .ZN(n8443)
         );
  MUX2_X2 U8383 ( .A(n8443), .B(\PCLOGIC/imm16_32 [18]), .S(net77276), .Z(
        aluA[18]) );
  NAND2_X2 U8384 ( .A1(\REGFILE/reg_out[30][17] ), .A2(net77564), .ZN(n7490)
         );
  NAND2_X2 U8385 ( .A1(\REGFILE/reg_out[31][17] ), .A2(net77492), .ZN(n7488)
         );
  NAND2_X2 U8386 ( .A1(\REGFILE/reg_out[29][17] ), .A2(net77456), .ZN(n7487)
         );
  NAND4_X2 U8387 ( .A1(n7490), .A2(n7489), .A3(n7488), .A4(n7487), .ZN(n7496)
         );
  NAND2_X2 U8388 ( .A1(\REGFILE/reg_out[28][17] ), .A2(net77384), .ZN(n7493)
         );
  NAND2_X2 U8389 ( .A1(\REGFILE/reg_out[26][17] ), .A2(net77348), .ZN(n7492)
         );
  NAND2_X2 U8390 ( .A1(\REGFILE/reg_out[24][17] ), .A2(net77312), .ZN(n7491)
         );
  NAND4_X2 U8391 ( .A1(n7494), .A2(n7493), .A3(n7492), .A4(n7491), .ZN(n7495)
         );
  NAND2_X2 U8392 ( .A1(\REGFILE/reg_out[22][17] ), .A2(net77564), .ZN(n7500)
         );
  NAND2_X2 U8393 ( .A1(\REGFILE/reg_out[17][17] ), .A2(net77528), .ZN(n7499)
         );
  NAND2_X2 U8394 ( .A1(\REGFILE/reg_out[23][17] ), .A2(net77492), .ZN(n7498)
         );
  NAND2_X2 U8395 ( .A1(\REGFILE/reg_out[21][17] ), .A2(net77456), .ZN(n7497)
         );
  NAND4_X2 U8396 ( .A1(n7500), .A2(n7499), .A3(n7498), .A4(n7497), .ZN(n7506)
         );
  NAND2_X2 U8397 ( .A1(\REGFILE/reg_out[19][17] ), .A2(net77420), .ZN(n7504)
         );
  NAND2_X2 U8398 ( .A1(\REGFILE/reg_out[20][17] ), .A2(net77384), .ZN(n7503)
         );
  NAND2_X2 U8399 ( .A1(\REGFILE/reg_out[18][17] ), .A2(net77348), .ZN(n7502)
         );
  NAND2_X2 U8400 ( .A1(\REGFILE/reg_out[16][17] ), .A2(net77312), .ZN(n7501)
         );
  NAND4_X2 U8401 ( .A1(n7504), .A2(n7503), .A3(n7502), .A4(n7501), .ZN(n7505)
         );
  NAND2_X2 U8402 ( .A1(\REGFILE/reg_out[14][17] ), .A2(net77564), .ZN(n7510)
         );
  NAND2_X2 U8403 ( .A1(\REGFILE/reg_out[9][17] ), .A2(net77528), .ZN(n7509) );
  NAND2_X2 U8404 ( .A1(\REGFILE/reg_out[15][17] ), .A2(net77492), .ZN(n7508)
         );
  NAND2_X2 U8405 ( .A1(\REGFILE/reg_out[13][17] ), .A2(net77456), .ZN(n7507)
         );
  NAND4_X2 U8406 ( .A1(n7510), .A2(n7509), .A3(n7508), .A4(n7507), .ZN(n7515)
         );
  NAND2_X2 U8407 ( .A1(\REGFILE/reg_out[11][17] ), .A2(net77420), .ZN(n7513)
         );
  NAND2_X2 U8408 ( .A1(\REGFILE/reg_out[12][17] ), .A2(net77384), .ZN(n7512)
         );
  NAND2_X2 U8409 ( .A1(\REGFILE/reg_out[8][17] ), .A2(net77312), .ZN(n7511) );
  NAND4_X2 U8410 ( .A1(n7513), .A2(n7512), .A3(net74808), .A4(n7511), .ZN(
        n7514) );
  NAND2_X2 U8411 ( .A1(\REGFILE/reg_out[6][17] ), .A2(net77564), .ZN(n7519) );
  NAND2_X2 U8412 ( .A1(\REGFILE/reg_out[1][17] ), .A2(net77528), .ZN(n7518) );
  NAND2_X2 U8413 ( .A1(\REGFILE/reg_out[7][17] ), .A2(net77492), .ZN(n7517) );
  NAND2_X2 U8414 ( .A1(\REGFILE/reg_out[5][17] ), .A2(net77456), .ZN(n7516) );
  NAND4_X2 U8415 ( .A1(n7519), .A2(n7518), .A3(n7517), .A4(n7516), .ZN(n7524)
         );
  NAND2_X2 U8416 ( .A1(\REGFILE/reg_out[3][17] ), .A2(net77420), .ZN(n7522) );
  NAND2_X2 U8417 ( .A1(\REGFILE/reg_out[4][17] ), .A2(net77384), .ZN(n7521) );
  NAND4_X2 U8418 ( .A1(n7522), .A2(n7521), .A3(n7520), .A4(net74799), .ZN(
        n7523) );
  NAND4_X2 U8419 ( .A1(n7528), .A2(n7527), .A3(n7526), .A4(n7525), .ZN(n8447)
         );
  MUX2_X2 U8420 ( .A(n8447), .B(\PCLOGIC/imm16_32 [17]), .S(net77276), .Z(
        aluA[17]) );
  NAND2_X2 U8421 ( .A1(\REGFILE/reg_out[30][16] ), .A2(net77564), .ZN(n7532)
         );
  NAND2_X2 U8422 ( .A1(\REGFILE/reg_out[31][16] ), .A2(net77492), .ZN(n7530)
         );
  NAND2_X2 U8423 ( .A1(\REGFILE/reg_out[29][16] ), .A2(net77456), .ZN(n7529)
         );
  NAND4_X2 U8424 ( .A1(n7532), .A2(n7531), .A3(n7530), .A4(n7529), .ZN(n7538)
         );
  NAND2_X2 U8425 ( .A1(\REGFILE/reg_out[28][16] ), .A2(net77384), .ZN(n7535)
         );
  NAND2_X2 U8426 ( .A1(\REGFILE/reg_out[26][16] ), .A2(net77348), .ZN(n7534)
         );
  NAND2_X2 U8427 ( .A1(\REGFILE/reg_out[24][16] ), .A2(net77312), .ZN(n7533)
         );
  NAND4_X2 U8428 ( .A1(n7536), .A2(n7535), .A3(n7534), .A4(n7533), .ZN(n7537)
         );
  NAND2_X2 U8429 ( .A1(\REGFILE/reg_out[22][16] ), .A2(net77562), .ZN(n7542)
         );
  NAND2_X2 U8430 ( .A1(\REGFILE/reg_out[17][16] ), .A2(net77526), .ZN(n7541)
         );
  NAND2_X2 U8431 ( .A1(\REGFILE/reg_out[23][16] ), .A2(net77490), .ZN(n7540)
         );
  NAND2_X2 U8432 ( .A1(\REGFILE/reg_out[21][16] ), .A2(net77454), .ZN(n7539)
         );
  NAND4_X2 U8433 ( .A1(n7542), .A2(n7541), .A3(n7540), .A4(n7539), .ZN(n7548)
         );
  NAND2_X2 U8434 ( .A1(\REGFILE/reg_out[19][16] ), .A2(net77418), .ZN(n7546)
         );
  NAND2_X2 U8435 ( .A1(\REGFILE/reg_out[20][16] ), .A2(net77382), .ZN(n7545)
         );
  NAND2_X2 U8436 ( .A1(\REGFILE/reg_out[16][16] ), .A2(net77310), .ZN(n7543)
         );
  NAND4_X2 U8437 ( .A1(n7546), .A2(n7545), .A3(n7544), .A4(n7543), .ZN(n7547)
         );
  NAND2_X2 U8438 ( .A1(\REGFILE/reg_out[14][16] ), .A2(net77562), .ZN(n7552)
         );
  NAND2_X2 U8439 ( .A1(\REGFILE/reg_out[9][16] ), .A2(net77526), .ZN(n7551) );
  NAND2_X2 U8440 ( .A1(\REGFILE/reg_out[15][16] ), .A2(net77490), .ZN(n7550)
         );
  NAND2_X2 U8441 ( .A1(\REGFILE/reg_out[13][16] ), .A2(net77454), .ZN(n7549)
         );
  NAND4_X2 U8442 ( .A1(n7552), .A2(n7551), .A3(n7550), .A4(n7549), .ZN(n7558)
         );
  NAND2_X2 U8443 ( .A1(\REGFILE/reg_out[11][16] ), .A2(net77418), .ZN(n7556)
         );
  NAND2_X2 U8444 ( .A1(\REGFILE/reg_out[10][16] ), .A2(net77346), .ZN(n7554)
         );
  NAND2_X2 U8445 ( .A1(\REGFILE/reg_out[8][16] ), .A2(net77310), .ZN(n7553) );
  NAND4_X2 U8446 ( .A1(n7556), .A2(n7555), .A3(n7554), .A4(n7553), .ZN(n7557)
         );
  NAND2_X2 U8447 ( .A1(\REGFILE/reg_out[7][16] ), .A2(net77490), .ZN(n7560) );
  NAND2_X2 U8448 ( .A1(\REGFILE/reg_out[5][16] ), .A2(net77454), .ZN(n7559) );
  NAND4_X2 U8449 ( .A1(n7562), .A2(n7561), .A3(n7560), .A4(n7559), .ZN(n7568)
         );
  NAND2_X2 U8450 ( .A1(\REGFILE/reg_out[3][16] ), .A2(net77418), .ZN(n7566) );
  NAND2_X2 U8451 ( .A1(\REGFILE/reg_out[4][16] ), .A2(net77382), .ZN(n7565) );
  NAND2_X2 U8452 ( .A1(\REGFILE/reg_out[2][16] ), .A2(net77346), .ZN(n7564) );
  NAND2_X2 U8453 ( .A1(\REGFILE/reg_out[0][16] ), .A2(net77310), .ZN(n7563) );
  NAND4_X2 U8454 ( .A1(n7566), .A2(n7565), .A3(n7564), .A4(n7563), .ZN(n7567)
         );
  NAND4_X2 U8455 ( .A1(n7572), .A2(n7571), .A3(n7570), .A4(n7569), .ZN(n8445)
         );
  MUX2_X2 U8456 ( .A(n8445), .B(\PCLOGIC/imm16_32 [16]), .S(net77276), .Z(
        aluA[16]) );
  NAND2_X2 U8457 ( .A1(\REGFILE/reg_out[30][15] ), .A2(net77562), .ZN(n7576)
         );
  NAND2_X2 U8458 ( .A1(\REGFILE/reg_out[31][15] ), .A2(net77490), .ZN(n7574)
         );
  NAND2_X2 U8459 ( .A1(\REGFILE/reg_out[29][15] ), .A2(net77454), .ZN(n7573)
         );
  NAND4_X2 U8460 ( .A1(n7576), .A2(n7575), .A3(n7574), .A4(n7573), .ZN(n7582)
         );
  NAND2_X2 U8461 ( .A1(\REGFILE/reg_out[26][15] ), .A2(net77346), .ZN(n7578)
         );
  NAND2_X2 U8462 ( .A1(\REGFILE/reg_out[24][15] ), .A2(net77310), .ZN(n7577)
         );
  NAND4_X2 U8463 ( .A1(n7580), .A2(n7579), .A3(n7578), .A4(n7577), .ZN(n7581)
         );
  NAND2_X2 U8464 ( .A1(\REGFILE/reg_out[17][15] ), .A2(net77526), .ZN(n7585)
         );
  NAND2_X2 U8465 ( .A1(\REGFILE/reg_out[23][15] ), .A2(net77490), .ZN(n7584)
         );
  NAND2_X2 U8466 ( .A1(\REGFILE/reg_out[21][15] ), .A2(net77454), .ZN(n7583)
         );
  NAND4_X2 U8467 ( .A1(n7586), .A2(n7585), .A3(n7584), .A4(n7583), .ZN(n7592)
         );
  NAND2_X2 U8468 ( .A1(\REGFILE/reg_out[19][15] ), .A2(net77418), .ZN(n7590)
         );
  NAND2_X2 U8469 ( .A1(\REGFILE/reg_out[20][15] ), .A2(net77382), .ZN(n7589)
         );
  NAND4_X2 U8470 ( .A1(n7590), .A2(n7589), .A3(n7588), .A4(n7587), .ZN(n7591)
         );
  NAND2_X2 U8471 ( .A1(\REGFILE/reg_out[14][15] ), .A2(net77562), .ZN(n7596)
         );
  NAND2_X2 U8472 ( .A1(\REGFILE/reg_out[9][15] ), .A2(net77526), .ZN(n7595) );
  NAND2_X2 U8473 ( .A1(\REGFILE/reg_out[15][15] ), .A2(net77490), .ZN(n7594)
         );
  NAND4_X2 U8474 ( .A1(n7596), .A2(n7595), .A3(n7594), .A4(n7593), .ZN(n7602)
         );
  NAND2_X2 U8475 ( .A1(\REGFILE/reg_out[11][15] ), .A2(net77418), .ZN(n7600)
         );
  NAND2_X2 U8476 ( .A1(\REGFILE/reg_out[10][15] ), .A2(net77346), .ZN(n7598)
         );
  NAND2_X2 U8477 ( .A1(\REGFILE/reg_out[8][15] ), .A2(net77310), .ZN(n7597) );
  NAND4_X2 U8478 ( .A1(n7600), .A2(n7599), .A3(n7598), .A4(n7597), .ZN(n7601)
         );
  NAND2_X2 U8479 ( .A1(\REGFILE/reg_out[6][15] ), .A2(net77562), .ZN(n7606) );
  NAND2_X2 U8480 ( .A1(\REGFILE/reg_out[7][15] ), .A2(net77490), .ZN(n7604) );
  NAND4_X2 U8481 ( .A1(n7606), .A2(n7605), .A3(n7604), .A4(n7603), .ZN(n7612)
         );
  NAND2_X2 U8482 ( .A1(\REGFILE/reg_out[4][15] ), .A2(net77382), .ZN(n7609) );
  NAND2_X2 U8483 ( .A1(\REGFILE/reg_out[0][15] ), .A2(net77310), .ZN(n7607) );
  NAND4_X2 U8484 ( .A1(n7610), .A2(n7609), .A3(n7608), .A4(n7607), .ZN(n7611)
         );
  NAND4_X2 U8485 ( .A1(n7616), .A2(n7615), .A3(n7614), .A4(n7613), .ZN(n8446)
         );
  NAND2_X2 U8486 ( .A1(n8446), .A2(net77272), .ZN(n10463) );
  INV_X4 U8487 ( .A(n10463), .ZN(\WIRE_ALU_A/MUX2TO1_32BIT[15].MUX/N1 ) );
  NAND2_X2 U8488 ( .A1(\REGFILE/reg_out[30][14] ), .A2(net77562), .ZN(n7620)
         );
  NAND2_X2 U8489 ( .A1(\REGFILE/reg_out[31][14] ), .A2(net77490), .ZN(n7618)
         );
  NAND2_X2 U8490 ( .A1(\REGFILE/reg_out[29][14] ), .A2(net77454), .ZN(n7617)
         );
  NAND4_X2 U8491 ( .A1(n7620), .A2(n7619), .A3(n7618), .A4(n7617), .ZN(n7626)
         );
  NAND2_X2 U8492 ( .A1(net77346), .A2(\REGFILE/reg_out[26][14] ), .ZN(n7622)
         );
  NAND2_X2 U8493 ( .A1(\REGFILE/reg_out[24][14] ), .A2(net77310), .ZN(n7621)
         );
  NAND4_X2 U8494 ( .A1(n7624), .A2(n7623), .A3(n7622), .A4(n7621), .ZN(n7625)
         );
  NAND2_X2 U8495 ( .A1(\REGFILE/reg_out[22][14] ), .A2(net77562), .ZN(n7630)
         );
  NAND2_X2 U8496 ( .A1(\REGFILE/reg_out[17][14] ), .A2(net77526), .ZN(n7629)
         );
  NAND2_X2 U8497 ( .A1(\REGFILE/reg_out[23][14] ), .A2(net77490), .ZN(n7628)
         );
  NAND2_X2 U8498 ( .A1(\REGFILE/reg_out[21][14] ), .A2(net77454), .ZN(n7627)
         );
  NAND4_X2 U8499 ( .A1(n7630), .A2(n7629), .A3(n7628), .A4(n7627), .ZN(n7636)
         );
  NAND2_X2 U8500 ( .A1(\REGFILE/reg_out[19][14] ), .A2(net77418), .ZN(n7634)
         );
  NAND2_X2 U8501 ( .A1(\REGFILE/reg_out[16][14] ), .A2(net77310), .ZN(n7631)
         );
  NAND4_X2 U8502 ( .A1(n7634), .A2(n7633), .A3(n7632), .A4(n7631), .ZN(n7635)
         );
  NAND2_X2 U8503 ( .A1(\REGFILE/reg_out[14][14] ), .A2(net77562), .ZN(n7640)
         );
  NAND2_X2 U8504 ( .A1(\REGFILE/reg_out[9][14] ), .A2(net77526), .ZN(n7639) );
  NAND2_X2 U8505 ( .A1(\REGFILE/reg_out[15][14] ), .A2(net77490), .ZN(n7638)
         );
  NAND2_X2 U8506 ( .A1(\REGFILE/reg_out[13][14] ), .A2(net77454), .ZN(n7637)
         );
  NAND4_X2 U8507 ( .A1(n7640), .A2(n7639), .A3(n7638), .A4(n7637), .ZN(n7646)
         );
  NAND2_X2 U8508 ( .A1(net77418), .A2(n5777), .ZN(n7644) );
  NAND4_X2 U8509 ( .A1(n7644), .A2(n7643), .A3(n7642), .A4(n7641), .ZN(n7645)
         );
  NAND2_X2 U8510 ( .A1(\REGFILE/reg_out[6][14] ), .A2(net77562), .ZN(n7650) );
  NAND2_X2 U8511 ( .A1(\REGFILE/reg_out[1][14] ), .A2(net77526), .ZN(n7649) );
  NAND2_X2 U8512 ( .A1(\REGFILE/reg_out[7][14] ), .A2(net77490), .ZN(n7648) );
  NAND2_X2 U8513 ( .A1(n5832), .A2(net77454), .ZN(n7647) );
  NAND4_X2 U8514 ( .A1(n7650), .A2(n7649), .A3(n7648), .A4(n7647), .ZN(n7656)
         );
  NAND2_X2 U8515 ( .A1(\REGFILE/reg_out[4][14] ), .A2(net77382), .ZN(n7653) );
  NAND4_X2 U8516 ( .A1(n7654), .A2(n7653), .A3(n7652), .A4(n7651), .ZN(n7655)
         );
  NAND4_X2 U8517 ( .A1(n7660), .A2(n7659), .A3(n7658), .A4(n7657), .ZN(n8438)
         );
  NAND2_X2 U8518 ( .A1(n8438), .A2(net77272), .ZN(n10247) );
  INV_X4 U8519 ( .A(n10247), .ZN(\WIRE_ALU_A/MUX2TO1_32BIT[14].MUX/N1 ) );
  NAND2_X2 U8520 ( .A1(\REGFILE/reg_out[25][13] ), .A2(net77524), .ZN(n7663)
         );
  NAND2_X2 U8521 ( .A1(\REGFILE/reg_out[31][13] ), .A2(net77488), .ZN(n7662)
         );
  NAND2_X2 U8522 ( .A1(\REGFILE/reg_out[29][13] ), .A2(net77452), .ZN(n7661)
         );
  NAND4_X2 U8523 ( .A1(n7664), .A2(n7663), .A3(n7662), .A4(n7661), .ZN(n7670)
         );
  NAND2_X2 U8524 ( .A1(\REGFILE/reg_out[27][13] ), .A2(net77416), .ZN(n7668)
         );
  NAND4_X2 U8525 ( .A1(n7668), .A2(n7667), .A3(n7666), .A4(n7665), .ZN(n7669)
         );
  NAND2_X2 U8526 ( .A1(\REGFILE/reg_out[22][13] ), .A2(net77560), .ZN(n7674)
         );
  NAND2_X2 U8527 ( .A1(\REGFILE/reg_out[17][13] ), .A2(net77524), .ZN(n7673)
         );
  NAND2_X2 U8528 ( .A1(\REGFILE/reg_out[23][13] ), .A2(net77488), .ZN(n7672)
         );
  NAND2_X2 U8529 ( .A1(\REGFILE/reg_out[21][13] ), .A2(net77452), .ZN(n7671)
         );
  NAND4_X2 U8530 ( .A1(n7674), .A2(n7673), .A3(n7672), .A4(n7671), .ZN(n7680)
         );
  NAND2_X2 U8531 ( .A1(\REGFILE/reg_out[19][13] ), .A2(net77416), .ZN(n7678)
         );
  NAND2_X2 U8532 ( .A1(\REGFILE/reg_out[20][13] ), .A2(net77380), .ZN(n7677)
         );
  NAND4_X2 U8533 ( .A1(n7678), .A2(n7677), .A3(n7676), .A4(n7675), .ZN(n7679)
         );
  NAND2_X2 U8534 ( .A1(\REGFILE/reg_out[9][13] ), .A2(net77524), .ZN(n7683) );
  NAND2_X2 U8535 ( .A1(\REGFILE/reg_out[15][13] ), .A2(net77488), .ZN(n7682)
         );
  NAND2_X2 U8536 ( .A1(\REGFILE/reg_out[13][13] ), .A2(net77452), .ZN(n7681)
         );
  NAND4_X2 U8537 ( .A1(n7684), .A2(n7683), .A3(n7682), .A4(n7681), .ZN(n7690)
         );
  NAND2_X2 U8538 ( .A1(net148736), .A2(net77416), .ZN(n7688) );
  NAND4_X2 U8539 ( .A1(n7688), .A2(n7687), .A3(n7686), .A4(n7685), .ZN(n7689)
         );
  NAND2_X2 U8540 ( .A1(\REGFILE/reg_out[7][13] ), .A2(net77488), .ZN(n7692) );
  NAND2_X2 U8541 ( .A1(\REGFILE/reg_out[5][13] ), .A2(net77452), .ZN(n7691) );
  NAND4_X2 U8542 ( .A1(n7694), .A2(n7693), .A3(n7692), .A4(n7691), .ZN(n7700)
         );
  NAND2_X2 U8543 ( .A1(\REGFILE/reg_out[3][13] ), .A2(net77416), .ZN(n7698) );
  NAND2_X2 U8544 ( .A1(\REGFILE/reg_out[4][13] ), .A2(net77380), .ZN(n7697) );
  NAND2_X2 U8545 ( .A1(\REGFILE/reg_out[0][13] ), .A2(net77308), .ZN(n7695) );
  NAND4_X2 U8546 ( .A1(n7698), .A2(n7697), .A3(n7696), .A4(n7695), .ZN(n7699)
         );
  NAND4_X2 U8547 ( .A1(n7704), .A2(n7703), .A3(n7702), .A4(n7701), .ZN(n8437)
         );
  NAND2_X2 U8548 ( .A1(n8437), .A2(net77272), .ZN(n10368) );
  INV_X4 U8549 ( .A(n10368), .ZN(\WIRE_ALU_A/MUX2TO1_32BIT[13].MUX/N1 ) );
  NAND2_X2 U8550 ( .A1(\REGFILE/reg_out[30][12] ), .A2(net77560), .ZN(n7708)
         );
  NAND2_X2 U8551 ( .A1(\REGFILE/reg_out[25][12] ), .A2(net77524), .ZN(n7707)
         );
  NAND2_X2 U8552 ( .A1(\REGFILE/reg_out[31][12] ), .A2(net77488), .ZN(n7706)
         );
  NAND2_X2 U8553 ( .A1(\REGFILE/reg_out[29][12] ), .A2(net77452), .ZN(n7705)
         );
  NAND4_X2 U8554 ( .A1(n7708), .A2(n7707), .A3(n7706), .A4(n7705), .ZN(n7714)
         );
  NAND2_X2 U8555 ( .A1(\REGFILE/reg_out[27][12] ), .A2(net77416), .ZN(n7712)
         );
  NAND2_X2 U8556 ( .A1(\REGFILE/reg_out[26][12] ), .A2(net77344), .ZN(n7710)
         );
  NAND2_X2 U8557 ( .A1(\REGFILE/reg_out[24][12] ), .A2(net77308), .ZN(n7709)
         );
  NAND4_X2 U8558 ( .A1(n7712), .A2(n7711), .A3(n7710), .A4(n7709), .ZN(n7713)
         );
  NAND2_X2 U8559 ( .A1(\REGFILE/reg_out[22][12] ), .A2(net77560), .ZN(n7718)
         );
  NAND2_X2 U8560 ( .A1(\REGFILE/reg_out[17][12] ), .A2(net77524), .ZN(n7717)
         );
  NAND2_X2 U8561 ( .A1(\REGFILE/reg_out[23][12] ), .A2(net77488), .ZN(n7716)
         );
  NAND2_X2 U8562 ( .A1(\REGFILE/reg_out[21][12] ), .A2(net77452), .ZN(n7715)
         );
  NAND4_X2 U8563 ( .A1(n7718), .A2(n7717), .A3(n7716), .A4(n7715), .ZN(n7724)
         );
  NAND2_X2 U8564 ( .A1(\REGFILE/reg_out[19][12] ), .A2(net77416), .ZN(n7722)
         );
  NAND2_X2 U8565 ( .A1(\REGFILE/reg_out[20][12] ), .A2(net77380), .ZN(n7721)
         );
  NAND2_X2 U8566 ( .A1(\REGFILE/reg_out[18][12] ), .A2(net77344), .ZN(n7720)
         );
  NAND2_X2 U8567 ( .A1(\REGFILE/reg_out[16][12] ), .A2(net77308), .ZN(n7719)
         );
  NAND4_X2 U8568 ( .A1(n7722), .A2(n7721), .A3(n7720), .A4(n7719), .ZN(n7723)
         );
  NAND2_X2 U8569 ( .A1(\REGFILE/reg_out[14][12] ), .A2(net77560), .ZN(n7728)
         );
  NAND2_X2 U8570 ( .A1(\REGFILE/reg_out[9][12] ), .A2(net77524), .ZN(n7727) );
  NAND4_X2 U8571 ( .A1(n7728), .A2(n7727), .A3(n7726), .A4(n7725), .ZN(n7734)
         );
  NAND2_X2 U8572 ( .A1(\REGFILE/reg_out[11][12] ), .A2(net77416), .ZN(n7732)
         );
  NAND2_X2 U8573 ( .A1(\REGFILE/reg_out[10][12] ), .A2(net77344), .ZN(n7730)
         );
  NAND4_X2 U8575 ( .A1(n7732), .A2(n7731), .A3(n7730), .A4(n7729), .ZN(n7733)
         );
  NAND2_X2 U8576 ( .A1(\REGFILE/reg_out[6][12] ), .A2(net77560), .ZN(n7738) );
  NAND2_X2 U8577 ( .A1(\REGFILE/reg_out[1][12] ), .A2(net77524), .ZN(n7737) );
  NAND2_X2 U8578 ( .A1(\REGFILE/reg_out[7][12] ), .A2(net77488), .ZN(n7736) );
  NAND2_X2 U8579 ( .A1(\REGFILE/reg_out[5][12] ), .A2(net77452), .ZN(n7735) );
  NAND4_X2 U8580 ( .A1(n7738), .A2(n7737), .A3(n7736), .A4(n7735), .ZN(n7744)
         );
  NAND2_X2 U8582 ( .A1(\REGFILE/reg_out[4][12] ), .A2(net77380), .ZN(n7741) );
  NAND2_X2 U8583 ( .A1(\REGFILE/reg_out[2][12] ), .A2(net77344), .ZN(n7740) );
  NAND2_X2 U8584 ( .A1(\REGFILE/reg_out[0][12] ), .A2(net77308), .ZN(n7739) );
  NAND4_X2 U8585 ( .A1(n7742), .A2(n7741), .A3(n7740), .A4(n7739), .ZN(n7743)
         );
  NAND4_X2 U8586 ( .A1(n7748), .A2(n7747), .A3(n7746), .A4(n7745), .ZN(n8436)
         );
  NAND2_X2 U8587 ( .A1(n8436), .A2(net77272), .ZN(n9075) );
  INV_X4 U8588 ( .A(n9075), .ZN(\WIRE_ALU_A/MUX2TO1_32BIT[12].MUX/N1 ) );
  NAND2_X2 U8589 ( .A1(\REGFILE/reg_out[30][11] ), .A2(net77560), .ZN(n7752)
         );
  NAND2_X2 U8590 ( .A1(\REGFILE/reg_out[25][11] ), .A2(net77524), .ZN(n7751)
         );
  NAND2_X2 U8591 ( .A1(\REGFILE/reg_out[31][11] ), .A2(net77488), .ZN(n7750)
         );
  NAND2_X2 U8592 ( .A1(\REGFILE/reg_out[29][11] ), .A2(net77452), .ZN(n7749)
         );
  NAND4_X2 U8593 ( .A1(n7752), .A2(n7751), .A3(n7750), .A4(n7749), .ZN(n7758)
         );
  NAND2_X2 U8594 ( .A1(\REGFILE/reg_out[26][11] ), .A2(net77344), .ZN(n7754)
         );
  NAND2_X2 U8595 ( .A1(\REGFILE/reg_out[24][11] ), .A2(net77308), .ZN(n7753)
         );
  NAND4_X2 U8596 ( .A1(n7756), .A2(n7755), .A3(n7754), .A4(n7753), .ZN(n7757)
         );
  NAND2_X2 U8597 ( .A1(\REGFILE/reg_out[22][11] ), .A2(net77560), .ZN(n7762)
         );
  NAND2_X2 U8598 ( .A1(\REGFILE/reg_out[17][11] ), .A2(net77524), .ZN(n7761)
         );
  NAND2_X2 U8599 ( .A1(\REGFILE/reg_out[23][11] ), .A2(net77488), .ZN(n7760)
         );
  NAND2_X2 U8600 ( .A1(\REGFILE/reg_out[21][11] ), .A2(net77452), .ZN(n7759)
         );
  NAND4_X2 U8601 ( .A1(n7762), .A2(n7761), .A3(n7760), .A4(n7759), .ZN(n7768)
         );
  NAND2_X2 U8602 ( .A1(\REGFILE/reg_out[19][11] ), .A2(net77416), .ZN(n7766)
         );
  NAND2_X2 U8603 ( .A1(\REGFILE/reg_out[20][11] ), .A2(net77380), .ZN(n7765)
         );
  NAND2_X2 U8604 ( .A1(\REGFILE/reg_out[18][11] ), .A2(net77344), .ZN(n7764)
         );
  NAND2_X2 U8605 ( .A1(\REGFILE/reg_out[16][11] ), .A2(net77308), .ZN(n7763)
         );
  NAND4_X2 U8606 ( .A1(n7766), .A2(n7765), .A3(n7764), .A4(n7763), .ZN(n7767)
         );
  NAND2_X2 U8607 ( .A1(\REGFILE/reg_out[14][11] ), .A2(net77560), .ZN(n7772)
         );
  NAND2_X2 U8608 ( .A1(\REGFILE/reg_out[9][11] ), .A2(net77524), .ZN(n7771) );
  NAND2_X2 U8609 ( .A1(\REGFILE/reg_out[15][11] ), .A2(net77488), .ZN(n7770)
         );
  NAND4_X2 U8610 ( .A1(n7772), .A2(n7771), .A3(n7770), .A4(n7769), .ZN(n7778)
         );
  NAND2_X2 U8611 ( .A1(\REGFILE/reg_out[11][11] ), .A2(net77416), .ZN(n7776)
         );
  NAND2_X2 U8612 ( .A1(n5907), .A2(net77344), .ZN(n7774) );
  NAND2_X2 U8613 ( .A1(\REGFILE/reg_out[8][11] ), .A2(net77308), .ZN(n7773) );
  NAND4_X2 U8614 ( .A1(n7776), .A2(n7775), .A3(n7774), .A4(n7773), .ZN(n7777)
         );
  NAND2_X2 U8615 ( .A1(\REGFILE/reg_out[6][11] ), .A2(net77560), .ZN(n7782) );
  NAND2_X2 U8616 ( .A1(\REGFILE/reg_out[1][11] ), .A2(net77524), .ZN(n7781) );
  NAND2_X2 U8617 ( .A1(\REGFILE/reg_out[7][11] ), .A2(net77488), .ZN(n7780) );
  NAND2_X2 U8618 ( .A1(\REGFILE/reg_out[5][11] ), .A2(net77452), .ZN(n7779) );
  NAND4_X2 U8619 ( .A1(n7782), .A2(n7781), .A3(n7780), .A4(n7779), .ZN(n7788)
         );
  NAND2_X2 U8620 ( .A1(\REGFILE/reg_out[3][11] ), .A2(net77416), .ZN(n7786) );
  NAND2_X2 U8621 ( .A1(\REGFILE/reg_out[4][11] ), .A2(net77380), .ZN(n7785) );
  NAND2_X2 U8622 ( .A1(net77344), .A2(\REGFILE/reg_out[2][11] ), .ZN(n7784) );
  NAND2_X2 U8623 ( .A1(\REGFILE/reg_out[0][11] ), .A2(net77308), .ZN(n7783) );
  NAND4_X2 U8624 ( .A1(n7786), .A2(n7785), .A3(n7784), .A4(n7783), .ZN(n7787)
         );
  NAND4_X2 U8625 ( .A1(n7792), .A2(n7791), .A3(n7790), .A4(n7789), .ZN(n8435)
         );
  NAND2_X2 U8626 ( .A1(n8435), .A2(net77272), .ZN(n10375) );
  INV_X4 U8627 ( .A(n10375), .ZN(\WIRE_ALU_A/MUX2TO1_32BIT[11].MUX/N1 ) );
  NAND2_X2 U8628 ( .A1(\REGFILE/reg_out[30][10] ), .A2(net77558), .ZN(n7796)
         );
  NAND2_X2 U8629 ( .A1(\REGFILE/reg_out[31][10] ), .A2(net77482), .ZN(n7794)
         );
  NAND2_X2 U8630 ( .A1(\REGFILE/reg_out[29][10] ), .A2(net77456), .ZN(n7793)
         );
  NAND4_X2 U8631 ( .A1(n7796), .A2(n7795), .A3(n7794), .A4(n7793), .ZN(n7802)
         );
  NAND2_X2 U8632 ( .A1(\REGFILE/reg_out[27][10] ), .A2(net77414), .ZN(n7800)
         );
  NAND2_X2 U8633 ( .A1(\REGFILE/reg_out[28][10] ), .A2(net77376), .ZN(n7799)
         );
  NAND2_X2 U8634 ( .A1(\REGFILE/reg_out[26][10] ), .A2(net77342), .ZN(n7798)
         );
  NAND2_X2 U8635 ( .A1(\REGFILE/reg_out[24][10] ), .A2(net77306), .ZN(n7797)
         );
  NAND4_X2 U8636 ( .A1(n7800), .A2(n7799), .A3(n7798), .A4(n7797), .ZN(n7801)
         );
  NAND2_X2 U8637 ( .A1(\REGFILE/reg_out[22][10] ), .A2(net77558), .ZN(n7806)
         );
  NAND2_X2 U8638 ( .A1(\REGFILE/reg_out[17][10] ), .A2(net77522), .ZN(n7805)
         );
  NAND2_X2 U8639 ( .A1(\REGFILE/reg_out[23][10] ), .A2(net77482), .ZN(n7804)
         );
  NAND2_X2 U8640 ( .A1(\REGFILE/reg_out[21][10] ), .A2(net77456), .ZN(n7803)
         );
  NAND4_X2 U8641 ( .A1(n7806), .A2(n7805), .A3(n7804), .A4(n7803), .ZN(n7812)
         );
  NAND2_X2 U8642 ( .A1(\REGFILE/reg_out[19][10] ), .A2(net77414), .ZN(n7810)
         );
  NAND2_X2 U8643 ( .A1(\REGFILE/reg_out[20][10] ), .A2(net77376), .ZN(n7809)
         );
  NAND2_X2 U8644 ( .A1(\REGFILE/reg_out[18][10] ), .A2(net77342), .ZN(n7808)
         );
  NAND2_X2 U8645 ( .A1(\REGFILE/reg_out[16][10] ), .A2(net77306), .ZN(n7807)
         );
  NAND4_X2 U8646 ( .A1(n7810), .A2(n7809), .A3(n7808), .A4(n7807), .ZN(n7811)
         );
  NAND2_X2 U8647 ( .A1(\REGFILE/reg_out[14][10] ), .A2(net77558), .ZN(n7816)
         );
  NAND2_X2 U8648 ( .A1(\REGFILE/reg_out[9][10] ), .A2(net77522), .ZN(n7815) );
  NAND4_X2 U8649 ( .A1(n7816), .A2(n7815), .A3(n7814), .A4(n7813), .ZN(n7822)
         );
  NAND2_X2 U8650 ( .A1(\REGFILE/reg_out[11][10] ), .A2(net77414), .ZN(n7820)
         );
  NAND2_X2 U8651 ( .A1(\REGFILE/reg_out[10][10] ), .A2(net77342), .ZN(n7818)
         );
  NAND2_X2 U8652 ( .A1(\REGFILE/reg_out[8][10] ), .A2(net77306), .ZN(n7817) );
  NAND4_X2 U8653 ( .A1(n7820), .A2(n7819), .A3(n7818), .A4(n7817), .ZN(n7821)
         );
  NAND2_X2 U8654 ( .A1(\REGFILE/reg_out[6][10] ), .A2(net77558), .ZN(n7826) );
  NAND2_X2 U8655 ( .A1(\REGFILE/reg_out[1][10] ), .A2(net77522), .ZN(n7825) );
  NAND2_X2 U8656 ( .A1(\REGFILE/reg_out[7][10] ), .A2(net77482), .ZN(n7824) );
  NAND2_X2 U8657 ( .A1(\REGFILE/reg_out[5][10] ), .A2(net77456), .ZN(n7823) );
  NAND4_X2 U8658 ( .A1(n7826), .A2(n7825), .A3(n7824), .A4(n7823), .ZN(n7832)
         );
  NAND2_X2 U8659 ( .A1(\REGFILE/reg_out[4][10] ), .A2(net77376), .ZN(n7829) );
  NAND2_X2 U8660 ( .A1(\REGFILE/reg_out[0][10] ), .A2(net77306), .ZN(n7827) );
  NAND4_X2 U8661 ( .A1(n7830), .A2(n7829), .A3(n7828), .A4(n7827), .ZN(n7831)
         );
  NAND4_X2 U8662 ( .A1(n7836), .A2(n7835), .A3(n7834), .A4(n7833), .ZN(n8434)
         );
  NAND2_X2 U8663 ( .A1(n8434), .A2(net77272), .ZN(n10125) );
  INV_X4 U8664 ( .A(n10125), .ZN(\WIRE_ALU_A/MUX2TO1_32BIT[10].MUX/N1 ) );
  NAND2_X2 U8665 ( .A1(\REGFILE/reg_out[30][9] ), .A2(net77558), .ZN(n7840) );
  NAND2_X2 U8666 ( .A1(\REGFILE/reg_out[31][9] ), .A2(net77482), .ZN(n7838) );
  NAND2_X2 U8667 ( .A1(\REGFILE/reg_out[29][9] ), .A2(net77456), .ZN(n7837) );
  NAND4_X2 U8668 ( .A1(n7840), .A2(n7839), .A3(n7838), .A4(n7837), .ZN(n7846)
         );
  NAND2_X2 U8669 ( .A1(\REGFILE/reg_out[27][9] ), .A2(net77414), .ZN(n7844) );
  NAND2_X2 U8670 ( .A1(\REGFILE/reg_out[28][9] ), .A2(net77376), .ZN(n7843) );
  NAND2_X2 U8671 ( .A1(\REGFILE/reg_out[26][9] ), .A2(net77342), .ZN(n7842) );
  NAND2_X2 U8672 ( .A1(\REGFILE/reg_out[24][9] ), .A2(net77306), .ZN(n7841) );
  NAND4_X2 U8673 ( .A1(n7844), .A2(n7843), .A3(n7842), .A4(n7841), .ZN(n7845)
         );
  NAND2_X2 U8674 ( .A1(\REGFILE/reg_out[22][9] ), .A2(net77558), .ZN(n7850) );
  NAND2_X2 U8675 ( .A1(\REGFILE/reg_out[17][9] ), .A2(net77522), .ZN(n7849) );
  NAND2_X2 U8676 ( .A1(\REGFILE/reg_out[23][9] ), .A2(net77482), .ZN(n7848) );
  NAND2_X2 U8677 ( .A1(\REGFILE/reg_out[21][9] ), .A2(net77456), .ZN(n7847) );
  NAND4_X2 U8678 ( .A1(n7850), .A2(n7849), .A3(n7848), .A4(n7847), .ZN(n7856)
         );
  NAND2_X2 U8679 ( .A1(\REGFILE/reg_out[19][9] ), .A2(net77414), .ZN(n7854) );
  NAND2_X2 U8680 ( .A1(\REGFILE/reg_out[20][9] ), .A2(net77376), .ZN(n7853) );
  NAND2_X2 U8681 ( .A1(\REGFILE/reg_out[18][9] ), .A2(net77342), .ZN(n7852) );
  NAND2_X2 U8682 ( .A1(\REGFILE/reg_out[16][9] ), .A2(net77306), .ZN(n7851) );
  NAND4_X2 U8683 ( .A1(n7854), .A2(n7853), .A3(n7852), .A4(n7851), .ZN(n7855)
         );
  NAND2_X2 U8684 ( .A1(\REGFILE/reg_out[14][9] ), .A2(net77558), .ZN(n7860) );
  NAND2_X2 U8685 ( .A1(\REGFILE/reg_out[9][9] ), .A2(net77522), .ZN(n7859) );
  NAND2_X2 U8686 ( .A1(\REGFILE/reg_out[15][9] ), .A2(net77482), .ZN(n7858) );
  NAND2_X2 U8687 ( .A1(\REGFILE/reg_out[13][9] ), .A2(net77456), .ZN(n7857) );
  NAND4_X2 U8688 ( .A1(n7860), .A2(n7859), .A3(n7858), .A4(n7857), .ZN(n7866)
         );
  NAND2_X2 U8689 ( .A1(\REGFILE/reg_out[11][9] ), .A2(net77414), .ZN(n7864) );
  NAND2_X2 U8690 ( .A1(net77376), .A2(\REGFILE/reg_out[12][9] ), .ZN(n7863) );
  NAND2_X2 U8691 ( .A1(\REGFILE/reg_out[10][9] ), .A2(net77342), .ZN(n7862) );
  NAND2_X2 U8692 ( .A1(\REGFILE/reg_out[8][9] ), .A2(net77306), .ZN(n7861) );
  NAND4_X2 U8693 ( .A1(n7864), .A2(n7863), .A3(n7862), .A4(n7861), .ZN(n7865)
         );
  NAND2_X2 U8694 ( .A1(\REGFILE/reg_out[6][9] ), .A2(net77558), .ZN(n7870) );
  NAND2_X2 U8695 ( .A1(\REGFILE/reg_out[1][9] ), .A2(net77522), .ZN(n7869) );
  NAND2_X2 U8696 ( .A1(\REGFILE/reg_out[7][9] ), .A2(net77482), .ZN(n7868) );
  NAND2_X2 U8697 ( .A1(\REGFILE/reg_out[5][9] ), .A2(net77456), .ZN(n7867) );
  NAND4_X2 U8698 ( .A1(n7870), .A2(n7869), .A3(n7868), .A4(n7867), .ZN(n7876)
         );
  NAND2_X2 U8699 ( .A1(\REGFILE/reg_out[3][9] ), .A2(net77414), .ZN(n7874) );
  NAND2_X2 U8700 ( .A1(\REGFILE/reg_out[4][9] ), .A2(net77376), .ZN(n7873) );
  NAND2_X2 U8701 ( .A1(\REGFILE/reg_out[0][9] ), .A2(net77306), .ZN(n7871) );
  NAND4_X2 U8702 ( .A1(n7874), .A2(n7873), .A3(n7872), .A4(n7871), .ZN(n7875)
         );
  NAND4_X2 U8703 ( .A1(n7880), .A2(n7879), .A3(n7878), .A4(n7877), .ZN(n8430)
         );
  NAND2_X2 U8704 ( .A1(n8430), .A2(net77272), .ZN(n10382) );
  INV_X4 U8705 ( .A(n10382), .ZN(\WIRE_ALU_A/MUX2TO1_32BIT[9].MUX/N1 ) );
  NAND2_X2 U8706 ( .A1(\REGFILE/reg_out[30][8] ), .A2(net77558), .ZN(n7884) );
  NAND2_X2 U8707 ( .A1(\REGFILE/reg_out[31][8] ), .A2(net77482), .ZN(n7882) );
  NAND2_X2 U8708 ( .A1(\REGFILE/reg_out[29][8] ), .A2(net77456), .ZN(n7881) );
  NAND4_X2 U8709 ( .A1(n7884), .A2(n7883), .A3(n7882), .A4(n7881), .ZN(n7890)
         );
  NAND2_X2 U8710 ( .A1(\REGFILE/reg_out[28][8] ), .A2(net77376), .ZN(n7887) );
  NAND2_X2 U8711 ( .A1(\REGFILE/reg_out[26][8] ), .A2(net77342), .ZN(n7886) );
  NAND2_X2 U8712 ( .A1(\REGFILE/reg_out[24][8] ), .A2(net77306), .ZN(n7885) );
  NAND4_X2 U8713 ( .A1(n7888), .A2(n7887), .A3(n7886), .A4(n7885), .ZN(n7889)
         );
  NAND2_X2 U8714 ( .A1(\REGFILE/reg_out[22][8] ), .A2(net77558), .ZN(n7894) );
  NAND2_X2 U8715 ( .A1(\REGFILE/reg_out[17][8] ), .A2(net77522), .ZN(n7893) );
  NAND2_X2 U8716 ( .A1(\REGFILE/reg_out[23][8] ), .A2(net77482), .ZN(n7892) );
  NAND2_X2 U8717 ( .A1(\REGFILE/reg_out[21][8] ), .A2(net77456), .ZN(n7891) );
  NAND4_X2 U8718 ( .A1(n7894), .A2(n7893), .A3(n7892), .A4(n7891), .ZN(n7900)
         );
  NAND2_X2 U8719 ( .A1(\REGFILE/reg_out[19][8] ), .A2(net77414), .ZN(n7898) );
  NAND2_X2 U8720 ( .A1(\REGFILE/reg_out[20][8] ), .A2(net77376), .ZN(n7897) );
  NAND2_X2 U8721 ( .A1(\REGFILE/reg_out[18][8] ), .A2(net77342), .ZN(n7896) );
  NAND2_X2 U8722 ( .A1(\REGFILE/reg_out[16][8] ), .A2(net77306), .ZN(n7895) );
  NAND4_X2 U8723 ( .A1(n7898), .A2(n7897), .A3(n7896), .A4(n7895), .ZN(n7899)
         );
  NAND2_X2 U8724 ( .A1(\REGFILE/reg_out[14][8] ), .A2(net77558), .ZN(n7904) );
  NAND2_X2 U8725 ( .A1(\REGFILE/reg_out[9][8] ), .A2(net77522), .ZN(n7903) );
  NAND2_X2 U8726 ( .A1(\REGFILE/reg_out[15][8] ), .A2(net77482), .ZN(n7902) );
  NAND2_X2 U8727 ( .A1(\REGFILE/reg_out[13][8] ), .A2(net77456), .ZN(n7901) );
  NAND4_X2 U8728 ( .A1(n7904), .A2(n7903), .A3(n7902), .A4(n7901), .ZN(n7910)
         );
  NAND2_X2 U8729 ( .A1(\REGFILE/reg_out[11][8] ), .A2(net77414), .ZN(n7908) );
  NAND2_X2 U8730 ( .A1(\REGFILE/reg_out[12][8] ), .A2(net77376), .ZN(n7907) );
  NAND2_X2 U8731 ( .A1(\REGFILE/reg_out[10][8] ), .A2(net77342), .ZN(n7906) );
  NAND2_X2 U8732 ( .A1(\REGFILE/reg_out[8][8] ), .A2(net77306), .ZN(n7905) );
  NAND4_X2 U8733 ( .A1(n7908), .A2(n7907), .A3(n7906), .A4(n7905), .ZN(n7909)
         );
  NAND2_X2 U8734 ( .A1(\REGFILE/reg_out[6][8] ), .A2(net77558), .ZN(n7914) );
  NAND2_X2 U8735 ( .A1(\REGFILE/reg_out[1][8] ), .A2(net77522), .ZN(n7913) );
  NAND2_X2 U8736 ( .A1(\REGFILE/reg_out[7][8] ), .A2(net77482), .ZN(n7912) );
  NAND2_X2 U8737 ( .A1(\REGFILE/reg_out[5][8] ), .A2(net77456), .ZN(n7911) );
  NAND4_X2 U8738 ( .A1(n7914), .A2(n7913), .A3(n7912), .A4(n7911), .ZN(n7920)
         );
  NAND2_X2 U8739 ( .A1(\REGFILE/reg_out[4][8] ), .A2(net77376), .ZN(n7917) );
  NAND2_X2 U8740 ( .A1(\REGFILE/reg_out[0][8] ), .A2(net77306), .ZN(n7915) );
  NAND4_X2 U8741 ( .A1(n7918), .A2(n7917), .A3(n7916), .A4(n7915), .ZN(n7919)
         );
  NAND4_X2 U8742 ( .A1(n7924), .A2(n7923), .A3(n7922), .A4(n7921), .ZN(n8431)
         );
  NAND2_X2 U8743 ( .A1(n8431), .A2(net77272), .ZN(n9535) );
  INV_X4 U8744 ( .A(n9535), .ZN(\WIRE_ALU_A/MUX2TO1_32BIT[8].MUX/N1 ) );
  NAND2_X2 U8745 ( .A1(\REGFILE/reg_out[30][7] ), .A2(net77556), .ZN(n7928) );
  NAND2_X2 U8746 ( .A1(\REGFILE/reg_out[31][7] ), .A2(net77484), .ZN(n7926) );
  NAND2_X2 U8747 ( .A1(\REGFILE/reg_out[29][7] ), .A2(net77456), .ZN(n7925) );
  NAND4_X2 U8748 ( .A1(n7928), .A2(n7927), .A3(n7926), .A4(n7925), .ZN(n7934)
         );
  NAND2_X2 U8749 ( .A1(\REGFILE/reg_out[28][7] ), .A2(net77376), .ZN(n7931) );
  NAND2_X2 U8750 ( .A1(\REGFILE/reg_out[26][7] ), .A2(net77338), .ZN(n7930) );
  NAND2_X2 U8751 ( .A1(\REGFILE/reg_out[24][7] ), .A2(net77304), .ZN(n7929) );
  NAND4_X2 U8752 ( .A1(n7932), .A2(n7931), .A3(n7930), .A4(n7929), .ZN(n7933)
         );
  NAND2_X2 U8753 ( .A1(\REGFILE/reg_out[22][7] ), .A2(net77556), .ZN(n7938) );
  NAND2_X2 U8754 ( .A1(\REGFILE/reg_out[17][7] ), .A2(net77520), .ZN(n7937) );
  NAND2_X2 U8755 ( .A1(\REGFILE/reg_out[23][7] ), .A2(net77484), .ZN(n7936) );
  NAND2_X2 U8756 ( .A1(\REGFILE/reg_out[21][7] ), .A2(net77456), .ZN(n7935) );
  NAND4_X2 U8757 ( .A1(n7938), .A2(n7937), .A3(n7936), .A4(n7935), .ZN(n7944)
         );
  NAND2_X2 U8758 ( .A1(\REGFILE/reg_out[19][7] ), .A2(net77410), .ZN(n7942) );
  NAND2_X2 U8759 ( .A1(\REGFILE/reg_out[20][7] ), .A2(net77376), .ZN(n7941) );
  NAND2_X2 U8760 ( .A1(\REGFILE/reg_out[18][7] ), .A2(net77338), .ZN(n7940) );
  NAND2_X2 U8761 ( .A1(\REGFILE/reg_out[16][7] ), .A2(net77304), .ZN(n7939) );
  NAND4_X2 U8762 ( .A1(n7942), .A2(n7941), .A3(n7940), .A4(n7939), .ZN(n7943)
         );
  NAND2_X2 U8763 ( .A1(\REGFILE/reg_out[14][7] ), .A2(net77556), .ZN(n7948) );
  NAND2_X2 U8764 ( .A1(\REGFILE/reg_out[9][7] ), .A2(net77520), .ZN(n7947) );
  NAND2_X2 U8765 ( .A1(\REGFILE/reg_out[15][7] ), .A2(net77484), .ZN(n7946) );
  NAND2_X2 U8766 ( .A1(\REGFILE/reg_out[13][7] ), .A2(net77456), .ZN(n7945) );
  NAND4_X2 U8767 ( .A1(n7948), .A2(n7947), .A3(n7946), .A4(n7945), .ZN(n7954)
         );
  NAND2_X2 U8768 ( .A1(\REGFILE/reg_out[11][7] ), .A2(net77410), .ZN(n7952) );
  NAND2_X2 U8769 ( .A1(\REGFILE/reg_out[12][7] ), .A2(net77376), .ZN(n7951) );
  NAND2_X2 U8770 ( .A1(\REGFILE/reg_out[8][7] ), .A2(net77304), .ZN(n7949) );
  NAND4_X2 U8771 ( .A1(n7952), .A2(n7951), .A3(n7950), .A4(n7949), .ZN(n7953)
         );
  NAND2_X2 U8772 ( .A1(\REGFILE/reg_out[1][7] ), .A2(net77520), .ZN(n7956) );
  NAND2_X2 U8773 ( .A1(\REGFILE/reg_out[5][7] ), .A2(net77456), .ZN(n7955) );
  NAND4_X2 U8774 ( .A1(net74359), .A2(n7956), .A3(net74361), .A4(n7955), .ZN(
        n7962) );
  NAND2_X2 U8775 ( .A1(\REGFILE/reg_out[3][7] ), .A2(net77410), .ZN(n7960) );
  NAND2_X2 U8776 ( .A1(\REGFILE/reg_out[4][7] ), .A2(net77376), .ZN(n7959) );
  NAND2_X2 U8777 ( .A1(\REGFILE/reg_out[0][7] ), .A2(net77304), .ZN(n7957) );
  NAND4_X2 U8778 ( .A1(n7960), .A2(n7959), .A3(n7958), .A4(n7957), .ZN(n7961)
         );
  NAND4_X2 U8779 ( .A1(n7966), .A2(n7965), .A3(n7964), .A4(n7963), .ZN(n8432)
         );
  NAND2_X2 U8780 ( .A1(n8432), .A2(net77272), .ZN(n10464) );
  INV_X4 U8781 ( .A(n10464), .ZN(\WIRE_ALU_A/MUX2TO1_32BIT[7].MUX/N1 ) );
  NAND2_X2 U8782 ( .A1(\REGFILE/reg_out[30][6] ), .A2(net77556), .ZN(n7970) );
  NAND2_X2 U8783 ( .A1(n5764), .A2(net77520), .ZN(n7969) );
  NAND2_X2 U8784 ( .A1(\REGFILE/reg_out[31][6] ), .A2(net77484), .ZN(n7968) );
  NAND2_X2 U8785 ( .A1(\REGFILE/reg_out[29][6] ), .A2(net77456), .ZN(n7967) );
  NAND4_X2 U8786 ( .A1(n7970), .A2(n7969), .A3(n7968), .A4(n7967), .ZN(n7976)
         );
  NAND2_X2 U8787 ( .A1(\REGFILE/reg_out[27][6] ), .A2(net77410), .ZN(n7974) );
  NAND2_X2 U8788 ( .A1(\REGFILE/reg_out[28][6] ), .A2(net77376), .ZN(n7973) );
  NAND2_X2 U8789 ( .A1(\REGFILE/reg_out[26][6] ), .A2(net77338), .ZN(n7972) );
  NAND2_X2 U8790 ( .A1(\REGFILE/reg_out[24][6] ), .A2(net77304), .ZN(n7971) );
  NAND4_X2 U8791 ( .A1(n7974), .A2(n7973), .A3(n7972), .A4(n7971), .ZN(n7975)
         );
  NAND2_X2 U8792 ( .A1(\REGFILE/reg_out[22][6] ), .A2(net77556), .ZN(n7980) );
  NAND2_X2 U8793 ( .A1(\REGFILE/reg_out[17][6] ), .A2(net77520), .ZN(n7979) );
  NAND2_X2 U8794 ( .A1(\REGFILE/reg_out[23][6] ), .A2(net77484), .ZN(n7978) );
  NAND2_X2 U8795 ( .A1(\REGFILE/reg_out[21][6] ), .A2(net77456), .ZN(n7977) );
  NAND4_X2 U8796 ( .A1(n7980), .A2(n7979), .A3(n7978), .A4(n7977), .ZN(n7986)
         );
  NAND2_X2 U8797 ( .A1(\REGFILE/reg_out[19][6] ), .A2(net77410), .ZN(n7984) );
  NAND2_X2 U8798 ( .A1(\REGFILE/reg_out[20][6] ), .A2(net77376), .ZN(n7983) );
  NAND2_X2 U8799 ( .A1(\REGFILE/reg_out[18][6] ), .A2(net77338), .ZN(n7982) );
  NAND2_X2 U8800 ( .A1(\REGFILE/reg_out[16][6] ), .A2(net77304), .ZN(n7981) );
  NAND4_X2 U8801 ( .A1(n7984), .A2(n7983), .A3(n7982), .A4(n7981), .ZN(n7985)
         );
  NAND2_X2 U8802 ( .A1(\REGFILE/reg_out[14][6] ), .A2(net77556), .ZN(n7990) );
  NAND2_X2 U8803 ( .A1(\REGFILE/reg_out[9][6] ), .A2(net77520), .ZN(n7989) );
  NAND2_X2 U8804 ( .A1(\REGFILE/reg_out[13][6] ), .A2(net77456), .ZN(n7987) );
  NAND4_X2 U8805 ( .A1(n7990), .A2(n7989), .A3(n7988), .A4(n7987), .ZN(n7996)
         );
  NAND2_X2 U8806 ( .A1(\REGFILE/reg_out[11][6] ), .A2(net77410), .ZN(n7994) );
  NAND2_X2 U8807 ( .A1(\REGFILE/reg_out[12][6] ), .A2(net77376), .ZN(n7993) );
  NAND2_X2 U8808 ( .A1(n5902), .A2(net77338), .ZN(n7992) );
  NAND2_X2 U8809 ( .A1(\REGFILE/reg_out[8][6] ), .A2(net77304), .ZN(n7991) );
  NAND4_X2 U8810 ( .A1(n7994), .A2(n7993), .A3(n7992), .A4(n7991), .ZN(n7995)
         );
  NAND2_X2 U8811 ( .A1(\REGFILE/reg_out[6][6] ), .A2(net77556), .ZN(n8000) );
  NAND2_X2 U8812 ( .A1(\REGFILE/reg_out[1][6] ), .A2(net77520), .ZN(n7999) );
  NAND2_X2 U8813 ( .A1(\REGFILE/reg_out[7][6] ), .A2(net77484), .ZN(n7998) );
  NAND2_X2 U8814 ( .A1(\REGFILE/reg_out[5][6] ), .A2(net77456), .ZN(n7997) );
  NAND4_X2 U8815 ( .A1(n8000), .A2(n7999), .A3(n7998), .A4(n7997), .ZN(n8006)
         );
  NAND2_X2 U8816 ( .A1(\REGFILE/reg_out[3][6] ), .A2(net77410), .ZN(n8004) );
  NAND2_X2 U8817 ( .A1(\REGFILE/reg_out[4][6] ), .A2(net77376), .ZN(n8003) );
  NAND2_X2 U8818 ( .A1(\REGFILE/reg_out[2][6] ), .A2(net77338), .ZN(n8002) );
  NAND2_X2 U8819 ( .A1(\REGFILE/reg_out[0][6] ), .A2(net77304), .ZN(n8001) );
  NAND4_X2 U8820 ( .A1(n8004), .A2(n8003), .A3(n8002), .A4(n8001), .ZN(n8005)
         );
  NAND4_X2 U8821 ( .A1(n8010), .A2(n8009), .A3(n8008), .A4(n8007), .ZN(n8433)
         );
  NAND2_X2 U8822 ( .A1(n8433), .A2(net77272), .ZN(n9656) );
  INV_X4 U8823 ( .A(n9656), .ZN(\WIRE_ALU_A/MUX2TO1_32BIT[6].MUX/N1 ) );
  NAND2_X2 U8824 ( .A1(\REGFILE/reg_out[30][5] ), .A2(net77556), .ZN(n8014) );
  NAND2_X2 U8825 ( .A1(\REGFILE/reg_out[25][5] ), .A2(net77520), .ZN(n8013) );
  NAND2_X2 U8826 ( .A1(\REGFILE/reg_out[31][5] ), .A2(net77484), .ZN(n8012) );
  NAND2_X2 U8827 ( .A1(\REGFILE/reg_out[29][5] ), .A2(net77456), .ZN(n8011) );
  NAND4_X2 U8828 ( .A1(n8014), .A2(n8013), .A3(n8012), .A4(n8011), .ZN(n8020)
         );
  NAND2_X2 U8829 ( .A1(\REGFILE/reg_out[27][5] ), .A2(net77410), .ZN(n8018) );
  NAND2_X2 U8830 ( .A1(\REGFILE/reg_out[28][5] ), .A2(net77376), .ZN(n8017) );
  NAND2_X2 U8831 ( .A1(\REGFILE/reg_out[26][5] ), .A2(net77338), .ZN(n8016) );
  NAND2_X2 U8832 ( .A1(\REGFILE/reg_out[24][5] ), .A2(net77304), .ZN(n8015) );
  NAND4_X2 U8833 ( .A1(n8018), .A2(n8017), .A3(n8016), .A4(n8015), .ZN(n8019)
         );
  NAND2_X2 U8834 ( .A1(\REGFILE/reg_out[22][5] ), .A2(net77556), .ZN(n8024) );
  NAND2_X2 U8835 ( .A1(\REGFILE/reg_out[17][5] ), .A2(net77520), .ZN(n8023) );
  NAND2_X2 U8836 ( .A1(\REGFILE/reg_out[23][5] ), .A2(net77484), .ZN(n8022) );
  NAND2_X2 U8837 ( .A1(\REGFILE/reg_out[21][5] ), .A2(net77456), .ZN(n8021) );
  NAND4_X2 U8838 ( .A1(n8024), .A2(n8023), .A3(n8022), .A4(n8021), .ZN(n8030)
         );
  NAND2_X2 U8839 ( .A1(\REGFILE/reg_out[19][5] ), .A2(net77410), .ZN(n8028) );
  NAND2_X2 U8840 ( .A1(\REGFILE/reg_out[20][5] ), .A2(net77376), .ZN(n8027) );
  NAND2_X2 U8841 ( .A1(\REGFILE/reg_out[18][5] ), .A2(net77338), .ZN(n8026) );
  NAND2_X2 U8842 ( .A1(\REGFILE/reg_out[16][5] ), .A2(net77304), .ZN(n8025) );
  NAND4_X2 U8843 ( .A1(n8028), .A2(n8027), .A3(n8026), .A4(n8025), .ZN(n8029)
         );
  NAND2_X2 U8844 ( .A1(\REGFILE/reg_out[14][5] ), .A2(net77556), .ZN(n8034) );
  NAND2_X2 U8845 ( .A1(\REGFILE/reg_out[9][5] ), .A2(net77520), .ZN(n8033) );
  NAND2_X2 U8846 ( .A1(\REGFILE/reg_out[15][5] ), .A2(net77484), .ZN(n8032) );
  NAND2_X2 U8847 ( .A1(\REGFILE/reg_out[13][5] ), .A2(net77456), .ZN(n8031) );
  NAND4_X2 U8848 ( .A1(n8034), .A2(n8033), .A3(n8032), .A4(n8031), .ZN(n8040)
         );
  NAND2_X2 U8849 ( .A1(\REGFILE/reg_out[11][5] ), .A2(net77410), .ZN(n8038) );
  NAND2_X2 U8850 ( .A1(\REGFILE/reg_out[12][5] ), .A2(net77376), .ZN(n8037) );
  NAND2_X2 U8851 ( .A1(\REGFILE/reg_out[8][5] ), .A2(net77304), .ZN(n8035) );
  NAND4_X2 U8852 ( .A1(n8038), .A2(n8037), .A3(n8036), .A4(n8035), .ZN(n8039)
         );
  NAND2_X2 U8853 ( .A1(\REGFILE/reg_out[6][5] ), .A2(net77556), .ZN(n8044) );
  NAND2_X2 U8854 ( .A1(\REGFILE/reg_out[1][5] ), .A2(net77520), .ZN(n8043) );
  NAND2_X2 U8855 ( .A1(\REGFILE/reg_out[7][5] ), .A2(net77484), .ZN(n8042) );
  NAND4_X2 U8856 ( .A1(n8044), .A2(n8043), .A3(n8042), .A4(n8041), .ZN(n8050)
         );
  NAND2_X2 U8857 ( .A1(\REGFILE/reg_out[3][5] ), .A2(net77410), .ZN(n8048) );
  NAND2_X2 U8858 ( .A1(\REGFILE/reg_out[4][5] ), .A2(net77376), .ZN(n8047) );
  NAND2_X2 U8859 ( .A1(\REGFILE/reg_out[0][5] ), .A2(net77304), .ZN(n8045) );
  NAND4_X2 U8860 ( .A1(n8048), .A2(n8047), .A3(n8046), .A4(n8045), .ZN(n8049)
         );
  NAND4_X2 U8861 ( .A1(n8054), .A2(n8053), .A3(n8052), .A4(n8051), .ZN(n8424)
         );
  NAND2_X2 U8862 ( .A1(n8424), .A2(n4866), .ZN(n10396) );
  INV_X4 U8863 ( .A(n10396), .ZN(\WIRE_ALU_A/MUX2TO1_32BIT[5].MUX/N1 ) );
  NAND2_X2 U8864 ( .A1(\REGFILE/reg_out[30][4] ), .A2(net77554), .ZN(n8058) );
  NAND2_X2 U8865 ( .A1(\REGFILE/reg_out[25][4] ), .A2(net77518), .ZN(n8057) );
  NAND2_X2 U8866 ( .A1(\REGFILE/reg_out[31][4] ), .A2(net77482), .ZN(n8056) );
  NAND2_X2 U8867 ( .A1(\REGFILE/reg_out[29][4] ), .A2(net77456), .ZN(n8055) );
  NAND4_X2 U8868 ( .A1(n8058), .A2(n8057), .A3(n8056), .A4(n8055), .ZN(n8064)
         );
  NAND2_X2 U8869 ( .A1(\REGFILE/reg_out[27][4] ), .A2(net77410), .ZN(n8062) );
  NAND2_X2 U8870 ( .A1(\REGFILE/reg_out[28][4] ), .A2(net77376), .ZN(n8061) );
  NAND2_X2 U8871 ( .A1(\REGFILE/reg_out[26][4] ), .A2(net77338), .ZN(n8060) );
  NAND2_X2 U8872 ( .A1(\REGFILE/reg_out[24][4] ), .A2(net77302), .ZN(n8059) );
  NAND4_X2 U8873 ( .A1(n8062), .A2(n8061), .A3(n8060), .A4(n8059), .ZN(n8063)
         );
  NAND2_X2 U8874 ( .A1(\REGFILE/reg_out[22][4] ), .A2(net77554), .ZN(n8068) );
  NAND2_X2 U8875 ( .A1(\REGFILE/reg_out[17][4] ), .A2(net77518), .ZN(n8067) );
  NAND2_X2 U8876 ( .A1(\REGFILE/reg_out[23][4] ), .A2(net77482), .ZN(n8066) );
  NAND2_X2 U8877 ( .A1(\REGFILE/reg_out[21][4] ), .A2(net77456), .ZN(n8065) );
  NAND4_X2 U8878 ( .A1(n8068), .A2(n8067), .A3(n8066), .A4(n8065), .ZN(n8074)
         );
  NAND2_X2 U8879 ( .A1(\REGFILE/reg_out[19][4] ), .A2(net77410), .ZN(n8072) );
  NAND2_X2 U8880 ( .A1(\REGFILE/reg_out[20][4] ), .A2(net77376), .ZN(n8071) );
  NAND2_X2 U8881 ( .A1(\REGFILE/reg_out[18][4] ), .A2(net77338), .ZN(n8070) );
  NAND2_X2 U8882 ( .A1(\REGFILE/reg_out[16][4] ), .A2(net77302), .ZN(n8069) );
  NAND4_X2 U8883 ( .A1(n8072), .A2(n8071), .A3(n8070), .A4(n8069), .ZN(n8073)
         );
  NAND2_X2 U8884 ( .A1(\REGFILE/reg_out[14][4] ), .A2(net77554), .ZN(n8078) );
  NAND2_X2 U8885 ( .A1(\REGFILE/reg_out[9][4] ), .A2(net77518), .ZN(n8077) );
  NAND2_X2 U8886 ( .A1(\REGFILE/reg_out[15][4] ), .A2(net77482), .ZN(n8076) );
  NAND2_X2 U8887 ( .A1(\REGFILE/reg_out[13][4] ), .A2(net77456), .ZN(n8075) );
  NAND4_X2 U8888 ( .A1(n8078), .A2(n8077), .A3(n8076), .A4(n8075), .ZN(n8084)
         );
  NAND2_X2 U8889 ( .A1(\REGFILE/reg_out[11][4] ), .A2(net77410), .ZN(n8082) );
  NAND2_X2 U8890 ( .A1(\REGFILE/reg_out[12][4] ), .A2(net77376), .ZN(n8081) );
  NAND2_X2 U8891 ( .A1(\REGFILE/reg_out[10][4] ), .A2(net77338), .ZN(n8080) );
  NAND2_X2 U8892 ( .A1(\REGFILE/reg_out[8][4] ), .A2(net77302), .ZN(n8079) );
  NAND4_X2 U8893 ( .A1(n8082), .A2(n8081), .A3(n8080), .A4(n8079), .ZN(n8083)
         );
  NAND2_X2 U8894 ( .A1(\REGFILE/reg_out[6][4] ), .A2(net77554), .ZN(n8088) );
  NAND2_X2 U8895 ( .A1(\REGFILE/reg_out[7][4] ), .A2(net77482), .ZN(n8086) );
  NAND2_X2 U8896 ( .A1(\REGFILE/reg_out[5][4] ), .A2(net77456), .ZN(n8085) );
  NAND4_X2 U8897 ( .A1(n8088), .A2(n8087), .A3(n8086), .A4(n8085), .ZN(n8094)
         );
  NAND2_X2 U8898 ( .A1(n5982), .A2(net77410), .ZN(n8092) );
  NAND2_X2 U8899 ( .A1(\REGFILE/reg_out[4][4] ), .A2(net77376), .ZN(n8091) );
  NAND2_X2 U8900 ( .A1(\REGFILE/reg_out[2][4] ), .A2(net77338), .ZN(n8090) );
  NAND2_X2 U8901 ( .A1(\REGFILE/reg_out[0][4] ), .A2(net77302), .ZN(n8089) );
  NAND4_X2 U8902 ( .A1(n8092), .A2(n8091), .A3(n8090), .A4(n8089), .ZN(n8093)
         );
  NAND4_X2 U8903 ( .A1(n8098), .A2(n8097), .A3(n8096), .A4(n8095), .ZN(n8425)
         );
  NAND2_X2 U8904 ( .A1(n8425), .A2(n4866), .ZN(n9954) );
  INV_X4 U8905 ( .A(n9954), .ZN(\WIRE_ALU_A/MUX2TO1_32BIT[4].MUX/N1 ) );
  NAND2_X2 U8906 ( .A1(\REGFILE/reg_out[30][3] ), .A2(net77554), .ZN(n8102) );
  NAND2_X2 U8907 ( .A1(n5957), .A2(net77518), .ZN(n8101) );
  NAND2_X2 U8908 ( .A1(\REGFILE/reg_out[31][3] ), .A2(net77482), .ZN(n8100) );
  NAND2_X2 U8909 ( .A1(\REGFILE/reg_out[29][3] ), .A2(net77460), .ZN(n8099) );
  NAND4_X2 U8910 ( .A1(n8102), .A2(n8101), .A3(n8100), .A4(n8099), .ZN(n8108)
         );
  NAND2_X2 U8911 ( .A1(\REGFILE/reg_out[27][3] ), .A2(net77410), .ZN(n8106) );
  NAND2_X2 U8912 ( .A1(\REGFILE/reg_out[28][3] ), .A2(net77376), .ZN(n8105) );
  NAND2_X2 U8913 ( .A1(\REGFILE/reg_out[26][3] ), .A2(net77338), .ZN(n8104) );
  NAND2_X2 U8914 ( .A1(\REGFILE/reg_out[24][3] ), .A2(net77302), .ZN(n8103) );
  NAND4_X2 U8915 ( .A1(n8106), .A2(n8105), .A3(n8104), .A4(n8103), .ZN(n8107)
         );
  NAND2_X2 U8916 ( .A1(\REGFILE/reg_out[22][3] ), .A2(net77554), .ZN(n8112) );
  NAND2_X2 U8917 ( .A1(\REGFILE/reg_out[17][3] ), .A2(net77518), .ZN(n8111) );
  NAND2_X2 U8918 ( .A1(\REGFILE/reg_out[23][3] ), .A2(net77482), .ZN(n8110) );
  NAND2_X2 U8919 ( .A1(\REGFILE/reg_out[21][3] ), .A2(net77456), .ZN(n8109) );
  NAND4_X2 U8920 ( .A1(n8112), .A2(n8111), .A3(n8110), .A4(n8109), .ZN(n8118)
         );
  NAND2_X2 U8921 ( .A1(\REGFILE/reg_out[19][3] ), .A2(net77410), .ZN(n8116) );
  NAND2_X2 U8922 ( .A1(\REGFILE/reg_out[20][3] ), .A2(net77376), .ZN(n8115) );
  NAND2_X2 U8923 ( .A1(\REGFILE/reg_out[18][3] ), .A2(net77338), .ZN(n8114) );
  NAND2_X2 U8924 ( .A1(\REGFILE/reg_out[16][3] ), .A2(net77302), .ZN(n8113) );
  NAND4_X2 U8925 ( .A1(n8116), .A2(n8115), .A3(n8114), .A4(n8113), .ZN(n8117)
         );
  NAND2_X2 U8926 ( .A1(\REGFILE/reg_out[14][3] ), .A2(net77554), .ZN(n8122) );
  NAND2_X2 U8927 ( .A1(\REGFILE/reg_out[9][3] ), .A2(net77518), .ZN(n8121) );
  NAND2_X2 U8928 ( .A1(\REGFILE/reg_out[15][3] ), .A2(net77482), .ZN(n8120) );
  NAND2_X2 U8929 ( .A1(\REGFILE/reg_out[13][3] ), .A2(net77456), .ZN(n8119) );
  NAND4_X2 U8930 ( .A1(n8122), .A2(n8121), .A3(n8120), .A4(n8119), .ZN(n8128)
         );
  NAND2_X2 U8931 ( .A1(\REGFILE/reg_out[11][3] ), .A2(net77410), .ZN(n8126) );
  NAND2_X2 U8932 ( .A1(\REGFILE/reg_out[12][3] ), .A2(net77376), .ZN(n8125) );
  NAND2_X2 U8933 ( .A1(\REGFILE/reg_out[10][3] ), .A2(net77338), .ZN(n8124) );
  NAND2_X2 U8934 ( .A1(\REGFILE/reg_out[8][3] ), .A2(net77302), .ZN(n8123) );
  NAND4_X2 U8935 ( .A1(n8126), .A2(n8125), .A3(n8124), .A4(n8123), .ZN(n8127)
         );
  NAND2_X2 U8936 ( .A1(\REGFILE/reg_out[6][3] ), .A2(net77554), .ZN(n8132) );
  NAND2_X2 U8937 ( .A1(\REGFILE/reg_out[1][3] ), .A2(net77518), .ZN(n8131) );
  NAND2_X2 U8938 ( .A1(\REGFILE/reg_out[7][3] ), .A2(net77482), .ZN(n8130) );
  NAND2_X2 U8939 ( .A1(\REGFILE/reg_out[5][3] ), .A2(net77456), .ZN(n8129) );
  NAND4_X2 U8940 ( .A1(n8132), .A2(n8131), .A3(n8130), .A4(n8129), .ZN(n8138)
         );
  NAND2_X2 U8941 ( .A1(\REGFILE/reg_out[4][3] ), .A2(net77376), .ZN(n8135) );
  NAND2_X2 U8942 ( .A1(\REGFILE/reg_out[0][3] ), .A2(net77302), .ZN(n8133) );
  NAND4_X2 U8943 ( .A1(n8136), .A2(n8135), .A3(n8134), .A4(n8133), .ZN(n8137)
         );
  NAND4_X2 U8944 ( .A1(n8142), .A2(n8141), .A3(n8140), .A4(n8139), .ZN(n8423)
         );
  NAND2_X2 U8945 ( .A1(n8423), .A2(n4866), .ZN(n10404) );
  INV_X4 U8946 ( .A(n10404), .ZN(\WIRE_ALU_A/MUX2TO1_32BIT[3].MUX/N1 ) );
  NAND2_X2 U8947 ( .A1(\REGFILE/reg_out[30][2] ), .A2(net77554), .ZN(n8146) );
  NAND2_X2 U8948 ( .A1(\REGFILE/reg_out[25][2] ), .A2(net77518), .ZN(n8145) );
  NAND2_X2 U8949 ( .A1(\REGFILE/reg_out[31][2] ), .A2(net77482), .ZN(n8144) );
  NAND2_X2 U8950 ( .A1(\REGFILE/reg_out[29][2] ), .A2(net77456), .ZN(n8143) );
  NAND4_X2 U8951 ( .A1(n8146), .A2(n8145), .A3(n8144), .A4(n8143), .ZN(n8152)
         );
  NAND2_X2 U8952 ( .A1(\REGFILE/reg_out[27][2] ), .A2(net77410), .ZN(n8150) );
  NAND2_X2 U8953 ( .A1(\REGFILE/reg_out[28][2] ), .A2(net77376), .ZN(n8149) );
  NAND2_X2 U8954 ( .A1(\REGFILE/reg_out[26][2] ), .A2(net77338), .ZN(n8148) );
  NAND2_X2 U8955 ( .A1(\REGFILE/reg_out[24][2] ), .A2(net77302), .ZN(n8147) );
  NAND4_X2 U8956 ( .A1(n8150), .A2(n8149), .A3(n8148), .A4(n8147), .ZN(n8151)
         );
  NAND2_X2 U8957 ( .A1(\REGFILE/reg_out[22][2] ), .A2(net77554), .ZN(n8156) );
  NAND2_X2 U8958 ( .A1(\REGFILE/reg_out[17][2] ), .A2(net77518), .ZN(n8155) );
  NAND2_X2 U8959 ( .A1(\REGFILE/reg_out[23][2] ), .A2(net77482), .ZN(n8154) );
  NAND2_X2 U8960 ( .A1(\REGFILE/reg_out[21][2] ), .A2(net77456), .ZN(n8153) );
  NAND4_X2 U8961 ( .A1(n8156), .A2(n8155), .A3(n8154), .A4(n8153), .ZN(n8162)
         );
  NAND2_X2 U8962 ( .A1(\REGFILE/reg_out[19][2] ), .A2(net77410), .ZN(n8160) );
  NAND2_X2 U8963 ( .A1(\REGFILE/reg_out[20][2] ), .A2(net77376), .ZN(n8159) );
  NAND2_X2 U8964 ( .A1(\REGFILE/reg_out[18][2] ), .A2(net77338), .ZN(n8158) );
  NAND2_X2 U8965 ( .A1(\REGFILE/reg_out[16][2] ), .A2(net77302), .ZN(n8157) );
  NAND4_X2 U8966 ( .A1(n8160), .A2(n8159), .A3(n8158), .A4(n8157), .ZN(n8161)
         );
  NAND2_X2 U8967 ( .A1(\REGFILE/reg_out[14][2] ), .A2(net77554), .ZN(n8166) );
  NAND2_X2 U8968 ( .A1(\REGFILE/reg_out[9][2] ), .A2(net77518), .ZN(n8165) );
  NAND2_X2 U8969 ( .A1(\REGFILE/reg_out[15][2] ), .A2(net77482), .ZN(n8164) );
  NAND2_X2 U8970 ( .A1(\REGFILE/reg_out[13][2] ), .A2(net77456), .ZN(n8163) );
  NAND4_X2 U8971 ( .A1(n8166), .A2(n8165), .A3(n8164), .A4(n8163), .ZN(n8172)
         );
  NAND2_X2 U8972 ( .A1(\REGFILE/reg_out[11][2] ), .A2(net77410), .ZN(n8170) );
  NAND2_X2 U8973 ( .A1(\REGFILE/reg_out[12][2] ), .A2(net77376), .ZN(n8169) );
  NAND2_X2 U8974 ( .A1(\REGFILE/reg_out[10][2] ), .A2(net77338), .ZN(n8168) );
  NAND2_X2 U8975 ( .A1(\REGFILE/reg_out[8][2] ), .A2(net77302), .ZN(n8167) );
  NAND4_X2 U8976 ( .A1(n8170), .A2(n8169), .A3(n8168), .A4(n8167), .ZN(n8171)
         );
  NAND2_X2 U8977 ( .A1(\REGFILE/reg_out[6][2] ), .A2(net77554), .ZN(n8176) );
  NAND2_X2 U8978 ( .A1(\REGFILE/reg_out[1][2] ), .A2(net77518), .ZN(n8175) );
  NAND2_X2 U8979 ( .A1(\REGFILE/reg_out[7][2] ), .A2(net77482), .ZN(n8174) );
  NAND2_X2 U8980 ( .A1(\REGFILE/reg_out[5][2] ), .A2(net77456), .ZN(n8173) );
  NAND4_X2 U8981 ( .A1(n8176), .A2(n8175), .A3(n8174), .A4(n8173), .ZN(n8182)
         );
  NAND2_X2 U8982 ( .A1(\REGFILE/reg_out[3][2] ), .A2(net77410), .ZN(n8180) );
  NAND2_X2 U8983 ( .A1(\REGFILE/reg_out[4][2] ), .A2(net77376), .ZN(n8179) );
  NAND2_X2 U8984 ( .A1(\REGFILE/reg_out[2][2] ), .A2(net77338), .ZN(n8178) );
  NAND2_X2 U8985 ( .A1(\REGFILE/reg_out[0][2] ), .A2(net77302), .ZN(n8177) );
  NAND4_X2 U8986 ( .A1(n8180), .A2(n8179), .A3(n8178), .A4(n8177), .ZN(n8181)
         );
  NAND4_X2 U8987 ( .A1(n8186), .A2(n8185), .A3(n8184), .A4(n8183), .ZN(n8421)
         );
  NAND2_X2 U8988 ( .A1(n8421), .A2(n4866), .ZN(n10109) );
  INV_X4 U8989 ( .A(n10109), .ZN(\WIRE_ALU_A/MUX2TO1_32BIT[2].MUX/N1 ) );
  NAND2_X2 U8990 ( .A1(\REGFILE/reg_out[25][1] ), .A2(net77516), .ZN(n8189) );
  NAND2_X2 U8991 ( .A1(\REGFILE/reg_out[31][1] ), .A2(net77480), .ZN(n8188) );
  NAND4_X2 U8992 ( .A1(n8190), .A2(n8189), .A3(n8188), .A4(n8187), .ZN(n8196)
         );
  NAND2_X2 U8993 ( .A1(\REGFILE/reg_out[27][1] ), .A2(net77410), .ZN(n8194) );
  NAND2_X2 U8994 ( .A1(\REGFILE/reg_out[28][1] ), .A2(net77376), .ZN(n8193) );
  NAND2_X2 U8995 ( .A1(\REGFILE/reg_out[26][1] ), .A2(net77336), .ZN(n8192) );
  NAND4_X2 U8997 ( .A1(n8194), .A2(n8193), .A3(n8192), .A4(n8191), .ZN(n8195)
         );
  NAND2_X2 U8998 ( .A1(\REGFILE/reg_out[17][1] ), .A2(net77516), .ZN(n8199) );
  NAND2_X2 U8999 ( .A1(\REGFILE/reg_out[23][1] ), .A2(net77480), .ZN(n8198) );
  NAND4_X2 U9000 ( .A1(n8200), .A2(n8199), .A3(n8198), .A4(n8197), .ZN(n8206)
         );
  NAND2_X2 U9001 ( .A1(\REGFILE/reg_out[19][1] ), .A2(net77410), .ZN(n8204) );
  NAND2_X2 U9002 ( .A1(\REGFILE/reg_out[18][1] ), .A2(net77336), .ZN(n8202) );
  NAND4_X2 U9004 ( .A1(n8204), .A2(n8203), .A3(n8202), .A4(n8201), .ZN(n8205)
         );
  NAND2_X2 U9005 ( .A1(\REGFILE/reg_out[9][1] ), .A2(net77516), .ZN(n8209) );
  NAND2_X2 U9006 ( .A1(\REGFILE/reg_out[15][1] ), .A2(net77480), .ZN(n8208) );
  NAND4_X2 U9007 ( .A1(n8210), .A2(n8209), .A3(n8208), .A4(n8207), .ZN(n8216)
         );
  NAND2_X2 U9008 ( .A1(\REGFILE/reg_out[11][1] ), .A2(net77410), .ZN(n8214) );
  NAND2_X2 U9009 ( .A1(\REGFILE/reg_out[12][1] ), .A2(net77376), .ZN(n8213) );
  NAND2_X2 U9010 ( .A1(\REGFILE/reg_out[10][1] ), .A2(net77336), .ZN(n8212) );
  NAND4_X2 U9012 ( .A1(n8214), .A2(n8213), .A3(n8212), .A4(n8211), .ZN(n8215)
         );
  NAND2_X2 U9013 ( .A1(\REGFILE/reg_out[1][1] ), .A2(net77516), .ZN(n8219) );
  NAND2_X2 U9014 ( .A1(\REGFILE/reg_out[7][1] ), .A2(net77480), .ZN(n8218) );
  NAND4_X2 U9015 ( .A1(n8220), .A2(n8219), .A3(n8218), .A4(n8217), .ZN(n8226)
         );
  NAND2_X2 U9016 ( .A1(\REGFILE/reg_out[3][1] ), .A2(net77410), .ZN(n8224) );
  NAND2_X2 U9017 ( .A1(\REGFILE/reg_out[4][1] ), .A2(net77376), .ZN(n8223) );
  NAND2_X2 U9018 ( .A1(\REGFILE/reg_out[2][1] ), .A2(net77336), .ZN(n8222) );
  NAND4_X2 U9020 ( .A1(n8224), .A2(n8223), .A3(n8222), .A4(n8221), .ZN(n8225)
         );
  NAND4_X2 U9021 ( .A1(n8230), .A2(n8229), .A3(n8228), .A4(n8227), .ZN(n8422)
         );
  NAND2_X2 U9022 ( .A1(n8422), .A2(n4866), .ZN(net71273) );
  NAND2_X2 U9023 ( .A1(\REGFILE/reg_out[25][0] ), .A2(net77516), .ZN(n8233) );
  NAND2_X2 U9024 ( .A1(\REGFILE/reg_out[31][0] ), .A2(net77480), .ZN(n8232) );
  NAND4_X2 U9025 ( .A1(n8234), .A2(n8233), .A3(n8232), .A4(n8231), .ZN(n8240)
         );
  NAND2_X2 U9026 ( .A1(\REGFILE/reg_out[27][0] ), .A2(net77410), .ZN(n8238) );
  NAND2_X2 U9028 ( .A1(\REGFILE/reg_out[26][0] ), .A2(net77336), .ZN(n8236) );
  NAND2_X2 U9029 ( .A1(\REGFILE/reg_out[24][0] ), .A2(net77300), .ZN(n8235) );
  NAND4_X2 U9030 ( .A1(n8238), .A2(n8237), .A3(n8236), .A4(n8235), .ZN(n8239)
         );
  NAND2_X2 U9031 ( .A1(\REGFILE/reg_out[17][0] ), .A2(net77516), .ZN(n8243) );
  NAND2_X2 U9032 ( .A1(\REGFILE/reg_out[23][0] ), .A2(net77480), .ZN(n8242) );
  NAND4_X2 U9033 ( .A1(n8244), .A2(n8243), .A3(n8242), .A4(n8241), .ZN(n8250)
         );
  NAND2_X2 U9034 ( .A1(\REGFILE/reg_out[19][0] ), .A2(net77410), .ZN(n8248) );
  NAND2_X2 U9035 ( .A1(\REGFILE/reg_out[18][0] ), .A2(net77336), .ZN(n8246) );
  NAND2_X2 U9036 ( .A1(\REGFILE/reg_out[16][0] ), .A2(net77300), .ZN(n8245) );
  NAND4_X2 U9037 ( .A1(n8248), .A2(n8247), .A3(n8246), .A4(n8245), .ZN(n8249)
         );
  NAND2_X2 U9038 ( .A1(\REGFILE/reg_out[9][0] ), .A2(net77516), .ZN(n8253) );
  NAND2_X2 U9039 ( .A1(\REGFILE/reg_out[15][0] ), .A2(net77480), .ZN(n8252) );
  NAND4_X2 U9040 ( .A1(n8254), .A2(n8253), .A3(n8252), .A4(n8251), .ZN(n8260)
         );
  NAND2_X2 U9041 ( .A1(\REGFILE/reg_out[11][0] ), .A2(net77410), .ZN(n8258) );
  NAND2_X2 U9042 ( .A1(\REGFILE/reg_out[12][0] ), .A2(net77376), .ZN(n8257) );
  NAND2_X2 U9043 ( .A1(\REGFILE/reg_out[10][0] ), .A2(net77336), .ZN(n8256) );
  NAND4_X2 U9045 ( .A1(n8258), .A2(n8257), .A3(n8256), .A4(n8255), .ZN(n8259)
         );
  NAND2_X2 U9046 ( .A1(\REGFILE/reg_out[6][0] ), .A2(net77562), .ZN(n8264) );
  NAND2_X2 U9047 ( .A1(\REGFILE/reg_out[1][0] ), .A2(net77526), .ZN(n8263) );
  NAND2_X2 U9048 ( .A1(\REGFILE/reg_out[7][0] ), .A2(net77490), .ZN(n8262) );
  NAND2_X2 U9049 ( .A1(\REGFILE/reg_out[5][0] ), .A2(net77454), .ZN(n8261) );
  NAND4_X2 U9050 ( .A1(n8264), .A2(n8263), .A3(n8262), .A4(n8261), .ZN(n8270)
         );
  NAND2_X2 U9051 ( .A1(\REGFILE/reg_out[3][0] ), .A2(net77418), .ZN(n8268) );
  NAND2_X2 U9052 ( .A1(\REGFILE/reg_out[4][0] ), .A2(net77382), .ZN(n8267) );
  NAND2_X2 U9053 ( .A1(\REGFILE/reg_out[2][0] ), .A2(net77346), .ZN(n8266) );
  NAND2_X2 U9054 ( .A1(\REGFILE/reg_out[0][0] ), .A2(net77310), .ZN(n8265) );
  NAND4_X2 U9055 ( .A1(n8268), .A2(n8267), .A3(n8266), .A4(n8265), .ZN(n8269)
         );
  NAND4_X2 U9056 ( .A1(n8274), .A2(n8273), .A3(n8272), .A4(n8271), .ZN(n8416)
         );
  NAND2_X2 U9057 ( .A1(n8416), .A2(n4866), .ZN(net70535) );
  NAND2_X2 U9058 ( .A1(instructionAddr_out[28]), .A2(instructionAddr_out[29]), 
        .ZN(n8337) );
  NOR2_X4 U9059 ( .A1(n8337), .A2(n4969), .ZN(n8344) );
  NAND2_X2 U9060 ( .A1(instructionAddr_out[26]), .A2(n8344), .ZN(n8343) );
  INV_X4 U9061 ( .A(n8343), .ZN(n8275) );
  NAND2_X2 U9062 ( .A1(instructionAddr_out[25]), .A2(n8275), .ZN(n8326) );
  NAND2_X2 U9063 ( .A1(instructionAddr_out[24]), .A2(n8328), .ZN(n8327) );
  INV_X4 U9064 ( .A(n8327), .ZN(n8276) );
  NAND2_X2 U9065 ( .A1(instructionAddr_out[23]), .A2(n8276), .ZN(n8321) );
  NAND2_X2 U9066 ( .A1(instructionAddr_out[22]), .A2(n8323), .ZN(n8322) );
  INV_X4 U9067 ( .A(n8322), .ZN(n8277) );
  NAND2_X2 U9068 ( .A1(instructionAddr_out[21]), .A2(n8277), .ZN(n8316) );
  NAND2_X2 U9069 ( .A1(instructionAddr_out[20]), .A2(n8318), .ZN(n8317) );
  INV_X4 U9070 ( .A(n8317), .ZN(n8278) );
  NAND2_X2 U9071 ( .A1(instructionAddr_out[19]), .A2(n8278), .ZN(n8315) );
  INV_X4 U9072 ( .A(n8315), .ZN(n8279) );
  NAND2_X2 U9073 ( .A1(instructionAddr_out[18]), .A2(n8279), .ZN(n8314) );
  INV_X4 U9074 ( .A(n8314), .ZN(n8280) );
  NAND2_X2 U9075 ( .A1(instructionAddr_out[17]), .A2(n8280), .ZN(n8312) );
  INV_X4 U9076 ( .A(n8312), .ZN(n8281) );
  NAND2_X2 U9077 ( .A1(instructionAddr_out[16]), .A2(n8281), .ZN(n8364) );
  INV_X4 U9078 ( .A(n8364), .ZN(n8282) );
  NAND2_X2 U9079 ( .A1(instructionAddr_out[15]), .A2(n8282), .ZN(n8362) );
  INV_X4 U9080 ( .A(n8362), .ZN(n8310) );
  NAND3_X4 U9081 ( .A1(instructionAddr_out[13]), .A2(instructionAddr_out[14]), 
        .A3(n8310), .ZN(n8308) );
  INV_X4 U9082 ( .A(n8308), .ZN(n8283) );
  NAND3_X4 U9083 ( .A1(instructionAddr_out[11]), .A2(instructionAddr_out[12]), 
        .A3(n8283), .ZN(n8303) );
  INV_X4 U9084 ( .A(n8303), .ZN(n8302) );
  NAND3_X4 U9085 ( .A1(instructionAddr_out[10]), .A2(instructionAddr_out[9]), 
        .A3(n8302), .ZN(n8379) );
  INV_X4 U9086 ( .A(n8379), .ZN(n8284) );
  NAND3_X4 U9087 ( .A1(instructionAddr_out[7]), .A2(instructionAddr_out[8]), 
        .A3(n8284), .ZN(n8296) );
  INV_X4 U9088 ( .A(n8296), .ZN(n8389) );
  NAND3_X4 U9089 ( .A1(instructionAddr_out[6]), .A2(instructionAddr_out[5]), 
        .A3(n8389), .ZN(n8391) );
  INV_X4 U9090 ( .A(n8391), .ZN(n8285) );
  NAND2_X2 U9091 ( .A1(instructionAddr_out[4]), .A2(n8285), .ZN(n8293) );
  INV_X4 U9092 ( .A(n8293), .ZN(n8291) );
  NAND2_X2 U9093 ( .A1(instructionAddr_out[3]), .A2(n8291), .ZN(n8290) );
  INV_X4 U9094 ( .A(n8290), .ZN(n8286) );
  NAND2_X2 U9095 ( .A1(instructionAddr_out[2]), .A2(n8286), .ZN(n8289) );
  INV_X4 U9096 ( .A(n8289), .ZN(n10538) );
  XNOR2_X2 U9097 ( .A(instructionAddr_out[1]), .B(n10538), .ZN(net73771) );
  NAND2_X2 U9098 ( .A1(instruction[3]), .A2(net74011), .ZN(net73519) );
  INV_X4 U9099 ( .A(net73519), .ZN(net74009) );
  NAND2_X2 U9100 ( .A1(net73878), .A2(n8287), .ZN(n8288) );
  NAND2_X2 U9101 ( .A1(net74009), .A2(net73878), .ZN(net73877) );
  NAND2_X2 U9102 ( .A1(n8288), .A2(net73877), .ZN(net70531) );
  INV_X4 U9103 ( .A(net73778), .ZN(net73855) );
  AOI21_X4 U9104 ( .B1(n8290), .B2(n4923), .A(n10538), .ZN(net71396) );
  XNOR2_X2 U9105 ( .A(net73858), .B(net71396), .ZN(n8470) );
  XNOR2_X2 U9106 ( .A(instructionAddr_out[3]), .B(n8291), .ZN(n8292) );
  INV_X4 U9107 ( .A(n8292), .ZN(n10043) );
  NAND2_X2 U9108 ( .A1(n10043), .A2(net73858), .ZN(n8397) );
  AOI21_X4 U9109 ( .B1(n8391), .B2(n4924), .A(n8291), .ZN(n9965) );
  XNOR2_X2 U9110 ( .A(net73858), .B(n9965), .ZN(n8479) );
  XNOR2_X2 U9111 ( .A(instructionAddr_out[6]), .B(n8389), .ZN(n8294) );
  INV_X4 U9112 ( .A(n8294), .ZN(n9671) );
  NAND2_X2 U9113 ( .A1(net73858), .A2(n9671), .ZN(n8388) );
  NAND2_X2 U9114 ( .A1(n8297), .A2(n8296), .ZN(n8298) );
  INV_X4 U9115 ( .A(n8298), .ZN(n9700) );
  XNOR2_X2 U9116 ( .A(n8385), .B(n9700), .ZN(n8493) );
  AOI21_X4 U9117 ( .B1(n8302), .B2(instructionAddr_out[10]), .A(
        instructionAddr_out[9]), .ZN(n8299) );
  INV_X4 U9118 ( .A(n8299), .ZN(n8300) );
  NAND2_X2 U9119 ( .A1(n8300), .A2(n8379), .ZN(n8499) );
  NAND2_X2 U9120 ( .A1(net73988), .A2(net73877), .ZN(n8378) );
  XNOR2_X2 U9121 ( .A(n8499), .B(n8378), .ZN(n8497) );
  XNOR2_X2 U9122 ( .A(instructionAddr_out[10]), .B(n8302), .ZN(n8376) );
  NAND2_X2 U9123 ( .A1(n8304), .A2(n8303), .ZN(n8305) );
  INV_X4 U9124 ( .A(n8305), .ZN(n9864) );
  XNOR2_X2 U9125 ( .A(n8374), .B(n9864), .ZN(n8516) );
  XNOR2_X2 U9126 ( .A(n8308), .B(n4908), .ZN(n9107) );
  NAND2_X2 U9127 ( .A1(n8306), .A2(net73877), .ZN(n8372) );
  AOI21_X4 U9128 ( .B1(n8310), .B2(instructionAddr_out[14]), .A(
        instructionAddr_out[13]), .ZN(n8307) );
  INV_X4 U9129 ( .A(n8307), .ZN(n8309) );
  NAND2_X2 U9130 ( .A1(n8309), .A2(n8308), .ZN(n8368) );
  NAND2_X2 U9131 ( .A1(net73974), .A2(net73877), .ZN(n8367) );
  XNOR2_X2 U9132 ( .A(n8368), .B(n8367), .ZN(n9389) );
  XNOR2_X2 U9133 ( .A(instructionAddr_out[14]), .B(n8310), .ZN(n8311) );
  INV_X4 U9134 ( .A(n8311), .ZN(n10261) );
  XNOR2_X2 U9135 ( .A(net73900), .B(n10261), .ZN(n8502) );
  INV_X4 U9136 ( .A(\PCLOGIC/imm16_32 [16]), .ZN(net73908) );
  OAI21_X4 U9137 ( .B1(instructionAddr_out[16]), .B2(n8281), .A(n8364), .ZN(
        n8512) );
  XNOR2_X2 U9138 ( .A(n8314), .B(n5084), .ZN(n8313) );
  INV_X4 U9139 ( .A(n8313), .ZN(n9041) );
  INV_X4 U9140 ( .A(\PCLOGIC/imm16_32 [17]), .ZN(n8650) );
  XNOR2_X2 U9141 ( .A(n8313), .B(n8650), .ZN(n8796) );
  INV_X4 U9142 ( .A(n8796), .ZN(n8360) );
  OAI21_X4 U9143 ( .B1(instructionAddr_out[18]), .B2(n8279), .A(n8314), .ZN(
        n8804) );
  AOI21_X4 U9144 ( .B1(n8317), .B2(n5063), .A(n8279), .ZN(n10003) );
  INV_X4 U9145 ( .A(n8316), .ZN(n8318) );
  OAI21_X4 U9146 ( .B1(instructionAddr_out[20]), .B2(n8318), .A(n8317), .ZN(
        n9279) );
  XNOR2_X2 U9147 ( .A(n8322), .B(n5085), .ZN(n8320) );
  INV_X4 U9148 ( .A(n8320), .ZN(n9569) );
  XNOR2_X2 U9149 ( .A(n8320), .B(n8319), .ZN(n9536) );
  INV_X4 U9150 ( .A(n9536), .ZN(n8357) );
  INV_X4 U9151 ( .A(\PCLOGIC/imm16_32 [22]), .ZN(n8356) );
  INV_X4 U9152 ( .A(n8321), .ZN(n8323) );
  OAI21_X4 U9153 ( .B1(instructionAddr_out[22]), .B2(n8323), .A(n8322), .ZN(
        n8950) );
  XNOR2_X2 U9154 ( .A(n8327), .B(n5086), .ZN(n8325) );
  INV_X4 U9155 ( .A(n8325), .ZN(n9316) );
  XNOR2_X2 U9156 ( .A(n8325), .B(n8324), .ZN(n9283) );
  INV_X4 U9157 ( .A(n9283), .ZN(n8353) );
  INV_X4 U9158 ( .A(\PCLOGIC/imm16_32 [24]), .ZN(n8352) );
  INV_X4 U9159 ( .A(n8326), .ZN(n8328) );
  OAI21_X4 U9160 ( .B1(instructionAddr_out[24]), .B2(n8328), .A(n8327), .ZN(
        n8530) );
  XNOR2_X2 U9161 ( .A(n8343), .B(n5087), .ZN(n8330) );
  INV_X4 U9162 ( .A(n8330), .ZN(n9000) );
  XNOR2_X2 U9163 ( .A(n8330), .B(n8329), .ZN(n8968) );
  INV_X4 U9164 ( .A(n8968), .ZN(n8349) );
  INV_X4 U9165 ( .A(n8331), .ZN(n8788) );
  NAND2_X2 U9166 ( .A1(n8788), .A2(\PCLOGIC/imm16_32 [28]), .ZN(n8336) );
  INV_X4 U9167 ( .A(\PCLOGIC/imm16_32 [28]), .ZN(net73670) );
  XNOR2_X2 U9168 ( .A(n8331), .B(net73670), .ZN(n8690) );
  INV_X4 U9169 ( .A(n8690), .ZN(n8335) );
  NAND2_X2 U9170 ( .A1(instructionAddr_out[31]), .A2(\PCLOGIC/imm16_32 [31]), 
        .ZN(n8699) );
  INV_X4 U9171 ( .A(n8699), .ZN(n8333) );
  XNOR2_X2 U9172 ( .A(instructionAddr_out[30]), .B(\PCLOGIC/imm16_32 [30]), 
        .ZN(n8700) );
  INV_X4 U9173 ( .A(n8700), .ZN(n8332) );
  NAND2_X2 U9174 ( .A1(n8333), .A2(n8332), .ZN(n8702) );
  INV_X4 U9175 ( .A(n8702), .ZN(n8334) );
  AOI21_X4 U9176 ( .B1(instructionAddr_out[30]), .B2(\PCLOGIC/imm16_32 [30]), 
        .A(n8334), .ZN(net73394) );
  XNOR2_X2 U9177 ( .A(instructionAddr_out[29]), .B(\PCLOGIC/imm16_32 [29]), 
        .ZN(net73395) );
  INV_X4 U9178 ( .A(net73395), .ZN(net73938) );
  NAND2_X2 U9179 ( .A1(n8335), .A2(net73400), .ZN(n8691) );
  NAND2_X2 U9180 ( .A1(n8336), .A2(n8691), .ZN(n8686) );
  INV_X4 U9181 ( .A(n8686), .ZN(n8342) );
  INV_X4 U9182 ( .A(n8337), .ZN(n8339) );
  INV_X4 U9183 ( .A(n8344), .ZN(n8338) );
  OAI21_X4 U9184 ( .B1(instructionAddr_out[27]), .B2(n8339), .A(n8338), .ZN(
        n8340) );
  INV_X4 U9185 ( .A(n8340), .ZN(n8908) );
  XNOR2_X2 U9186 ( .A(\PCLOGIC/imm16_32 [27]), .B(n8908), .ZN(n8685) );
  NAND2_X2 U9187 ( .A1(n8908), .A2(\PCLOGIC/imm16_32 [27]), .ZN(n8341) );
  OAI21_X4 U9188 ( .B1(n8342), .B2(n8685), .A(n8341), .ZN(n8681) );
  INV_X4 U9189 ( .A(n8681), .ZN(n8348) );
  OAI21_X4 U9190 ( .B1(instructionAddr_out[26]), .B2(n8344), .A(n8343), .ZN(
        n8346) );
  INV_X4 U9191 ( .A(\PCLOGIC/imm16_32 [26]), .ZN(n8345) );
  XNOR2_X2 U9192 ( .A(n8346), .B(n8345), .ZN(n8680) );
  INV_X4 U9193 ( .A(n8346), .ZN(n9791) );
  NAND2_X2 U9194 ( .A1(n9791), .A2(\PCLOGIC/imm16_32 [26]), .ZN(n8347) );
  OAI21_X4 U9195 ( .B1(n8348), .B2(n8680), .A(n8347), .ZN(n8970) );
  NAND2_X2 U9196 ( .A1(n8349), .A2(n8970), .ZN(n8969) );
  INV_X4 U9197 ( .A(n8969), .ZN(n8350) );
  AOI21_X4 U9198 ( .B1(n9000), .B2(\PCLOGIC/imm16_32 [25]), .A(n8350), .ZN(
        n8528) );
  XNOR2_X2 U9199 ( .A(n8530), .B(n8351), .ZN(n8529) );
  OAI22_X2 U9200 ( .A1(n8352), .A2(n8530), .B1(n8528), .B2(n8529), .ZN(n9285)
         );
  NAND2_X2 U9201 ( .A1(n8353), .A2(n9285), .ZN(n9284) );
  INV_X4 U9202 ( .A(n9284), .ZN(n8354) );
  AOI21_X4 U9203 ( .B1(n9316), .B2(\PCLOGIC/imm16_32 [23]), .A(n8354), .ZN(
        n8963) );
  XNOR2_X2 U9204 ( .A(n8950), .B(n8355), .ZN(n8962) );
  OAI22_X2 U9205 ( .A1(n8356), .A2(n8950), .B1(n8963), .B2(n8962), .ZN(n9538)
         );
  NAND2_X2 U9206 ( .A1(n8357), .A2(n9538), .ZN(n9537) );
  INV_X4 U9207 ( .A(n9537), .ZN(n8358) );
  AOI21_X4 U9208 ( .B1(n9569), .B2(\PCLOGIC/imm16_32 [21]), .A(n8358), .ZN(
        n9278) );
  INV_X4 U9209 ( .A(\PCLOGIC/imm16_32 [20]), .ZN(net73512) );
  XNOR2_X2 U9210 ( .A(n9279), .B(net73512), .ZN(n9277) );
  OAI22_X2 U9211 ( .A1(net73512), .A2(n9279), .B1(n9278), .B2(n9277), .ZN(
        n9271) );
  NAND2_X2 U9212 ( .A1(n4968), .A2(n9271), .ZN(n9272) );
  INV_X4 U9213 ( .A(n9272), .ZN(n8359) );
  AOI21_X4 U9214 ( .B1(n10003), .B2(\PCLOGIC/imm16_32 [19]), .A(n8359), .ZN(
        n8803) );
  INV_X4 U9215 ( .A(\PCLOGIC/imm16_32 [18]), .ZN(net73529) );
  XNOR2_X2 U9216 ( .A(n8804), .B(net73529), .ZN(n8802) );
  OAI22_X2 U9217 ( .A1(net73529), .A2(n8804), .B1(n8803), .B2(n8802), .ZN(
        n8798) );
  NAND2_X2 U9218 ( .A1(n8360), .A2(n8798), .ZN(n8797) );
  INV_X4 U9219 ( .A(n8797), .ZN(n8361) );
  AOI21_X4 U9220 ( .B1(n9041), .B2(\PCLOGIC/imm16_32 [17]), .A(n8361), .ZN(
        n8511) );
  XNOR2_X2 U9221 ( .A(n8512), .B(net73908), .ZN(n8510) );
  OAI22_X2 U9222 ( .A1(net73908), .A2(n8512), .B1(n8511), .B2(n8510), .ZN(
        n8506) );
  INV_X4 U9223 ( .A(n8362), .ZN(n8363) );
  AOI21_X4 U9224 ( .B1(n8364), .B2(n5064), .A(n8363), .ZN(n10294) );
  XNOR2_X2 U9225 ( .A(net73902), .B(n10294), .ZN(n8507) );
  INV_X4 U9226 ( .A(n8507), .ZN(n8365) );
  AOI22_X2 U9227 ( .A1(n8506), .A2(n8365), .B1(net73902), .B2(n10294), .ZN(
        n8503) );
  NAND2_X2 U9228 ( .A1(net73900), .A2(n10261), .ZN(n8366) );
  INV_X4 U9229 ( .A(n9388), .ZN(n8371) );
  INV_X4 U9230 ( .A(n8367), .ZN(n8369) );
  INV_X4 U9231 ( .A(n8368), .ZN(n9422) );
  NAND2_X2 U9232 ( .A1(n8369), .A2(n9422), .ZN(n8370) );
  OAI21_X4 U9233 ( .B1(n9389), .B2(n8371), .A(n8370), .ZN(n8521) );
  XNOR2_X2 U9234 ( .A(n9107), .B(n8372), .ZN(n8520) );
  NAND2_X2 U9235 ( .A1(n8521), .A2(n8522), .ZN(n8523) );
  INV_X4 U9236 ( .A(n8373), .ZN(n8517) );
  NAND2_X2 U9237 ( .A1(n8374), .A2(n9864), .ZN(n8375) );
  OAI21_X4 U9238 ( .B1(n8516), .B2(n8517), .A(n8375), .ZN(n9384) );
  INV_X4 U9239 ( .A(n8376), .ZN(n10139) );
  XNOR2_X2 U9240 ( .A(n4921), .B(n10139), .ZN(n8377) );
  INV_X4 U9241 ( .A(n8377), .ZN(n9385) );
  AOI22_X2 U9242 ( .A1(n4921), .A2(n10139), .B1(n9384), .B2(n9385), .ZN(n8498)
         );
  OAI22_X2 U9243 ( .A1(n8499), .A2(n8378), .B1(n8497), .B2(n8498), .ZN(n9529)
         );
  XNOR2_X2 U9244 ( .A(n8379), .B(n4909), .ZN(n8382) );
  NAND2_X2 U9245 ( .A1(n8380), .A2(net73877), .ZN(n8381) );
  XNOR2_X2 U9246 ( .A(n8382), .B(n8381), .ZN(n9530) );
  INV_X4 U9247 ( .A(n9530), .ZN(n8384) );
  INV_X4 U9248 ( .A(n8381), .ZN(n8383) );
  INV_X4 U9249 ( .A(n8382), .ZN(n9531) );
  AOI22_X2 U9250 ( .A1(n9529), .A2(n8384), .B1(n8383), .B2(n9531), .ZN(n8494)
         );
  NAND2_X2 U9251 ( .A1(n8385), .A2(n9700), .ZN(n8386) );
  XNOR2_X2 U9252 ( .A(net73858), .B(n9671), .ZN(n8387) );
  INV_X4 U9253 ( .A(n8387), .ZN(n8488) );
  NAND2_X2 U9254 ( .A1(n8487), .A2(n8488), .ZN(n8489) );
  NAND2_X2 U9255 ( .A1(n8388), .A2(n8489), .ZN(n8483) );
  AOI21_X4 U9256 ( .B1(n8389), .B2(instructionAddr_out[6]), .A(
        instructionAddr_out[5]), .ZN(n8390) );
  INV_X4 U9257 ( .A(n8390), .ZN(n8392) );
  NAND2_X2 U9258 ( .A1(n8392), .A2(n8391), .ZN(n8393) );
  XNOR2_X2 U9259 ( .A(n8393), .B(net70531), .ZN(n8484) );
  INV_X4 U9260 ( .A(n8484), .ZN(n8394) );
  INV_X4 U9261 ( .A(n8393), .ZN(n9634) );
  AOI22_X2 U9262 ( .A1(n8483), .A2(n8394), .B1(n9634), .B2(net73858), .ZN(
        n8480) );
  NAND2_X2 U9263 ( .A1(n9965), .A2(net73858), .ZN(n8395) );
  XNOR2_X2 U9264 ( .A(net73858), .B(n10043), .ZN(n8396) );
  INV_X4 U9265 ( .A(n8396), .ZN(n8474) );
  NAND2_X2 U9266 ( .A1(n8473), .A2(n8474), .ZN(n8475) );
  NAND2_X2 U9267 ( .A1(n8397), .A2(n8475), .ZN(n8469) );
  INV_X4 U9268 ( .A(n8469), .ZN(n8399) );
  NAND2_X2 U9269 ( .A1(net71396), .A2(net73858), .ZN(n8398) );
  OAI21_X4 U9270 ( .B1(n8470), .B2(n8399), .A(n8398), .ZN(n8462) );
  INV_X4 U9271 ( .A(n10650), .ZN(n8464) );
  INV_X4 U9272 ( .A(net73842), .ZN(net73838) );
  INV_X4 U9273 ( .A(n8409), .ZN(n8411) );
  NAND4_X2 U9274 ( .A1(n8415), .A2(n8414), .A3(n8413), .A4(n8412), .ZN(n8459)
         );
  NAND4_X2 U9275 ( .A1(n8429), .A2(n8428), .A3(n8427), .A4(n8426), .ZN(n8458)
         );
  NAND4_X2 U9276 ( .A1(n8442), .A2(n8441), .A3(n8440), .A4(n8439), .ZN(n8457)
         );
  NOR4_X2 U9277 ( .A1(n8446), .A2(n8445), .A3(n8444), .A4(n8443), .ZN(n8455)
         );
  INV_X4 U9278 ( .A(n8447), .ZN(n8454) );
  NAND4_X2 U9279 ( .A1(n8455), .A2(n8454), .A3(n8453), .A4(n8452), .ZN(n8456)
         );
  NOR4_X2 U9280 ( .A1(n8459), .A2(n8458), .A3(n8457), .A4(n8456), .ZN(n8460)
         );
  XNOR2_X2 U9281 ( .A(n8460), .B(instruction[5]), .ZN(n8461) );
  NAND2_X2 U9282 ( .A1(n8462), .A2(net73855), .ZN(n10640) );
  NAND2_X2 U9283 ( .A1(n10649), .A2(n10640), .ZN(n8467) );
  INV_X4 U9284 ( .A(n8463), .ZN(n8465) );
  NAND2_X2 U9285 ( .A1(n8465), .A2(n8464), .ZN(n8527) );
  NAND2_X2 U9286 ( .A1(n6190), .A2(n5592), .ZN(n8466) );
  OAI221_X2 U9287 ( .B1(net71273), .B2(n4962), .C1(n8468), .C2(n8467), .A(
        n8466), .ZN(\PCLOGIC/PC_REG/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  XOR2_X2 U9288 ( .A(n8470), .B(n8469), .Z(n8472) );
  NAND2_X2 U9289 ( .A1(n6190), .A2(net71396), .ZN(n8471) );
  OAI221_X2 U9290 ( .B1(n10109), .B2(n4962), .C1(n8472), .C2(n6008), .A(n8471), 
        .ZN(\PCLOGIC/PC_REG/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9291 ( .A1(n10649), .A2(n8475), .ZN(n8477) );
  NAND2_X2 U9292 ( .A1(n6190), .A2(n10043), .ZN(n8476) );
  OAI221_X2 U9293 ( .B1(n10404), .B2(n4962), .C1(n8478), .C2(n8477), .A(n8476), 
        .ZN(\PCLOGIC/PC_REG/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  XNOR2_X2 U9294 ( .A(n8480), .B(n8479), .ZN(n8482) );
  NAND2_X2 U9295 ( .A1(n6190), .A2(n9965), .ZN(n8481) );
  OAI221_X2 U9296 ( .B1(n9954), .B2(n4962), .C1(n6008), .C2(n8482), .A(n8481), 
        .ZN(\PCLOGIC/PC_REG/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  XOR2_X2 U9297 ( .A(n8484), .B(n8483), .Z(n8486) );
  NAND2_X2 U9298 ( .A1(n6190), .A2(n9634), .ZN(n8485) );
  OAI221_X2 U9299 ( .B1(n10396), .B2(n4962), .C1(n8486), .C2(n9533), .A(n8485), 
        .ZN(\PCLOGIC/PC_REG/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9300 ( .A1(n10649), .A2(n8489), .ZN(n8491) );
  NAND2_X2 U9301 ( .A1(n6190), .A2(n9671), .ZN(n8490) );
  OAI221_X2 U9302 ( .B1(n9656), .B2(n4962), .C1(n8492), .C2(n8491), .A(n8490), 
        .ZN(\PCLOGIC/PC_REG/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  XNOR2_X2 U9303 ( .A(n8494), .B(n8493), .ZN(n8496) );
  NAND2_X2 U9304 ( .A1(n6190), .A2(n9700), .ZN(n8495) );
  OAI221_X2 U9305 ( .B1(n10464), .B2(n4962), .C1(n9533), .C2(n8496), .A(n8495), 
        .ZN(\PCLOGIC/PC_REG/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  XNOR2_X2 U9306 ( .A(n8498), .B(n8497), .ZN(n8501) );
  INV_X4 U9307 ( .A(n8499), .ZN(n9375) );
  NAND2_X2 U9308 ( .A1(n6190), .A2(n9375), .ZN(n8500) );
  OAI221_X2 U9309 ( .B1(n10382), .B2(n4962), .C1(n6008), .C2(n8501), .A(n8500), 
        .ZN(\PCLOGIC/PC_REG/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  XNOR2_X2 U9310 ( .A(n8503), .B(n8502), .ZN(n8505) );
  NAND2_X2 U9311 ( .A1(n6190), .A2(n10261), .ZN(n8504) );
  OAI221_X2 U9312 ( .B1(n10247), .B2(n4962), .C1(n9533), .C2(n8505), .A(n8504), 
        .ZN(\PCLOGIC/PC_REG/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  XOR2_X2 U9313 ( .A(n8507), .B(n8506), .Z(n8509) );
  NAND2_X2 U9314 ( .A1(n6190), .A2(n10294), .ZN(n8508) );
  OAI221_X2 U9315 ( .B1(n10463), .B2(n4962), .C1(n8509), .C2(n6008), .A(n8508), 
        .ZN(\PCLOGIC/PC_REG/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  XNOR2_X2 U9316 ( .A(n8511), .B(n8510), .ZN(n8515) );
  INV_X4 U9317 ( .A(n8512), .ZN(n9203) );
  NAND2_X2 U9318 ( .A1(n6190), .A2(n9203), .ZN(n8514) );
  NAND2_X2 U9319 ( .A1(net73708), .A2(aluA[16]), .ZN(n8513) );
  OAI211_X2 U9320 ( .C1(n8515), .C2(n9533), .A(n8514), .B(n8513), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  XNOR2_X2 U9321 ( .A(n8517), .B(n8516), .ZN(n8519) );
  NAND2_X2 U9322 ( .A1(n6190), .A2(n9864), .ZN(n8518) );
  OAI221_X2 U9323 ( .B1(n10375), .B2(n4962), .C1(n6008), .C2(n8519), .A(n8518), 
        .ZN(\PCLOGIC/PC_REG/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9324 ( .A(n8520), .ZN(n8522) );
  NAND2_X2 U9325 ( .A1(n8523), .A2(n10649), .ZN(n8525) );
  INV_X4 U9326 ( .A(n4962), .ZN(net73708) );
  NAND2_X2 U9327 ( .A1(net73708), .A2(\WIRE_ALU_A/MUX2TO1_32BIT[12].MUX/N1 ), 
        .ZN(n8524) );
  OAI221_X2 U9328 ( .B1(n9107), .B2(n8527), .C1(n8526), .C2(n8525), .A(n8524), 
        .ZN(\PCLOGIC/PC_REG/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  XNOR2_X2 U9329 ( .A(n8529), .B(n8528), .ZN(n8533) );
  NAND2_X2 U9330 ( .A1(net73708), .A2(net36391), .ZN(n8532) );
  INV_X4 U9331 ( .A(n8530), .ZN(n8664) );
  NAND2_X2 U9332 ( .A1(n6190), .A2(n8664), .ZN(n8531) );
  OAI211_X2 U9333 ( .C1(n8533), .C2(n6008), .A(n8532), .B(n8531), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9335 ( .A(net73620), .ZN(net73684) );
  INV_X4 U9336 ( .A(net73695), .ZN(net73638) );
  NAND2_X2 U9337 ( .A1(net73638), .A2(net73619), .ZN(n8558) );
  INV_X4 U9338 ( .A(instruction[4]), .ZN(net73694) );
  NAND2_X2 U9339 ( .A1(n8576), .A2(net73694), .ZN(n8557) );
  INV_X4 U9340 ( .A(n8565), .ZN(n8576) );
  INV_X4 U9341 ( .A(\PCLOGIC/imm16_32 [31]), .ZN(net73652) );
  NAND3_X2 U9342 ( .A1(net73638), .A2(net73652), .A3(net73619), .ZN(n8534) );
  NAND2_X2 U9343 ( .A1(n8535), .A2(n8534), .ZN(n8582) );
  INV_X4 U9344 ( .A(n8582), .ZN(n8548) );
  NAND2_X2 U9345 ( .A1(instruction[4]), .A2(net73503), .ZN(n8655) );
  INV_X4 U9346 ( .A(n8655), .ZN(n8536) );
  NAND2_X2 U9347 ( .A1(n8536), .A2(instruction[3]), .ZN(n8538) );
  NAND2_X2 U9348 ( .A1(\PCLOGIC/imm16_32 [30]), .A2(net73652), .ZN(net73630)
         );
  NAND4_X2 U9349 ( .A1(net73646), .A2(\PCLOGIC/imm16_32 [29]), .A3(net73670), 
        .A4(net73684), .ZN(n8537) );
  OAI21_X4 U9350 ( .B1(net73622), .B2(n8538), .A(n8537), .ZN(n8574) );
  INV_X4 U9351 ( .A(n8574), .ZN(n8547) );
  NAND3_X4 U9352 ( .A1(n8539), .A2(instruction[3]), .A3(net73498), .ZN(n8540)
         );
  INV_X4 U9353 ( .A(n8540), .ZN(n8564) );
  NAND3_X2 U9354 ( .A1(n4967), .A2(\PCLOGIC/imm16_32 [31]), .A3(net73670), 
        .ZN(n8541) );
  NAND2_X2 U9355 ( .A1(n8542), .A2(n8541), .ZN(n8543) );
  INV_X4 U9356 ( .A(n8543), .ZN(n8579) );
  NOR2_X4 U9357 ( .A1(\PCLOGIC/imm16_32 [26]), .A2(\PCLOGIC/imm16_32 [27]), 
        .ZN(n8544) );
  NAND4_X2 U9358 ( .A1(net73509), .A2(\PCLOGIC/imm16_32 [29]), .A3(net73670), 
        .A4(n8544), .ZN(n8563) );
  INV_X4 U9359 ( .A(n8563), .ZN(n8545) );
  NAND2_X2 U9360 ( .A1(instruction[1]), .A2(instruction[3]), .ZN(n8559) );
  NAND4_X2 U9361 ( .A1(n8548), .A2(n8547), .A3(n8579), .A4(n8546), .ZN(n8549)
         );
  INV_X4 U9362 ( .A(n8549), .ZN(n8572) );
  NAND3_X2 U9363 ( .A1(n4967), .A2(net73670), .A3(net73652), .ZN(n8550) );
  NAND2_X2 U9364 ( .A1(n8551), .A2(n8550), .ZN(n8575) );
  NAND2_X2 U9365 ( .A1(n8552), .A2(net73619), .ZN(n8555) );
  NAND3_X2 U9366 ( .A1(n8555), .A2(n8554), .A3(net77272), .ZN(n8581) );
  NAND4_X2 U9367 ( .A1(n8558), .A2(n8557), .A3(n8572), .A4(n8556), .ZN(
        net73543) );
  INV_X4 U9368 ( .A(net73543), .ZN(net70821) );
  NAND2_X2 U9369 ( .A1(\PCLOGIC/imm16_32 [31]), .A2(\PCLOGIC/imm16_32 [30]), 
        .ZN(n8562) );
  INV_X4 U9370 ( .A(n8559), .ZN(n8560) );
  NAND3_X2 U9371 ( .A1(n4966), .A2(instruction[5]), .A3(n8560), .ZN(n8561) );
  OAI21_X4 U9372 ( .B1(n8563), .B2(n8562), .A(n8561), .ZN(n8573) );
  INV_X4 U9373 ( .A(n8573), .ZN(n8571) );
  NAND2_X2 U9374 ( .A1(n4967), .A2(\PCLOGIC/imm16_32 [28]), .ZN(net73653) );
  INV_X4 U9375 ( .A(net73653), .ZN(net73616) );
  NAND2_X2 U9376 ( .A1(net73616), .A2(net73652), .ZN(n8570) );
  NAND2_X2 U9377 ( .A1(n8564), .A2(instruction[1]), .ZN(net73612) );
  INV_X4 U9378 ( .A(net73612), .ZN(net73637) );
  AOI21_X4 U9379 ( .B1(net73637), .B2(net73503), .A(n8566), .ZN(n8567) );
  INV_X4 U9380 ( .A(n8567), .ZN(n8568) );
  NOR3_X4 U9381 ( .A1(n8575), .A2(n8574), .A3(n8573), .ZN(net73611) );
  NAND4_X2 U9382 ( .A1(net73611), .A2(n8579), .A3(n8578), .A4(n8577), .ZN(
        net73541) );
  NOR2_X4 U9383 ( .A1(n8582), .A2(n8581), .ZN(net73613) );
  NOR2_X4 U9384 ( .A1(net73498), .A2(net73622), .ZN(net73615) );
  XNOR2_X2 U9385 ( .A(n10315), .B(net77042), .ZN(n8591) );
  INV_X4 U9386 ( .A(n8591), .ZN(n8593) );
  XNOR2_X2 U9387 ( .A(n10099), .B(net77042), .ZN(n8587) );
  INV_X4 U9388 ( .A(n9809), .ZN(n8590) );
  XNOR2_X2 U9389 ( .A(net71026), .B(net77042), .ZN(n8585) );
  XNOR2_X2 U9390 ( .A(n10928), .B(net77038), .ZN(n8584) );
  INV_X4 U9391 ( .A(n8583), .ZN(n10490) );
  OAI22_X2 U9392 ( .A1(net73608), .A2(n8584), .B1(net77042), .B2(n10490), .ZN(
        n8707) );
  INV_X4 U9393 ( .A(n8585), .ZN(n8586) );
  AOI22_X2 U9394 ( .A1(n8706), .A2(n8707), .B1(n8586), .B2(n5798), .ZN(n9810)
         );
  INV_X4 U9395 ( .A(n8587), .ZN(n8588) );
  OAI21_X4 U9396 ( .B1(n8590), .B2(n9810), .A(n8589), .ZN(n8772) );
  NAND2_X2 U9397 ( .A1(n8772), .A2(n8773), .ZN(n8771) );
  INV_X4 U9398 ( .A(n8771), .ZN(n8592) );
  XNOR2_X2 U9399 ( .A(n8594), .B(n5761), .ZN(n8883) );
  NAND2_X2 U9400 ( .A1(n8594), .A2(n5761), .ZN(n8595) );
  NAND2_X2 U9401 ( .A1(n9776), .A2(n9777), .ZN(n9774) );
  OAI21_X4 U9402 ( .B1(n8597), .B2(n8596), .A(n9774), .ZN(n8987) );
  INV_X4 U9403 ( .A(n8988), .ZN(n8598) );
  AOI22_X2 U9404 ( .A1(n8987), .A2(n8598), .B1(n10930), .B2(n4808), .ZN(n8809)
         );
  INV_X4 U9405 ( .A(n8808), .ZN(n8600) );
  XNOR2_X2 U9406 ( .A(n8809), .B(n8600), .ZN(n8603) );
  XNOR2_X2 U9407 ( .A(net36391), .B(n10331), .ZN(n10430) );
  NAND2_X2 U9408 ( .A1(n10494), .A2(net73541), .ZN(net70845) );
  NAND2_X2 U9409 ( .A1(multOut[24]), .A2(net81873), .ZN(n8648) );
  NAND2_X2 U9410 ( .A1(n10928), .A2(n10494), .ZN(n10474) );
  INV_X4 U9411 ( .A(n10474), .ZN(n8854) );
  INV_X4 U9412 ( .A(net73541), .ZN(net70826) );
  NAND2_X2 U9413 ( .A1(net77042), .A2(n10494), .ZN(n10304) );
  INV_X4 U9414 ( .A(n10494), .ZN(n10457) );
  NAND2_X2 U9415 ( .A1(n10457), .A2(net77040), .ZN(n8642) );
  NAND2_X2 U9416 ( .A1(n10304), .A2(n8642), .ZN(n10475) );
  NAND2_X2 U9417 ( .A1(net70826), .A2(n10475), .ZN(n8604) );
  MUX2_X2 U9418 ( .A(n8604), .B(net70845), .S(net70821), .Z(net72163) );
  NAND2_X2 U9419 ( .A1(n8854), .A2(net70697), .ZN(n9803) );
  NAND2_X2 U9420 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[5].MUX/N1 ), .A2(net70720), 
        .ZN(n8607) );
  INV_X4 U9421 ( .A(n9581), .ZN(n9330) );
  NAND2_X2 U9422 ( .A1(n10933), .A2(n6041), .ZN(n8821) );
  NAND2_X2 U9423 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[13].MUX/N1 ), .A2(n9065), 
        .ZN(n9597) );
  INV_X4 U9424 ( .A(n9597), .ZN(n8605) );
  NAND2_X2 U9425 ( .A1(net70534), .A2(net73541), .ZN(net71300) );
  NAND2_X2 U9426 ( .A1(net70719), .A2(net70696), .ZN(n8855) );
  INV_X4 U9427 ( .A(n8855), .ZN(n8624) );
  NOR2_X4 U9428 ( .A1(n8605), .A2(n8624), .ZN(n8606) );
  NAND3_X4 U9429 ( .A1(n8607), .A2(n8821), .A3(n8606), .ZN(n8977) );
  NAND2_X2 U9430 ( .A1(n10102), .A2(n8977), .ZN(n8619) );
  NAND2_X2 U9431 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[7].MUX/N1 ), .A2(net70720), 
        .ZN(n8610) );
  NAND2_X2 U9432 ( .A1(n10931), .A2(n6041), .ZN(n8826) );
  NAND2_X2 U9433 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[15].MUX/N1 ), .A2(n9065), 
        .ZN(n9593) );
  INV_X4 U9434 ( .A(n9593), .ZN(n8608) );
  NOR2_X4 U9435 ( .A1(n8608), .A2(n8624), .ZN(n8609) );
  NAND3_X4 U9436 ( .A1(n8610), .A2(n8826), .A3(n8609), .ZN(n8976) );
  NAND2_X2 U9437 ( .A1(net77086), .A2(n8976), .ZN(n8618) );
  NAND2_X2 U9438 ( .A1(n6040), .A2(aluA[19]), .ZN(n8828) );
  NAND2_X2 U9439 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[11].MUX/N1 ), .A2(n9065), 
        .ZN(n10018) );
  INV_X4 U9440 ( .A(n10018), .ZN(n8612) );
  NOR2_X4 U9441 ( .A1(n8612), .A2(n8611), .ZN(n8613) );
  NAND3_X4 U9442 ( .A1(n8855), .A2(n8828), .A3(n8613), .ZN(n9976) );
  NAND2_X2 U9443 ( .A1(n6040), .A2(aluA[17]), .ZN(n9017) );
  NAND2_X2 U9444 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[9].MUX/N1 ), .A2(n9065), .ZN(
        n10155) );
  INV_X4 U9445 ( .A(n10155), .ZN(n8615) );
  NOR2_X4 U9446 ( .A1(n8615), .A2(n8614), .ZN(n8616) );
  NAND3_X4 U9447 ( .A1(n8855), .A2(n9017), .A3(n8616), .ZN(n9975) );
  AOI22_X2 U9448 ( .A1(n6082), .A2(n9976), .B1(n6083), .B2(n9975), .ZN(n8617)
         );
  NAND2_X2 U9449 ( .A1(n10058), .A2(n9294), .ZN(n8633) );
  INV_X4 U9450 ( .A(n10928), .ZN(n10470) );
  INV_X4 U9451 ( .A(n10472), .ZN(n8861) );
  INV_X4 U9452 ( .A(n9854), .ZN(n10060) );
  NAND2_X2 U9453 ( .A1(n6040), .A2(aluA[18]), .ZN(n8842) );
  NAND2_X2 U9454 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[10].MUX/N1 ), .A2(n9065), 
        .ZN(n10095) );
  INV_X4 U9455 ( .A(n10095), .ZN(n8621) );
  NOR2_X4 U9456 ( .A1(n8621), .A2(n8620), .ZN(n8622) );
  NAND3_X4 U9457 ( .A1(n8855), .A2(n8842), .A3(n8622), .ZN(n9546) );
  NAND2_X2 U9458 ( .A1(n6083), .A2(n9546), .ZN(n8631) );
  NAND2_X2 U9459 ( .A1(n6040), .A2(aluA[20]), .ZN(n8836) );
  NAND2_X2 U9460 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[12].MUX/N1 ), .A2(n9065), 
        .ZN(n9938) );
  NAND3_X4 U9461 ( .A1(n8836), .A2(n9938), .A3(n8625), .ZN(n9547) );
  NAND2_X2 U9462 ( .A1(n6082), .A2(n9547), .ZN(n8630) );
  NAND2_X2 U9463 ( .A1(n10932), .A2(n6041), .ZN(n8840) );
  NAND2_X2 U9464 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[14].MUX/N1 ), .A2(n9065), 
        .ZN(n9617) );
  NAND2_X2 U9465 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[6].MUX/N1 ), .A2(net70720), 
        .ZN(n8626) );
  NAND4_X2 U9466 ( .A1(n8840), .A2(n9617), .A3(n8626), .A4(n8855), .ZN(n8928)
         );
  NAND2_X2 U9467 ( .A1(n8728), .A2(n8928), .ZN(n8629) );
  NAND2_X2 U9468 ( .A1(net36391), .A2(n6041), .ZN(n8637) );
  NAND2_X2 U9469 ( .A1(n9065), .A2(aluA[16]), .ZN(n9499) );
  AOI22_X2 U9470 ( .A1(net70719), .A2(net70534), .B1(net70720), .B2(
        \WIRE_ALU_A/MUX2TO1_32BIT[8].MUX/N1 ), .ZN(n8627) );
  NAND2_X2 U9471 ( .A1(net77084), .A2(n8892), .ZN(n8628) );
  NAND4_X2 U9472 ( .A1(n8631), .A2(n8630), .A3(n8629), .A4(n8628), .ZN(n8975)
         );
  NAND2_X2 U9473 ( .A1(n10060), .A2(n8975), .ZN(n8632) );
  NAND2_X2 U9474 ( .A1(n8633), .A2(n8632), .ZN(n8646) );
  NAND2_X2 U9475 ( .A1(n10457), .A2(n10928), .ZN(n9770) );
  INV_X4 U9476 ( .A(n9770), .ZN(n10303) );
  NAND2_X2 U9477 ( .A1(n6040), .A2(n6005), .ZN(n8823) );
  INV_X4 U9478 ( .A(n5761), .ZN(n10319) );
  NAND2_X2 U9479 ( .A1(n6040), .A2(n10099), .ZN(n8634) );
  NAND2_X2 U9480 ( .A1(n10064), .A2(n8974), .ZN(n8636) );
  NAND2_X2 U9481 ( .A1(n10457), .A2(n10470), .ZN(n9802) );
  NAND2_X2 U9482 ( .A1(n10066), .A2(n9297), .ZN(n8635) );
  NAND2_X2 U9483 ( .A1(n8636), .A2(n8635), .ZN(n8641) );
  NAND2_X2 U9484 ( .A1(n10930), .A2(n6041), .ZN(n8724) );
  OAI22_X2 U9485 ( .A1(n10312), .A2(n8823), .B1(n6005), .B2(n8724), .ZN(n9298)
         );
  NAND2_X2 U9486 ( .A1(n10064), .A2(n9298), .ZN(n8640) );
  OAI22_X2 U9487 ( .A1(n8638), .A2(n8823), .B1(n6005), .B2(n8637), .ZN(n9301)
         );
  NAND2_X2 U9488 ( .A1(n10066), .A2(n9301), .ZN(n8639) );
  NAND2_X2 U9489 ( .A1(n8640), .A2(n8639), .ZN(n8942) );
  MUX2_X2 U9490 ( .A(n8641), .B(n8942), .S(net71026), .Z(n8645) );
  INV_X4 U9491 ( .A(n8642), .ZN(n10491) );
  NAND2_X2 U9492 ( .A1(n10491), .A2(net73543), .ZN(n8643) );
  NAND2_X2 U9493 ( .A1(n8643), .A2(n10304), .ZN(net70706) );
  NAND3_X2 U9494 ( .A1(n8649), .A2(n8648), .A3(n8647), .ZN(dmem_addr_out[24])
         );
  MUX2_X2 U9495 ( .A(net88253), .B(n8650), .S(net73509), .Z(n8651) );
  NAND2_X2 U9496 ( .A1(n8651), .A2(net70738), .ZN(net73443) );
  NAND2_X2 U9497 ( .A1(net73527), .A2(net70738), .ZN(net73429) );
  MUX2_X2 U9498 ( .A(n4820), .B(net73908), .S(net73509), .Z(n8652) );
  NAND2_X2 U9499 ( .A1(n8652), .A2(net70738), .ZN(net73468) );
  NAND2_X2 U9500 ( .A1(instruction[0]), .A2(instruction[2]), .ZN(n8653) );
  NAND2_X2 U9501 ( .A1(net73510), .A2(net70738), .ZN(n8671) );
  INV_X4 U9502 ( .A(n8671), .ZN(n8669) );
  INV_X4 U9503 ( .A(\PCLOGIC/imm16_32 [19]), .ZN(n8656) );
  MUX2_X2 U9504 ( .A(net86793), .B(n8656), .S(net73509), .Z(n8657) );
  NAND2_X2 U9505 ( .A1(n8657), .A2(net70738), .ZN(n8670) );
  INV_X4 U9506 ( .A(n8670), .ZN(n8672) );
  INV_X4 U9507 ( .A(dmem_addr_out[24]), .ZN(n8667) );
  INV_X4 U9508 ( .A(n8870), .ZN(dmem_dsize[1]) );
  INV_X4 U9509 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [24]), .ZN(n9516) );
  NAND2_X2 U9510 ( .A1(n4899), .A2(n8870), .ZN(net70811) );
  INV_X4 U9511 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [16]), .ZN(n10540) );
  INV_X4 U9512 ( .A(dmem_read_in[24]), .ZN(n8662) );
  OAI211_X2 U9513 ( .C1(n8667), .C2(net76646), .A(n8666), .B(n8665), .ZN(n8668) );
  OAI22_X2 U9514 ( .A1(n5128), .A2(n6088), .B1(net76660), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9515 ( .A1(n8669), .A2(n8670), .ZN(net73436) );
  INV_X4 U9516 ( .A(net73436), .ZN(net73423) );
  NAND2_X2 U9517 ( .A1(net76270), .A2(n6156), .ZN(n10512) );
  OAI22_X2 U9518 ( .A1(n5253), .A2(n6091), .B1(n6156), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9519 ( .A1(n8670), .A2(n8671), .ZN(net73434) );
  INV_X4 U9520 ( .A(net73434), .ZN(net73421) );
  OAI22_X2 U9521 ( .A1(n6192), .A2(n5563), .B1(n6195), .B2(n8679), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9522 ( .A1(n6196), .A2(n5564), .B1(n6199), .B2(n8679), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9523 ( .A1(n8672), .A2(n8671), .ZN(net73439) );
  NAND2_X2 U9524 ( .A1(n4894), .A2(net73416), .ZN(n10516) );
  NAND2_X2 U9525 ( .A1(net76270), .A2(n10516), .ZN(n10517) );
  OAI22_X2 U9526 ( .A1(n4946), .A2(n6097), .B1(n6095), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9527 ( .A1(n4894), .A2(net73423), .ZN(n10519) );
  OAI22_X2 U9528 ( .A1(n5129), .A2(n6103), .B1(n6102), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9529 ( .A1(n4894), .A2(net73421), .ZN(n10521) );
  OAI22_X2 U9530 ( .A1(n4947), .A2(n6108), .B1(n6106), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9531 ( .A1(n5130), .A2(n6112), .B1(n6158), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9532 ( .A1(n5131), .A2(n6115), .B1(n6160), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9533 ( .A1(n5254), .A2(n6118), .B1(n6162), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9534 ( .A1(n6200), .A2(n5363), .B1(n6204), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9535 ( .A1(n5255), .A2(net76862), .B1(net76616), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9536 ( .A1(n6205), .A2(n5398), .B1(n6208), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9537 ( .A1(n5132), .A2(n6121), .B1(n6164), .B2(n8679), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9538 ( .A1(n5256), .A2(n6124), .B1(n6166), .B2(n8679), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9539 ( .A1(n5133), .A2(n6127), .B1(n6168), .B2(n8679), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9540 ( .A1(n5134), .A2(n6129), .B1(n6170), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9541 ( .A1(n5257), .A2(n6132), .B1(n6172), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9542 ( .A1(n5135), .A2(n6136), .B1(n6174), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9543 ( .A1(n6209), .A2(n5399), .B1(n6212), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9544 ( .A(n8677), .ZN(n8673) );
  NAND2_X2 U9545 ( .A1(\REGFILE/reg_out[28][24] ), .A2(n6177), .ZN(n8674) );
  OAI21_X4 U9546 ( .B1(n6213), .B2(n6021), .A(n8674), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9547 ( .A(n10607), .ZN(n10532) );
  NAND2_X2 U9548 ( .A1(n6178), .A2(\REGFILE/reg_out[29][24] ), .ZN(n8675) );
  OAI21_X4 U9549 ( .B1(n6138), .B2(n6021), .A(n8675), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9550 ( .A1(n5258), .A2(n6139), .B1(net76550), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9551 ( .A(n10614), .ZN(n10534) );
  NAND2_X2 U9552 ( .A1(n6180), .A2(\REGFILE/reg_out[30][24] ), .ZN(n8676) );
  OAI21_X4 U9553 ( .B1(n6142), .B2(n6021), .A(n8676), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9554 ( .A(net70574), .ZN(net70509) );
  NAND2_X2 U9555 ( .A1(net76488), .A2(\REGFILE/reg_out[31][24] ), .ZN(n8678)
         );
  OAI21_X4 U9556 ( .B1(net76480), .B2(n6021), .A(n8678), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9557 ( .A1(n6215), .A2(n5400), .B1(net76320), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9558 ( .A1(n6217), .A2(n5364), .B1(n6220), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9559 ( .A1(n5259), .A2(n6144), .B1(n6183), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9560 ( .A1(net73423), .A2(n4895), .ZN(n10535) );
  OAI22_X2 U9561 ( .A1(n5260), .A2(net76706), .B1(n6147), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9562 ( .A1(n5136), .A2(net76692), .B1(n6185), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9563 ( .A1(n5261), .A2(n6150), .B1(n6187), .B2(n6021), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9564 ( .A1(n5137), .A2(n6153), .B1(n6189), .B2(n8679), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[24].REGISTER1/STORE_DATA/N3 ) );
  XOR2_X2 U9565 ( .A(n8681), .B(n8680), .Z(n8684) );
  NAND2_X2 U9566 ( .A1(n6190), .A2(n9791), .ZN(n8682) );
  OAI211_X2 U9567 ( .C1(n8684), .C2(n9533), .A(n8683), .B(n8682), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  XOR2_X2 U9568 ( .A(n8686), .B(n8685), .Z(n8689) );
  NAND2_X2 U9569 ( .A1(net73708), .A2(n5761), .ZN(n8688) );
  NAND2_X2 U9570 ( .A1(n6190), .A2(n8908), .ZN(n8687) );
  OAI211_X2 U9571 ( .C1(n8689), .C2(n6008), .A(n8688), .B(n8687), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI211_X2 U9572 ( .C1(n8335), .C2(net73400), .A(n8691), .B(n10649), .ZN(
        n8693) );
  NAND2_X2 U9573 ( .A1(n6190), .A2(n8788), .ZN(n8692) );
  XOR2_X2 U9574 ( .A(net73394), .B(net73395), .Z(n8697) );
  NAND2_X2 U9575 ( .A1(n6190), .A2(n5016), .ZN(n8695) );
  OAI211_X2 U9576 ( .C1(n8697), .C2(n9533), .A(n8696), .B(n8695), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9578 ( .A1(n6190), .A2(instructionAddr_out[30]), .ZN(n8705) );
  NAND2_X2 U9579 ( .A1(n8700), .A2(n8699), .ZN(n8701) );
  XOR2_X2 U9580 ( .A(n8707), .B(n8706), .Z(n8719) );
  NAND2_X2 U9581 ( .A1(net77084), .A2(n6041), .ZN(n10159) );
  INV_X4 U9582 ( .A(n10159), .ZN(n10542) );
  NAND2_X2 U9583 ( .A1(n10542), .A2(n5798), .ZN(n9805) );
  NAND2_X2 U9584 ( .A1(n10932), .A2(n9065), .ZN(n9076) );
  OAI21_X4 U9585 ( .B1(n8709), .B2(n8708), .A(net77084), .ZN(n8717) );
  NAND2_X2 U9586 ( .A1(n9065), .A2(aluA[20]), .ZN(n9079) );
  AOI22_X2 U9587 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[4].MUX/N1 ), .A2(net70719), 
        .B1(\WIRE_ALU_A/MUX2TO1_32BIT[12].MUX/N1 ), .B2(net70720), .ZN(n8710)
         );
  NAND3_X2 U9588 ( .A1(n9079), .A2(n8711), .A3(n8710), .ZN(n8712) );
  MUX2_X2 U9589 ( .A(n8892), .B(n8712), .S(n10099), .Z(n8758) );
  NAND2_X2 U9590 ( .A1(n8758), .A2(net78051), .ZN(n8716) );
  NAND2_X2 U9591 ( .A1(n9065), .A2(aluA[18]), .ZN(n9360) );
  AOI22_X2 U9592 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[2].MUX/N1 ), .A2(net70719), 
        .B1(\WIRE_ALU_A/MUX2TO1_32BIT[10].MUX/N1 ), .B2(net70720), .ZN(n8713)
         );
  NAND3_X4 U9593 ( .A1(n9360), .A2(n8714), .A3(n8713), .ZN(n8891) );
  NAND2_X2 U9594 ( .A1(n6081), .A2(n8891), .ZN(n8715) );
  AOI21_X4 U9595 ( .B1(n4910), .B2(n8719), .A(n8718), .ZN(n8734) );
  XNOR2_X2 U9596 ( .A(n5798), .B(net78051), .ZN(n10433) );
  INV_X4 U9597 ( .A(n10433), .ZN(n10310) );
  NAND2_X2 U9598 ( .A1(net70701), .A2(n10310), .ZN(n8733) );
  INV_X4 U9599 ( .A(n10094), .ZN(n8728) );
  NAND2_X2 U9600 ( .A1(n6040), .A2(n5761), .ZN(n8722) );
  NAND2_X2 U9601 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[11].MUX/N1 ), .A2(net70720), 
        .ZN(n8721) );
  NAND2_X2 U9602 ( .A1(n9065), .A2(aluA[19]), .ZN(n9340) );
  NAND2_X2 U9603 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[3].MUX/N1 ), .A2(net70719), 
        .ZN(n8720) );
  NAND4_X2 U9604 ( .A1(n8722), .A2(n8721), .A3(n9340), .A4(n8720), .ZN(n10466)
         );
  NAND2_X2 U9605 ( .A1(n9065), .A2(aluA[17]), .ZN(n9343) );
  AOI22_X2 U9606 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[1].MUX/N1 ), .A2(net70719), 
        .B1(\WIRE_ALU_A/MUX2TO1_32BIT[9].MUX/N1 ), .B2(net70720), .ZN(n8723)
         );
  NAND2_X2 U9607 ( .A1(n10933), .A2(n9065), .ZN(n9068) );
  AOI22_X2 U9608 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[5].MUX/N1 ), .A2(net70719), 
        .B1(\WIRE_ALU_A/MUX2TO1_32BIT[13].MUX/N1 ), .B2(net70720), .ZN(n8725)
         );
  NAND3_X2 U9609 ( .A1(n9068), .A2(n8726), .A3(n8725), .ZN(n8727) );
  MUX2_X2 U9610 ( .A(n8978), .B(n8727), .S(n10099), .Z(n10465) );
  NAND2_X2 U9611 ( .A1(n8854), .A2(net70697), .ZN(n9012) );
  OAI22_X2 U9612 ( .A1(n9801), .A2(n9012), .B1(n9606), .B2(n9805), .ZN(n8731)
         );
  NOR3_X4 U9613 ( .A1(n8731), .A2(n8730), .A3(n5062), .ZN(n8732) );
  MUX2_X2 U9614 ( .A(n8735), .B(multOut[30]), .S(net76452), .Z(
        dmem_addr_out[30]) );
  INV_X4 U9615 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [22]), .ZN(n9669) );
  INV_X4 U9616 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [30]), .ZN(n10259) );
  OAI22_X2 U9617 ( .A1(net70811), .A2(n9669), .B1(net77999), .B2(n10259), .ZN(
        n8736) );
  AOI21_X4 U9618 ( .B1(net76650), .B2(dmem_addr_out[30]), .A(n8736), .ZN(n8741) );
  INV_X4 U9619 ( .A(dmem_read_in[30]), .ZN(n8737) );
  NAND2_X2 U9620 ( .A1(n8741), .A2(n8740), .ZN(n8742) );
  OAI22_X2 U9621 ( .A1(n4975), .A2(n6088), .B1(n6223), .B2(net76658), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9622 ( .A(\REGFILE/reg_out[10][30] ), .ZN(n8743) );
  OAI22_X2 U9623 ( .A1(n8743), .A2(n6091), .B1(n6223), .B2(n6155), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9624 ( .A1(n5958), .A2(n6097), .B1(n6223), .B2(n6094), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9625 ( .A(\REGFILE/reg_out[14][30] ), .ZN(n8744) );
  OAI22_X2 U9626 ( .A1(n8744), .A2(n6103), .B1(n6223), .B2(n6102), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9627 ( .A1(n5918), .A2(n6108), .B1(n6223), .B2(n6105), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9628 ( .A1(n8745), .A2(n6112), .B1(n6223), .B2(n6157), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9629 ( .A(\REGFILE/reg_out[17][30] ), .ZN(n8746) );
  OAI22_X2 U9630 ( .A1(n8746), .A2(n6115), .B1(n6223), .B2(n6159), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9631 ( .A(\REGFILE/reg_out[18][30] ), .ZN(n8747) );
  OAI22_X2 U9632 ( .A1(n8747), .A2(n6118), .B1(n6223), .B2(n6161), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9633 ( .A1(n5124), .A2(net76862), .B1(n6223), .B2(net76614), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9634 ( .A(\REGFILE/reg_out[21][30] ), .ZN(n8748) );
  OAI22_X2 U9635 ( .A1(n8748), .A2(n6121), .B1(n6223), .B2(n6163), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9636 ( .A(\REGFILE/reg_out[22][30] ), .ZN(n8749) );
  OAI22_X2 U9637 ( .A1(n8749), .A2(n6124), .B1(n6223), .B2(n6165), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9638 ( .A(\REGFILE/reg_out[23][30] ), .ZN(n8750) );
  OAI22_X2 U9639 ( .A1(n8750), .A2(n6127), .B1(n6223), .B2(n6167), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9640 ( .A(\REGFILE/reg_out[24][30] ), .ZN(n8751) );
  OAI22_X2 U9641 ( .A1(n8751), .A2(n6129), .B1(n6223), .B2(n6169), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9642 ( .A1(n5924), .A2(n6132), .B1(n6223), .B2(n6171), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9643 ( .A(\REGFILE/reg_out[26][30] ), .ZN(n8752) );
  OAI22_X2 U9644 ( .A1(n8752), .A2(n6136), .B1(n6223), .B2(n6173), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9645 ( .A1(n6178), .A2(\REGFILE/reg_out[29][30] ), .ZN(n8753) );
  OAI22_X2 U9646 ( .A1(n5680), .A2(n6139), .B1(n6223), .B2(net76548), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9647 ( .A1(n5070), .A2(n6144), .B1(n6223), .B2(n6182), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9648 ( .A1(n5440), .A2(net76706), .B1(n6223), .B2(n6146), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9649 ( .A1(n5507), .A2(net76692), .B1(n6223), .B2(n6184), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9650 ( .A1(n8756), .A2(n6150), .B1(n6223), .B2(n6186), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9651 ( .A1(n8757), .A2(n6153), .B1(n6223), .B2(n6188), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9652 ( .A1(multOut[28]), .A2(net92392), .ZN(n8783) );
  INV_X4 U9653 ( .A(n10094), .ZN(n8759) );
  NAND2_X2 U9654 ( .A1(net77084), .A2(n10466), .ZN(n8763) );
  NAND2_X2 U9655 ( .A1(n8759), .A2(n8978), .ZN(n8762) );
  NAND2_X2 U9656 ( .A1(n6083), .A2(n8977), .ZN(n8761) );
  NAND2_X2 U9657 ( .A1(n6082), .A2(n8976), .ZN(n8760) );
  NAND4_X2 U9658 ( .A1(n8763), .A2(n8762), .A3(n8761), .A4(n8760), .ZN(n8890)
         );
  NAND2_X2 U9659 ( .A1(n8854), .A2(n8890), .ZN(n8764) );
  OAI22_X2 U9660 ( .A1(n4896), .A2(n9802), .B1(n4922), .B2(n9770), .ZN(n8769)
         );
  INV_X4 U9661 ( .A(n8772), .ZN(n8775) );
  INV_X4 U9662 ( .A(n8773), .ZN(n8774) );
  NAND2_X2 U9663 ( .A1(n8775), .A2(n8774), .ZN(n8779) );
  INV_X4 U9664 ( .A(n10441), .ZN(n10317) );
  NAND2_X2 U9665 ( .A1(net70701), .A2(n10317), .ZN(n8777) );
  NAND2_X2 U9666 ( .A1(n8777), .A2(n8776), .ZN(n8778) );
  AOI21_X4 U9667 ( .B1(n8780), .B2(n8779), .A(n8778), .ZN(n8781) );
  NAND3_X2 U9668 ( .A1(n8783), .A2(n8782), .A3(n8781), .ZN(dmem_addr_out[28])
         );
  INV_X4 U9669 ( .A(dmem_addr_out[28]), .ZN(n8791) );
  INV_X4 U9670 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [28]), .ZN(n9108) );
  INV_X4 U9671 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [20]), .ZN(n10083) );
  INV_X4 U9672 ( .A(dmem_read_in[28]), .ZN(n8786) );
  OAI211_X2 U9673 ( .C1(n8791), .C2(net76646), .A(n8790), .B(n8789), .ZN(n8792) );
  OAI22_X2 U9674 ( .A1(n5047), .A2(n6088), .B1(n6221), .B2(net76658), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9675 ( .A1(n5484), .A2(n6091), .B1(n6221), .B2(n6155), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9676 ( .A1(n5494), .A2(n6097), .B1(n6221), .B2(n6094), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9677 ( .A1(n5491), .A2(n6103), .B1(n6221), .B2(n6102), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9678 ( .A1(n5485), .A2(n6108), .B1(n6221), .B2(n6105), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9679 ( .A1(n5568), .A2(n6112), .B1(n6221), .B2(n6157), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9680 ( .A1(n5544), .A2(n6115), .B1(n6221), .B2(n6159), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9681 ( .A1(n5486), .A2(n6118), .B1(n6221), .B2(n6161), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9682 ( .A1(n5357), .A2(net76862), .B1(n6221), .B2(net76614), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9683 ( .A1(n5069), .A2(n6121), .B1(n6221), .B2(n6163), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9684 ( .A1(n5495), .A2(n6124), .B1(n6221), .B2(n6165), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9685 ( .A1(n5351), .A2(n6127), .B1(n6221), .B2(n6167), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9686 ( .A1(n5569), .A2(n6129), .B1(n6221), .B2(n6169), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9687 ( .A1(n5487), .A2(n6132), .B1(n6221), .B2(n6171), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9688 ( .A1(n5545), .A2(n6136), .B1(n6221), .B2(n6173), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9689 ( .A1(n6178), .A2(\REGFILE/reg_out[29][28] ), .ZN(n8793) );
  OAI22_X2 U9690 ( .A1(n5488), .A2(n6139), .B1(n6221), .B2(net76548), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9691 ( .A1(n6180), .A2(\REGFILE/reg_out[30][28] ), .ZN(n8794) );
  NAND2_X2 U9692 ( .A1(net76488), .A2(\REGFILE/reg_out[31][28] ), .ZN(n8795)
         );
  OAI22_X2 U9693 ( .A1(n5358), .A2(n6144), .B1(n6221), .B2(n6182), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9694 ( .A1(n5565), .A2(net76706), .B1(n6221), .B2(n6146), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9695 ( .A1(n5546), .A2(net76692), .B1(n6221), .B2(n6184), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9696 ( .A1(n5032), .A2(n6150), .B1(n6221), .B2(n6186), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9697 ( .A1(n5547), .A2(n6153), .B1(n6221), .B2(n6188), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[28].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9698 ( .A1(net73708), .A2(aluA[17]), .ZN(n8801) );
  OAI211_X2 U9699 ( .C1(n8360), .C2(n8798), .A(n8797), .B(n10649), .ZN(n8800)
         );
  NAND2_X2 U9700 ( .A1(n6190), .A2(n9041), .ZN(n8799) );
  NAND3_X4 U9701 ( .A1(n8801), .A2(n8800), .A3(n8799), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  XNOR2_X2 U9702 ( .A(n8803), .B(n8802), .ZN(n8807) );
  INV_X4 U9703 ( .A(n8804), .ZN(n8873) );
  NAND2_X2 U9704 ( .A1(n6190), .A2(n8873), .ZN(n8806) );
  NAND2_X2 U9705 ( .A1(net73708), .A2(aluA[18]), .ZN(n8805) );
  OAI211_X2 U9706 ( .C1(n8807), .C2(n6008), .A(n8806), .B(n8805), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9707 ( .A(n10053), .ZN(n8818) );
  OAI22_X2 U9708 ( .A1(n8810), .A2(net72312), .B1(n8809), .B2(n8808), .ZN(
        n9289) );
  XNOR2_X2 U9709 ( .A(n10931), .B(n4814), .ZN(n9290) );
  INV_X4 U9710 ( .A(n9290), .ZN(n8811) );
  AOI22_X2 U9711 ( .A1(n9289), .A2(n8811), .B1(n10931), .B2(n4814), .ZN(n8920)
         );
  INV_X4 U9712 ( .A(n8813), .ZN(n8812) );
  XNOR2_X2 U9713 ( .A(n10932), .B(n8812), .ZN(n8918) );
  OAI22_X2 U9714 ( .A1(n8813), .A2(n8967), .B1(n8920), .B2(n8918), .ZN(n9542)
         );
  INV_X4 U9715 ( .A(n9543), .ZN(n8814) );
  AOI22_X2 U9716 ( .A1(n9542), .A2(n8814), .B1(n10933), .B2(n4810), .ZN(n10054) );
  AOI22_X2 U9717 ( .A1(n9992), .A2(n9993), .B1(n8820), .B2(aluA[19]), .ZN(
        n9033) );
  XNOR2_X2 U9718 ( .A(n9033), .B(n9028), .ZN(n8835) );
  NAND2_X2 U9719 ( .A1(n8822), .A2(n8821), .ZN(n10241) );
  INV_X4 U9720 ( .A(n10241), .ZN(n8825) );
  INV_X4 U9721 ( .A(n8823), .ZN(n8937) );
  NAND2_X2 U9722 ( .A1(n8937), .A2(n10930), .ZN(n8824) );
  OAI21_X4 U9723 ( .B1(n6005), .B2(n8825), .A(n8824), .ZN(n10063) );
  INV_X4 U9724 ( .A(n10063), .ZN(n8832) );
  NAND2_X2 U9725 ( .A1(n8827), .A2(n8826), .ZN(n9018) );
  NAND2_X2 U9726 ( .A1(n6082), .A2(n9018), .ZN(n8831) );
  NAND2_X2 U9727 ( .A1(n9065), .A2(n5761), .ZN(n8829) );
  NAND2_X2 U9728 ( .A1(n8829), .A2(n8828), .ZN(n10240) );
  NAND2_X2 U9729 ( .A1(net77084), .A2(n10240), .ZN(n8830) );
  OAI211_X2 U9730 ( .C1(net71026), .C2(n8832), .A(n8831), .B(n8830), .ZN(n9986) );
  INV_X4 U9731 ( .A(n9986), .ZN(n8833) );
  NAND2_X2 U9732 ( .A1(multOut[18]), .A2(net81873), .ZN(n8868) );
  NAND2_X2 U9733 ( .A1(n8837), .A2(n8836), .ZN(n9397) );
  INV_X4 U9734 ( .A(n9397), .ZN(n8839) );
  NAND2_X2 U9735 ( .A1(n8937), .A2(net36391), .ZN(n8838) );
  OAI21_X4 U9736 ( .B1(n6005), .B2(n8839), .A(n8838), .ZN(n10065) );
  INV_X4 U9737 ( .A(n10065), .ZN(n8846) );
  NAND2_X2 U9738 ( .A1(n8841), .A2(n8840), .ZN(n9183) );
  NAND2_X2 U9739 ( .A1(n6082), .A2(n9183), .ZN(n8845) );
  NAND2_X2 U9740 ( .A1(n8843), .A2(n8842), .ZN(n9396) );
  NAND2_X2 U9741 ( .A1(net77084), .A2(n9396), .ZN(n8844) );
  OAI211_X2 U9742 ( .C1(net71026), .C2(n8846), .A(n8845), .B(n8844), .ZN(n9010) );
  INV_X4 U9743 ( .A(n9010), .ZN(n8848) );
  INV_X4 U9744 ( .A(n10445), .ZN(n10354) );
  NAND2_X2 U9745 ( .A1(net70701), .A2(n10354), .ZN(n8847) );
  INV_X4 U9746 ( .A(aluA[18]), .ZN(n8849) );
  NAND2_X2 U9747 ( .A1(net77084), .A2(n9975), .ZN(n8853) );
  NAND2_X2 U9748 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[11].MUX/N1 ), .A2(n6041), 
        .ZN(n9341) );
  OAI211_X2 U9749 ( .C1(n9094), .C2(n10404), .A(n9093), .B(n9341), .ZN(n9408)
         );
  NAND2_X2 U9750 ( .A1(n6083), .A2(n9408), .ZN(n8852) );
  NAND2_X2 U9751 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[15].MUX/N1 ), .A2(n6041), 
        .ZN(n9066) );
  NAND2_X2 U9752 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[7].MUX/N1 ), .A2(n9065), .ZN(
        n8850) );
  NAND2_X2 U9753 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[13].MUX/N1 ), .A2(n6041), 
        .ZN(n9069) );
  OAI211_X2 U9754 ( .C1(n9094), .C2(n10396), .A(n9093), .B(n9069), .ZN(n9977)
         );
  AOI22_X2 U9755 ( .A1(n8728), .A2(n9978), .B1(n6081), .B2(n9977), .ZN(n8851)
         );
  NAND2_X2 U9756 ( .A1(n8854), .A2(n9011), .ZN(n8863) );
  NAND2_X2 U9757 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[14].MUX/N1 ), .A2(n6041), 
        .ZN(n9077) );
  OAI211_X2 U9758 ( .C1(n9094), .C2(n9656), .A(n9093), .B(n9077), .ZN(n10233)
         );
  NAND2_X2 U9759 ( .A1(n6081), .A2(n10233), .ZN(n8860) );
  NAND2_X2 U9760 ( .A1(n6040), .A2(aluA[16]), .ZN(n9082) );
  NAND2_X2 U9761 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[8].MUX/N1 ), .A2(n9065), .ZN(
        net70717) );
  NAND2_X2 U9762 ( .A1(net70720), .A2(net70534), .ZN(n8856) );
  NAND4_X2 U9763 ( .A1(n9082), .A2(net70717), .A3(n8856), .A4(n8855), .ZN(
        n9548) );
  NAND2_X2 U9764 ( .A1(n8728), .A2(n9548), .ZN(n8859) );
  NAND2_X2 U9765 ( .A1(net77084), .A2(n9546), .ZN(n8858) );
  NAND2_X2 U9766 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[12].MUX/N1 ), .A2(n6040), 
        .ZN(n9080) );
  OAI211_X2 U9767 ( .C1(n9094), .C2(n9954), .A(n9093), .B(n9080), .ZN(n10232)
         );
  NAND2_X2 U9768 ( .A1(n6083), .A2(n10232), .ZN(n8857) );
  NAND4_X2 U9769 ( .A1(n8860), .A2(n8859), .A3(n8858), .A4(n8857), .ZN(n9984)
         );
  NAND2_X2 U9770 ( .A1(n8861), .A2(n9984), .ZN(n8862) );
  NOR3_X4 U9771 ( .A1(n8866), .A2(n8865), .A3(n8864), .ZN(n8867) );
  NAND3_X2 U9772 ( .A1(n8869), .A2(n8868), .A3(n8867), .ZN(dmem_addr_out[18])
         );
  INV_X4 U9773 ( .A(dmem_addr_out[18]), .ZN(n8876) );
  INV_X4 U9774 ( .A(net70740), .ZN(net73167) );
  NAND2_X2 U9775 ( .A1(net73167), .A2(n8870), .ZN(n10079) );
  INV_X4 U9776 ( .A(n10079), .ZN(n10000) );
  INV_X4 U9777 ( .A(dmem_read_in[18]), .ZN(n8871) );
  OAI211_X2 U9778 ( .C1(n8876), .C2(net76646), .A(n8875), .B(n8874), .ZN(n8877) );
  NAND2_X2 U9779 ( .A1(net76270), .A2(n8877), .ZN(n8882) );
  OAI22_X2 U9780 ( .A1(n5088), .A2(n6088), .B1(net76660), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9781 ( .A1(n5886), .A2(n6091), .B1(n6156), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9782 ( .A1(n6192), .A2(n5115), .B1(n6195), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9783 ( .A1(n6196), .A2(n4980), .B1(n6199), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9784 ( .A1(n4925), .A2(n6097), .B1(n6095), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9785 ( .A1(n5089), .A2(n6103), .B1(n6102), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9786 ( .A1(n5878), .A2(n6108), .B1(n6106), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9787 ( .A1(n5138), .A2(n6112), .B1(n6158), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9788 ( .A1(n5139), .A2(n6115), .B1(n6160), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9789 ( .A1(n5262), .A2(n6118), .B1(n6162), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9790 ( .A1(n6200), .A2(n5365), .B1(n6204), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9791 ( .A1(n5263), .A2(net76862), .B1(net76616), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9792 ( .A1(n6205), .A2(n5401), .B1(n6208), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9793 ( .A1(n5140), .A2(n6121), .B1(n6164), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9794 ( .A1(n5071), .A2(n6124), .B1(n6166), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9795 ( .A1(n5090), .A2(n6127), .B1(n6168), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9796 ( .A1(n5141), .A2(n6129), .B1(n6170), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9797 ( .A1(n5857), .A2(n6132), .B1(n6172), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9798 ( .A1(n5142), .A2(n6136), .B1(n6174), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9799 ( .A1(n6209), .A2(n5913), .B1(n6212), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9800 ( .A1(\REGFILE/reg_out[28][18] ), .A2(n6177), .ZN(n8878) );
  NAND2_X2 U9801 ( .A1(n6178), .A2(\REGFILE/reg_out[29][18] ), .ZN(n8879) );
  OAI22_X2 U9802 ( .A1(n5785), .A2(n6139), .B1(net76550), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9803 ( .A1(n6180), .A2(\REGFILE/reg_out[30][18] ), .ZN(n8880) );
  NAND2_X2 U9804 ( .A1(net76488), .A2(\REGFILE/reg_out[31][18] ), .ZN(n8881)
         );
  OAI22_X2 U9805 ( .A1(n6215), .A2(n5685), .B1(net76320), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9806 ( .A1(n6217), .A2(n5366), .B1(n6220), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9807 ( .A1(n5030), .A2(n6144), .B1(n6183), .B2(n8882), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9808 ( .A1(n5264), .A2(net76706), .B1(n6147), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9809 ( .A1(n5143), .A2(net76692), .B1(n6185), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9810 ( .A1(n5072), .A2(n6150), .B1(n6187), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9811 ( .A1(n5091), .A2(n6153), .B1(n6189), .B2(n6023), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[18].REGISTER1/STORE_DATA/N3 ) );
  XOR2_X2 U9812 ( .A(n8884), .B(n8883), .Z(n8889) );
  NAND2_X2 U9813 ( .A1(net70701), .A2(n10436), .ZN(n8887) );
  NAND2_X2 U9814 ( .A1(n8887), .A2(n8886), .ZN(n8888) );
  INV_X4 U9815 ( .A(n8890), .ZN(n8898) );
  NAND2_X2 U9816 ( .A1(n6083), .A2(n9547), .ZN(n8896) );
  NAND2_X2 U9817 ( .A1(net77084), .A2(n8891), .ZN(n8895) );
  NAND2_X2 U9818 ( .A1(n6082), .A2(n8928), .ZN(n8894) );
  NAND2_X2 U9819 ( .A1(n8759), .A2(n8892), .ZN(n8893) );
  NAND4_X2 U9820 ( .A1(n8896), .A2(n8895), .A3(n8894), .A4(n8893), .ZN(n8897)
         );
  INV_X4 U9821 ( .A(n8897), .ZN(n9768) );
  OAI22_X2 U9822 ( .A1(n10472), .A2(n8898), .B1(n9768), .B2(n10474), .ZN(n8900) );
  OAI22_X2 U9823 ( .A1(n4896), .A2(n9770), .B1(n9771), .B2(n9802), .ZN(n8899)
         );
  NAND2_X2 U9824 ( .A1(multOut[27]), .A2(net92392), .ZN(n8901) );
  NAND3_X4 U9825 ( .A1(n8903), .A2(n8902), .A3(n8901), .ZN(dmem_addr_out[27])
         );
  INV_X4 U9826 ( .A(dmem_addr_out[27]), .ZN(n8911) );
  INV_X4 U9827 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [27]), .ZN(n9862) );
  INV_X4 U9828 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [19]), .ZN(n10041) );
  INV_X4 U9829 ( .A(dmem_read_in[27]), .ZN(n8906) );
  OAI211_X2 U9830 ( .C1(n8911), .C2(net76646), .A(n8910), .B(n8909), .ZN(n8912) );
  NAND2_X2 U9831 ( .A1(net76270), .A2(n8912), .ZN(n8917) );
  OAI22_X2 U9832 ( .A1(n5548), .A2(n6088), .B1(net76660), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9833 ( .A1(n5489), .A2(n6091), .B1(n6156), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9834 ( .A1(n6192), .A2(n5562), .B1(n6195), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9835 ( .A1(n6196), .A2(n5567), .B1(n6199), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9836 ( .A1(n4955), .A2(n6097), .B1(n6095), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9837 ( .A1(n5492), .A2(n6103), .B1(n6102), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9838 ( .A1(n4949), .A2(n6108), .B1(n6106), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9839 ( .A1(n5493), .A2(n6112), .B1(n6158), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9840 ( .A1(n5549), .A2(n6115), .B1(n6160), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9841 ( .A1(n5490), .A2(n6118), .B1(n6162), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9842 ( .A1(n6200), .A2(n5432), .B1(n6204), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9843 ( .A1(n5359), .A2(net76862), .B1(net76616), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9844 ( .A1(n6205), .A2(n5434), .B1(n6208), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9845 ( .A1(n5352), .A2(n6121), .B1(n6164), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9846 ( .A1(n5496), .A2(n6124), .B1(n6166), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9847 ( .A1(n5353), .A2(n6127), .B1(n6168), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9848 ( .A1(n5354), .A2(n6129), .B1(n6170), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9849 ( .A1(n5360), .A2(n6132), .B1(n6172), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9850 ( .A1(n5355), .A2(n6136), .B1(n6174), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9851 ( .A1(n6209), .A2(n5435), .B1(n6212), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9852 ( .A1(\REGFILE/reg_out[28][27] ), .A2(n6177), .ZN(n8913) );
  NAND2_X2 U9853 ( .A1(n6178), .A2(\REGFILE/reg_out[29][27] ), .ZN(n8914) );
  OAI22_X2 U9854 ( .A1(n5361), .A2(n6139), .B1(net76550), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9855 ( .A1(n6180), .A2(\REGFILE/reg_out[30][27] ), .ZN(n8915) );
  NAND2_X2 U9856 ( .A1(net76488), .A2(\REGFILE/reg_out[31][27] ), .ZN(n8916)
         );
  OAI22_X2 U9857 ( .A1(n6215), .A2(n5436), .B1(net76320), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9858 ( .A1(n6217), .A2(n5542), .B1(n6220), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9859 ( .A1(n5497), .A2(n6144), .B1(n6183), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9860 ( .A1(n5566), .A2(net76706), .B1(n6147), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9861 ( .A1(n5550), .A2(net76692), .B1(n6185), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9862 ( .A1(n5362), .A2(n6150), .B1(n6187), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9863 ( .A1(n5356), .A2(n6153), .B1(n6189), .B2(n6025), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U9864 ( .A(n8918), .ZN(n8919) );
  XNOR2_X2 U9865 ( .A(n8920), .B(n8919), .ZN(n8923) );
  XNOR2_X2 U9866 ( .A(n10932), .B(n10338), .ZN(n10432) );
  INV_X4 U9867 ( .A(n10432), .ZN(n8921) );
  NAND2_X2 U9868 ( .A1(multOut[22]), .A2(net92392), .ZN(n8947) );
  NAND2_X2 U9869 ( .A1(n10102), .A2(n9976), .ZN(n8927) );
  NAND2_X2 U9870 ( .A1(n9978), .A2(n4880), .ZN(n8926) );
  NAND2_X2 U9871 ( .A1(n6081), .A2(n9975), .ZN(n8925) );
  NAND2_X2 U9872 ( .A1(net77084), .A2(n8977), .ZN(n8924) );
  NAND4_X2 U9873 ( .A1(n8927), .A2(n8926), .A3(n8925), .A4(n8924), .ZN(n9552)
         );
  NAND2_X2 U9874 ( .A1(n10058), .A2(n9552), .ZN(n8934) );
  NAND2_X2 U9875 ( .A1(n8728), .A2(n9547), .ZN(n8932) );
  NAND2_X2 U9876 ( .A1(n4880), .A2(n9548), .ZN(n8931) );
  NAND2_X2 U9877 ( .A1(net77084), .A2(n8928), .ZN(n8930) );
  NAND2_X2 U9878 ( .A1(n6081), .A2(n9546), .ZN(n8929) );
  NAND4_X2 U9879 ( .A1(n8932), .A2(n8931), .A3(n8930), .A4(n8929), .ZN(n9293)
         );
  NAND2_X2 U9880 ( .A1(n10060), .A2(n9293), .ZN(n8933) );
  NAND2_X2 U9881 ( .A1(n8934), .A2(n8933), .ZN(n8945) );
  INV_X4 U9882 ( .A(n9018), .ZN(n8936) );
  NAND2_X2 U9883 ( .A1(n8937), .A2(n5761), .ZN(n8935) );
  NAND2_X2 U9884 ( .A1(n10064), .A2(n9302), .ZN(n8941) );
  INV_X4 U9885 ( .A(n9183), .ZN(n8939) );
  OAI21_X4 U9886 ( .B1(n6005), .B2(n8939), .A(n8938), .ZN(n9982) );
  NAND2_X2 U9887 ( .A1(n10066), .A2(n9982), .ZN(n8940) );
  NAND2_X2 U9888 ( .A1(n8941), .A2(n8940), .ZN(n10070) );
  MUX2_X2 U9889 ( .A(n8942), .B(n10070), .S(net71026), .Z(n8944) );
  NOR3_X4 U9890 ( .A1(n8945), .A2(n8944), .A3(n8943), .ZN(n8946) );
  NAND3_X2 U9891 ( .A1(n8948), .A2(n8947), .A3(n8946), .ZN(dmem_addr_out[22])
         );
  INV_X4 U9892 ( .A(dmem_addr_out[22]), .ZN(n8955) );
  INV_X4 U9893 ( .A(n8950), .ZN(n8964) );
  INV_X4 U9894 ( .A(dmem_read_in[22]), .ZN(n8951) );
  OAI211_X2 U9895 ( .C1(n8955), .C2(net76646), .A(n8954), .B(n8953), .ZN(n8956) );
  OAI22_X2 U9896 ( .A1(n5144), .A2(n6088), .B1(net76660), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9897 ( .A1(n4983), .A2(n6091), .B1(n6156), .B2(n8961), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9898 ( .A1(n6192), .A2(n5367), .B1(n6195), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9899 ( .A1(n6196), .A2(n5621), .B1(n6199), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9900 ( .A1(n5265), .A2(n6097), .B1(n6095), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9901 ( .A1(n5145), .A2(n6103), .B1(n6102), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9902 ( .A1(n5017), .A2(n6108), .B1(n6106), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9903 ( .A1(n5092), .A2(n6112), .B1(n6158), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9904 ( .A1(n5146), .A2(n6115), .B1(n6160), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9905 ( .A1(n5266), .A2(n6118), .B1(n6162), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9906 ( .A1(n6200), .A2(n5368), .B1(n6204), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9907 ( .A1(n5267), .A2(net76862), .B1(net76616), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9908 ( .A1(n6205), .A2(n5504), .B1(n6208), .B2(n8961), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9909 ( .A1(n5147), .A2(n6121), .B1(n6164), .B2(n8961), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9910 ( .A1(n5268), .A2(n6124), .B1(n6166), .B2(n8961), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9911 ( .A1(n5148), .A2(n6127), .B1(n6168), .B2(n8961), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9912 ( .A1(n5149), .A2(n6129), .B1(n6170), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9913 ( .A1(n5269), .A2(n6132), .B1(n6172), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9914 ( .A1(n5150), .A2(n6136), .B1(n6174), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9915 ( .A1(n6209), .A2(n5402), .B1(n6212), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9916 ( .A1(\REGFILE/reg_out[28][22] ), .A2(n6177), .ZN(n8957) );
  OAI21_X4 U9917 ( .B1(n6213), .B2(n6027), .A(n8957), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9918 ( .A1(n6178), .A2(\REGFILE/reg_out[29][22] ), .ZN(n8958) );
  OAI21_X4 U9919 ( .B1(n6138), .B2(n6027), .A(n8958), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9920 ( .A1(n5270), .A2(n6139), .B1(net76550), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9921 ( .A1(n6180), .A2(\REGFILE/reg_out[30][22] ), .ZN(n8959) );
  OAI21_X4 U9922 ( .B1(n6142), .B2(n6027), .A(n8959), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9923 ( .A1(net76488), .A2(\REGFILE/reg_out[31][22] ), .ZN(n8960)
         );
  OAI21_X4 U9924 ( .B1(net76480), .B2(n6027), .A(n8960), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9925 ( .A1(n6215), .A2(n5403), .B1(net76320), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9926 ( .A1(n6217), .A2(n5498), .B1(n6220), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9927 ( .A1(n5271), .A2(n6144), .B1(n6183), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9928 ( .A1(n5272), .A2(net76706), .B1(n6147), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9929 ( .A1(n5151), .A2(net76692), .B1(n6185), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9930 ( .A1(n5273), .A2(n6150), .B1(n6187), .B2(n6027), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9931 ( .A1(n5152), .A2(n6153), .B1(n6189), .B2(n8961), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  XNOR2_X2 U9932 ( .A(n8963), .B(n8962), .ZN(n8966) );
  NAND2_X2 U9933 ( .A1(n6190), .A2(n8964), .ZN(n8965) );
  OAI221_X2 U9934 ( .B1(n8967), .B2(n4962), .C1(n9533), .C2(n8966), .A(n8965), 
        .ZN(\PCLOGIC/PC_REG/REG_32BIT[22].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9935 ( .A1(net73708), .A2(n10930), .ZN(n8973) );
  OAI211_X2 U9936 ( .C1(n8349), .C2(n8970), .A(n8969), .B(n10649), .ZN(n8972)
         );
  NAND2_X2 U9937 ( .A1(n6190), .A2(n9000), .ZN(n8971) );
  MUX2_X2 U9938 ( .A(n8974), .B(n9298), .S(net71026), .Z(n8986) );
  INV_X4 U9939 ( .A(n9802), .ZN(n8985) );
  INV_X4 U9940 ( .A(n8975), .ZN(n8982) );
  NAND2_X2 U9941 ( .A1(n8728), .A2(n8976), .ZN(n8981) );
  NAND2_X2 U9942 ( .A1(n6081), .A2(n8977), .ZN(n8980) );
  AOI22_X2 U9943 ( .A1(net77084), .A2(n8978), .B1(n6083), .B2(n9976), .ZN(
        n8979) );
  OAI22_X2 U9944 ( .A1(n10474), .A2(n8982), .B1(n5061), .B2(n10472), .ZN(n8984) );
  AOI211_X4 U9945 ( .C1(n8986), .C2(n8985), .A(n8984), .B(n8983), .ZN(n8996)
         );
  XNOR2_X2 U9946 ( .A(n8988), .B(n8987), .ZN(n8993) );
  NAND2_X2 U9947 ( .A1(n8991), .A2(n8990), .ZN(n8992) );
  NAND2_X2 U9948 ( .A1(multOut[25]), .A2(net92392), .ZN(n8994) );
  OAI211_X2 U9949 ( .C1(n8996), .C2(net72163), .A(n8995), .B(n8994), .ZN(
        dmem_addr_out[25]) );
  INV_X4 U9950 ( .A(dmem_addr_out[25]), .ZN(n9003) );
  INV_X4 U9951 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [25]), .ZN(n9373) );
  INV_X4 U9952 ( .A(dmem_read_in[25]), .ZN(n8998) );
  OAI211_X2 U9953 ( .C1(n9003), .C2(net76646), .A(n9002), .B(n9001), .ZN(n9004) );
  NAND2_X2 U9954 ( .A1(net76270), .A2(n9004), .ZN(n9009) );
  OAI22_X2 U9955 ( .A1(n5153), .A2(n6088), .B1(net76660), .B2(n6029), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9956 ( .A1(n5274), .A2(n6091), .B1(n6156), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9957 ( .A1(n6192), .A2(n5551), .B1(n6195), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9958 ( .A1(n6196), .A2(n5501), .B1(n6199), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9959 ( .A1(n5275), .A2(n6097), .B1(n6095), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9960 ( .A1(n5154), .A2(n6103), .B1(n6102), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9961 ( .A1(n5276), .A2(n6108), .B1(n6106), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9962 ( .A1(n5155), .A2(n6112), .B1(n6158), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9963 ( .A1(n5508), .A2(n6115), .B1(n6160), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9964 ( .A1(n5441), .A2(n6118), .B1(n6162), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9965 ( .A1(n6200), .A2(n5552), .B1(n6204), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9966 ( .A1(n5442), .A2(net76862), .B1(net76616), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9967 ( .A1(n6205), .A2(n5404), .B1(n6208), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9968 ( .A1(n5156), .A2(n6121), .B1(n6164), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9969 ( .A1(n5277), .A2(n6124), .B1(n6166), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9970 ( .A1(n5157), .A2(n6127), .B1(n6168), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9971 ( .A1(n5158), .A2(n6129), .B1(n6170), .B2(n6029), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9972 ( .A1(n5278), .A2(n6132), .B1(n6172), .B2(n6029), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9973 ( .A1(n5159), .A2(n6136), .B1(n6174), .B2(n6029), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9974 ( .A1(n6209), .A2(n5405), .B1(n6212), .B2(n6029), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9975 ( .A1(\REGFILE/reg_out[28][25] ), .A2(n6177), .ZN(n9005) );
  OAI21_X4 U9976 ( .B1(n6213), .B2(n6029), .A(n9005), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9977 ( .A1(n6178), .A2(\REGFILE/reg_out[29][25] ), .ZN(n9006) );
  OAI21_X4 U9978 ( .B1(n6138), .B2(n6029), .A(n9006), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9979 ( .A1(n5443), .A2(n6139), .B1(net76550), .B2(n6029), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9980 ( .A1(n6180), .A2(\REGFILE/reg_out[30][25] ), .ZN(n9007) );
  OAI21_X4 U9981 ( .B1(n6142), .B2(n6029), .A(n9007), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U9982 ( .A1(net76488), .A2(\REGFILE/reg_out[31][25] ), .ZN(n9008)
         );
  OAI21_X4 U9983 ( .B1(net76480), .B2(n6029), .A(n9008), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9984 ( .A1(n6215), .A2(n5406), .B1(net76320), .B2(n6029), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9985 ( .A1(n6217), .A2(n5369), .B1(n6220), .B2(n6029), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9986 ( .A1(n5279), .A2(n6144), .B1(n6183), .B2(n6029), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9987 ( .A1(n5444), .A2(net76706), .B1(n6147), .B2(n6029), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9988 ( .A1(n5509), .A2(net76692), .B1(n6185), .B2(n6029), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9989 ( .A1(n5445), .A2(n6150), .B1(n6187), .B2(n6029), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U9990 ( .A1(n5510), .A2(n6153), .B1(n6189), .B2(n6030), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ) );
  AOI22_X2 U9991 ( .A1(net71092), .A2(n9011), .B1(net71094), .B2(n9010), .ZN(
        n9026) );
  NAND2_X2 U9992 ( .A1(net77084), .A2(n9548), .ZN(n9016) );
  NAND2_X2 U9993 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[10].MUX/N1 ), .A2(n6041), 
        .ZN(n9361) );
  OAI211_X2 U9994 ( .C1(n9094), .C2(n10109), .A(n9093), .B(n9361), .ZN(n10230)
         );
  NAND2_X2 U9995 ( .A1(n6083), .A2(n10230), .ZN(n9015) );
  NAND2_X2 U9996 ( .A1(n6081), .A2(n10232), .ZN(n9014) );
  NAND2_X2 U9997 ( .A1(n8728), .A2(n10233), .ZN(n9013) );
  NAND4_X2 U9998 ( .A1(n9016), .A2(n9015), .A3(n9014), .A4(n9013), .ZN(n9194)
         );
  NAND2_X2 U9999 ( .A1(n10280), .A2(n9194), .ZN(n9025) );
  INV_X4 U10000 ( .A(n9606), .ZN(net71085) );
  NAND2_X2 U10001 ( .A1(n6081), .A2(n10241), .ZN(n9022) );
  NAND2_X2 U10002 ( .A1(net77086), .A2(n10238), .ZN(n9021) );
  NAND2_X2 U10003 ( .A1(n8728), .A2(n10240), .ZN(n9020) );
  NAND2_X2 U10004 ( .A1(n6083), .A2(n9018), .ZN(n9019) );
  NAND4_X2 U10005 ( .A1(n9022), .A2(n9021), .A3(n9020), .A4(n9019), .ZN(n9182)
         );
  NAND3_X2 U10006 ( .A1(n9026), .A2(n9025), .A3(n9024), .ZN(n9027) );
  MUX2_X2 U10007 ( .A(n9027), .B(multOut[17]), .S(net76452), .Z(n9038) );
  INV_X4 U10008 ( .A(n9028), .ZN(n9032) );
  NAND2_X2 U10009 ( .A1(n9030), .A2(aluA[18]), .ZN(n9031) );
  XNOR2_X2 U10010 ( .A(n9052), .B(n9053), .ZN(n9036) );
  NAND2_X2 U10011 ( .A1(net71078), .A2(aluA[17]), .ZN(n9034) );
  OAI22_X2 U10012 ( .A1(n9036), .A2(net70691), .B1(n9035), .B2(n9034), .ZN(
        n9037) );
  NOR2_X4 U10013 ( .A1(n9038), .A2(n9037), .ZN(n9044) );
  INV_X4 U10014 ( .A(n9044), .ZN(dmem_addr_out[17]) );
  INV_X4 U10015 ( .A(dmem_read_in[17]), .ZN(n9039) );
  OAI211_X2 U10016 ( .C1(n9044), .C2(net76646), .A(n9043), .B(n9042), .ZN(
        n9045) );
  OAI22_X2 U10017 ( .A1(n5093), .A2(n6088), .B1(net76660), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10018 ( .A1(n5073), .A2(n6091), .B1(n6156), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10019 ( .A1(n6192), .A2(n5370), .B1(n6194), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10020 ( .A1(n6196), .A2(n5620), .B1(n6198), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10021 ( .A1(n5280), .A2(n6097), .B1(n6095), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10022 ( .A1(n5160), .A2(n6103), .B1(n6102), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10023 ( .A1(n5018), .A2(n6108), .B1(n6106), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10024 ( .A1(n5094), .A2(n6112), .B1(n6158), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10025 ( .A1(n5095), .A2(n6115), .B1(n6160), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10026 ( .A1(n5074), .A2(n6118), .B1(n6162), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10027 ( .A1(n6200), .A2(n5116), .B1(n6203), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10028 ( .A1(n5075), .A2(net76862), .B1(net76616), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10029 ( .A1(n6205), .A2(n5407), .B1(n6207), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10030 ( .A1(n5161), .A2(n6121), .B1(n6164), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10031 ( .A1(n5281), .A2(n6124), .B1(n6166), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10032 ( .A1(n5162), .A2(n6127), .B1(n6168), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10033 ( .A1(n5096), .A2(n6129), .B1(n6170), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10034 ( .A1(n5019), .A2(n6132), .B1(n6172), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10035 ( .A1(n5097), .A2(n6136), .B1(n6174), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10036 ( .A1(n6209), .A2(n5027), .B1(n6211), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10037 ( .A1(\REGFILE/reg_out[28][17] ), .A2(n6177), .ZN(n9046) );
  NAND2_X2 U10038 ( .A1(n6178), .A2(\REGFILE/reg_out[29][17] ), .ZN(n9047) );
  OAI22_X2 U10039 ( .A1(n5020), .A2(n6139), .B1(net76550), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10040 ( .A1(n6180), .A2(\REGFILE/reg_out[30][17] ), .ZN(n9048) );
  NAND2_X2 U10041 ( .A1(net76488), .A2(\REGFILE/reg_out[31][17] ), .ZN(n9049)
         );
  OAI22_X2 U10042 ( .A1(n6215), .A2(n5111), .B1(net76318), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10043 ( .A1(n6217), .A2(n5117), .B1(n6219), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10044 ( .A1(n5076), .A2(n6144), .B1(n6183), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10045 ( .A1(n5077), .A2(net76706), .B1(n6147), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10046 ( .A1(n5098), .A2(net76692), .B1(n6185), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10047 ( .A1(n5078), .A2(n6150), .B1(n6187), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10048 ( .A1(n5099), .A2(n6153), .B1(n6189), .B2(n6032), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[17].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10049 ( .A1(multOut[12]), .A2(net92392), .ZN(n9106) );
  XNOR2_X2 U10050 ( .A(n9351), .B(n9075), .ZN(n9352) );
  INV_X4 U10051 ( .A(n9352), .ZN(n9063) );
  AOI22_X2 U10052 ( .A1(n9053), .A2(n9052), .B1(n9051), .B2(aluA[17]), .ZN(
        n9179) );
  INV_X4 U10053 ( .A(n9179), .ZN(n9056) );
  AOI22_X2 U10054 ( .A1(n9178), .A2(n9056), .B1(n9055), .B2(aluA[16]), .ZN(
        n10287) );
  OAI22_X2 U10055 ( .A1(n9058), .A2(n10463), .B1(n10287), .B2(n4807), .ZN(
        n10253) );
  XNOR2_X2 U10056 ( .A(n9059), .B(n10247), .ZN(n10254) );
  AOI22_X2 U10057 ( .A1(n10253), .A2(n10254), .B1(
        \WIRE_ALU_A/MUX2TO1_32BIT[14].MUX/N1 ), .B2(n9059), .ZN(n9393) );
  XNOR2_X2 U10058 ( .A(n9060), .B(n10368), .ZN(n9392) );
  INV_X4 U10059 ( .A(n9392), .ZN(n9062) );
  NAND2_X2 U10060 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[13].MUX/N1 ), .A2(n9060), 
        .ZN(n9061) );
  XNOR2_X2 U10061 ( .A(n9063), .B(n9353), .ZN(n9064) );
  NAND2_X2 U10062 ( .A1(net71271), .A2(n9064), .ZN(n9105) );
  NAND2_X2 U10063 ( .A1(net70720), .A2(net80189), .ZN(n9067) );
  NAND2_X2 U10064 ( .A1(n10931), .A2(n9065), .ZN(n10462) );
  NAND2_X2 U10065 ( .A1(n10102), .A2(n10239), .ZN(n9074) );
  NAND2_X2 U10066 ( .A1(net77086), .A2(n9838), .ZN(n9073) );
  NAND2_X2 U10067 ( .A1(n6083), .A2(n10240), .ZN(n9072) );
  NAND2_X2 U10068 ( .A1(n6081), .A2(n10238), .ZN(n9071) );
  NAND4_X2 U10069 ( .A1(n9074), .A2(n9073), .A3(n9072), .A4(n9071), .ZN(n9403)
         );
  INV_X4 U10070 ( .A(n10423), .ZN(n10373) );
  NAND2_X2 U10071 ( .A1(n8759), .A2(n9500), .ZN(n9086) );
  NAND2_X2 U10072 ( .A1(net77086), .A2(n9621), .ZN(n9085) );
  NAND2_X2 U10073 ( .A1(n6083), .A2(n9396), .ZN(n9084) );
  NAND2_X2 U10074 ( .A1(n6081), .A2(n9395), .ZN(n9083) );
  NAND4_X2 U10075 ( .A1(n9086), .A2(n9085), .A3(n9084), .A4(n9083), .ZN(n9837)
         );
  NAND2_X2 U10076 ( .A1(n10066), .A2(n9837), .ZN(n9092) );
  NAND2_X2 U10077 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[7].MUX/N1 ), .A2(n6040), 
        .ZN(n9594) );
  NAND2_X2 U10078 ( .A1(net70696), .A2(n9581), .ZN(n9580) );
  NAND2_X2 U10079 ( .A1(n9594), .A2(n9580), .ZN(n9493) );
  NAND2_X2 U10080 ( .A1(n6081), .A2(n9493), .ZN(n9090) );
  NAND2_X2 U10081 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[9].MUX/N1 ), .A2(n6041), 
        .ZN(n9342) );
  OAI211_X2 U10082 ( .C1(n9094), .C2(net71273), .A(n9093), .B(n9342), .ZN(
        n9407) );
  NAND2_X2 U10083 ( .A1(n8759), .A2(n9407), .ZN(n9089) );
  NAND2_X2 U10084 ( .A1(net77086), .A2(n9408), .ZN(n9088) );
  NAND2_X2 U10085 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[5].MUX/N1 ), .A2(n6041), 
        .ZN(n9598) );
  NAND2_X2 U10086 ( .A1(n9598), .A2(n9580), .ZN(n9585) );
  NAND2_X2 U10087 ( .A1(n4880), .A2(n9585), .ZN(n9087) );
  NAND4_X2 U10088 ( .A1(n9090), .A2(n9089), .A3(n9088), .A4(n9087), .ZN(n9852)
         );
  NAND2_X2 U10089 ( .A1(n10058), .A2(n9852), .ZN(n9091) );
  NAND2_X2 U10090 ( .A1(n9092), .A2(n9091), .ZN(n9102) );
  NAND2_X2 U10091 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[6].MUX/N1 ), .A2(n6040), 
        .ZN(n9618) );
  NAND2_X2 U10092 ( .A1(n9618), .A2(n9580), .ZN(n9845) );
  NAND2_X2 U10093 ( .A1(n4880), .A2(n9845), .ZN(n9098) );
  NAND2_X2 U10094 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[8].MUX/N1 ), .A2(n6040), 
        .ZN(n9498) );
  OAI211_X2 U10095 ( .C1(net70535), .C2(n9094), .A(n9498), .B(n9093), .ZN(
        n10231) );
  NAND2_X2 U10096 ( .A1(n6081), .A2(n10231), .ZN(n9097) );
  NAND2_X2 U10097 ( .A1(net77086), .A2(n10232), .ZN(n9096) );
  NAND2_X2 U10098 ( .A1(n8728), .A2(n10230), .ZN(n9095) );
  NAND4_X2 U10099 ( .A1(n9098), .A2(n9097), .A3(n9096), .A4(n9095), .ZN(n9404)
         );
  INV_X4 U10100 ( .A(n9404), .ZN(n9100) );
  NOR2_X4 U10101 ( .A1(n9102), .A2(n9101), .ZN(n9103) );
  NAND4_X2 U10102 ( .A1(n9106), .A2(n9105), .A3(n9104), .A4(n9103), .ZN(
        dmem_addr_out[12]) );
  NAND2_X2 U10103 ( .A1(net76650), .A2(dmem_addr_out[12]), .ZN(n9112) );
  INV_X4 U10104 ( .A(n9107), .ZN(n9110) );
  AOI21_X4 U10105 ( .B1(n9110), .B2(net77030), .A(n9109), .ZN(n9111) );
  NAND3_X2 U10106 ( .A1(n9112), .A2(net70740), .A3(n9111), .ZN(n9113) );
  NAND2_X2 U10107 ( .A1(n6034), .A2(n4992), .ZN(n9115) );
  NAND2_X2 U10108 ( .A1(n4867), .A2(\REGFILE/reg_out[0][12] ), .ZN(n9114) );
  NAND2_X2 U10109 ( .A1(n9115), .A2(n9114), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10110 ( .A1(n6034), .A2(n4990), .ZN(n9117) );
  NAND2_X2 U10111 ( .A1(n6093), .A2(\REGFILE/reg_out[10][12] ), .ZN(n9116) );
  NAND2_X2 U10112 ( .A1(n9117), .A2(n9116), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10113 ( .A1(n6034), .A2(n4998), .ZN(n9119) );
  NAND2_X2 U10114 ( .A1(\REGFILE/reg_out[11][12] ), .A2(n4869), .ZN(n9118) );
  NAND2_X2 U10115 ( .A1(n9119), .A2(n9118), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10116 ( .A1(n6034), .A2(n4993), .ZN(n9121) );
  NAND2_X2 U10117 ( .A1(n9121), .A2(n9120), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10118 ( .A1(n6034), .A2(n6096), .ZN(n9123) );
  NAND2_X2 U10119 ( .A1(n9123), .A2(n9122), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10120 ( .A1(n6034), .A2(n6101), .ZN(n9125) );
  NAND2_X2 U10121 ( .A1(n4805), .A2(\REGFILE/reg_out[14][12] ), .ZN(n9124) );
  NAND2_X2 U10122 ( .A1(n9125), .A2(n9124), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10123 ( .A1(n6034), .A2(n6107), .ZN(n9127) );
  NAND2_X2 U10124 ( .A1(n9127), .A2(n9126), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10125 ( .A1(n6034), .A2(n4994), .ZN(n9129) );
  NAND2_X2 U10126 ( .A1(n4891), .A2(\REGFILE/reg_out[16][12] ), .ZN(n9128) );
  NAND2_X2 U10127 ( .A1(n9129), .A2(n9128), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10128 ( .A1(n6034), .A2(n4999), .ZN(n9131) );
  NAND2_X2 U10129 ( .A1(n4892), .A2(\REGFILE/reg_out[17][12] ), .ZN(n9130) );
  NAND2_X2 U10130 ( .A1(n9131), .A2(n9130), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10131 ( .A1(n6034), .A2(n5000), .ZN(n9133) );
  NAND2_X2 U10132 ( .A1(n4884), .A2(\REGFILE/reg_out[18][12] ), .ZN(n9132) );
  NAND2_X2 U10133 ( .A1(n9133), .A2(n9132), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10134 ( .A1(n6033), .A2(n5001), .ZN(n9135) );
  NAND2_X2 U10135 ( .A1(\REGFILE/reg_out[19][12] ), .A2(n4876), .ZN(n9134) );
  NAND2_X2 U10136 ( .A1(n9135), .A2(n9134), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10137 ( .A1(n6033), .A2(n4997), .ZN(n9137) );
  NAND2_X2 U10138 ( .A1(n4877), .A2(\REGFILE/reg_out[1][12] ), .ZN(n9136) );
  NAND2_X2 U10139 ( .A1(n9137), .A2(n9136), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10140 ( .A1(n6033), .A2(n4903), .ZN(n9139) );
  NAND2_X2 U10141 ( .A1(\REGFILE/reg_out[20][12] ), .A2(n4868), .ZN(n9138) );
  NAND2_X2 U10142 ( .A1(n9139), .A2(n9138), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10143 ( .A1(n6033), .A2(n4904), .ZN(n9141) );
  NAND2_X2 U10144 ( .A1(n4882), .A2(\REGFILE/reg_out[21][12] ), .ZN(n9140) );
  NAND2_X2 U10145 ( .A1(n9141), .A2(n9140), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10146 ( .A1(n6033), .A2(n4905), .ZN(n9143) );
  NAND2_X2 U10147 ( .A1(n4888), .A2(\REGFILE/reg_out[22][12] ), .ZN(n9142) );
  NAND2_X2 U10148 ( .A1(n9143), .A2(n9142), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10149 ( .A1(n6033), .A2(n4906), .ZN(n9145) );
  NAND2_X2 U10150 ( .A1(n4883), .A2(\REGFILE/reg_out[23][12] ), .ZN(n9144) );
  NAND2_X2 U10151 ( .A1(n9145), .A2(n9144), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10152 ( .A1(n6033), .A2(n4995), .ZN(n9147) );
  NAND2_X2 U10153 ( .A1(n4875), .A2(\REGFILE/reg_out[24][12] ), .ZN(n9146) );
  NAND2_X2 U10154 ( .A1(n9147), .A2(n9146), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10155 ( .A1(n6033), .A2(n5002), .ZN(n9149) );
  NAND2_X2 U10156 ( .A1(n4878), .A2(\REGFILE/reg_out[25][12] ), .ZN(n9148) );
  NAND2_X2 U10157 ( .A1(n9149), .A2(n9148), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10158 ( .A1(n6033), .A2(n5003), .ZN(n9151) );
  NAND2_X2 U10159 ( .A1(n4893), .A2(\REGFILE/reg_out[26][12] ), .ZN(n9150) );
  NAND2_X2 U10160 ( .A1(n9151), .A2(n9150), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10161 ( .A1(n6033), .A2(n5004), .ZN(n9153) );
  NAND2_X2 U10162 ( .A1(\REGFILE/reg_out[27][12] ), .A2(n4872), .ZN(n9152) );
  NAND2_X2 U10163 ( .A1(n9153), .A2(n9152), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10164 ( .A1(n6033), .A2(n4806), .ZN(n9155) );
  NAND2_X2 U10165 ( .A1(n9155), .A2(n9154), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10166 ( .A1(n6033), .A2(n10607), .ZN(n9157) );
  NAND2_X2 U10167 ( .A1(n6178), .A2(\REGFILE/reg_out[29][12] ), .ZN(n9156) );
  NAND2_X2 U10168 ( .A1(n9157), .A2(n9156), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10169 ( .A1(n6033), .A2(n5005), .ZN(n9159) );
  NAND2_X2 U10170 ( .A1(n4879), .A2(\REGFILE/reg_out[2][12] ), .ZN(n9158) );
  NAND2_X2 U10171 ( .A1(n9159), .A2(n9158), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10172 ( .A1(n6033), .A2(n10614), .ZN(n9161) );
  NAND2_X2 U10173 ( .A1(n6180), .A2(\REGFILE/reg_out[30][12] ), .ZN(n9160) );
  NAND2_X2 U10174 ( .A1(n9161), .A2(n9160), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10175 ( .A1(n6034), .A2(net70574), .ZN(n9163) );
  NAND2_X2 U10176 ( .A1(net76488), .A2(\REGFILE/reg_out[31][12] ), .ZN(n9162)
         );
  NAND2_X2 U10177 ( .A1(n9163), .A2(n9162), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10178 ( .A1(n6034), .A2(n5009), .ZN(n9165) );
  NAND2_X2 U10180 ( .A1(n9165), .A2(n9164), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10181 ( .A1(n6034), .A2(n4996), .ZN(n9167) );
  NAND2_X2 U10182 ( .A1(\REGFILE/reg_out[4][12] ), .A2(n4870), .ZN(n9166) );
  NAND2_X2 U10183 ( .A1(n9167), .A2(n9166), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10184 ( .A1(n6034), .A2(n5006), .ZN(n9169) );
  NAND2_X2 U10185 ( .A1(n4885), .A2(\REGFILE/reg_out[5][12] ), .ZN(n9168) );
  NAND2_X2 U10186 ( .A1(n9169), .A2(n9168), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10187 ( .A1(n6034), .A2(n6148), .ZN(n9171) );
  NAND2_X2 U10188 ( .A1(n4889), .A2(\REGFILE/reg_out[6][12] ), .ZN(n9170) );
  NAND2_X2 U10189 ( .A1(n9171), .A2(n9170), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10190 ( .A1(n6033), .A2(n5007), .ZN(n9173) );
  NAND2_X2 U10191 ( .A1(n4886), .A2(\REGFILE/reg_out[7][12] ), .ZN(n9172) );
  NAND2_X2 U10192 ( .A1(n9173), .A2(n9172), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10193 ( .A1(n6033), .A2(n4991), .ZN(n9175) );
  NAND2_X2 U10195 ( .A1(n9175), .A2(n9174), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10196 ( .A1(n6034), .A2(n5008), .ZN(n9177) );
  NAND2_X2 U10197 ( .A1(n4887), .A2(\REGFILE/reg_out[9][12] ), .ZN(n9176) );
  NAND2_X2 U10198 ( .A1(n9177), .A2(n9176), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10199 ( .A1(multOut[16]), .A2(net92392), .ZN(n9202) );
  XNOR2_X2 U10200 ( .A(n9179), .B(n9178), .ZN(n9180) );
  NAND2_X2 U10201 ( .A1(net71271), .A2(n9180), .ZN(n9201) );
  NAND2_X2 U10202 ( .A1(n6081), .A2(n9397), .ZN(n9187) );
  NAND2_X2 U10203 ( .A1(net77086), .A2(n9395), .ZN(n9186) );
  NAND2_X2 U10204 ( .A1(n8759), .A2(n9396), .ZN(n9185) );
  NAND2_X2 U10205 ( .A1(n6083), .A2(n9183), .ZN(n9184) );
  NAND4_X2 U10206 ( .A1(n9187), .A2(n9186), .A3(n9185), .A4(n9184), .ZN(n10277) );
  NAND2_X2 U10207 ( .A1(n10066), .A2(n10277), .ZN(n9193) );
  NAND2_X2 U10208 ( .A1(net77086), .A2(n9978), .ZN(n9191) );
  NAND2_X2 U10209 ( .A1(n6083), .A2(n9407), .ZN(n9190) );
  NAND2_X2 U10210 ( .A1(n6081), .A2(n9408), .ZN(n9189) );
  NAND2_X2 U10211 ( .A1(n8759), .A2(n9977), .ZN(n9188) );
  NAND4_X2 U10212 ( .A1(n9191), .A2(n9190), .A3(n9189), .A4(n9188), .ZN(n10278) );
  NAND2_X2 U10213 ( .A1(n10058), .A2(n10278), .ZN(n9192) );
  NAND2_X2 U10214 ( .A1(n9193), .A2(n9192), .ZN(n9198) );
  INV_X4 U10215 ( .A(n9194), .ZN(n9196) );
  NAND4_X2 U10216 ( .A1(n9202), .A2(n9201), .A3(n9200), .A4(n9199), .ZN(
        dmem_addr_out[16]) );
  AOI21_X4 U10217 ( .B1(n9205), .B2(n9204), .A(net76278), .ZN(n9268) );
  NAND2_X2 U10218 ( .A1(n6036), .A2(n4992), .ZN(n9207) );
  NAND2_X2 U10219 ( .A1(n4867), .A2(\REGFILE/reg_out[0][16] ), .ZN(n9206) );
  NAND2_X2 U10220 ( .A1(n9207), .A2(n9206), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10221 ( .A1(n6036), .A2(n4990), .ZN(n9209) );
  NAND2_X2 U10222 ( .A1(n6093), .A2(\REGFILE/reg_out[10][16] ), .ZN(n9208) );
  NAND2_X2 U10223 ( .A1(n9209), .A2(n9208), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10224 ( .A1(n6036), .A2(n4998), .ZN(n9211) );
  NAND2_X2 U10225 ( .A1(\REGFILE/reg_out[11][16] ), .A2(n4869), .ZN(n9210) );
  NAND2_X2 U10226 ( .A1(n9211), .A2(n9210), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10227 ( .A1(n6036), .A2(n4993), .ZN(n9213) );
  NAND2_X2 U10228 ( .A1(n9213), .A2(n9212), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10229 ( .A1(n6036), .A2(n6096), .ZN(n9215) );
  NAND2_X2 U10230 ( .A1(n6100), .A2(\REGFILE/reg_out[13][16] ), .ZN(n9214) );
  NAND2_X2 U10231 ( .A1(n9215), .A2(n9214), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10232 ( .A1(n6036), .A2(n6101), .ZN(n9217) );
  NAND2_X2 U10233 ( .A1(n4805), .A2(\REGFILE/reg_out[14][16] ), .ZN(n9216) );
  NAND2_X2 U10234 ( .A1(n9217), .A2(n9216), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10235 ( .A1(n6036), .A2(n6107), .ZN(n9219) );
  NAND2_X2 U10236 ( .A1(n9219), .A2(n9218), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10237 ( .A1(n6036), .A2(n4994), .ZN(n9221) );
  NAND2_X2 U10238 ( .A1(n4891), .A2(\REGFILE/reg_out[16][16] ), .ZN(n9220) );
  NAND2_X2 U10239 ( .A1(n9221), .A2(n9220), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10240 ( .A1(n6036), .A2(n4999), .ZN(n9223) );
  NAND2_X2 U10241 ( .A1(n4892), .A2(\REGFILE/reg_out[17][16] ), .ZN(n9222) );
  NAND2_X2 U10242 ( .A1(n9223), .A2(n9222), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10243 ( .A1(n6036), .A2(n5000), .ZN(n9225) );
  NAND2_X2 U10244 ( .A1(n9225), .A2(n9224), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10245 ( .A1(n6035), .A2(n5001), .ZN(n9227) );
  NAND2_X2 U10246 ( .A1(\REGFILE/reg_out[19][16] ), .A2(n4876), .ZN(n9226) );
  NAND2_X2 U10247 ( .A1(n9227), .A2(n9226), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10248 ( .A1(n6035), .A2(n4997), .ZN(n9229) );
  NAND2_X2 U10249 ( .A1(n4877), .A2(\REGFILE/reg_out[1][16] ), .ZN(n9228) );
  NAND2_X2 U10250 ( .A1(n9229), .A2(n9228), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10251 ( .A1(n6035), .A2(n4903), .ZN(n9231) );
  NAND2_X2 U10252 ( .A1(\REGFILE/reg_out[20][16] ), .A2(n4868), .ZN(n9230) );
  NAND2_X2 U10253 ( .A1(n9231), .A2(n9230), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10254 ( .A1(n6035), .A2(n4904), .ZN(n9233) );
  NAND2_X2 U10255 ( .A1(n4882), .A2(\REGFILE/reg_out[21][16] ), .ZN(n9232) );
  NAND2_X2 U10256 ( .A1(n9233), .A2(n9232), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10257 ( .A1(n6035), .A2(n4905), .ZN(n9235) );
  NAND2_X2 U10258 ( .A1(n9235), .A2(n9234), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10259 ( .A1(n6035), .A2(n4906), .ZN(n9237) );
  NAND2_X2 U10260 ( .A1(n4883), .A2(\REGFILE/reg_out[23][16] ), .ZN(n9236) );
  NAND2_X2 U10261 ( .A1(n9237), .A2(n9236), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10262 ( .A1(n6035), .A2(n4995), .ZN(n9239) );
  NAND2_X2 U10263 ( .A1(n4875), .A2(\REGFILE/reg_out[24][16] ), .ZN(n9238) );
  NAND2_X2 U10264 ( .A1(n9239), .A2(n9238), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10265 ( .A1(n6035), .A2(n5002), .ZN(n9241) );
  NAND2_X2 U10266 ( .A1(n9241), .A2(n9240), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10267 ( .A1(n6035), .A2(n5003), .ZN(n9243) );
  NAND2_X2 U10268 ( .A1(n4893), .A2(\REGFILE/reg_out[26][16] ), .ZN(n9242) );
  NAND2_X2 U10269 ( .A1(n9243), .A2(n9242), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10270 ( .A1(n6035), .A2(n5004), .ZN(n9245) );
  NAND2_X2 U10271 ( .A1(n9245), .A2(n9244), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10272 ( .A1(n6035), .A2(n4806), .ZN(n9247) );
  NAND2_X2 U10273 ( .A1(\REGFILE/reg_out[28][16] ), .A2(n6177), .ZN(n9246) );
  NAND2_X2 U10274 ( .A1(n9247), .A2(n9246), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10275 ( .A1(n6035), .A2(n10607), .ZN(n9249) );
  NAND2_X2 U10276 ( .A1(n6178), .A2(\REGFILE/reg_out[29][16] ), .ZN(n9248) );
  NAND2_X2 U10277 ( .A1(n9249), .A2(n9248), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10278 ( .A1(n6035), .A2(n5005), .ZN(n9251) );
  NAND2_X2 U10279 ( .A1(n4879), .A2(\REGFILE/reg_out[2][16] ), .ZN(n9250) );
  NAND2_X2 U10280 ( .A1(n9251), .A2(n9250), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10281 ( .A1(n6035), .A2(n10614), .ZN(n9253) );
  NAND2_X2 U10282 ( .A1(n6180), .A2(\REGFILE/reg_out[30][16] ), .ZN(n9252) );
  NAND2_X2 U10283 ( .A1(n9253), .A2(n9252), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10284 ( .A1(n6036), .A2(net70574), .ZN(n9255) );
  NAND2_X2 U10285 ( .A1(net76488), .A2(\REGFILE/reg_out[31][16] ), .ZN(n9254)
         );
  NAND2_X2 U10286 ( .A1(n9255), .A2(n9254), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10287 ( .A1(n6036), .A2(n5009), .ZN(n9257) );
  NAND2_X2 U10288 ( .A1(n9257), .A2(n9256), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10289 ( .A1(n6036), .A2(n4996), .ZN(n9259) );
  NAND2_X2 U10290 ( .A1(\REGFILE/reg_out[4][16] ), .A2(n4870), .ZN(n9258) );
  NAND2_X2 U10291 ( .A1(n9259), .A2(n9258), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10292 ( .A1(n6036), .A2(n5006), .ZN(n9261) );
  NAND2_X2 U10293 ( .A1(n4885), .A2(\REGFILE/reg_out[5][16] ), .ZN(n9260) );
  NAND2_X2 U10294 ( .A1(n9261), .A2(n9260), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10295 ( .A1(n6036), .A2(n6148), .ZN(n9263) );
  NAND2_X2 U10296 ( .A1(n9263), .A2(n9262), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10297 ( .A1(n6036), .A2(n5007), .ZN(n9265) );
  NAND2_X2 U10298 ( .A1(n4886), .A2(\REGFILE/reg_out[7][16] ), .ZN(n9264) );
  NAND2_X2 U10299 ( .A1(n9265), .A2(n9264), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10300 ( .A1(n6035), .A2(n4991), .ZN(n9267) );
  NAND2_X2 U10301 ( .A1(n4890), .A2(\REGFILE/reg_out[8][16] ), .ZN(n9266) );
  NAND2_X2 U10302 ( .A1(n9267), .A2(n9266), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10303 ( .A1(n6035), .A2(n5008), .ZN(n9270) );
  NAND2_X2 U10304 ( .A1(n4887), .A2(\REGFILE/reg_out[9][16] ), .ZN(n9269) );
  NAND2_X2 U10305 ( .A1(n9270), .A2(n9269), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[16].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10306 ( .A1(n10649), .A2(n9272), .ZN(n9275) );
  NAND2_X2 U10307 ( .A1(n6190), .A2(n10003), .ZN(n9274) );
  NAND2_X2 U10308 ( .A1(net73708), .A2(aluA[19]), .ZN(n9273) );
  OAI211_X2 U10309 ( .C1(n9276), .C2(n9275), .A(n9274), .B(n9273), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  XNOR2_X2 U10310 ( .A(n9278), .B(n9277), .ZN(n9282) );
  INV_X4 U10311 ( .A(n9279), .ZN(n10080) );
  NAND2_X2 U10312 ( .A1(n6190), .A2(n10080), .ZN(n9281) );
  NAND2_X2 U10313 ( .A1(net73708), .A2(aluA[20]), .ZN(n9280) );
  OAI211_X2 U10314 ( .C1(n9282), .C2(n9533), .A(n9281), .B(n9280), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10315 ( .A1(net73708), .A2(n10931), .ZN(n9288) );
  OAI211_X2 U10316 ( .C1(n8353), .C2(n9285), .A(n9284), .B(n10649), .ZN(n9287)
         );
  NAND2_X2 U10317 ( .A1(n6190), .A2(n9316), .ZN(n9286) );
  XNOR2_X2 U10318 ( .A(n9290), .B(n9289), .ZN(n9292) );
  XNOR2_X2 U10319 ( .A(n10931), .B(n9306), .ZN(n10429) );
  INV_X4 U10320 ( .A(n10429), .ZN(n10336) );
  NAND2_X2 U10321 ( .A1(multOut[23]), .A2(net92392), .ZN(n9311) );
  NAND2_X2 U10322 ( .A1(n10058), .A2(n9293), .ZN(n9296) );
  NAND2_X2 U10323 ( .A1(n10060), .A2(n9294), .ZN(n9295) );
  NAND2_X2 U10324 ( .A1(n9296), .A2(n9295), .ZN(n9309) );
  NAND2_X2 U10325 ( .A1(n10064), .A2(n9297), .ZN(n9300) );
  NAND2_X2 U10326 ( .A1(n10066), .A2(n9298), .ZN(n9299) );
  NAND2_X2 U10327 ( .A1(n9300), .A2(n9299), .ZN(n9305) );
  NAND2_X2 U10328 ( .A1(n10064), .A2(n9301), .ZN(n9304) );
  NAND2_X2 U10329 ( .A1(n10066), .A2(n9302), .ZN(n9303) );
  NAND2_X2 U10330 ( .A1(n9304), .A2(n9303), .ZN(n9558) );
  MUX2_X2 U10331 ( .A(n9305), .B(n9558), .S(net71026), .Z(n9308) );
  NOR3_X4 U10332 ( .A1(n9309), .A2(n9308), .A3(n9307), .ZN(n9310) );
  NAND3_X2 U10333 ( .A1(n9312), .A2(n9311), .A3(n9310), .ZN(dmem_addr_out[23])
         );
  INV_X4 U10334 ( .A(dmem_addr_out[23]), .ZN(n9319) );
  INV_X4 U10335 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [23]), .ZN(n10505) );
  INV_X4 U10336 ( .A(dmem_read_in[23]), .ZN(n9314) );
  OAI211_X2 U10337 ( .C1(n9319), .C2(net76646), .A(n9318), .B(n9317), .ZN(
        n9320) );
  OAI22_X2 U10338 ( .A1(n5511), .A2(n6088), .B1(net76660), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10339 ( .A1(n5446), .A2(n6091), .B1(n6156), .B2(n9325), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10340 ( .A1(n6192), .A2(n5553), .B1(n6195), .B2(n9325), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10341 ( .A1(n6196), .A2(n5502), .B1(n6199), .B2(n9325), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10342 ( .A1(n5282), .A2(n6097), .B1(n6095), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10343 ( .A1(n5163), .A2(n6103), .B1(n6102), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10344 ( .A1(n5283), .A2(n6108), .B1(n6106), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10345 ( .A1(n5164), .A2(n6112), .B1(n6158), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10346 ( .A1(n5512), .A2(n6115), .B1(n6160), .B2(n9325), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10347 ( .A1(n5447), .A2(n6118), .B1(n6162), .B2(n9325), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10348 ( .A1(n6200), .A2(n5371), .B1(n6204), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10349 ( .A1(n5284), .A2(net76862), .B1(net76616), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10350 ( .A1(n6206), .A2(n5408), .B1(n6208), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10351 ( .A1(n5165), .A2(n6121), .B1(n6164), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10352 ( .A1(n5285), .A2(n6124), .B1(n6166), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10353 ( .A1(n5166), .A2(n6127), .B1(n6168), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10354 ( .A1(n5513), .A2(n6129), .B1(n6170), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10355 ( .A1(n5448), .A2(n6132), .B1(n6172), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10356 ( .A1(n5167), .A2(n6136), .B1(n6174), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10357 ( .A1(n6209), .A2(n5409), .B1(n6212), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10358 ( .A1(\REGFILE/reg_out[28][23] ), .A2(n6177), .ZN(n9321) );
  OAI21_X4 U10359 ( .B1(n6213), .B2(n6038), .A(n9321), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10360 ( .A1(n6178), .A2(\REGFILE/reg_out[29][23] ), .ZN(n9322) );
  OAI21_X4 U10361 ( .B1(n6138), .B2(n6038), .A(n9322), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10362 ( .A1(n5449), .A2(n6139), .B1(net76550), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10363 ( .A1(n6180), .A2(\REGFILE/reg_out[30][23] ), .ZN(n9323) );
  OAI21_X4 U10364 ( .B1(n6142), .B2(n6038), .A(n9323), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10365 ( .A1(net76488), .A2(\REGFILE/reg_out[31][23] ), .ZN(n9324)
         );
  OAI21_X4 U10366 ( .B1(net76480), .B2(n6038), .A(n9324), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10367 ( .A1(n6215), .A2(n5410), .B1(net76320), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10368 ( .A1(n6218), .A2(n5372), .B1(n6220), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10369 ( .A1(n5286), .A2(n6144), .B1(n6183), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10370 ( .A1(n5450), .A2(net76706), .B1(n6147), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10371 ( .A1(n5514), .A2(net76692), .B1(n6185), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10372 ( .A1(n5287), .A2(n6150), .B1(n6187), .B2(n6038), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10373 ( .A1(n5168), .A2(n6153), .B1(n6189), .B2(n9325), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10374 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[2].MUX/N1 ), .A2(n6040), 
        .ZN(n10096) );
  NAND2_X2 U10375 ( .A1(n10096), .A2(n9580), .ZN(n10013) );
  NAND2_X2 U10376 ( .A1(n4880), .A2(n10013), .ZN(n9329) );
  NAND2_X2 U10377 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[4].MUX/N1 ), .A2(n6040), 
        .ZN(n9939) );
  NAND2_X2 U10378 ( .A1(n9939), .A2(n9580), .ZN(n9844) );
  NAND2_X2 U10379 ( .A1(n9844), .A2(n6082), .ZN(n9328) );
  NAND2_X2 U10380 ( .A1(net77086), .A2(n10231), .ZN(n9327) );
  NAND2_X2 U10381 ( .A1(n8759), .A2(n9845), .ZN(n9326) );
  NAND4_X2 U10382 ( .A1(n9329), .A2(n9328), .A3(n9327), .A4(n9326), .ZN(n9492)
         );
  INV_X4 U10383 ( .A(n9492), .ZN(n9336) );
  NAND2_X2 U10384 ( .A1(net77086), .A2(n9407), .ZN(n9334) );
  NAND2_X2 U10385 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[3].MUX/N1 ), .A2(n6041), 
        .ZN(n10019) );
  NAND2_X2 U10386 ( .A1(n10019), .A2(n9580), .ZN(n9935) );
  NAND2_X2 U10387 ( .A1(n4880), .A2(n9935), .ZN(n9333) );
  NAND2_X2 U10388 ( .A1(n6082), .A2(n9585), .ZN(n9332) );
  NAND2_X2 U10389 ( .A1(n10102), .A2(n9493), .ZN(n9331) );
  NAND4_X2 U10390 ( .A1(n9334), .A2(n9333), .A3(n9332), .A4(n9331), .ZN(n10124) );
  INV_X4 U10391 ( .A(n10124), .ZN(n9335) );
  OAI22_X2 U10392 ( .A1(n10474), .A2(n9336), .B1(n10472), .B2(n9335), .ZN(
        n9338) );
  NAND2_X2 U10393 ( .A1(net70720), .A2(n5761), .ZN(n9339) );
  NAND2_X2 U10394 ( .A1(n10102), .A2(n9839), .ZN(n9347) );
  OAI211_X2 U10395 ( .C1(net70868), .C2(n10327), .A(n9343), .B(n9342), .ZN(
        n10024) );
  NAND2_X2 U10396 ( .A1(net77086), .A2(n10024), .ZN(n9346) );
  NAND2_X2 U10397 ( .A1(n6083), .A2(n10239), .ZN(n9345) );
  NAND2_X2 U10398 ( .A1(n6082), .A2(n9838), .ZN(n9344) );
  NAND4_X2 U10399 ( .A1(n9347), .A2(n9346), .A3(n9345), .A4(n9344), .ZN(n9491)
         );
  INV_X4 U10400 ( .A(n9491), .ZN(n9348) );
  NOR2_X4 U10401 ( .A1(n9350), .A2(n9349), .ZN(n9371) );
  AOI22_X2 U10402 ( .A1(n9353), .A2(n9352), .B1(
        \WIRE_ALU_A/MUX2TO1_32BIT[12].MUX/N1 ), .B2(n9351), .ZN(n9833) );
  XNOR2_X2 U10403 ( .A(n9354), .B(n10375), .ZN(n9832) );
  INV_X4 U10404 ( .A(n9832), .ZN(n9356) );
  XNOR2_X2 U10405 ( .A(n9357), .B(n10125), .ZN(n10132) );
  AOI22_X2 U10406 ( .A1(n10131), .A2(n10132), .B1(
        \WIRE_ALU_A/MUX2TO1_32BIT[10].MUX/N1 ), .B2(n9357), .ZN(n9511) );
  XNOR2_X2 U10407 ( .A(n9508), .B(n10382), .ZN(n9507) );
  XNOR2_X2 U10408 ( .A(n9511), .B(n9507), .ZN(n9368) );
  NAND2_X2 U10409 ( .A1(n8759), .A2(n9621), .ZN(n9365) );
  NAND2_X2 U10410 ( .A1(net77086), .A2(n9945), .ZN(n9364) );
  NAND2_X2 U10411 ( .A1(n6083), .A2(n9395), .ZN(n9363) );
  NAND2_X2 U10412 ( .A1(n6082), .A2(n9500), .ZN(n9362) );
  NAND4_X2 U10413 ( .A1(n9365), .A2(n9364), .A3(n9363), .A4(n9362), .ZN(n10126) );
  INV_X4 U10414 ( .A(n10126), .ZN(n9366) );
  INV_X4 U10415 ( .A(dmem_addr_out[9]), .ZN(n9377) );
  OAI22_X2 U10416 ( .A1(n5169), .A2(n6088), .B1(net76660), .B2(n6043), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10417 ( .A1(n5616), .A2(n6091), .B1(n6156), .B2(n6044), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10418 ( .A1(n6193), .A2(n5373), .B1(n6195), .B2(n6044), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10419 ( .A1(n6196), .A2(n5653), .B1(n6199), .B2(n6044), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10420 ( .A1(n5288), .A2(n6097), .B1(n6095), .B2(n6044), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10421 ( .A1(n5170), .A2(n6103), .B1(n6102), .B2(n6044), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10422 ( .A1(n4976), .A2(n6108), .B1(n6106), .B2(n6044), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10423 ( .A1(n5171), .A2(n6112), .B1(n6044), .B2(n6158), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10424 ( .A1(n5172), .A2(n6115), .B1(n6160), .B2(n6044), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10425 ( .A1(n5289), .A2(n6118), .B1(n6162), .B2(n6044), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10426 ( .A1(n6200), .A2(n5374), .B1(n6204), .B2(n6044), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10427 ( .A1(n5290), .A2(net76862), .B1(net76616), .B2(n6044), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10428 ( .A1(n6206), .A2(n5411), .B1(n6208), .B2(n6044), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10429 ( .A1(n5173), .A2(n6121), .B1(n6164), .B2(n6044), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10430 ( .A1(n5291), .A2(n6124), .B1(n6166), .B2(n6044), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10431 ( .A1(n5174), .A2(n6127), .B1(n6168), .B2(n6044), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10432 ( .A1(n5100), .A2(n6129), .B1(n6170), .B2(n6043), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10433 ( .A1(n5021), .A2(n6132), .B1(n6172), .B2(n6043), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10434 ( .A1(n5175), .A2(n6136), .B1(n6174), .B2(n6043), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10435 ( .A1(n6210), .A2(n5412), .B1(n6212), .B2(n6043), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10436 ( .A1(\REGFILE/reg_out[28][9] ), .A2(n6177), .ZN(n9379) );
  NAND2_X2 U10437 ( .A1(n6178), .A2(\REGFILE/reg_out[29][9] ), .ZN(n9380) );
  OAI22_X2 U10438 ( .A1(n5022), .A2(n6139), .B1(net76550), .B2(n6043), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10439 ( .A1(n6180), .A2(\REGFILE/reg_out[30][9] ), .ZN(n9381) );
  NAND2_X2 U10440 ( .A1(n5688), .A2(\REGFILE/reg_out[31][9] ), .ZN(n9382) );
  OAI22_X2 U10441 ( .A1(n6216), .A2(n5112), .B1(net76320), .B2(n6043), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10442 ( .A1(n6218), .A2(n5375), .B1(n6220), .B2(n6043), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10443 ( .A1(n5292), .A2(n6144), .B1(n6183), .B2(n6043), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10444 ( .A1(n5293), .A2(net76706), .B1(n6147), .B2(n6043), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10445 ( .A1(n5176), .A2(net76692), .B1(n6185), .B2(n6043), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10446 ( .A1(n5294), .A2(n6150), .B1(n6187), .B2(n6043), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10447 ( .A1(n5177), .A2(n6153), .B1(n6189), .B2(n6044), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[9].REGISTER1/STORE_DATA/N3 ) );
  XNOR2_X2 U10448 ( .A(n9385), .B(n9384), .ZN(n9387) );
  NAND2_X2 U10449 ( .A1(n6190), .A2(n10139), .ZN(n9386) );
  OAI221_X2 U10450 ( .B1(n10125), .B2(n4962), .C1(n6008), .C2(n9387), .A(n9386), .ZN(\PCLOGIC/PC_REG/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  XOR2_X2 U10451 ( .A(n9389), .B(n9388), .Z(n9391) );
  NAND2_X2 U10452 ( .A1(n6190), .A2(n9422), .ZN(n9390) );
  OAI221_X2 U10453 ( .B1(n10368), .B2(n4962), .C1(n9391), .C2(n9533), .A(n9390), .ZN(\PCLOGIC/PC_REG/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10454 ( .A1(multOut[13]), .A2(net92392), .ZN(n9420) );
  XNOR2_X2 U10455 ( .A(n9393), .B(n9392), .ZN(n9394) );
  NAND2_X2 U10456 ( .A1(net71271), .A2(n9394), .ZN(n9419) );
  NAND2_X2 U10457 ( .A1(n10102), .A2(n9395), .ZN(n9401) );
  NAND2_X2 U10458 ( .A1(net77086), .A2(n9500), .ZN(n9400) );
  NAND2_X2 U10459 ( .A1(n6082), .A2(n9396), .ZN(n9399) );
  NAND2_X2 U10460 ( .A1(n6083), .A2(n9397), .ZN(n9398) );
  NAND4_X2 U10461 ( .A1(n9401), .A2(n9400), .A3(n9399), .A4(n9398), .ZN(n10248) );
  NAND2_X2 U10462 ( .A1(n10066), .A2(n9403), .ZN(n9406) );
  NAND2_X2 U10463 ( .A1(n10058), .A2(n9404), .ZN(n9405) );
  NAND2_X2 U10464 ( .A1(n9406), .A2(n9405), .ZN(n9416) );
  NAND2_X2 U10465 ( .A1(n4880), .A2(n9493), .ZN(n9412) );
  NAND2_X2 U10466 ( .A1(n6082), .A2(n9407), .ZN(n9411) );
  NAND2_X2 U10467 ( .A1(n8759), .A2(n9408), .ZN(n9410) );
  NAND2_X2 U10468 ( .A1(net77086), .A2(n9977), .ZN(n9409) );
  NAND4_X2 U10469 ( .A1(n9412), .A2(n9411), .A3(n9410), .A4(n9409), .ZN(n10246) );
  INV_X4 U10470 ( .A(n10246), .ZN(n9414) );
  NOR2_X4 U10471 ( .A1(n9416), .A2(n9415), .ZN(n9417) );
  NAND4_X2 U10472 ( .A1(n9420), .A2(n9419), .A3(n9418), .A4(n9417), .ZN(
        dmem_addr_out[13]) );
  NAND2_X2 U10473 ( .A1(net76650), .A2(dmem_addr_out[13]), .ZN(n9424) );
  INV_X4 U10474 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [29]), .ZN(n9816) );
  NAND3_X2 U10475 ( .A1(n9424), .A2(net70740), .A3(n9423), .ZN(n9425) );
  NAND2_X2 U10476 ( .A1(n6047), .A2(n4992), .ZN(n9428) );
  NAND2_X2 U10477 ( .A1(n4867), .A2(\REGFILE/reg_out[0][13] ), .ZN(n9427) );
  NAND2_X2 U10478 ( .A1(n9428), .A2(n9427), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10479 ( .A1(n6047), .A2(n4990), .ZN(n9430) );
  NAND2_X2 U10480 ( .A1(n9430), .A2(n9429), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10481 ( .A1(n6047), .A2(n4998), .ZN(n9432) );
  NAND2_X2 U10482 ( .A1(net148736), .A2(n4869), .ZN(n9431) );
  NAND2_X2 U10483 ( .A1(n9432), .A2(n9431), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10484 ( .A1(n6047), .A2(n4993), .ZN(n9434) );
  NAND2_X2 U10485 ( .A1(n9434), .A2(n9433), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10486 ( .A1(n6047), .A2(n6096), .ZN(n9436) );
  NAND2_X2 U10487 ( .A1(n6100), .A2(\REGFILE/reg_out[13][13] ), .ZN(n9435) );
  NAND2_X2 U10488 ( .A1(n9436), .A2(n9435), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10489 ( .A1(n6047), .A2(n6101), .ZN(n9438) );
  NAND2_X2 U10490 ( .A1(n9438), .A2(n9437), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10491 ( .A1(n6047), .A2(n6107), .ZN(n9440) );
  NAND2_X2 U10492 ( .A1(n4804), .A2(\REGFILE/reg_out[15][13] ), .ZN(n9439) );
  NAND2_X2 U10493 ( .A1(n9440), .A2(n9439), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10494 ( .A1(n6047), .A2(n4994), .ZN(n9442) );
  NAND2_X2 U10495 ( .A1(n9442), .A2(n9441), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10496 ( .A1(n6047), .A2(n4999), .ZN(n9444) );
  NAND2_X2 U10497 ( .A1(n4892), .A2(\REGFILE/reg_out[17][13] ), .ZN(n9443) );
  NAND2_X2 U10498 ( .A1(n9444), .A2(n9443), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10499 ( .A1(n6047), .A2(n5000), .ZN(n9446) );
  NAND2_X2 U10500 ( .A1(n4884), .A2(\REGFILE/reg_out[18][13] ), .ZN(n9445) );
  NAND2_X2 U10501 ( .A1(n9446), .A2(n9445), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10502 ( .A1(n6046), .A2(n5001), .ZN(n9448) );
  NAND2_X2 U10503 ( .A1(\REGFILE/reg_out[19][13] ), .A2(n4876), .ZN(n9447) );
  NAND2_X2 U10504 ( .A1(n9448), .A2(n9447), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10505 ( .A1(n6046), .A2(n4997), .ZN(n9450) );
  NAND2_X2 U10506 ( .A1(n9450), .A2(n9449), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10507 ( .A1(n6046), .A2(n4903), .ZN(n9452) );
  NAND2_X2 U10508 ( .A1(\REGFILE/reg_out[20][13] ), .A2(n4868), .ZN(n9451) );
  NAND2_X2 U10509 ( .A1(n9452), .A2(n9451), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10510 ( .A1(n6046), .A2(n4904), .ZN(n9454) );
  NAND2_X2 U10511 ( .A1(n4882), .A2(\REGFILE/reg_out[21][13] ), .ZN(n9453) );
  NAND2_X2 U10512 ( .A1(n9454), .A2(n9453), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10513 ( .A1(n6046), .A2(n4905), .ZN(n9456) );
  NAND2_X2 U10514 ( .A1(n4888), .A2(\REGFILE/reg_out[22][13] ), .ZN(n9455) );
  NAND2_X2 U10515 ( .A1(n9456), .A2(n9455), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10516 ( .A1(n6046), .A2(n4906), .ZN(n9458) );
  NAND2_X2 U10517 ( .A1(n4883), .A2(\REGFILE/reg_out[23][13] ), .ZN(n9457) );
  NAND2_X2 U10518 ( .A1(n9458), .A2(n9457), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10519 ( .A1(n6046), .A2(n4995), .ZN(n9460) );
  NAND2_X2 U10520 ( .A1(n9460), .A2(n9459), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10521 ( .A1(n6046), .A2(n5002), .ZN(n9462) );
  NAND2_X2 U10522 ( .A1(n4878), .A2(\REGFILE/reg_out[25][13] ), .ZN(n9461) );
  NAND2_X2 U10523 ( .A1(n9462), .A2(n9461), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10524 ( .A1(n6046), .A2(n5003), .ZN(n9464) );
  NAND2_X2 U10525 ( .A1(n9464), .A2(n9463), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10526 ( .A1(n6046), .A2(n5004), .ZN(n9466) );
  NAND2_X2 U10527 ( .A1(\REGFILE/reg_out[27][13] ), .A2(n4872), .ZN(n9465) );
  NAND2_X2 U10528 ( .A1(n9466), .A2(n9465), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10529 ( .A1(n6046), .A2(n4806), .ZN(n9468) );
  NAND2_X2 U10530 ( .A1(n9468), .A2(n9467), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10531 ( .A1(n6046), .A2(n10607), .ZN(n9470) );
  NAND2_X2 U10532 ( .A1(n6178), .A2(\REGFILE/reg_out[29][13] ), .ZN(n9469) );
  NAND2_X2 U10533 ( .A1(n9470), .A2(n9469), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10534 ( .A1(n6047), .A2(n5005), .ZN(n9472) );
  NAND2_X2 U10535 ( .A1(n9472), .A2(n9471), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10536 ( .A1(n6046), .A2(n10614), .ZN(n9474) );
  NAND2_X2 U10537 ( .A1(n9474), .A2(n9473), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10538 ( .A1(n6047), .A2(net70574), .ZN(n9476) );
  NAND2_X2 U10539 ( .A1(n5688), .A2(\REGFILE/reg_out[31][13] ), .ZN(n9475) );
  NAND2_X2 U10540 ( .A1(n9476), .A2(n9475), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10541 ( .A1(n6047), .A2(n5009), .ZN(n9478) );
  NAND2_X2 U10542 ( .A1(\REGFILE/reg_out[3][13] ), .A2(n4871), .ZN(n9477) );
  NAND2_X2 U10543 ( .A1(n9478), .A2(n9477), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10544 ( .A1(n6046), .A2(n4996), .ZN(n9480) );
  NAND2_X2 U10545 ( .A1(\REGFILE/reg_out[4][13] ), .A2(n4870), .ZN(n9479) );
  NAND2_X2 U10546 ( .A1(n9480), .A2(n9479), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10547 ( .A1(n6046), .A2(n5006), .ZN(n9482) );
  NAND2_X2 U10548 ( .A1(n4885), .A2(\REGFILE/reg_out[5][13] ), .ZN(n9481) );
  NAND2_X2 U10549 ( .A1(n9482), .A2(n9481), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10550 ( .A1(n6047), .A2(n6148), .ZN(n9484) );
  NAND2_X2 U10551 ( .A1(n4889), .A2(\REGFILE/reg_out[6][13] ), .ZN(n9483) );
  NAND2_X2 U10552 ( .A1(n9484), .A2(n9483), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10553 ( .A1(n6046), .A2(n5007), .ZN(n9486) );
  NAND2_X2 U10554 ( .A1(n4886), .A2(\REGFILE/reg_out[7][13] ), .ZN(n9485) );
  NAND2_X2 U10555 ( .A1(n9486), .A2(n9485), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10556 ( .A1(n6047), .A2(n4991), .ZN(n9488) );
  NAND2_X2 U10557 ( .A1(n9488), .A2(n9487), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10558 ( .A1(n6047), .A2(n5008), .ZN(n9490) );
  NAND2_X2 U10559 ( .A1(n4887), .A2(\REGFILE/reg_out[9][13] ), .ZN(n9489) );
  NAND2_X2 U10560 ( .A1(n9490), .A2(n9489), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[13].REGISTER1/STORE_DATA/N3 ) );
  AOI22_X2 U10561 ( .A1(net71092), .A2(n9492), .B1(net71094), .B2(n9491), .ZN(
        n9505) );
  NAND2_X2 U10562 ( .A1(n6082), .A2(n9935), .ZN(n9497) );
  NAND2_X2 U10563 ( .A1(n4880), .A2(n10091), .ZN(n9496) );
  NAND2_X2 U10564 ( .A1(n10102), .A2(n9585), .ZN(n9495) );
  NAND2_X2 U10565 ( .A1(net77086), .A2(n9493), .ZN(n9494) );
  NAND4_X2 U10566 ( .A1(n9497), .A2(n9496), .A3(n9495), .A4(n9494), .ZN(n9690)
         );
  NAND2_X2 U10567 ( .A1(n10280), .A2(n9690), .ZN(n9504) );
  OAI211_X2 U10568 ( .C1(net72312), .C2(net70868), .A(n9499), .B(n9498), .ZN(
        n10103) );
  AOI22_X2 U10569 ( .A1(net77084), .A2(n10103), .B1(n8728), .B2(n9945), .ZN(
        n9502) );
  AOI22_X2 U10570 ( .A1(n6082), .A2(n9621), .B1(n6083), .B2(n9500), .ZN(n9501)
         );
  NAND2_X2 U10571 ( .A1(n9502), .A2(n9501), .ZN(n9685) );
  INV_X4 U10572 ( .A(n10419), .ZN(n10387) );
  NAND3_X2 U10573 ( .A1(n9505), .A2(n9504), .A3(n9503), .ZN(n9506) );
  INV_X4 U10575 ( .A(n9507), .ZN(n9510) );
  NAND2_X2 U10576 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[9].MUX/N1 ), .A2(n9508), 
        .ZN(n9509) );
  XNOR2_X2 U10577 ( .A(n9610), .B(n9611), .ZN(n9513) );
  NAND2_X2 U10578 ( .A1(net71078), .A2(\WIRE_ALU_A/MUX2TO1_32BIT[8].MUX/N1 ), 
        .ZN(n9512) );
  NOR2_X4 U10579 ( .A1(n9515), .A2(n9514), .ZN(n9519) );
  OAI22_X2 U10581 ( .A1(n5977), .A2(n6091), .B1(n6156), .B2(n6049), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10582 ( .A1(n6193), .A2(n5376), .B1(n6195), .B2(n6049), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U10583 ( .A(\REGFILE/reg_out[12][8] ), .ZN(n9521) );
  OAI22_X2 U10584 ( .A1(n6196), .A2(n9521), .B1(n6199), .B2(n6049), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10585 ( .A1(n5295), .A2(n6097), .B1(n6095), .B2(n6049), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10586 ( .A1(n5178), .A2(n6103), .B1(n6102), .B2(n6049), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10587 ( .A1(n5910), .A2(n6108), .B1(n6106), .B2(n6049), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10588 ( .A1(n5179), .A2(n6112), .B1(n6158), .B2(n6048), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10589 ( .A1(n5180), .A2(n6115), .B1(n6160), .B2(n4801), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10590 ( .A1(n5296), .A2(n6118), .B1(n6162), .B2(n6048), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10591 ( .A1(n6200), .A2(n5377), .B1(n6204), .B2(n6049), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10592 ( .A1(n5297), .A2(net76862), .B1(net76616), .B2(n4801), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10593 ( .A1(n6206), .A2(n5413), .B1(n6208), .B2(n6049), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10594 ( .A1(n5181), .A2(n6121), .B1(n6164), .B2(n6048), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10595 ( .A1(n5298), .A2(n6124), .B1(n6166), .B2(n4801), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10596 ( .A1(n5182), .A2(n6127), .B1(n6168), .B2(n6049), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10597 ( .A1(n5183), .A2(n6129), .B1(n6170), .B2(n6048), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10598 ( .A1(n5869), .A2(n6132), .B1(n6172), .B2(n6048), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10599 ( .A1(n5184), .A2(n6136), .B1(n6174), .B2(n6048), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10600 ( .A1(n6210), .A2(n5978), .B1(n6212), .B2(n4801), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10601 ( .A1(\REGFILE/reg_out[28][8] ), .A2(n6175), .ZN(n9522) );
  NAND2_X2 U10602 ( .A1(n6178), .A2(\REGFILE/reg_out[29][8] ), .ZN(n9523) );
  OAI22_X2 U10603 ( .A1(n9524), .A2(n6139), .B1(net76550), .B2(n4801), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10604 ( .A1(n6180), .A2(\REGFILE/reg_out[30][8] ), .ZN(n9525) );
  NAND2_X2 U10605 ( .A1(n5688), .A2(\REGFILE/reg_out[31][8] ), .ZN(n9526) );
  OAI22_X2 U10606 ( .A1(n6216), .A2(n5028), .B1(net76320), .B2(n4801), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10607 ( .A1(n6218), .A2(n5378), .B1(n6220), .B2(n6048), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U10608 ( .A(\REGFILE/reg_out[5][8] ), .ZN(n9527) );
  OAI22_X2 U10609 ( .A1(n9527), .A2(n6144), .B1(n6183), .B2(n6048), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10610 ( .A1(n5079), .A2(net76706), .B1(n6147), .B2(n4801), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10611 ( .A1(n5101), .A2(net76692), .B1(n6185), .B2(n4801), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10612 ( .A1(n4972), .A2(n6150), .B1(n6187), .B2(n4801), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10613 ( .A1(n5102), .A2(n6153), .B1(n6189), .B2(n6049), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  XOR2_X2 U10614 ( .A(n9530), .B(n9529), .Z(n9534) );
  NAND2_X2 U10615 ( .A1(n6190), .A2(n9531), .ZN(n9532) );
  OAI221_X2 U10616 ( .B1(n9535), .B2(n4962), .C1(n9534), .C2(n6008), .A(n9532), 
        .ZN(\PCLOGIC/PC_REG/REG_32BIT[8].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10617 ( .A1(net73708), .A2(n10933), .ZN(n9541) );
  OAI211_X2 U10618 ( .C1(n8357), .C2(n9538), .A(n9537), .B(n10649), .ZN(n9540)
         );
  NAND2_X2 U10619 ( .A1(n6190), .A2(n9569), .ZN(n9539) );
  XNOR2_X2 U10620 ( .A(n9543), .B(n9542), .ZN(n9545) );
  INV_X4 U10621 ( .A(n10431), .ZN(n10343) );
  NAND2_X2 U10622 ( .A1(multOut[21]), .A2(net92392), .ZN(n9564) );
  NAND2_X2 U10623 ( .A1(n10102), .A2(n9546), .ZN(n9551) );
  NAND2_X2 U10624 ( .A1(net77086), .A2(n9547), .ZN(n9550) );
  AOI22_X2 U10625 ( .A1(n6082), .A2(n9548), .B1(n6083), .B2(n10233), .ZN(n9549) );
  NAND2_X2 U10626 ( .A1(n10058), .A2(n10059), .ZN(n9554) );
  NAND2_X2 U10627 ( .A1(n10060), .A2(n9552), .ZN(n9553) );
  NAND2_X2 U10628 ( .A1(n9554), .A2(n9553), .ZN(n9562) );
  NAND2_X2 U10629 ( .A1(n10064), .A2(n9982), .ZN(n9556) );
  NAND2_X2 U10630 ( .A1(n10066), .A2(n10063), .ZN(n9555) );
  NAND2_X2 U10631 ( .A1(n9556), .A2(n9555), .ZN(n9557) );
  MUX2_X2 U10632 ( .A(n9558), .B(n9557), .S(net71026), .Z(n9561) );
  NAND3_X2 U10633 ( .A1(n9565), .A2(n9564), .A3(n9563), .ZN(dmem_addr_out[21])
         );
  INV_X4 U10634 ( .A(dmem_addr_out[21]), .ZN(n9572) );
  INV_X4 U10635 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [21]), .ZN(n9817) );
  INV_X4 U10636 ( .A(dmem_read_in[21]), .ZN(n9567) );
  OAI211_X2 U10637 ( .C1(n9572), .C2(net76646), .A(n9571), .B(n9570), .ZN(
        n9573) );
  OAI22_X2 U10638 ( .A1(n5185), .A2(n6089), .B1(net76658), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U10639 ( .A(\REGFILE/reg_out[10][21] ), .ZN(n9574) );
  OAI22_X2 U10640 ( .A1(n9574), .A2(n6092), .B1(n6155), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10641 ( .A1(n6192), .A2(n5379), .B1(n6195), .B2(n9579), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10642 ( .A1(n6196), .A2(n5810), .B1(n6199), .B2(n9579), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10643 ( .A1(n5299), .A2(n6098), .B1(n6095), .B2(n9579), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10644 ( .A1(n5186), .A2(n6104), .B1(n6102), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10645 ( .A1(n5300), .A2(n6109), .B1(n6106), .B2(n9579), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10646 ( .A1(n5187), .A2(n6113), .B1(n6157), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10647 ( .A1(n5188), .A2(n6116), .B1(n6159), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10648 ( .A1(n5301), .A2(n6119), .B1(n6161), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10649 ( .A1(n6200), .A2(n5380), .B1(n6204), .B2(n9579), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10650 ( .A1(n5302), .A2(net76864), .B1(net76614), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10651 ( .A1(n6205), .A2(n5505), .B1(n6208), .B2(n9579), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10652 ( .A1(n5189), .A2(n6122), .B1(n6163), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10653 ( .A1(n5303), .A2(n6125), .B1(n6165), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10654 ( .A1(n5190), .A2(n6128), .B1(n6167), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10655 ( .A1(n5191), .A2(n6130), .B1(n6169), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10656 ( .A1(n5807), .A2(n6133), .B1(n6171), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10657 ( .A1(n5192), .A2(n6137), .B1(n6173), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10658 ( .A1(n6209), .A2(n5034), .B1(n6212), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10659 ( .A1(\REGFILE/reg_out[28][21] ), .A2(n6175), .ZN(n9575) );
  OAI21_X4 U10660 ( .B1(n6213), .B2(n6051), .A(n9575), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10661 ( .A1(n6178), .A2(\REGFILE/reg_out[29][21] ), .ZN(n9576) );
  OAI21_X4 U10662 ( .B1(n6138), .B2(n6051), .A(n9576), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10663 ( .A1(n5304), .A2(n6140), .B1(net76548), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10664 ( .A1(n6180), .A2(\REGFILE/reg_out[30][21] ), .ZN(n9577) );
  OAI21_X4 U10665 ( .B1(n6142), .B2(n6051), .A(n9577), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10666 ( .A1(n5688), .A2(\REGFILE/reg_out[31][21] ), .ZN(n9578) );
  OAI21_X4 U10667 ( .B1(net76480), .B2(n6051), .A(n9578), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10668 ( .A1(n6215), .A2(n5414), .B1(net76320), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10669 ( .A1(n6217), .A2(n5499), .B1(n6220), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10670 ( .A1(n5305), .A2(n6145), .B1(n6182), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10671 ( .A1(n5306), .A2(net76708), .B1(n6147), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10672 ( .A1(n5193), .A2(net76694), .B1(n6184), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10673 ( .A1(n5307), .A2(n6151), .B1(n6186), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10674 ( .A1(n5194), .A2(n6154), .B1(n6188), .B2(n6051), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[21].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10675 ( .A1(net77086), .A2(n9844), .ZN(n9584) );
  NAND2_X2 U10676 ( .A1(n6082), .A2(net70727), .ZN(n9583) );
  INV_X4 U10677 ( .A(n9934), .ZN(n9590) );
  NAND2_X2 U10678 ( .A1(n8759), .A2(n9935), .ZN(n9588) );
  NAND2_X2 U10679 ( .A1(n6082), .A2(n10091), .ZN(n9587) );
  INV_X4 U10680 ( .A(n9655), .ZN(n9589) );
  OAI22_X2 U10681 ( .A1(n10474), .A2(n9590), .B1(n10472), .B2(n9589), .ZN(
        n9592) );
  NAND2_X2 U10682 ( .A1(n10931), .A2(net70720), .ZN(n9596) );
  NAND2_X2 U10683 ( .A1(net70719), .A2(net80189), .ZN(n9595) );
  NAND4_X2 U10684 ( .A1(n9596), .A2(n9595), .A3(n9594), .A4(n9593), .ZN(n10023) );
  NAND2_X2 U10685 ( .A1(n10102), .A2(n10023), .ZN(n9604) );
  NAND2_X2 U10686 ( .A1(n10933), .A2(net70720), .ZN(n9600) );
  NAND4_X2 U10687 ( .A1(n9600), .A2(n9599), .A3(n9598), .A4(n9597), .ZN(n10158) );
  NAND2_X2 U10688 ( .A1(net77086), .A2(n10158), .ZN(n9603) );
  NAND2_X2 U10689 ( .A1(n6083), .A2(n9839), .ZN(n9602) );
  NAND2_X2 U10690 ( .A1(n6082), .A2(n10024), .ZN(n9601) );
  NAND4_X2 U10691 ( .A1(n9604), .A2(n9603), .A3(n9602), .A4(n9601), .ZN(n9933)
         );
  INV_X4 U10692 ( .A(n9933), .ZN(n9605) );
  NOR2_X4 U10693 ( .A1(n9608), .A2(n9607), .ZN(n9631) );
  AOI22_X2 U10695 ( .A1(n9611), .A2(n9610), .B1(
        \WIRE_ALU_A/MUX2TO1_32BIT[8].MUX/N1 ), .B2(n9609), .ZN(n9683) );
  XNOR2_X2 U10696 ( .A(n9612), .B(n10464), .ZN(n9682) );
  INV_X4 U10697 ( .A(n9682), .ZN(n9614) );
  NAND2_X2 U10698 ( .A1(\WIRE_ALU_A/MUX2TO1_32BIT[7].MUX/N1 ), .A2(n9612), 
        .ZN(n9613) );
  AOI22_X2 U10699 ( .A1(n9663), .A2(n9664), .B1(
        \WIRE_ALU_A/MUX2TO1_32BIT[6].MUX/N1 ), .B2(n9615), .ZN(n9959) );
  XNOR2_X2 U10700 ( .A(n9956), .B(n10396), .ZN(n9955) );
  XNOR2_X2 U10701 ( .A(n9959), .B(n9955), .ZN(n9628) );
  NAND2_X2 U10702 ( .A1(n8759), .A2(n10103), .ZN(n9625) );
  NAND2_X2 U10703 ( .A1(n10932), .A2(net70720), .ZN(n9620) );
  NAND4_X2 U10704 ( .A1(n9620), .A2(n9619), .A3(n9618), .A4(n9617), .ZN(n10101) );
  NAND2_X2 U10705 ( .A1(net77086), .A2(n10101), .ZN(n9624) );
  NAND2_X2 U10706 ( .A1(n4880), .A2(n9621), .ZN(n9623) );
  NAND2_X2 U10707 ( .A1(n6082), .A2(n9945), .ZN(n9622) );
  NAND4_X2 U10708 ( .A1(n9625), .A2(n9624), .A3(n9623), .A4(n9622), .ZN(n9658)
         );
  INV_X4 U10709 ( .A(n9658), .ZN(n9626) );
  OAI22_X2 U10712 ( .A1(n5515), .A2(n6089), .B1(n6053), .B2(net76658), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10713 ( .A1(n5043), .A2(n6092), .B1(n6054), .B2(n6155), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10716 ( .A1(n6196), .A2(n5660), .B1(n6054), .B2(n6199), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10717 ( .A1(n5308), .A2(n6098), .B1(n6054), .B2(n6095), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10720 ( .A1(n5309), .A2(n6109), .B1(n6054), .B2(n6106), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10722 ( .A1(n5196), .A2(n6116), .B1(n6054), .B2(n6159), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10723 ( .A1(n5310), .A2(n6119), .B1(n6054), .B2(n6161), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10724 ( .A1(n6200), .A2(n5381), .B1(n6054), .B2(n6204), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10725 ( .A1(n5311), .A2(net76864), .B1(n6054), .B2(net76614), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10726 ( .A1(n6205), .A2(n5415), .B1(n6054), .B2(n6208), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10727 ( .A1(n5197), .A2(n6122), .B1(n6054), .B2(n6163), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10728 ( .A1(n5312), .A2(n6125), .B1(n6054), .B2(n6165), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10729 ( .A1(n5198), .A2(n6128), .B1(n6054), .B2(n6167), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10732 ( .A1(n5313), .A2(n6133), .B1(n6053), .B2(n6171), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10734 ( .A1(n9641), .A2(n6137), .B1(n6053), .B2(n6173), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10735 ( .A1(n6210), .A2(n5416), .B1(n6053), .B2(n6212), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10736 ( .A1(\REGFILE/reg_out[28][5] ), .A2(n6175), .ZN(n9642) );
  NAND2_X2 U10737 ( .A1(n6178), .A2(\REGFILE/reg_out[29][5] ), .ZN(n9643) );
  OAI22_X2 U10738 ( .A1(n4984), .A2(n6140), .B1(n6053), .B2(net76548), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10739 ( .A1(n6180), .A2(\REGFILE/reg_out[30][5] ), .ZN(n9644) );
  NAND2_X2 U10740 ( .A1(n5688), .A2(\REGFILE/reg_out[31][5] ), .ZN(n9645) );
  OAI22_X2 U10741 ( .A1(n6216), .A2(n4985), .B1(n6053), .B2(net76320), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10742 ( .A1(n6217), .A2(n5554), .B1(n6053), .B2(n6220), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10743 ( .A1(n5044), .A2(n6145), .B1(n6053), .B2(n6182), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10744 ( .A1(n5451), .A2(net76708), .B1(n6053), .B2(n6147), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10745 ( .A1(n5516), .A2(net76694), .B1(n6053), .B2(n6184), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10746 ( .A1(n5314), .A2(n6151), .B1(n6053), .B2(n6186), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10747 ( .A1(n5199), .A2(n6154), .B1(n6054), .B2(n6188), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10748 ( .A1(n10102), .A2(n9844), .ZN(n9650) );
  NAND2_X2 U10749 ( .A1(n4880), .A2(net70727), .ZN(n9649) );
  NAND2_X2 U10750 ( .A1(net77086), .A2(n9845), .ZN(n9648) );
  NAND2_X2 U10751 ( .A1(n6082), .A2(n10013), .ZN(n9647) );
  NAND4_X2 U10752 ( .A1(n9650), .A2(n9649), .A3(n9648), .A4(n9647), .ZN(n9687)
         );
  NAND2_X2 U10753 ( .A1(n8759), .A2(n10024), .ZN(n9654) );
  NAND2_X2 U10754 ( .A1(net77086), .A2(n10023), .ZN(n9653) );
  NAND2_X2 U10755 ( .A1(n6083), .A2(n9838), .ZN(n9652) );
  NAND2_X2 U10756 ( .A1(n6082), .A2(n9839), .ZN(n9651) );
  NAND4_X2 U10757 ( .A1(n9654), .A2(n9653), .A3(n9652), .A4(n9651), .ZN(n9686)
         );
  AOI22_X2 U10758 ( .A1(net71092), .A2(n9687), .B1(net71094), .B2(n9686), .ZN(
        n9661) );
  NAND2_X2 U10759 ( .A1(n10280), .A2(n9655), .ZN(n9660) );
  INV_X4 U10760 ( .A(n9657), .ZN(n10394) );
  AOI21_X4 U10761 ( .B1(net71085), .B2(n9658), .A(n5052), .ZN(n9659) );
  NAND3_X2 U10762 ( .A1(n9661), .A2(n9660), .A3(n9659), .ZN(n9662) );
  XNOR2_X2 U10763 ( .A(n9664), .B(n9663), .ZN(n9666) );
  NAND2_X2 U10764 ( .A1(net71078), .A2(\WIRE_ALU_A/MUX2TO1_32BIT[6].MUX/N1 ), 
        .ZN(n9665) );
  NOR2_X4 U10765 ( .A1(n9668), .A2(n9667), .ZN(n9673) );
  OAI22_X2 U10766 ( .A1(n5437), .A2(n6089), .B1(n4802), .B2(net76658), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10768 ( .A1(n9675), .A2(n6092), .B1(n4802), .B2(n6155), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10769 ( .A1(n6193), .A2(n5382), .B1(n4802), .B2(n6194), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10770 ( .A1(n6197), .A2(n5417), .B1(n6057), .B2(n6198), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10771 ( .A1(n5315), .A2(n6098), .B1(n6056), .B2(n6095), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10772 ( .A1(n5200), .A2(n6104), .B1(n6102), .B2(n6057), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10773 ( .A1(n4982), .A2(n6109), .B1(n6057), .B2(n6106), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10774 ( .A1(n5517), .A2(n6113), .B1(n6057), .B2(n6157), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10775 ( .A1(n5201), .A2(n6116), .B1(n6057), .B2(n6159), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10776 ( .A1(n5316), .A2(n6119), .B1(n6056), .B2(n6161), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10777 ( .A1(n6201), .A2(n5383), .B1(n6056), .B2(n6203), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10778 ( .A1(n5317), .A2(net76864), .B1(n4802), .B2(net76614), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10779 ( .A1(n6206), .A2(n5418), .B1(n4802), .B2(n6207), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10780 ( .A1(n5202), .A2(n6122), .B1(n6057), .B2(n6163), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10781 ( .A1(n5318), .A2(n6125), .B1(n6056), .B2(n6165), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10782 ( .A1(n5203), .A2(n6128), .B1(n6056), .B2(n6167), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10783 ( .A1(n5204), .A2(n6130), .B1(n6057), .B2(n6169), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U10784 ( .A(n5764), .ZN(n9676) );
  OAI22_X2 U10785 ( .A1(n9676), .A2(n6133), .B1(n6056), .B2(n6171), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10786 ( .A1(n5103), .A2(n6137), .B1(n6056), .B2(n6173), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10787 ( .A1(n6210), .A2(n5113), .B1(n4802), .B2(n6211), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10788 ( .A1(\REGFILE/reg_out[28][6] ), .A2(n6175), .ZN(n9677) );
  NAND2_X2 U10789 ( .A1(n6178), .A2(\REGFILE/reg_out[29][6] ), .ZN(n9678) );
  OAI22_X2 U10790 ( .A1(n5319), .A2(n6140), .B1(n4802), .B2(net76548), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10791 ( .A1(n6180), .A2(\REGFILE/reg_out[30][6] ), .ZN(n9679) );
  NAND2_X2 U10792 ( .A1(n5688), .A2(\REGFILE/reg_out[31][6] ), .ZN(n9680) );
  OAI22_X2 U10793 ( .A1(n6216), .A2(n5419), .B1(n6056), .B2(net76318), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10794 ( .A1(n6218), .A2(n5384), .B1(n6057), .B2(n6219), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10795 ( .A1(n5320), .A2(n6145), .B1(n6057), .B2(n6182), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10796 ( .A1(n5321), .A2(net76708), .B1(n4802), .B2(n6147), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10797 ( .A1(n5205), .A2(net76694), .B1(n6056), .B2(n6184), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10798 ( .A1(n5322), .A2(n6151), .B1(n4802), .B2(n6186), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10799 ( .A1(n5206), .A2(n6154), .B1(n6057), .B2(n6188), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ) );
  XNOR2_X2 U10801 ( .A(n9683), .B(n9682), .ZN(n9684) );
  NAND2_X2 U10802 ( .A1(net71271), .A2(n9684), .ZN(n9697) );
  INV_X4 U10803 ( .A(n10391), .ZN(n10307) );
  NAND2_X2 U10804 ( .A1(n10066), .A2(n9686), .ZN(n9689) );
  NAND2_X2 U10805 ( .A1(n10058), .A2(n9687), .ZN(n9688) );
  NAND2_X2 U10806 ( .A1(n9689), .A2(n9688), .ZN(n9694) );
  INV_X4 U10807 ( .A(n9690), .ZN(n9692) );
  NAND2_X2 U10808 ( .A1(n6060), .A2(n4992), .ZN(n9706) );
  NAND2_X2 U10809 ( .A1(n4867), .A2(\REGFILE/reg_out[0][7] ), .ZN(n9705) );
  NAND2_X2 U10810 ( .A1(n9706), .A2(n9705), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10811 ( .A1(n6060), .A2(n4990), .ZN(n9708) );
  NAND2_X2 U10812 ( .A1(n9708), .A2(n9707), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10813 ( .A1(n6059), .A2(n4998), .ZN(n9710) );
  NAND2_X2 U10814 ( .A1(\REGFILE/reg_out[11][7] ), .A2(n4869), .ZN(n9709) );
  NAND2_X2 U10815 ( .A1(n9710), .A2(n9709), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10816 ( .A1(n6060), .A2(n4993), .ZN(n9712) );
  NAND2_X2 U10817 ( .A1(\REGFILE/reg_out[12][7] ), .A2(n4873), .ZN(n9711) );
  NAND2_X2 U10818 ( .A1(n9712), .A2(n9711), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10819 ( .A1(n6060), .A2(n6096), .ZN(n9714) );
  NAND2_X2 U10820 ( .A1(n6100), .A2(\REGFILE/reg_out[13][7] ), .ZN(n9713) );
  NAND2_X2 U10821 ( .A1(n9714), .A2(n9713), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10822 ( .A1(n9765), .A2(n6101), .ZN(n9716) );
  NAND2_X2 U10823 ( .A1(n4805), .A2(\REGFILE/reg_out[14][7] ), .ZN(n9715) );
  NAND2_X2 U10824 ( .A1(n9716), .A2(n9715), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10825 ( .A1(n6059), .A2(n6107), .ZN(n9718) );
  NAND2_X2 U10826 ( .A1(n4804), .A2(\REGFILE/reg_out[15][7] ), .ZN(n9717) );
  NAND2_X2 U10827 ( .A1(n9718), .A2(n9717), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10828 ( .A1(n6060), .A2(n4994), .ZN(n9720) );
  NAND2_X2 U10829 ( .A1(n4891), .A2(\REGFILE/reg_out[16][7] ), .ZN(n9719) );
  NAND2_X2 U10830 ( .A1(n9720), .A2(n9719), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10831 ( .A1(n6060), .A2(n4999), .ZN(n9722) );
  NAND2_X2 U10832 ( .A1(n4892), .A2(\REGFILE/reg_out[17][7] ), .ZN(n9721) );
  NAND2_X2 U10833 ( .A1(n9722), .A2(n9721), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10834 ( .A1(n6060), .A2(n5000), .ZN(n9724) );
  NAND2_X2 U10835 ( .A1(n4884), .A2(\REGFILE/reg_out[18][7] ), .ZN(n9723) );
  NAND2_X2 U10836 ( .A1(n9724), .A2(n9723), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10837 ( .A1(n6060), .A2(n5001), .ZN(n9726) );
  NAND2_X2 U10838 ( .A1(\REGFILE/reg_out[19][7] ), .A2(n4876), .ZN(n9725) );
  NAND2_X2 U10839 ( .A1(n9726), .A2(n9725), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10840 ( .A1(n6060), .A2(n4997), .ZN(n9728) );
  NAND2_X2 U10841 ( .A1(n4877), .A2(\REGFILE/reg_out[1][7] ), .ZN(n9727) );
  NAND2_X2 U10842 ( .A1(n9728), .A2(n9727), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10843 ( .A1(n6060), .A2(n4903), .ZN(n9730) );
  NAND2_X2 U10844 ( .A1(\REGFILE/reg_out[20][7] ), .A2(n4868), .ZN(n9729) );
  NAND2_X2 U10845 ( .A1(n9730), .A2(n9729), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10846 ( .A1(n6060), .A2(n4904), .ZN(n9732) );
  NAND2_X2 U10847 ( .A1(n4882), .A2(\REGFILE/reg_out[21][7] ), .ZN(n9731) );
  NAND2_X2 U10848 ( .A1(n9732), .A2(n9731), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10849 ( .A1(n6060), .A2(n4905), .ZN(n9734) );
  NAND2_X2 U10850 ( .A1(n4888), .A2(\REGFILE/reg_out[22][7] ), .ZN(n9733) );
  NAND2_X2 U10851 ( .A1(n9734), .A2(n9733), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10852 ( .A1(n6060), .A2(n4906), .ZN(n9736) );
  NAND2_X2 U10853 ( .A1(n4883), .A2(\REGFILE/reg_out[23][7] ), .ZN(n9735) );
  NAND2_X2 U10854 ( .A1(n9736), .A2(n9735), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10855 ( .A1(n6060), .A2(n4995), .ZN(n9738) );
  NAND2_X2 U10856 ( .A1(n4875), .A2(\REGFILE/reg_out[24][7] ), .ZN(n9737) );
  NAND2_X2 U10857 ( .A1(n9738), .A2(n9737), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10858 ( .A1(n6060), .A2(n5002), .ZN(n9740) );
  NAND2_X2 U10859 ( .A1(n9740), .A2(n9739), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10860 ( .A1(n6060), .A2(n5003), .ZN(n9742) );
  NAND2_X2 U10861 ( .A1(n4893), .A2(\REGFILE/reg_out[26][7] ), .ZN(n9741) );
  NAND2_X2 U10862 ( .A1(n9742), .A2(n9741), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10863 ( .A1(n6060), .A2(n5004), .ZN(n9744) );
  NAND2_X2 U10864 ( .A1(n9744), .A2(n9743), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10865 ( .A1(n6060), .A2(n4806), .ZN(n9746) );
  NAND2_X2 U10866 ( .A1(\REGFILE/reg_out[28][7] ), .A2(n10604), .ZN(n9745) );
  NAND2_X2 U10867 ( .A1(n9746), .A2(n9745), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10868 ( .A1(n6059), .A2(n10607), .ZN(n9748) );
  NAND2_X2 U10869 ( .A1(n6178), .A2(\REGFILE/reg_out[29][7] ), .ZN(n9747) );
  NAND2_X2 U10870 ( .A1(n9748), .A2(n9747), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10871 ( .A1(n6059), .A2(n5005), .ZN(n9750) );
  NAND2_X2 U10872 ( .A1(n9750), .A2(n9749), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10873 ( .A1(n6059), .A2(n10614), .ZN(n9752) );
  NAND2_X2 U10874 ( .A1(n6180), .A2(\REGFILE/reg_out[30][7] ), .ZN(n9751) );
  NAND2_X2 U10875 ( .A1(n9752), .A2(n9751), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10876 ( .A1(n6059), .A2(net70574), .ZN(n9754) );
  NAND2_X2 U10877 ( .A1(n5688), .A2(\REGFILE/reg_out[31][7] ), .ZN(n9753) );
  NAND2_X2 U10878 ( .A1(n9754), .A2(n9753), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10879 ( .A1(n6059), .A2(n5009), .ZN(n9756) );
  NAND2_X2 U10880 ( .A1(\REGFILE/reg_out[3][7] ), .A2(n4871), .ZN(n9755) );
  NAND2_X2 U10881 ( .A1(n9756), .A2(n9755), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10882 ( .A1(n6059), .A2(n4996), .ZN(n9758) );
  NAND2_X2 U10883 ( .A1(\REGFILE/reg_out[4][7] ), .A2(n4870), .ZN(n9757) );
  NAND2_X2 U10884 ( .A1(n9758), .A2(n9757), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10885 ( .A1(n6059), .A2(n5006), .ZN(n9760) );
  NAND2_X2 U10886 ( .A1(n4885), .A2(\REGFILE/reg_out[5][7] ), .ZN(n9759) );
  NAND2_X2 U10887 ( .A1(n9760), .A2(n9759), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10888 ( .A1(n6059), .A2(n6148), .ZN(n9761) );
  NAND2_X2 U10889 ( .A1(n9761), .A2(net71936), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10890 ( .A1(n6059), .A2(n5007), .ZN(n9762) );
  NAND2_X2 U10891 ( .A1(n9762), .A2(net71934), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10892 ( .A1(n6059), .A2(n4991), .ZN(n9764) );
  NAND2_X2 U10893 ( .A1(n4890), .A2(\REGFILE/reg_out[8][7] ), .ZN(n9763) );
  NAND2_X2 U10894 ( .A1(n9764), .A2(n9763), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10895 ( .A1(n6059), .A2(n5008), .ZN(n9767) );
  NAND2_X2 U10896 ( .A1(n4887), .A2(\REGFILE/reg_out[9][7] ), .ZN(n9766) );
  NAND2_X2 U10897 ( .A1(n9767), .A2(n9766), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[7].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10898 ( .A1(multOut[26]), .A2(net92392), .ZN(n9787) );
  OAI22_X2 U10899 ( .A1(n9768), .A2(n10472), .B1(n5061), .B2(n10474), .ZN(
        n9773) );
  INV_X4 U10900 ( .A(n9774), .ZN(n9775) );
  NOR2_X4 U10901 ( .A1(n9775), .A2(net70691), .ZN(n9784) );
  INV_X4 U10902 ( .A(n9776), .ZN(n9779) );
  INV_X4 U10903 ( .A(n9777), .ZN(n9778) );
  NAND2_X2 U10904 ( .A1(n9779), .A2(n9778), .ZN(n9783) );
  INV_X4 U10905 ( .A(n10444), .ZN(n10325) );
  NAND2_X2 U10906 ( .A1(net70701), .A2(n10325), .ZN(n9781) );
  NAND2_X2 U10907 ( .A1(n9781), .A2(n9780), .ZN(n9782) );
  NAND3_X2 U10908 ( .A1(n9787), .A2(n9786), .A3(n9785), .ZN(dmem_addr_out[26])
         );
  INV_X4 U10909 ( .A(dmem_addr_out[26]), .ZN(n9794) );
  INV_X4 U10910 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [26]), .ZN(n10137) );
  INV_X4 U10911 ( .A(dmem_read_in[26]), .ZN(n9789) );
  OAI211_X2 U10912 ( .C1(n9794), .C2(net76646), .A(n9793), .B(n9792), .ZN(
        n9795) );
  NAND2_X2 U10913 ( .A1(net76270), .A2(n9795), .ZN(n9800) );
  OAI22_X2 U10914 ( .A1(n5518), .A2(n6089), .B1(net76658), .B2(n6062), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10915 ( .A1(n5452), .A2(n6092), .B1(n6155), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10916 ( .A1(n6193), .A2(n5555), .B1(n6194), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10917 ( .A1(n6197), .A2(n5503), .B1(n6198), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10918 ( .A1(n5323), .A2(n6098), .B1(n6095), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10919 ( .A1(n5207), .A2(n6104), .B1(n6102), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10920 ( .A1(n5324), .A2(n6109), .B1(n6106), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10921 ( .A1(n5208), .A2(n6113), .B1(n6157), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10922 ( .A1(n5519), .A2(n6116), .B1(n6159), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10923 ( .A1(n5453), .A2(n6119), .B1(n6161), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10924 ( .A1(n6201), .A2(n5385), .B1(n6203), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10925 ( .A1(n5325), .A2(net76864), .B1(net76614), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10926 ( .A1(n6206), .A2(n5420), .B1(n6207), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10927 ( .A1(n5209), .A2(n6122), .B1(n6163), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10928 ( .A1(n5326), .A2(n6125), .B1(n6165), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10929 ( .A1(n5210), .A2(n6128), .B1(n6167), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10930 ( .A1(n5211), .A2(n6130), .B1(n6169), .B2(n6062), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10931 ( .A1(n5327), .A2(n6133), .B1(n6171), .B2(n6062), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10932 ( .A1(n5212), .A2(n6137), .B1(n6173), .B2(n6062), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10933 ( .A1(n6210), .A2(n5421), .B1(n6211), .B2(n6062), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10934 ( .A1(\REGFILE/reg_out[28][26] ), .A2(n6175), .ZN(n9796) );
  OAI21_X4 U10935 ( .B1(n6214), .B2(n6062), .A(n9796), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10936 ( .A1(n6178), .A2(\REGFILE/reg_out[29][26] ), .ZN(n9797) );
  OAI21_X4 U10937 ( .B1(n10532), .B2(n6062), .A(n9797), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10938 ( .A1(n5454), .A2(n6140), .B1(net76548), .B2(n6062), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10939 ( .A1(n6180), .A2(\REGFILE/reg_out[30][26] ), .ZN(n9798) );
  OAI21_X4 U10940 ( .B1(n10534), .B2(n6062), .A(n9798), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10941 ( .A1(n5688), .A2(\REGFILE/reg_out[31][26] ), .ZN(n9799) );
  OAI21_X4 U10942 ( .B1(net70509), .B2(n6062), .A(n9799), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10943 ( .A1(n6216), .A2(n5422), .B1(net76318), .B2(n6062), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10944 ( .A1(n6218), .A2(n5556), .B1(n6219), .B2(n6062), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10945 ( .A1(n5455), .A2(n6145), .B1(n6182), .B2(n6062), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10946 ( .A1(n5456), .A2(net76708), .B1(n6147), .B2(n6062), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10947 ( .A1(n5520), .A2(net76694), .B1(n6184), .B2(n6062), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10948 ( .A1(n5457), .A2(n6151), .B1(n6186), .B2(n6062), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10949 ( .A1(n5521), .A2(n6154), .B1(n6188), .B2(n6063), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10950 ( .A1(n4922), .A2(n9802), .B1(n9801), .B2(n10472), .ZN(n9808) );
  OAI22_X2 U10951 ( .A1(net70710), .A2(n9805), .B1(n9804), .B2(n9803), .ZN(
        n9807) );
  AOI211_X4 U10952 ( .C1(n9808), .C2(net70697), .A(n9807), .B(n9806), .ZN(
        n9815) );
  NAND2_X2 U10953 ( .A1(multOut[29]), .A2(net92392), .ZN(n9814) );
  XNOR2_X2 U10954 ( .A(n9810), .B(n9809), .ZN(n9812) );
  INV_X4 U10955 ( .A(dmem_addr_out[29]), .ZN(n9825) );
  INV_X4 U10956 ( .A(dmem_read_in[29]), .ZN(n9820) );
  OAI211_X2 U10957 ( .C1(n9825), .C2(net76646), .A(n9824), .B(n9823), .ZN(
        n9826) );
  OAI22_X2 U10958 ( .A1(n5522), .A2(n6089), .B1(n6222), .B2(net76658), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10959 ( .A1(n5458), .A2(n6092), .B1(n6222), .B2(n6155), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10960 ( .A1(n5328), .A2(n6098), .B1(n6222), .B2(n6094), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U10961 ( .A(\REGFILE/reg_out[14][29] ), .ZN(n9827) );
  OAI22_X2 U10962 ( .A1(n9827), .A2(n6104), .B1(n6222), .B2(n6102), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10963 ( .A1(n9828), .A2(n6109), .B1(n6222), .B2(n6105), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10964 ( .A1(n5213), .A2(n6113), .B1(n6222), .B2(n6157), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10965 ( .A1(n5126), .A2(n6116), .B1(n6222), .B2(n6159), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10966 ( .A1(n5459), .A2(n6119), .B1(n6222), .B2(n6161), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10967 ( .A1(n4977), .A2(net76864), .B1(n6222), .B2(net76614), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10968 ( .A1(n4988), .A2(n6122), .B1(n6222), .B2(n6163), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10969 ( .A1(n5460), .A2(n6125), .B1(n6222), .B2(n6165), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10970 ( .A1(net71824), .A2(n6128), .B1(n6222), .B2(n6167), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10971 ( .A1(n5123), .A2(n6130), .B1(n6222), .B2(n6169), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10972 ( .A1(n4974), .A2(n6133), .B1(n6222), .B2(n6171), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10973 ( .A1(n5214), .A2(n6137), .B1(n6222), .B2(n6173), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10974 ( .A1(n6178), .A2(\REGFILE/reg_out[29][29] ), .ZN(n9829) );
  OAI22_X2 U10975 ( .A1(n5461), .A2(n6140), .B1(n6222), .B2(net76548), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10976 ( .A1(n6180), .A2(\REGFILE/reg_out[30][29] ), .ZN(n9830) );
  OAI22_X2 U10977 ( .A1(n5125), .A2(n6145), .B1(n6222), .B2(n6182), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10978 ( .A1(n5462), .A2(net76708), .B1(n6222), .B2(n6146), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10979 ( .A1(n5523), .A2(net76694), .B1(n6222), .B2(n6184), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10980 ( .A1(n5463), .A2(n6151), .B1(n6222), .B2(n6186), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U10981 ( .A1(n5987), .A2(n6154), .B1(n6222), .B2(n6188), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U10982 ( .A1(multOut[11]), .A2(net92392), .ZN(n9861) );
  XNOR2_X2 U10983 ( .A(n9833), .B(n9832), .ZN(n9834) );
  NAND2_X2 U10984 ( .A1(net71271), .A2(n9834), .ZN(n9860) );
  NAND2_X2 U10985 ( .A1(n8759), .A2(n9838), .ZN(n9843) );
  NAND2_X2 U10986 ( .A1(net105360), .A2(n9839), .ZN(n9842) );
  NAND2_X2 U10987 ( .A1(n6083), .A2(n10238), .ZN(n9841) );
  NAND2_X2 U10988 ( .A1(n6082), .A2(n10239), .ZN(n9840) );
  NAND4_X2 U10989 ( .A1(n9843), .A2(n9842), .A3(n9841), .A4(n9840), .ZN(n10122) );
  NAND2_X2 U10990 ( .A1(n10066), .A2(n10122), .ZN(n9851) );
  NAND2_X2 U10991 ( .A1(n8759), .A2(n10231), .ZN(n9849) );
  NAND2_X2 U10992 ( .A1(n6083), .A2(n9844), .ZN(n9848) );
  NAND2_X2 U10993 ( .A1(net105360), .A2(n10230), .ZN(n9847) );
  NAND2_X2 U10994 ( .A1(n6082), .A2(n9845), .ZN(n9846) );
  NAND4_X2 U10995 ( .A1(n9849), .A2(n9848), .A3(n9847), .A4(n9846), .ZN(n10123) );
  NAND2_X2 U10996 ( .A1(n10058), .A2(n10123), .ZN(n9850) );
  NAND2_X2 U10997 ( .A1(n9851), .A2(n9850), .ZN(n9857) );
  INV_X4 U10998 ( .A(n9852), .ZN(n9855) );
  NAND4_X2 U10999 ( .A1(n9861), .A2(n9860), .A3(n9859), .A4(n9858), .ZN(
        dmem_addr_out[11]) );
  NAND2_X2 U11000 ( .A1(net76650), .A2(dmem_addr_out[11]), .ZN(n9866) );
  NAND3_X2 U11001 ( .A1(n9866), .A2(net70740), .A3(n9865), .ZN(n9867) );
  NAND2_X2 U11002 ( .A1(n6066), .A2(n4992), .ZN(n9870) );
  NAND2_X2 U11003 ( .A1(n4867), .A2(\REGFILE/reg_out[0][11] ), .ZN(n9869) );
  NAND2_X2 U11004 ( .A1(n9870), .A2(n9869), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11005 ( .A1(n6066), .A2(n4990), .ZN(n9872) );
  NAND2_X2 U11006 ( .A1(n6093), .A2(n5907), .ZN(n9871) );
  NAND2_X2 U11007 ( .A1(n9872), .A2(n9871), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11008 ( .A1(n6066), .A2(n4998), .ZN(n9874) );
  NAND2_X2 U11009 ( .A1(\REGFILE/reg_out[11][11] ), .A2(n4869), .ZN(n9873) );
  NAND2_X2 U11010 ( .A1(n9874), .A2(n9873), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11011 ( .A1(n6066), .A2(n4993), .ZN(n9876) );
  NAND2_X2 U11012 ( .A1(n9876), .A2(n9875), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11013 ( .A1(n6066), .A2(n6096), .ZN(n9878) );
  NAND2_X2 U11014 ( .A1(n9878), .A2(n9877), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11015 ( .A1(n6066), .A2(n6101), .ZN(n9880) );
  NAND2_X2 U11016 ( .A1(n4805), .A2(\REGFILE/reg_out[14][11] ), .ZN(n9879) );
  NAND2_X2 U11017 ( .A1(n9880), .A2(n9879), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11018 ( .A1(n6066), .A2(n6107), .ZN(n9882) );
  NAND2_X2 U11019 ( .A1(n4804), .A2(\REGFILE/reg_out[15][11] ), .ZN(n9881) );
  NAND2_X2 U11020 ( .A1(n9882), .A2(n9881), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11021 ( .A1(n6066), .A2(n4994), .ZN(n9884) );
  NAND2_X2 U11022 ( .A1(n4891), .A2(\REGFILE/reg_out[16][11] ), .ZN(n9883) );
  NAND2_X2 U11023 ( .A1(n9884), .A2(n9883), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11024 ( .A1(n6066), .A2(n4999), .ZN(n9886) );
  NAND2_X2 U11025 ( .A1(n4892), .A2(\REGFILE/reg_out[17][11] ), .ZN(n9885) );
  NAND2_X2 U11026 ( .A1(n9886), .A2(n9885), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11027 ( .A1(n6066), .A2(n5000), .ZN(n9888) );
  NAND2_X2 U11028 ( .A1(n4884), .A2(\REGFILE/reg_out[18][11] ), .ZN(n9887) );
  NAND2_X2 U11029 ( .A1(n9888), .A2(n9887), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11030 ( .A1(n6065), .A2(n5001), .ZN(n9890) );
  NAND2_X2 U11031 ( .A1(\REGFILE/reg_out[19][11] ), .A2(n4876), .ZN(n9889) );
  NAND2_X2 U11032 ( .A1(n9890), .A2(n9889), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11033 ( .A1(n6065), .A2(n4997), .ZN(n9892) );
  NAND2_X2 U11034 ( .A1(n4877), .A2(\REGFILE/reg_out[1][11] ), .ZN(n9891) );
  NAND2_X2 U11035 ( .A1(n9892), .A2(n9891), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11036 ( .A1(n6065), .A2(n4903), .ZN(n9894) );
  NAND2_X2 U11037 ( .A1(\REGFILE/reg_out[20][11] ), .A2(n4868), .ZN(n9893) );
  NAND2_X2 U11038 ( .A1(n9894), .A2(n9893), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11039 ( .A1(n6065), .A2(n4904), .ZN(n9896) );
  NAND2_X2 U11040 ( .A1(n4882), .A2(\REGFILE/reg_out[21][11] ), .ZN(n9895) );
  NAND2_X2 U11041 ( .A1(n9896), .A2(n9895), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11042 ( .A1(n6065), .A2(n4905), .ZN(n9898) );
  NAND2_X2 U11043 ( .A1(n4888), .A2(\REGFILE/reg_out[22][11] ), .ZN(n9897) );
  NAND2_X2 U11044 ( .A1(n9898), .A2(n9897), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11045 ( .A1(n6065), .A2(n4906), .ZN(n9900) );
  NAND2_X2 U11046 ( .A1(n4883), .A2(\REGFILE/reg_out[23][11] ), .ZN(n9899) );
  NAND2_X2 U11047 ( .A1(n9900), .A2(n9899), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11048 ( .A1(n6065), .A2(n4995), .ZN(n9902) );
  NAND2_X2 U11049 ( .A1(n4875), .A2(\REGFILE/reg_out[24][11] ), .ZN(n9901) );
  NAND2_X2 U11050 ( .A1(n9902), .A2(n9901), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11051 ( .A1(n6065), .A2(n5002), .ZN(n9904) );
  NAND2_X2 U11052 ( .A1(n4878), .A2(\REGFILE/reg_out[25][11] ), .ZN(n9903) );
  NAND2_X2 U11053 ( .A1(n9904), .A2(n9903), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11054 ( .A1(n6065), .A2(n5003), .ZN(n9906) );
  NAND2_X2 U11055 ( .A1(n4893), .A2(\REGFILE/reg_out[26][11] ), .ZN(n9905) );
  NAND2_X2 U11056 ( .A1(n9906), .A2(n9905), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11057 ( .A1(n6065), .A2(n5004), .ZN(n9908) );
  NAND2_X2 U11058 ( .A1(n9908), .A2(n9907), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11059 ( .A1(n6065), .A2(n4806), .ZN(n9910) );
  NAND2_X2 U11060 ( .A1(n9910), .A2(n9909), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11061 ( .A1(n6065), .A2(n10607), .ZN(n9912) );
  NAND2_X2 U11062 ( .A1(n6178), .A2(\REGFILE/reg_out[29][11] ), .ZN(n9911) );
  NAND2_X2 U11063 ( .A1(n9912), .A2(n9911), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11064 ( .A1(n6065), .A2(n5005), .ZN(n9914) );
  NAND2_X2 U11065 ( .A1(n4879), .A2(\REGFILE/reg_out[2][11] ), .ZN(n9913) );
  NAND2_X2 U11066 ( .A1(n9914), .A2(n9913), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11067 ( .A1(n6066), .A2(n10614), .ZN(n9916) );
  NAND2_X2 U11068 ( .A1(n6180), .A2(\REGFILE/reg_out[30][11] ), .ZN(n9915) );
  NAND2_X2 U11069 ( .A1(n9916), .A2(n9915), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11070 ( .A1(n6065), .A2(net70574), .ZN(n9918) );
  NAND2_X2 U11071 ( .A1(n5688), .A2(\REGFILE/reg_out[31][11] ), .ZN(n9917) );
  NAND2_X2 U11072 ( .A1(n9918), .A2(n9917), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11073 ( .A1(n6066), .A2(n5009), .ZN(n9920) );
  NAND2_X2 U11074 ( .A1(\REGFILE/reg_out[3][11] ), .A2(n4871), .ZN(n9919) );
  NAND2_X2 U11075 ( .A1(n9920), .A2(n9919), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11076 ( .A1(n6066), .A2(n4996), .ZN(n9922) );
  NAND2_X2 U11077 ( .A1(\REGFILE/reg_out[4][11] ), .A2(n4870), .ZN(n9921) );
  NAND2_X2 U11078 ( .A1(n9922), .A2(n9921), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11079 ( .A1(n6066), .A2(n5006), .ZN(n9924) );
  NAND2_X2 U11080 ( .A1(n4885), .A2(\REGFILE/reg_out[5][11] ), .ZN(n9923) );
  NAND2_X2 U11081 ( .A1(n9924), .A2(n9923), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11082 ( .A1(n6066), .A2(n6148), .ZN(n9926) );
  NAND2_X2 U11083 ( .A1(n4889), .A2(\REGFILE/reg_out[6][11] ), .ZN(n9925) );
  NAND2_X2 U11084 ( .A1(n9926), .A2(n9925), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11085 ( .A1(n6065), .A2(n5007), .ZN(n9928) );
  NAND2_X2 U11086 ( .A1(n4886), .A2(\REGFILE/reg_out[7][11] ), .ZN(n9927) );
  NAND2_X2 U11087 ( .A1(n9928), .A2(n9927), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11088 ( .A1(n6065), .A2(n4991), .ZN(n9930) );
  NAND2_X2 U11089 ( .A1(n4890), .A2(\REGFILE/reg_out[8][11] ), .ZN(n9929) );
  NAND2_X2 U11090 ( .A1(n9930), .A2(n9929), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11091 ( .A1(n6066), .A2(n5008), .ZN(n9932) );
  NAND2_X2 U11092 ( .A1(n4887), .A2(\REGFILE/reg_out[9][11] ), .ZN(n9931) );
  NAND2_X2 U11093 ( .A1(n9932), .A2(n9931), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ) );
  AOI22_X2 U11094 ( .A1(net71092), .A2(n9934), .B1(net71094), .B2(n9933), .ZN(
        n9952) );
  INV_X4 U11095 ( .A(n10091), .ZN(n9937) );
  INV_X4 U11096 ( .A(n9935), .ZN(n9936) );
  NAND2_X2 U11097 ( .A1(net70696), .A2(n6005), .ZN(n10014) );
  OAI221_X2 U11098 ( .B1(n9937), .B2(n10094), .C1(n9936), .C2(net70718), .A(
        n10014), .ZN(n10017) );
  NAND2_X2 U11099 ( .A1(n10280), .A2(n10017), .ZN(n9951) );
  NAND2_X2 U11100 ( .A1(n10102), .A2(n10101), .ZN(n9949) );
  NAND2_X2 U11101 ( .A1(net70720), .A2(aluA[20]), .ZN(n9944) );
  INV_X4 U11102 ( .A(n9938), .ZN(n9941) );
  INV_X4 U11103 ( .A(n9939), .ZN(n9940) );
  NAND2_X2 U11104 ( .A1(net105360), .A2(n10541), .ZN(n9948) );
  NAND2_X2 U11105 ( .A1(n4880), .A2(n9945), .ZN(n9947) );
  NAND2_X2 U11106 ( .A1(n6082), .A2(n10103), .ZN(n9946) );
  NAND4_X2 U11107 ( .A1(n9949), .A2(n9948), .A3(n9947), .A4(n9946), .ZN(n10016) );
  INV_X4 U11108 ( .A(n10306), .ZN(n10402) );
  NAND3_X2 U11109 ( .A1(n9952), .A2(n9951), .A3(n9950), .ZN(n9953) );
  MUX2_X2 U11110 ( .A(n9953), .B(multOut[4]), .S(net76452), .Z(n9963) );
  XNOR2_X2 U11111 ( .A(n10033), .B(n9954), .ZN(n10034) );
  INV_X4 U11112 ( .A(n9955), .ZN(n9958) );
  XNOR2_X2 U11113 ( .A(n10034), .B(n10035), .ZN(n9961) );
  NAND2_X2 U11114 ( .A1(net71078), .A2(\WIRE_ALU_A/MUX2TO1_32BIT[4].MUX/N1 ), 
        .ZN(n9960) );
  OAI22_X2 U11115 ( .A1(n5524), .A2(n6089), .B1(net76658), .B2(n4803), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11116 ( .A1(n5464), .A2(n6092), .B1(n6155), .B2(n6068), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11117 ( .A1(n6193), .A2(n5557), .B1(n6194), .B2(n4803), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11118 ( .A1(n6197), .A2(n5033), .B1(n6198), .B2(n6067), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11119 ( .A1(n5465), .A2(n6098), .B1(n6094), .B2(n6067), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11120 ( .A1(n5525), .A2(n6104), .B1(n10519), .B2(n6067), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11121 ( .A1(n5329), .A2(n6109), .B1(n6105), .B2(n6067), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11122 ( .A1(n5215), .A2(n6113), .B1(n6157), .B2(n6067), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11123 ( .A1(n5526), .A2(n6116), .B1(n6159), .B2(n6067), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11124 ( .A1(n5466), .A2(n6119), .B1(n6161), .B2(n4803), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11125 ( .A1(n6201), .A2(n5438), .B1(n6203), .B2(n6068), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11126 ( .A1(n5048), .A2(net76864), .B1(net76614), .B2(n4803), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11127 ( .A1(n6206), .A2(n5423), .B1(n6207), .B2(n4803), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11128 ( .A1(n5216), .A2(n6122), .B1(n6163), .B2(n6067), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11129 ( .A1(n5467), .A2(n6125), .B1(n6165), .B2(n6068), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11130 ( .A1(n5527), .A2(n6128), .B1(n6167), .B2(n6068), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11131 ( .A1(n5528), .A2(n6130), .B1(n6169), .B2(n6068), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11132 ( .A1(n5468), .A2(n6133), .B1(n6171), .B2(n4803), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11133 ( .A1(n5217), .A2(n6137), .B1(n6067), .B2(n6173), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11134 ( .A1(n6210), .A2(n5424), .B1(n6211), .B2(n6068), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11135 ( .A1(\REGFILE/reg_out[28][4] ), .A2(n10604), .ZN(n9969) );
  NAND2_X2 U11136 ( .A1(n10608), .A2(\REGFILE/reg_out[29][4] ), .ZN(n9970) );
  OAI22_X2 U11137 ( .A1(n5770), .A2(n6140), .B1(net76548), .B2(n6068), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11138 ( .A1(n10615), .A2(\REGFILE/reg_out[30][4] ), .ZN(n9971) );
  NAND2_X2 U11139 ( .A1(net76488), .A2(\REGFILE/reg_out[31][4] ), .ZN(n9972)
         );
  OAI22_X2 U11141 ( .A1(n6216), .A2(n9973), .B1(net76318), .B2(n4803), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11142 ( .A1(n6218), .A2(n5386), .B1(n6219), .B2(n6067), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11143 ( .A1(n5330), .A2(n6145), .B1(n6182), .B2(n4803), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11144 ( .A1(n5469), .A2(net76708), .B1(n6146), .B2(n6068), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11145 ( .A1(n5529), .A2(net76694), .B1(n6184), .B2(n4803), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11146 ( .A1(n5331), .A2(n6151), .B1(n6186), .B2(n6068), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11147 ( .A1(n5218), .A2(n6154), .B1(n6188), .B2(n6067), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11148 ( .A1(n8759), .A2(n9975), .ZN(n9981) );
  NAND2_X2 U11149 ( .A1(net77086), .A2(n9976), .ZN(n9980) );
  AOI22_X2 U11150 ( .A1(n6082), .A2(n9978), .B1(n6083), .B2(n9977), .ZN(n9979)
         );
  NAND2_X2 U11151 ( .A1(net71092), .A2(n10057), .ZN(n9990) );
  MUX2_X2 U11152 ( .A(n9982), .B(n10065), .S(net71026), .Z(n9983) );
  NAND2_X2 U11153 ( .A1(net71094), .A2(n9983), .ZN(n9989) );
  NAND2_X2 U11154 ( .A1(n10280), .A2(n9984), .ZN(n9988) );
  AOI21_X4 U11155 ( .B1(net71085), .B2(n9986), .A(n9985), .ZN(n9987) );
  NAND4_X2 U11156 ( .A1(n9990), .A2(n9989), .A3(n9988), .A4(n9987), .ZN(n9991)
         );
  MUX2_X2 U11157 ( .A(n9991), .B(multOut[19]), .S(net76452), .Z(n9998) );
  XNOR2_X2 U11158 ( .A(n9993), .B(n9992), .ZN(n9996) );
  NAND2_X2 U11159 ( .A1(net71078), .A2(aluA[19]), .ZN(n9994) );
  OAI22_X2 U11160 ( .A1(n9996), .A2(net70691), .B1(n9995), .B2(n9994), .ZN(
        n9997) );
  NOR2_X4 U11161 ( .A1(n9998), .A2(n9997), .ZN(n10006) );
  INV_X4 U11162 ( .A(n10006), .ZN(dmem_addr_out[19]) );
  INV_X4 U11163 ( .A(dmem_read_in[19]), .ZN(n10001) );
  OAI211_X2 U11164 ( .C1(n10006), .C2(net76646), .A(n10005), .B(n10004), .ZN(
        n10007) );
  NAND2_X2 U11165 ( .A1(net76270), .A2(n10007), .ZN(n10012) );
  OAI22_X2 U11166 ( .A1(n5219), .A2(n6089), .B1(net76658), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11167 ( .A1(n5031), .A2(n6092), .B1(n6155), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11168 ( .A1(n6193), .A2(n5387), .B1(n6194), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11169 ( .A1(n6197), .A2(n5035), .B1(n6198), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11170 ( .A1(n5332), .A2(n6098), .B1(n6094), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11171 ( .A1(n5220), .A2(n6104), .B1(n6102), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11172 ( .A1(n4978), .A2(n6109), .B1(n6105), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11173 ( .A1(n5221), .A2(n6113), .B1(n6157), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11174 ( .A1(n5222), .A2(n6116), .B1(n6159), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11175 ( .A1(n5333), .A2(n6119), .B1(n6161), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11176 ( .A1(n6201), .A2(n5118), .B1(n6203), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11177 ( .A1(n5080), .A2(net76864), .B1(net76614), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11178 ( .A1(n6206), .A2(n5425), .B1(n6207), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11179 ( .A1(n5223), .A2(n6122), .B1(n6163), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11180 ( .A1(n5334), .A2(n6125), .B1(n6165), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11181 ( .A1(n5224), .A2(n6128), .B1(n6167), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11182 ( .A1(n5104), .A2(n6130), .B1(n6169), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11183 ( .A1(n4973), .A2(n6133), .B1(n6171), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11184 ( .A1(n5225), .A2(n6137), .B1(n6173), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11185 ( .A1(n6210), .A2(n5036), .B1(n6211), .B2(n10012), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11186 ( .A1(\REGFILE/reg_out[28][19] ), .A2(n10604), .ZN(n10008)
         );
  NAND2_X2 U11187 ( .A1(n10608), .A2(\REGFILE/reg_out[29][19] ), .ZN(n10009)
         );
  OAI22_X2 U11188 ( .A1(n5651), .A2(n6140), .B1(net76548), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11189 ( .A1(n10615), .A2(\REGFILE/reg_out[30][19] ), .ZN(n10010)
         );
  NAND2_X2 U11190 ( .A1(net76488), .A2(\REGFILE/reg_out[31][19] ), .ZN(n10011)
         );
  OAI22_X2 U11191 ( .A1(n6216), .A2(n5426), .B1(net76318), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11192 ( .A1(n6218), .A2(n5388), .B1(n6219), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11193 ( .A1(n5335), .A2(n6145), .B1(n6182), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11194 ( .A1(n5336), .A2(net76708), .B1(n6146), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11195 ( .A1(n5226), .A2(net76694), .B1(n6184), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11196 ( .A1(n5337), .A2(n6151), .B1(n6186), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11197 ( .A1(n5227), .A2(n6154), .B1(n6188), .B2(n6070), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[19].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11198 ( .A(net70727), .ZN(net71299) );
  INV_X4 U11199 ( .A(n10013), .ZN(n10015) );
  OAI221_X2 U11200 ( .B1(net71299), .B2(n10094), .C1(n10015), .C2(net70718), 
        .A(n10014), .ZN(n10092) );
  AOI222_X2 U11201 ( .A1(n10280), .A2(n10092), .B1(net71092), .B2(n10017), 
        .C1(net71094), .C2(n10016), .ZN(n10031) );
  NAND2_X2 U11202 ( .A1(net70720), .A2(aluA[19]), .ZN(n10021) );
  NAND2_X2 U11203 ( .A1(net70719), .A2(n5761), .ZN(n10020) );
  NAND4_X2 U11204 ( .A1(n10021), .A2(n10020), .A3(n10019), .A4(n10018), .ZN(
        n10022) );
  MUX2_X2 U11205 ( .A(n10023), .B(n10022), .S(n10099), .Z(n10156) );
  INV_X4 U11206 ( .A(n10156), .ZN(n10027) );
  NAND2_X2 U11207 ( .A1(n8759), .A2(n10158), .ZN(n10026) );
  NAND2_X2 U11208 ( .A1(n6083), .A2(n10024), .ZN(n10025) );
  OAI211_X2 U11209 ( .C1(net78051), .C2(n10027), .A(n10026), .B(n10025), .ZN(
        n10028) );
  INV_X4 U11210 ( .A(n10028), .ZN(n10093) );
  INV_X4 U11211 ( .A(n10407), .ZN(n10415) );
  NOR2_X4 U11212 ( .A1(n10029), .A2(n5040), .ZN(n10030) );
  NAND2_X2 U11213 ( .A1(n10031), .A2(n10030), .ZN(n10032) );
  AOI22_X2 U11214 ( .A1(n10035), .A2(n10034), .B1(
        \WIRE_ALU_A/MUX2TO1_32BIT[4].MUX/N1 ), .B2(n10033), .ZN(n10111) );
  XNOR2_X2 U11215 ( .A(n10111), .B(n4813), .ZN(n10038) );
  NAND2_X2 U11216 ( .A1(net71078), .A2(\WIRE_ALU_A/MUX2TO1_32BIT[3].MUX/N1 ), 
        .ZN(n10037) );
  OAI22_X2 U11217 ( .A1(n5530), .A2(n6089), .B1(net76658), .B2(n6072), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11218 ( .A1(n5470), .A2(n6092), .B1(n6073), .B2(n6155), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11219 ( .A1(n6193), .A2(n5389), .B1(n6194), .B2(n6073), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11220 ( .A1(n6197), .A2(n5427), .B1(n6073), .B2(n6198), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11221 ( .A1(n5471), .A2(n6098), .B1(n6095), .B2(n6072), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11222 ( .A1(n5531), .A2(n6104), .B1(n6073), .B2(n6102), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11223 ( .A1(n5338), .A2(n6109), .B1(n6073), .B2(n6106), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11224 ( .A1(n5228), .A2(n6113), .B1(n6073), .B2(n6157), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11225 ( .A1(n5532), .A2(n6116), .B1(n6073), .B2(n6159), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11226 ( .A1(n5472), .A2(n6119), .B1(n6073), .B2(n6161), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11227 ( .A1(n6201), .A2(n5558), .B1(n6073), .B2(n6203), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11228 ( .A1(n5473), .A2(net76864), .B1(n6073), .B2(net76614), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11229 ( .A1(n6206), .A2(n5428), .B1(n6073), .B2(n6207), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11230 ( .A1(n5229), .A2(n6122), .B1(n6073), .B2(n6163), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11231 ( .A1(n5339), .A2(n6125), .B1(n6073), .B2(n6165), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11232 ( .A1(n5230), .A2(n6128), .B1(n6073), .B2(n6167), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11233 ( .A1(n5533), .A2(n6130), .B1(n6169), .B2(n6072), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11234 ( .A(n5957), .ZN(n10047) );
  OAI22_X2 U11235 ( .A1(n10047), .A2(n6133), .B1(n6171), .B2(n6072), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11236 ( .A1(n5231), .A2(n6137), .B1(n6173), .B2(n6072), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11237 ( .A1(n6210), .A2(n5429), .B1(n6211), .B2(n6072), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11238 ( .A1(\REGFILE/reg_out[28][3] ), .A2(n6175), .ZN(n10048) );
  OAI22_X2 U11239 ( .A1(n5045), .A2(n6140), .B1(net76548), .B2(n6072), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11240 ( .A1(n10615), .A2(\REGFILE/reg_out[30][3] ), .ZN(n10050) );
  NAND2_X2 U11241 ( .A1(net76488), .A2(\REGFILE/reg_out[31][3] ), .ZN(n10051)
         );
  OAI22_X2 U11242 ( .A1(n6216), .A2(n5046), .B1(net76318), .B2(n6072), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11243 ( .A1(n6218), .A2(n5559), .B1(n6219), .B2(n6072), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11244 ( .A1(n5474), .A2(n6145), .B1(n6182), .B2(n6072), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11245 ( .A1(n5475), .A2(net76708), .B1(n6147), .B2(n6072), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11246 ( .A1(n5534), .A2(net76694), .B1(n6184), .B2(n6072), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11247 ( .A1(n5476), .A2(n6151), .B1(n6186), .B2(n6072), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11248 ( .A1(n5535), .A2(n6154), .B1(n6073), .B2(n6188), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  XNOR2_X2 U11249 ( .A(n10054), .B(n10053), .ZN(n10056) );
  NAND2_X2 U11250 ( .A1(multOut[20]), .A2(net92392), .ZN(n10076) );
  NAND2_X2 U11251 ( .A1(n10058), .A2(n10057), .ZN(n10062) );
  NAND2_X2 U11252 ( .A1(n10060), .A2(n10059), .ZN(n10061) );
  NAND2_X2 U11253 ( .A1(n10062), .A2(n10061), .ZN(n10074) );
  NAND2_X2 U11254 ( .A1(n10064), .A2(n10063), .ZN(n10068) );
  NAND2_X2 U11255 ( .A1(n10066), .A2(n10065), .ZN(n10067) );
  NAND2_X2 U11256 ( .A1(n10068), .A2(n10067), .ZN(n10069) );
  MUX2_X2 U11257 ( .A(n10070), .B(n10069), .S(net71026), .Z(n10073) );
  INV_X4 U11258 ( .A(aluA[20]), .ZN(n10071) );
  NAND3_X2 U11259 ( .A1(n10077), .A2(n10076), .A3(n10075), .ZN(
        dmem_addr_out[20]) );
  INV_X4 U11260 ( .A(dmem_read_in[20]), .ZN(n10078) );
  NAND2_X2 U11261 ( .A1(n5573), .A2(n10079), .ZN(n10085) );
  INV_X4 U11262 ( .A(dmem_addr_out[20]), .ZN(n10082) );
  NAND2_X2 U11263 ( .A1(n10080), .A2(net77030), .ZN(n10081) );
  OAI221_X2 U11264 ( .B1(net77999), .B2(n10083), .C1(n10082), .C2(net76646), 
        .A(n10081), .ZN(n10084) );
  OAI21_X4 U11265 ( .B1(n10085), .B2(n10084), .A(reset), .ZN(n10090) );
  OAI22_X2 U11266 ( .A1(n5232), .A2(n6089), .B1(net76658), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11267 ( .A1(n5821), .A2(n6092), .B1(n6155), .B2(n6075), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11268 ( .A1(n6193), .A2(n5390), .B1(n6194), .B2(n6075), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11269 ( .A1(n6197), .A2(n5682), .B1(n6198), .B2(n6075), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11270 ( .A1(n5340), .A2(n6098), .B1(n6094), .B2(n6075), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11271 ( .A1(n5233), .A2(n6104), .B1(n6102), .B2(n6075), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11272 ( .A1(n5081), .A2(n6109), .B1(n6105), .B2(n6075), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11273 ( .A1(n5105), .A2(n6113), .B1(n6157), .B2(n6075), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11274 ( .A1(n5234), .A2(n6116), .B1(n6159), .B2(n6075), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11275 ( .A1(n5341), .A2(n6119), .B1(n6161), .B2(n6075), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11276 ( .A1(n6201), .A2(n5391), .B1(n6203), .B2(n6075), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11277 ( .A1(n5342), .A2(net76864), .B1(net76614), .B2(n6075), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11278 ( .A1(n6206), .A2(n5506), .B1(n6207), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11279 ( .A1(n5235), .A2(n6122), .B1(n6163), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11280 ( .A1(n5343), .A2(n6125), .B1(n6165), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11281 ( .A1(n5236), .A2(n6128), .B1(n6167), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11282 ( .A1(n5237), .A2(n6130), .B1(n6169), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11283 ( .A1(n5661), .A2(n6133), .B1(n6171), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11284 ( .A1(n5238), .A2(n6137), .B1(n6173), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11285 ( .A1(n6210), .A2(n5681), .B1(n6211), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11286 ( .A1(\REGFILE/reg_out[28][20] ), .A2(n10604), .ZN(n10086)
         );
  OAI21_X4 U11287 ( .B1(n6214), .B2(n6075), .A(n10086), .ZN(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11288 ( .A1(n10608), .A2(\REGFILE/reg_out[29][20] ), .ZN(n10087)
         );
  OAI21_X4 U11289 ( .B1(n10532), .B2(n6075), .A(n10087), .ZN(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11290 ( .A1(n5023), .A2(n6140), .B1(net76548), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11291 ( .A1(n10615), .A2(\REGFILE/reg_out[30][20] ), .ZN(n10088)
         );
  OAI21_X4 U11292 ( .B1(n10534), .B2(n6075), .A(n10088), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11293 ( .A1(net76488), .A2(\REGFILE/reg_out[31][20] ), .ZN(n10089)
         );
  OAI21_X4 U11294 ( .B1(net70509), .B2(n6075), .A(n10089), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11295 ( .A1(n6216), .A2(n5037), .B1(net76318), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11296 ( .A1(n6218), .A2(n5500), .B1(n6219), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11297 ( .A1(n5344), .A2(n6145), .B1(n6182), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11298 ( .A1(n5345), .A2(net76708), .B1(n6146), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11299 ( .A1(n5239), .A2(net76694), .B1(n6184), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11300 ( .A1(n5346), .A2(n6151), .B1(n6186), .B2(n6076), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11301 ( .A1(n5240), .A2(n6154), .B1(n6188), .B2(n6075), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[20].REGISTER1/STORE_DATA/N3 ) );
  MUX2_X2 U11302 ( .A(net70696), .B(n10091), .S(net77084), .Z(n10150) );
  AOI22_X2 U11303 ( .A1(n10280), .A2(n10150), .B1(net71092), .B2(n10092), .ZN(
        n10107) );
  INV_X4 U11304 ( .A(n10094), .ZN(n10102) );
  NAND2_X2 U11305 ( .A1(net70720), .A2(aluA[18]), .ZN(n10098) );
  NAND4_X2 U11306 ( .A1(n10098), .A2(n10097), .A3(n10096), .A4(n10095), .ZN(
        n10100) );
  MUX2_X2 U11307 ( .A(n10101), .B(n10100), .S(n10099), .Z(net70713) );
  INV_X4 U11308 ( .A(n10104), .ZN(n10414) );
  NOR2_X4 U11309 ( .A1(n10105), .A2(n5041), .ZN(n10106) );
  XNOR2_X2 U11310 ( .A(n10165), .B(n10109), .ZN(n10166) );
  INV_X4 U11311 ( .A(n10110), .ZN(n10112) );
  OAI22_X2 U11312 ( .A1(n10112), .A2(n10404), .B1(n10111), .B2(n4813), .ZN(
        n10167) );
  XNOR2_X2 U11313 ( .A(n10166), .B(n10167), .ZN(n10114) );
  NAND2_X2 U11314 ( .A1(net71078), .A2(\WIRE_ALU_A/MUX2TO1_32BIT[2].MUX/N1 ), 
        .ZN(n10113) );
  OAI22_X2 U11315 ( .A1(n5536), .A2(n6089), .B1(net76658), .B2(net77116), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11316 ( .A1(n5477), .A2(n6092), .B1(n6155), .B2(net77114), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11317 ( .A1(n6193), .A2(n5560), .B1(n6194), .B2(net77116), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11318 ( .A1(n6197), .A2(n4989), .B1(net77116), .B2(n6198), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11319 ( .A1(n5478), .A2(n6098), .B1(n6094), .B2(net77116), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11320 ( .A1(n5537), .A2(n6104), .B1(n10519), .B2(net77114), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11321 ( .A1(n5347), .A2(n6109), .B1(n6105), .B2(net77114), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11322 ( .A1(n5241), .A2(n6113), .B1(n6157), .B2(net77116), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11323 ( .A1(n5538), .A2(n6116), .B1(n6159), .B2(net77114), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11324 ( .A1(n5479), .A2(n6119), .B1(n6161), .B2(net77114), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11325 ( .A1(n6201), .A2(n5392), .B1(n6203), .B2(net77116), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11327 ( .A1(n10116), .A2(net76864), .B1(net76614), .B2(net77114), 
        .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11328 ( .A1(n6206), .A2(n4986), .B1(net77116), .B2(n6207), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11329 ( .A1(n5242), .A2(n6122), .B1(n6163), .B2(net77114), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11330 ( .A1(n5348), .A2(n6125), .B1(n6165), .B2(net77114), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11331 ( .A1(n5243), .A2(n6128), .B1(n6167), .B2(net77116), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11332 ( .A1(n5539), .A2(n6130), .B1(n6169), .B2(net77114), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11334 ( .A1(n10117), .A2(n6133), .B1(n6171), .B2(net77116), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11335 ( .A1(n5244), .A2(n6137), .B1(n6173), .B2(net77114), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11336 ( .A1(n6210), .A2(n4987), .B1(n6211), .B2(net77116), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11337 ( .A1(\REGFILE/reg_out[28][2] ), .A2(n6175), .ZN(n10118) );
  NAND2_X2 U11338 ( .A1(n10608), .A2(\REGFILE/reg_out[29][2] ), .ZN(n10119) );
  OAI22_X2 U11339 ( .A1(n5480), .A2(n6140), .B1(net76548), .B2(net77116), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11340 ( .A1(n6180), .A2(\REGFILE/reg_out[30][2] ), .ZN(n10120) );
  OAI22_X2 U11342 ( .A1(n6216), .A2(n10121), .B1(net76318), .B2(net77114), 
        .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11343 ( .A1(n6218), .A2(n5561), .B1(n6219), .B2(net77116), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11344 ( .A1(n5481), .A2(n6145), .B1(n6182), .B2(net77114), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11345 ( .A1(n5482), .A2(net76708), .B1(n6146), .B2(net77114), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11346 ( .A1(n5540), .A2(net76694), .B1(n6184), .B2(net77116), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11347 ( .A1(n5483), .A2(n6151), .B1(n6186), .B2(net77114), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11348 ( .A1(n5541), .A2(n6154), .B1(n6188), .B2(net77116), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  AOI22_X2 U11349 ( .A1(net71092), .A2(n10123), .B1(net71094), .B2(n10122), 
        .ZN(n10129) );
  NAND2_X2 U11350 ( .A1(n10280), .A2(n10124), .ZN(n10128) );
  INV_X4 U11351 ( .A(n10421), .ZN(n10380) );
  NAND3_X2 U11352 ( .A1(n10129), .A2(n10128), .A3(n10127), .ZN(n10130) );
  XNOR2_X2 U11353 ( .A(n10132), .B(n10131), .ZN(n10134) );
  NAND2_X2 U11354 ( .A1(net71078), .A2(\WIRE_ALU_A/MUX2TO1_32BIT[10].MUX/N1 ), 
        .ZN(n10133) );
  NOR2_X4 U11355 ( .A1(n10136), .A2(n10135), .ZN(n10141) );
  OAI22_X2 U11356 ( .A1(n5106), .A2(n6089), .B1(net76658), .B2(n6078), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11357 ( .A(\REGFILE/reg_out[10][10] ), .ZN(n10143) );
  OAI22_X2 U11358 ( .A1(n10143), .A2(n6092), .B1(n6155), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11359 ( .A1(n6193), .A2(n5119), .B1(n6194), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11360 ( .A1(n6197), .A2(n5775), .B1(n6198), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11361 ( .A1(n5024), .A2(n6098), .B1(n6094), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11362 ( .A1(n5107), .A2(n6104), .B1(n6102), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11363 ( .A1(n10144), .A2(n6109), .B1(n6105), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11364 ( .A1(n5245), .A2(n6113), .B1(n6157), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11365 ( .A1(n5108), .A2(n6116), .B1(n6159), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11366 ( .A1(n5774), .A2(n6119), .B1(n6161), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11367 ( .A1(n6201), .A2(n5393), .B1(n6203), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11368 ( .A1(n4979), .A2(net76864), .B1(net76614), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11369 ( .A1(n6206), .A2(n5430), .B1(n6207), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11370 ( .A1(n5246), .A2(n6122), .B1(n6163), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11371 ( .A1(n5082), .A2(n6125), .B1(n6165), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11372 ( .A1(n5109), .A2(n6128), .B1(n6167), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11373 ( .A1(n5110), .A2(n6130), .B1(n6169), .B2(n6078), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11374 ( .A1(n5025), .A2(n6133), .B1(n6171), .B2(n6078), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11375 ( .A1(n5247), .A2(n6137), .B1(n6173), .B2(n6078), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11376 ( .A1(n6210), .A2(n5877), .B1(n6211), .B2(n6078), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11377 ( .A1(\REGFILE/reg_out[28][10] ), .A2(n6177), .ZN(n10145) );
  NAND2_X2 U11378 ( .A1(n10608), .A2(\REGFILE/reg_out[29][10] ), .ZN(n10146)
         );
  OAI22_X2 U11379 ( .A1(n5773), .A2(n6140), .B1(net76548), .B2(n6078), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11380 ( .A1(n10615), .A2(\REGFILE/reg_out[30][10] ), .ZN(n10147)
         );
  NAND2_X2 U11381 ( .A1(net76488), .A2(\REGFILE/reg_out[31][10] ), .ZN(n10148)
         );
  OAI22_X2 U11382 ( .A1(n6216), .A2(n5114), .B1(net76318), .B2(n6078), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11383 ( .A1(n6218), .A2(n5120), .B1(n6219), .B2(n6078), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11384 ( .A1(n5083), .A2(n6145), .B1(n6182), .B2(n6078), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11385 ( .A1(n5349), .A2(net76708), .B1(n6146), .B2(n6078), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11386 ( .A1(n5248), .A2(net76694), .B1(n6184), .B2(n6078), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11387 ( .A1(n5350), .A2(n6151), .B1(n6186), .B2(n6078), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11388 ( .A1(n5249), .A2(n6154), .B1(n6188), .B2(n6079), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[10].REGISTER1/STORE_DATA/N3 ) );
  AOI22_X2 U11389 ( .A1(n10280), .A2(n10151), .B1(net71092), .B2(n10150), .ZN(
        net71277) );
  NAND2_X2 U11390 ( .A1(n10930), .A2(net70719), .ZN(n10154) );
  NAND2_X2 U11391 ( .A1(net70720), .A2(aluA[17]), .ZN(n10153) );
  NAND3_X4 U11392 ( .A1(n10155), .A2(n10154), .A3(n10153), .ZN(n10163) );
  NAND2_X2 U11393 ( .A1(n10156), .A2(net78051), .ZN(n10157) );
  INV_X4 U11394 ( .A(n10157), .ZN(n10162) );
  INV_X4 U11395 ( .A(n10158), .ZN(n10160) );
  OAI22_X2 U11396 ( .A1(n10160), .A2(n10544), .B1(n10159), .B2(net71273), .ZN(
        n10161) );
  AOI211_X4 U11397 ( .C1(net77084), .C2(n10163), .A(n10162), .B(n10161), .ZN(
        net70709) );
  INV_X4 U11398 ( .A(n10164), .ZN(n10416) );
  AOI22_X2 U11399 ( .A1(n10167), .A2(n10166), .B1(
        \WIRE_ALU_A/MUX2TO1_32BIT[2].MUX/N1 ), .B2(n10165), .ZN(net70731) );
  XNOR2_X2 U11400 ( .A(net70734), .B(net71273), .ZN(net70735) );
  NAND2_X2 U11401 ( .A1(net77104), .A2(n4992), .ZN(n10169) );
  NAND2_X2 U11402 ( .A1(n4867), .A2(\REGFILE/reg_out[0][1] ), .ZN(n10168) );
  NAND2_X2 U11403 ( .A1(n6093), .A2(\REGFILE/reg_out[10][1] ), .ZN(n10170) );
  NAND2_X2 U11404 ( .A1(net77102), .A2(n4998), .ZN(n10173) );
  NAND2_X2 U11405 ( .A1(\REGFILE/reg_out[11][1] ), .A2(n4869), .ZN(n10172) );
  NAND2_X2 U11406 ( .A1(n10173), .A2(n10172), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11407 ( .A1(net77102), .A2(n4993), .ZN(n10175) );
  NAND2_X2 U11408 ( .A1(\REGFILE/reg_out[12][1] ), .A2(n4873), .ZN(n10174) );
  NAND2_X2 U11409 ( .A1(n10175), .A2(n10174), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11410 ( .A1(net77104), .A2(n6096), .ZN(n10177) );
  NAND2_X2 U11411 ( .A1(n10177), .A2(n10176), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11412 ( .A1(net77104), .A2(n6101), .ZN(n10179) );
  NAND2_X2 U11413 ( .A1(n4805), .A2(\REGFILE/reg_out[14][1] ), .ZN(n10178) );
  NAND2_X2 U11414 ( .A1(n10179), .A2(n10178), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11415 ( .A1(net77100), .A2(n6107), .ZN(n10181) );
  NAND2_X2 U11416 ( .A1(n4804), .A2(\REGFILE/reg_out[15][1] ), .ZN(n10180) );
  NAND2_X2 U11417 ( .A1(n10181), .A2(n10180), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11418 ( .A1(net77104), .A2(n4994), .ZN(n10183) );
  NAND2_X2 U11419 ( .A1(n4891), .A2(\REGFILE/reg_out[16][1] ), .ZN(n10182) );
  NAND2_X2 U11420 ( .A1(n10183), .A2(n10182), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11421 ( .A1(net77102), .A2(n4999), .ZN(n10185) );
  NAND2_X2 U11422 ( .A1(n4892), .A2(\REGFILE/reg_out[17][1] ), .ZN(n10184) );
  NAND2_X2 U11423 ( .A1(net77104), .A2(n5000), .ZN(n10187) );
  NAND2_X2 U11424 ( .A1(n4884), .A2(\REGFILE/reg_out[18][1] ), .ZN(n10186) );
  NAND2_X2 U11425 ( .A1(net77100), .A2(n5001), .ZN(n10189) );
  NAND2_X2 U11426 ( .A1(\REGFILE/reg_out[19][1] ), .A2(n4876), .ZN(n10188) );
  NAND2_X2 U11427 ( .A1(n10189), .A2(n10188), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11428 ( .A1(net77100), .A2(n4903), .ZN(n10191) );
  NAND2_X2 U11429 ( .A1(\REGFILE/reg_out[20][1] ), .A2(n4868), .ZN(n10190) );
  NAND2_X2 U11430 ( .A1(net77100), .A2(n4904), .ZN(n10193) );
  NAND2_X2 U11431 ( .A1(n4882), .A2(\REGFILE/reg_out[21][1] ), .ZN(n10192) );
  NAND2_X2 U11432 ( .A1(n10193), .A2(n10192), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11433 ( .A1(n10947), .A2(n4905), .ZN(n10195) );
  NAND2_X2 U11435 ( .A1(n10195), .A2(n10194), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11436 ( .A1(net77102), .A2(n4906), .ZN(n10197) );
  NAND2_X2 U11437 ( .A1(n4883), .A2(\REGFILE/reg_out[23][1] ), .ZN(n10196) );
  NAND2_X2 U11438 ( .A1(net77102), .A2(n4995), .ZN(n10199) );
  NAND2_X2 U11439 ( .A1(n4875), .A2(\REGFILE/reg_out[24][1] ), .ZN(n10198) );
  NAND2_X2 U11440 ( .A1(n10199), .A2(n10198), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11441 ( .A1(net77100), .A2(n5002), .ZN(n10201) );
  NAND2_X2 U11442 ( .A1(n4878), .A2(\REGFILE/reg_out[25][1] ), .ZN(n10200) );
  NAND2_X2 U11443 ( .A1(n10201), .A2(n10200), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11444 ( .A1(net77100), .A2(n5003), .ZN(n10203) );
  NAND2_X2 U11445 ( .A1(n4893), .A2(\REGFILE/reg_out[26][1] ), .ZN(n10202) );
  NAND2_X2 U11446 ( .A1(net77104), .A2(n5004), .ZN(n10205) );
  NAND2_X2 U11447 ( .A1(\REGFILE/reg_out[27][1] ), .A2(n4872), .ZN(n10204) );
  NAND2_X2 U11448 ( .A1(\REGFILE/reg_out[28][1] ), .A2(n6175), .ZN(n10206) );
  NAND2_X2 U11449 ( .A1(n10608), .A2(\REGFILE/reg_out[29][1] ), .ZN(n10208) );
  NAND2_X2 U11450 ( .A1(net77102), .A2(n5005), .ZN(n10211) );
  NAND2_X2 U11451 ( .A1(n4879), .A2(\REGFILE/reg_out[2][1] ), .ZN(n10210) );
  NAND2_X2 U11452 ( .A1(n10211), .A2(n10210), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11453 ( .A1(n10615), .A2(\REGFILE/reg_out[30][1] ), .ZN(n10212) );
  NAND2_X2 U11454 ( .A1(net76488), .A2(\REGFILE/reg_out[31][1] ), .ZN(n10214)
         );
  NAND2_X2 U11455 ( .A1(\REGFILE/reg_out[3][1] ), .A2(n4871), .ZN(n10216) );
  NAND2_X2 U11456 ( .A1(n10217), .A2(n10216), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11457 ( .A1(net77100), .A2(n4996), .ZN(n10219) );
  NAND2_X2 U11458 ( .A1(\REGFILE/reg_out[4][1] ), .A2(n4870), .ZN(n10218) );
  NAND2_X2 U11459 ( .A1(net77102), .A2(n5006), .ZN(n10221) );
  NAND2_X2 U11460 ( .A1(n4885), .A2(\REGFILE/reg_out[5][1] ), .ZN(n10220) );
  NAND2_X2 U11461 ( .A1(net77102), .A2(n6148), .ZN(n10223) );
  NAND2_X2 U11462 ( .A1(n4889), .A2(\REGFILE/reg_out[6][1] ), .ZN(n10222) );
  NAND2_X2 U11463 ( .A1(n10223), .A2(n10222), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11464 ( .A1(net77100), .A2(n5007), .ZN(n10225) );
  NAND2_X2 U11465 ( .A1(n4886), .A2(\REGFILE/reg_out[7][1] ), .ZN(n10224) );
  NAND2_X2 U11466 ( .A1(n10225), .A2(n10224), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11467 ( .A1(net77104), .A2(n4991), .ZN(n10227) );
  NAND2_X2 U11468 ( .A1(n4890), .A2(\REGFILE/reg_out[8][1] ), .ZN(n10226) );
  NAND2_X2 U11469 ( .A1(n10227), .A2(n10226), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11470 ( .A1(net77102), .A2(n5008), .ZN(n10229) );
  NAND2_X2 U11471 ( .A1(n4887), .A2(\REGFILE/reg_out[9][1] ), .ZN(n10228) );
  NAND2_X2 U11472 ( .A1(n10229), .A2(n10228), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[1].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11473 ( .A1(n6082), .A2(n10230), .ZN(n10237) );
  NAND2_X2 U11474 ( .A1(n6083), .A2(n10231), .ZN(n10236) );
  NAND2_X2 U11475 ( .A1(n8759), .A2(n10232), .ZN(n10235) );
  NAND2_X2 U11476 ( .A1(net105360), .A2(n10233), .ZN(n10234) );
  NAND4_X2 U11477 ( .A1(n10237), .A2(n10236), .A3(n10235), .A4(n10234), .ZN(
        n10279) );
  NAND2_X2 U11478 ( .A1(n8728), .A2(n10238), .ZN(n10245) );
  NAND2_X2 U11479 ( .A1(net77084), .A2(n10239), .ZN(n10244) );
  NAND2_X2 U11480 ( .A1(n6082), .A2(n10240), .ZN(n10243) );
  NAND2_X2 U11481 ( .A1(n6083), .A2(n10241), .ZN(n10242) );
  NAND4_X2 U11482 ( .A1(n10245), .A2(n10244), .A3(n10243), .A4(n10242), .ZN(
        n10282) );
  AOI22_X2 U11483 ( .A1(net71092), .A2(n10279), .B1(net71094), .B2(n10282), 
        .ZN(n10251) );
  NAND2_X2 U11484 ( .A1(n10280), .A2(n10246), .ZN(n10250) );
  INV_X4 U11485 ( .A(n10425), .ZN(n10366) );
  NAND3_X2 U11486 ( .A1(n10251), .A2(n10250), .A3(n10249), .ZN(n10252) );
  MUX2_X2 U11487 ( .A(n10252), .B(multOut[14]), .S(net76452), .Z(n10258) );
  XNOR2_X2 U11488 ( .A(n10254), .B(n10253), .ZN(n10256) );
  NAND2_X2 U11489 ( .A1(net71078), .A2(\WIRE_ALU_A/MUX2TO1_32BIT[14].MUX/N1 ), 
        .ZN(n10255) );
  NOR2_X4 U11490 ( .A1(n10258), .A2(n10257), .ZN(n10263) );
  INV_X4 U11491 ( .A(n10263), .ZN(dmem_addr_out[14]) );
  OAI211_X2 U11492 ( .C1(n10263), .C2(net76646), .A(net70740), .B(n10262), 
        .ZN(n10264) );
  NAND2_X2 U11493 ( .A1(reset), .A2(n10264), .ZN(n10276) );
  OAI22_X2 U11494 ( .A1(n5029), .A2(n6090), .B1(net76658), .B2(n10276), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11495 ( .A1(n5844), .A2(n10512), .B1(n6155), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11496 ( .A(n5777), .ZN(n10265) );
  OAI22_X2 U11497 ( .A1(n6193), .A2(n10265), .B1(n6194), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11498 ( .A1(n6197), .A2(n10266), .B1(n6198), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11499 ( .A1(n5843), .A2(n6099), .B1(n6094), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11500 ( .A1(n4928), .A2(n6104), .B1(n10519), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11501 ( .A(\REGFILE/reg_out[15][14] ), .ZN(n10267) );
  OAI22_X2 U11502 ( .A1(n10267), .A2(n6110), .B1(n6105), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11503 ( .A1(n5819), .A2(n6111), .B1(n6157), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11504 ( .A1(n4929), .A2(n6114), .B1(n6159), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11505 ( .A1(n5842), .A2(n6117), .B1(n6161), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11506 ( .A1(n6201), .A2(n5394), .B1(n6203), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11507 ( .A1(n5841), .A2(net76866), .B1(net76614), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11508 ( .A(n5781), .ZN(n10268) );
  OAI22_X2 U11509 ( .A1(n6206), .A2(n10268), .B1(n6207), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11510 ( .A1(n4930), .A2(n6120), .B1(n6163), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11511 ( .A1(n5837), .A2(n6123), .B1(n6165), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11512 ( .A1(n4931), .A2(n6126), .B1(n6167), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11513 ( .A1(n5662), .A2(n6131), .B1(n6169), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11514 ( .A1(n10269), .A2(n6134), .B1(n6171), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11515 ( .A1(n4936), .A2(n6135), .B1(n6173), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11516 ( .A1(n6210), .A2(n10270), .B1(n6211), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11517 ( .A1(n10608), .A2(\REGFILE/reg_out[29][14] ), .ZN(n10272)
         );
  OAI22_X2 U11518 ( .A1(n5838), .A2(n6141), .B1(net76548), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11519 ( .A1(n10615), .A2(\REGFILE/reg_out[30][14] ), .ZN(n10273)
         );
  NAND2_X2 U11520 ( .A1(net76488), .A2(\REGFILE/reg_out[31][14] ), .ZN(n10274)
         );
  OAI22_X2 U11521 ( .A1(n6216), .A2(n4981), .B1(net76318), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11522 ( .A1(n6218), .A2(n5395), .B1(n6219), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11523 ( .A(n5832), .ZN(n10275) );
  OAI22_X2 U11524 ( .A1(n10275), .A2(n6143), .B1(n6182), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11525 ( .A1(n4926), .A2(net76716), .B1(n6146), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11526 ( .A1(n4932), .A2(net76702), .B1(n6184), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11527 ( .A1(n4918), .A2(n6149), .B1(n6186), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11528 ( .A1(n4933), .A2(n6152), .B1(n6188), .B2(n6085), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[14].REGISTER1/STORE_DATA/N3 ) );
  AOI22_X2 U11529 ( .A1(net71092), .A2(n10278), .B1(net71094), .B2(n10277), 
        .ZN(n10285) );
  NAND2_X2 U11530 ( .A1(n10280), .A2(n10279), .ZN(n10284) );
  NAND3_X2 U11531 ( .A1(n10285), .A2(n10284), .A3(n10283), .ZN(n10286) );
  MUX2_X2 U11532 ( .A(n10286), .B(multOut[15]), .S(net76452), .Z(n10292) );
  XNOR2_X2 U11533 ( .A(n10287), .B(n4807), .ZN(n10290) );
  NAND2_X2 U11534 ( .A1(net71078), .A2(\WIRE_ALU_A/MUX2TO1_32BIT[15].MUX/N1 ), 
        .ZN(n10289) );
  NOR2_X4 U11535 ( .A1(n10292), .A2(n10291), .ZN(n10296) );
  INV_X4 U11536 ( .A(n10296), .ZN(dmem_addr_out[15]) );
  INV_X4 U11537 ( .A(\SELECT_CORRECT_SEGMENTS/selHalf [31]), .ZN(n10504) );
  OAI211_X2 U11538 ( .C1(n10296), .C2(net76646), .A(net70740), .B(n10295), 
        .ZN(n10297) );
  OAI22_X2 U11539 ( .A1(n5250), .A2(n6090), .B1(net76658), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11540 ( .A1(n10298), .A2(n10512), .B1(n6155), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11541 ( .A1(n6193), .A2(n5121), .B1(n6194), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11542 ( .A1(n6197), .A2(n5856), .B1(n6198), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11543 ( .A1(n5714), .A2(n6099), .B1(n6094), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11544 ( .A1(n4941), .A2(n6103), .B1(n10519), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11545 ( .A1(n5866), .A2(n6110), .B1(n6105), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11546 ( .A1(n4954), .A2(n6111), .B1(n6157), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11547 ( .A1(n4942), .A2(n6114), .B1(n6159), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11548 ( .A1(n4901), .A2(n6117), .B1(n6161), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11549 ( .A1(n6201), .A2(n5122), .B1(n6203), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11550 ( .A1(n5656), .A2(net76866), .B1(net76614), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11551 ( .A1(n6206), .A2(n5431), .B1(n6207), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11552 ( .A1(n4943), .A2(n6120), .B1(n6163), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11553 ( .A1(n4919), .A2(n6123), .B1(n6165), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11554 ( .A1(n4934), .A2(n6126), .B1(n6167), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11555 ( .A1(n5251), .A2(n6131), .B1(n6169), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11556 ( .A1(n5784), .A2(n6134), .B1(n6171), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11557 ( .A1(n4944), .A2(n6135), .B1(n6173), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11558 ( .A1(n6210), .A2(n5683), .B1(n6211), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11559 ( .A1(n10608), .A2(\REGFILE/reg_out[29][15] ), .ZN(n10300)
         );
  OAI22_X2 U11560 ( .A1(n5917), .A2(n6141), .B1(net76548), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11561 ( .A1(n10615), .A2(\REGFILE/reg_out[30][15] ), .ZN(n10301)
         );
  NAND2_X2 U11562 ( .A1(net76488), .A2(\REGFILE/reg_out[31][15] ), .ZN(n10302)
         );
  OAI22_X2 U11563 ( .A1(n6216), .A2(n5038), .B1(net76318), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11564 ( .A1(n6218), .A2(n5396), .B1(n6219), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11565 ( .A1(n4902), .A2(n6143), .B1(n6182), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11566 ( .A1(n4948), .A2(net76716), .B1(n6146), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11567 ( .A1(n4945), .A2(net76702), .B1(n6184), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11568 ( .A1(n4927), .A2(n6149), .B1(n6186), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11569 ( .A1(n4935), .A2(n6152), .B1(n6188), .B2(n6087), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11570 ( .A1(n10303), .A2(net77040), .ZN(n10305) );
  XNOR2_X2 U11571 ( .A(net80189), .B(n10928), .ZN(n10434) );
  INV_X4 U11572 ( .A(n10434), .ZN(n10459) );
  NAND2_X2 U11573 ( .A1(n10306), .A2(n10399), .ZN(n10308) );
  XNOR2_X2 U11574 ( .A(net71027), .B(net70535), .ZN(net70703) );
  NOR2_X4 U11575 ( .A1(n10470), .A2(n10434), .ZN(n10311) );
  OAI21_X4 U11576 ( .B1(n10311), .B2(n10310), .A(n10309), .ZN(n10314) );
  AOI21_X4 U11577 ( .B1(n10442), .B2(n10314), .A(n10313), .ZN(n10318) );
  OAI21_X4 U11578 ( .B1(n10318), .B2(n10317), .A(n10316), .ZN(n10322) );
  INV_X4 U11579 ( .A(n10436), .ZN(n10321) );
  AOI21_X4 U11580 ( .B1(n10322), .B2(n10321), .A(n10320), .ZN(n10326) );
  NAND2_X2 U11581 ( .A1(aluA[26]), .A2(n10323), .ZN(n10324) );
  OAI21_X4 U11582 ( .B1(n10326), .B2(n10325), .A(n10324), .ZN(n10330) );
  INV_X4 U11583 ( .A(n10435), .ZN(n10329) );
  AOI21_X4 U11584 ( .B1(n10330), .B2(n10329), .A(n10328), .ZN(n10333) );
  OAI21_X4 U11585 ( .B1(n10430), .B2(n10333), .A(n10332), .ZN(n10337) );
  AOI21_X4 U11586 ( .B1(n10337), .B2(n10336), .A(n10335), .ZN(n10340) );
  NAND2_X2 U11587 ( .A1(n10932), .A2(n10338), .ZN(n10339) );
  OAI21_X4 U11588 ( .B1(n10432), .B2(n10340), .A(n10339), .ZN(n10344) );
  INV_X4 U11589 ( .A(n10443), .ZN(n10347) );
  INV_X4 U11590 ( .A(aluA[19]), .ZN(n10349) );
  INV_X4 U11591 ( .A(aluA[17]), .ZN(n10356) );
  INV_X4 U11592 ( .A(n10447), .ZN(n10360) );
  OAI21_X4 U11593 ( .B1(n10361), .B2(n10360), .A(n10359), .ZN(n10363) );
  OAI21_X4 U11594 ( .B1(n10374), .B2(n10373), .A(n10372), .ZN(n10377) );
  INV_X4 U11595 ( .A(n10411), .ZN(n10413) );
  OAI21_X4 U11596 ( .B1(n10413), .B2(n10416), .A(n10412), .ZN(n10486) );
  NAND2_X2 U11597 ( .A1(net70703), .A2(n10486), .ZN(net70838) );
  OAI21_X4 U11598 ( .B1(net70703), .B2(n10486), .A(net70838), .ZN(n10485) );
  INV_X4 U11599 ( .A(n10485), .ZN(n10417) );
  NOR4_X2 U11600 ( .A1(n10417), .A2(n10416), .A3(n10415), .A4(n10414), .ZN(
        n10454) );
  NAND2_X2 U11601 ( .A1(n10425), .A2(n10424), .ZN(n10426) );
  NOR3_X4 U11602 ( .A1(n10428), .A2(n10427), .A3(n10426), .ZN(n10453) );
  NAND2_X2 U11603 ( .A1(n10434), .A2(n10433), .ZN(n10437) );
  NAND4_X2 U11604 ( .A1(n10455), .A2(n10454), .A3(n10453), .A4(n10452), .ZN(
        n10456) );
  INV_X4 U11605 ( .A(n10456), .ZN(n10484) );
  MUX2_X2 U11606 ( .A(n10459), .B(n10458), .S(n10457), .Z(n10460) );
  NOR2_X4 U11607 ( .A1(n10461), .A2(n10460), .ZN(n10477) );
  OAI221_X2 U11608 ( .B1(net70866), .B2(n10464), .C1(net70868), .C2(n10463), 
        .A(n10462), .ZN(n10469) );
  INV_X4 U11609 ( .A(n10466), .ZN(n10467) );
  NOR2_X4 U11610 ( .A1(n10467), .A2(n10544), .ZN(n10468) );
  AOI211_X4 U11611 ( .C1(n10469), .C2(net105360), .A(n4811), .B(n10468), .ZN(
        n10473) );
  OAI221_X2 U11612 ( .B1(n4812), .B2(n10474), .C1(n10473), .C2(n10472), .A(
        n10471), .ZN(n10480) );
  NAND2_X2 U11613 ( .A1(n10480), .A2(n10475), .ZN(n10476) );
  MUX2_X2 U11614 ( .A(n10477), .B(n10476), .S(net70826), .Z(n10478) );
  NAND4_X2 U11615 ( .A1(net77040), .A2(n10494), .A3(net70826), .A4(n10484), 
        .ZN(n10479) );
  NAND2_X2 U11616 ( .A1(n10478), .A2(n10479), .ZN(n10501) );
  INV_X4 U11617 ( .A(n10479), .ZN(n10483) );
  INV_X4 U11618 ( .A(n10480), .ZN(n10481) );
  NOR2_X4 U11619 ( .A1(n10481), .A2(net70845), .ZN(n10482) );
  NOR2_X4 U11620 ( .A1(n10483), .A2(n10482), .ZN(n10499) );
  XNOR2_X2 U11621 ( .A(n10486), .B(n10485), .ZN(n10487) );
  XNOR2_X2 U11622 ( .A(n10487), .B(net70837), .ZN(n10489) );
  NAND2_X2 U11623 ( .A1(n10488), .A2(n10489), .ZN(n10497) );
  INV_X4 U11624 ( .A(n10489), .ZN(n10495) );
  MUX2_X2 U11625 ( .A(n10492), .B(n10491), .S(n10490), .Z(n10493) );
  MUX2_X2 U11626 ( .A(n10497), .B(n10496), .S(net70826), .Z(n10498) );
  NAND2_X2 U11627 ( .A1(n10499), .A2(n10498), .ZN(n10500) );
  MUX2_X2 U11628 ( .A(n10501), .B(n10500), .S(net70821), .Z(n10502) );
  MUX2_X2 U11629 ( .A(n10502), .B(multOut[31]), .S(net76452), .Z(
        dmem_addr_out[31]) );
  AOI22_X2 U11630 ( .A1(dmem_read_in[31]), .A2(net76468), .B1(
        instructionAddr_out[31]), .B2(net77030), .ZN(n10510) );
  INV_X4 U11631 ( .A(dmem_addr_out[31]), .ZN(n10503) );
  NOR3_X4 U11632 ( .A1(n10508), .A2(n10507), .A3(n10506), .ZN(n10509) );
  AOI21_X4 U11633 ( .B1(n10510), .B2(n10509), .A(net76278), .ZN(n10511) );
  OAI22_X2 U11634 ( .A1(n10513), .A2(n10512), .B1(n6191), .B2(n6155), .ZN(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11635 ( .A(\REGFILE/reg_out[11][31] ), .ZN(n10514) );
  OAI22_X2 U11636 ( .A1(n6193), .A2(n10514), .B1(n6194), .B2(n6191), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11637 ( .A1(n6197), .A2(n10515), .B1(n6198), .B2(n6191), .ZN(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11638 ( .A1(n10518), .A2(n6099), .B1(n6191), .B2(n6094), .ZN(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11639 ( .A1(n10520), .A2(n6103), .B1(n6191), .B2(n6102), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11640 ( .A1(n10522), .A2(n6110), .B1(n6191), .B2(n6105), .ZN(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11641 ( .A1(n10523), .A2(n6111), .B1(n6191), .B2(n6157), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11642 ( .A1(n4917), .A2(n6114), .B1(n6191), .B2(n6159), .ZN(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11643 ( .A1(n10524), .A2(n6117), .B1(n6191), .B2(n6161), .ZN(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11644 ( .A1(n6201), .A2(n5026), .B1(n6203), .B2(n6191), .ZN(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11645 ( .A1(net70780), .A2(net76866), .B1(n6191), .B2(net76614), 
        .ZN(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11646 ( .A1(n6206), .A2(n10525), .B1(n6207), .B2(n6191), .ZN(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11647 ( .A1(n4939), .A2(n6120), .B1(n6191), .B2(n6163), .ZN(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11648 ( .A(\REGFILE/reg_out[22][31] ), .ZN(n10526) );
  OAI22_X2 U11649 ( .A1(n10526), .A2(n6123), .B1(n6191), .B2(n6165), .ZN(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11650 ( .A1(n4953), .A2(n6126), .B1(n6191), .B2(n6167), .ZN(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11651 ( .A1(n5999), .A2(n6131), .B1(n6191), .B2(n6169), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11652 ( .A(\REGFILE/reg_out[25][31] ), .ZN(n10527) );
  OAI22_X2 U11653 ( .A1(n10527), .A2(n6134), .B1(n6191), .B2(n6171), .ZN(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11654 ( .A(\REGFILE/reg_out[26][31] ), .ZN(n10528) );
  OAI22_X2 U11655 ( .A1(n10528), .A2(n6135), .B1(n6191), .B2(n6173), .ZN(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11656 ( .A(\REGFILE/reg_out[27][31] ), .ZN(n10529) );
  OAI22_X2 U11657 ( .A1(n6210), .A2(n10529), .B1(n6211), .B2(n6191), .ZN(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11658 ( .A1(\REGFILE/reg_out[28][31] ), .A2(n6175), .ZN(n10530) );
  NAND2_X2 U11659 ( .A1(n6178), .A2(\REGFILE/reg_out[29][31] ), .ZN(n10531) );
  OAI22_X2 U11660 ( .A1(net70761), .A2(n6141), .B1(n6191), .B2(net76548), .ZN(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11661 ( .A1(n6180), .A2(\REGFILE/reg_out[30][31] ), .ZN(n10533) );
  INV_X4 U11662 ( .A(\REGFILE/reg_out[3][31] ), .ZN(net70758) );
  OAI22_X2 U11663 ( .A1(n6216), .A2(net70758), .B1(net76318), .B2(n6191), .ZN(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11664 ( .A1(n6218), .A2(net70757), .B1(n6219), .B2(n6191), .ZN(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11665 ( .A(\REGFILE/reg_out[5][31] ), .ZN(net70755) );
  OAI22_X2 U11666 ( .A1(net70755), .A2(n6143), .B1(n6191), .B2(n6182), .ZN(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11667 ( .A(\REGFILE/reg_out[6][31] ), .ZN(net70752) );
  OAI22_X2 U11668 ( .A1(net70752), .A2(net76716), .B1(n6191), .B2(n6146), .ZN(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11669 ( .A(\REGFILE/reg_out[7][31] ), .ZN(net70750) );
  OAI22_X2 U11670 ( .A1(net70750), .A2(net76702), .B1(n6191), .B2(n6184), .ZN(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  INV_X4 U11671 ( .A(\REGFILE/reg_out[8][31] ), .ZN(n10536) );
  OAI22_X2 U11672 ( .A1(n10536), .A2(n6149), .B1(n6191), .B2(n6186), .ZN(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U11673 ( .A1(n10537), .A2(n6152), .B1(n6191), .B2(n6188), .ZN(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11674 ( .A1(instructionAddr_out[1]), .A2(n10538), .ZN(n10539) );
  XNOR2_X2 U11675 ( .A(n10539), .B(n5439), .ZN(n10644) );
  OAI211_X2 U11676 ( .C1(net70738), .C2(n10644), .A(n5572), .B(net70740), .ZN(
        net70737) );
  INV_X4 U11677 ( .A(net70737), .ZN(net70685) );
  INV_X4 U11678 ( .A(n10541), .ZN(n10545) );
  NAND2_X2 U11679 ( .A1(n10542), .A2(net70534), .ZN(n10543) );
  OAI21_X4 U11680 ( .B1(n10545), .B2(n10544), .A(n10543), .ZN(net70714) );
  INV_X4 U11681 ( .A(net70687), .ZN(net70684) );
  NAND2_X2 U11682 ( .A1(n10546), .A2(net76510), .ZN(n10548) );
  NAND2_X2 U11683 ( .A1(n10549), .A2(net76510), .ZN(n10551) );
  NAND2_X2 U11684 ( .A1(n6093), .A2(\REGFILE/reg_out[10][0] ), .ZN(n10550) );
  NAND2_X2 U11685 ( .A1(n10552), .A2(net76510), .ZN(n10554) );
  NAND2_X2 U11686 ( .A1(\REGFILE/reg_out[11][0] ), .A2(n4869), .ZN(n10553) );
  NAND2_X2 U11687 ( .A1(n10555), .A2(net76510), .ZN(n10557) );
  NAND2_X2 U11688 ( .A1(\REGFILE/reg_out[12][0] ), .A2(n4873), .ZN(n10556) );
  NAND2_X2 U11690 ( .A1(n4805), .A2(\REGFILE/reg_out[14][0] ), .ZN(n10560) );
  NAND2_X2 U11691 ( .A1(n4804), .A2(\REGFILE/reg_out[15][0] ), .ZN(n10562) );
  NAND2_X2 U11692 ( .A1(n10564), .A2(net76510), .ZN(n10566) );
  NAND2_X2 U11693 ( .A1(n4891), .A2(\REGFILE/reg_out[16][0] ), .ZN(n10565) );
  NAND2_X2 U11694 ( .A1(n10567), .A2(net76510), .ZN(n10569) );
  NAND2_X2 U11695 ( .A1(n10570), .A2(net76510), .ZN(n10572) );
  NAND2_X2 U11696 ( .A1(n4884), .A2(\REGFILE/reg_out[18][0] ), .ZN(n10571) );
  NAND2_X2 U11697 ( .A1(n10573), .A2(net76510), .ZN(n10575) );
  NAND2_X2 U11698 ( .A1(\REGFILE/reg_out[19][0] ), .A2(n4876), .ZN(n10574) );
  NAND2_X2 U11699 ( .A1(n10576), .A2(net76510), .ZN(n10578) );
  NAND2_X2 U11700 ( .A1(n4877), .A2(\REGFILE/reg_out[1][0] ), .ZN(n10577) );
  NAND2_X2 U11701 ( .A1(n10579), .A2(net76510), .ZN(n10581) );
  NAND2_X2 U11703 ( .A1(n10582), .A2(net76510), .ZN(n10584) );
  NAND2_X2 U11704 ( .A1(n4882), .A2(\REGFILE/reg_out[21][0] ), .ZN(n10583) );
  NAND2_X2 U11705 ( .A1(n10585), .A2(net76510), .ZN(n10587) );
  NAND2_X2 U11706 ( .A1(n4888), .A2(\REGFILE/reg_out[22][0] ), .ZN(n10586) );
  NAND2_X2 U11707 ( .A1(n10588), .A2(net76510), .ZN(n10590) );
  NAND2_X2 U11709 ( .A1(n10591), .A2(net76510), .ZN(n10593) );
  NAND2_X2 U11710 ( .A1(n4875), .A2(\REGFILE/reg_out[24][0] ), .ZN(n10592) );
  NAND2_X2 U11711 ( .A1(n10594), .A2(net76510), .ZN(n10596) );
  NAND2_X2 U11712 ( .A1(n4878), .A2(\REGFILE/reg_out[25][0] ), .ZN(n10595) );
  NAND2_X2 U11713 ( .A1(n10597), .A2(net76510), .ZN(n10599) );
  NAND2_X2 U11714 ( .A1(n4893), .A2(\REGFILE/reg_out[26][0] ), .ZN(n10598) );
  NAND2_X2 U11715 ( .A1(n10600), .A2(net76510), .ZN(n10602) );
  NAND2_X2 U11716 ( .A1(\REGFILE/reg_out[27][0] ), .A2(n4872), .ZN(n10601) );
  NAND2_X2 U11717 ( .A1(n10603), .A2(net76510), .ZN(n10606) );
  NAND2_X2 U11718 ( .A1(\REGFILE/reg_out[28][0] ), .A2(n6175), .ZN(n10605) );
  NAND2_X2 U11719 ( .A1(n10608), .A2(\REGFILE/reg_out[29][0] ), .ZN(n10609) );
  NAND2_X2 U11720 ( .A1(n10611), .A2(net76510), .ZN(n10613) );
  NAND2_X2 U11722 ( .A1(n10615), .A2(\REGFILE/reg_out[30][0] ), .ZN(n10616) );
  NAND2_X2 U11724 ( .A1(n10620), .A2(net76510), .ZN(n10622) );
  NAND2_X2 U11725 ( .A1(\REGFILE/reg_out[3][0] ), .A2(n4871), .ZN(n10621) );
  NAND2_X2 U11726 ( .A1(n10623), .A2(net76510), .ZN(n10625) );
  NAND2_X2 U11727 ( .A1(\REGFILE/reg_out[4][0] ), .A2(n4870), .ZN(n10624) );
  NAND2_X2 U11728 ( .A1(n10626), .A2(net76510), .ZN(n10628) );
  NAND2_X2 U11729 ( .A1(n4885), .A2(\REGFILE/reg_out[5][0] ), .ZN(n10627) );
  NAND2_X2 U11731 ( .A1(n10631), .A2(net76510), .ZN(n10633) );
  NAND2_X2 U11733 ( .A1(n10634), .A2(net76510), .ZN(n10636) );
  NAND2_X2 U11735 ( .A1(net76510), .A2(n10637), .ZN(n10639) );
  INV_X4 U11737 ( .A(net70535), .ZN(net70534) );
  NAND2_X2 U11738 ( .A1(net73708), .A2(net70534), .ZN(n10648) );
  INV_X4 U11739 ( .A(n10640), .ZN(n10641) );
  XNOR2_X2 U11740 ( .A(n10641), .B(net70529), .ZN(n10642) );
  INV_X4 U11741 ( .A(n10642), .ZN(n10643) );
  NAND2_X2 U11742 ( .A1(n10649), .A2(n10643), .ZN(n10645) );
  MUX2_X2 U11743 ( .A(n10646), .B(n10645), .S(n10644), .Z(n10647) );
  NAND2_X2 U11744 ( .A1(n10648), .A2(n10647), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11745 ( .A1(n10649), .A2(\PCLOGIC/imm16_32 [31]), .ZN(n10653) );
  MUX2_X2 U11746 ( .A(n10653), .B(n10652), .S(instructionAddr_out[31]), .Z(
        n10654) );
  NAND2_X2 U11747 ( .A1(n10655), .A2(n10654), .ZN(
        \PCLOGIC/PC_REG/REG_32BIT[31].REGISTER1/STORE_DATA/N3 ) );
  NAND2_X2 U11748 ( .A1(net76488), .A2(\REGFILE/reg_out[31][31] ), .ZN(n10656)
         );
  INV_X4 U11749 ( .A(net70506), .ZN(dmem_writeEnable_out) );
  INV_X4 U11750 ( .A(\REGFILE/reg_out[20][29] ), .ZN(n10935) );
  INV_X4 U11751 ( .A(\REGFILE/reg_out[28][30] ), .ZN(n10937) );
  INV_X4 U11752 ( .A(\REGFILE/reg_out[27][30] ), .ZN(n10938) );
  INV_X4 U11753 ( .A(\REGFILE/reg_out[20][30] ), .ZN(n10939) );
  INV_X4 U11754 ( .A(\REGFILE/reg_out[12][30] ), .ZN(n10940) );
  INV_X4 U11755 ( .A(\REGFILE/reg_out[11][30] ), .ZN(n10941) );
  single_cycle_DW02_mult_0 \MULT/mult_6  ( .A({net70534, 
        \WIRE_ALU_A/MUX2TO1_32BIT[1].MUX/N1 , 
        \WIRE_ALU_A/MUX2TO1_32BIT[2].MUX/N1 , 
        \WIRE_ALU_A/MUX2TO1_32BIT[3].MUX/N1 , 
        \WIRE_ALU_A/MUX2TO1_32BIT[4].MUX/N1 , 
        \WIRE_ALU_A/MUX2TO1_32BIT[5].MUX/N1 , 
        \WIRE_ALU_A/MUX2TO1_32BIT[6].MUX/N1 , 
        \WIRE_ALU_A/MUX2TO1_32BIT[7].MUX/N1 , 
        \WIRE_ALU_A/MUX2TO1_32BIT[8].MUX/N1 , 
        \WIRE_ALU_A/MUX2TO1_32BIT[9].MUX/N1 , 
        \WIRE_ALU_A/MUX2TO1_32BIT[10].MUX/N1 , 
        \WIRE_ALU_A/MUX2TO1_32BIT[11].MUX/N1 , 
        \WIRE_ALU_A/MUX2TO1_32BIT[12].MUX/N1 , 
        \WIRE_ALU_A/MUX2TO1_32BIT[13].MUX/N1 , 
        \WIRE_ALU_A/MUX2TO1_32BIT[14].MUX/N1 , 
        \WIRE_ALU_A/MUX2TO1_32BIT[15].MUX/N1 , aluA[16:20], n10933, n10932, 
        n10931, net36391, n10930, aluA[26], n5761, n6007, aluA[29:31]}), .B({
        net36488, net36466, n10907, n10908, n10909, n10910, n10911, net36479, 
        n10912, n10913, n10914, n10915, n5943, net36470, n10916, n5851, n10917, 
        net36463, n5759, n10918, n10919, n10920, n10921, n10922, n10923, 
        n10924, n10925, n10929, n10926, n6005, net78051, n10928}), .TC(1'b0), 
        .PRODUCT({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, multOut}) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][0] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][0] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][5] ), .QN(n5415) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][5] ), .QN(n5312) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][5] ), .QN(n5311) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][4] ), .QN(n5465) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][4] ), .QN(n5329) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][4] ), .QN(n5526) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][4] ), .QN(n5525) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][4] ), .QN(n5438) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][4] ), .QN(n5524) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][4] ), .QN(n5528) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][4] ), .QN(n5467) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][4] ), .QN(n5466) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][4] ), .QN(n5331) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][4] ), .QN(n5469) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][4] ), .QN(n5048) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][4] ), .QN(n5527) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][4] ), .QN(n5529) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][4] ), .QN(n5330) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][4] ), .QN(n5424) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][4] ), .QN(n5423) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][4] ), .QN(n5557) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][2] ), .QN(n4989) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][2] ), .QN(n5347) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][2] ), .QN(n5482) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][2] ), .QN(n5537) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][2] ), .QN(n5539) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][2] ), .QN(n5348) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][2] ), .QN(n5479) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][2] ), .QN(n5538) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][2] ), .QN(n5477) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][2] ), .QN(n5483) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][2] ), .QN(n5481) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][2] ), .QN(n5478) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][2] ), .QN(n5560) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][2] ), .QN(n5561) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][2] ), .QN(n5541) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][2] ), .QN(n5540) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][2] ), .QN(n5480) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][2] ), .QN(n5536) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][3] ), .QN(n5338) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][3] ), .QN(n5558) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][3] ), .QN(n5427) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][3] ), .QN(n5230) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][3] ), .QN(n5339) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][3] ), .QN(n5229) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][3] ), .QN(n5472) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][3] ), .QN(n5532) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][3] ), .QN(n5228) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][3] ), .QN(n5470) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][3] ), .QN(n5535) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][3] ), .QN(n5473) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][3] ), .QN(n5531) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][3] ), .QN(n5471) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[30].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[30].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[30]), .QN(n5014) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[29].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[29].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[29]), .QN(n5016) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[27]), .QN(n4969) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][27] ), .QN(n5492) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][26] ), .QN(n5519) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][26] ), .QN(n5520) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[15].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[15].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[15]), .QN(n5064) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[12].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[12].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[12]), .QN(n4908) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][25] ), .QN(n5510) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][25] ), .QN(n5552) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][25] ), .QN(n5509) );
  DFF_X2 \PCLOGIC/PC_REG/REG_32BIT[11].REGISTER1/STORE_DATA/q_reg  ( .D(
        \PCLOGIC/PC_REG/REG_32BIT[11].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(
        instructionAddr_out[11]), .QN(n5060) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][23] ), .QN(n5512) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][23] ), .QN(n5511) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[27].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][27] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[26].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][26] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][25] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[25].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][25] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[23].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][23] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(n5902), .QN(n9675) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][2] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][2] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][3] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][3] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][2] ), .QN(n10121) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][2] ), .QN(n10116) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][2] ), .QN(n10117) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[13].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[13][0] ) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(n5982), .QN(n9973) );
  DFF_X1 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][5] ), .QN(n9641) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[6].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(n5764) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[15].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[15][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[0].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[0][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[27].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[27][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[26].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[26][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[25].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[25][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[22].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[22][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[21].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[21][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[19].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[19][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[18].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[18][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[16][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[12].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[12][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[4].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[4][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[3].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[3][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[1].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[1][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[10].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[10][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[6].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[6][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[17].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[17][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[2].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[2][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[23].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[23][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[20].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[20][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[9].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[9][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[8].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[8][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[7].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[7][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[5].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[5][0] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][2] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][3] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][2] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[28].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[28][4] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[31][4] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[30][4] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[4].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][4] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][5] ), .QN(n9639) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[11][5] ), .QN(n9638) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[24][5] ), .QN(n9640) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[29].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[29][5] ) );
  DFF_X2 \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/q_reg  ( 
        .D(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[0].REGISTER1/STORE_DATA/N3 ), .CK(clk), .Q(\REGFILE/reg_out[14][0] ) );
  INV_X8 U4890 ( .A(n4881), .ZN(n10945) );
  INV_X8 U4892 ( .A(n4881), .ZN(net78042) );
  AOI22_X2 U4900 ( .A1(\REGFILE/reg_out[26][18] ), .A2(net75439), .B1(n4818), 
        .B2(net75440), .ZN(n6545) );
  AOI22_X2 U4901 ( .A1(\REGFILE/reg_out[30][20] ), .A2(net84761), .B1(
        \REGFILE/reg_out[2][20] ), .B2(net82613), .ZN(n6498) );
  AOI22_X1 U4914 ( .A1(\REGFILE/reg_out[30][27] ), .A2(net77638), .B1(
        \REGFILE/reg_out[2][27] ), .B2(net75442), .ZN(n6337) );
  INV_X8 U4917 ( .A(n10947), .ZN(n10946) );
  AOI21_X4 U4929 ( .B1(net81874), .B2(n4970), .A(net76274), .ZN(n10947) );
  NAND2_X2 U4930 ( .A1(net73838), .A2(net77272), .ZN(n4830) );
  INV_X8 U4934 ( .A(net77856), .ZN(net77854) );
  INV_X1 U5036 ( .A(net73837), .ZN(n10948) );
  INV_X4 U5043 ( .A(n10948), .ZN(n10949) );
  INV_X2 U5049 ( .A(n10950), .ZN(n10951) );
  NAND2_X1 U5060 ( .A1(\REGFILE/reg_out[28][0] ), .A2(net77388), .ZN(n8237) );
  NAND2_X1 U5066 ( .A1(\REGFILE/reg_out[28][22] ), .A2(net77388), .ZN(n7267)
         );
  NAND2_X1 U5083 ( .A1(\REGFILE/reg_out[28][23] ), .A2(net77388), .ZN(n7222)
         );
  NAND2_X1 U5094 ( .A1(\REGFILE/reg_out[4][23] ), .A2(net77388), .ZN(n7232) );
  NAND2_X1 U5168 ( .A1(\REGFILE/reg_out[12][23] ), .A2(net77388), .ZN(n7242)
         );
  NAND2_X1 U5171 ( .A1(\REGFILE/reg_out[20][23] ), .A2(net77388), .ZN(n7252)
         );
  NAND2_X1 U5175 ( .A1(\REGFILE/reg_out[28][24] ), .A2(net77388), .ZN(n7177)
         );
  NAND2_X1 U5185 ( .A1(\REGFILE/reg_out[4][24] ), .A2(net77388), .ZN(n7187) );
  NAND2_X1 U5291 ( .A1(\REGFILE/reg_out[12][24] ), .A2(net77388), .ZN(n7197)
         );
  NAND2_X1 U5919 ( .A1(\REGFILE/reg_out[20][24] ), .A2(net77388), .ZN(n7207)
         );
  NAND2_X1 U6111 ( .A1(\REGFILE/reg_out[4][25] ), .A2(net77388), .ZN(n7142) );
  NAND2_X1 U6117 ( .A1(\REGFILE/reg_out[12][25] ), .A2(net77388), .ZN(n7152)
         );
  NAND2_X1 U6118 ( .A1(\REGFILE/reg_out[20][25] ), .A2(net77388), .ZN(n7162)
         );
  NAND2_X1 U6380 ( .A1(net77388), .A2(\REGFILE/reg_out[20][27] ), .ZN(n7058)
         );
  AOI22_X2 U6493 ( .A1(\REGFILE/reg_out[21][31] ), .A2(net77458), .B1(n5766), 
        .B2(net77388), .ZN(n6923) );
  NAND2_X1 U6537 ( .A1(net77298), .A2(\REGFILE/reg_out[0][28] ), .ZN(n7032) );
  NAND2_X1 U6546 ( .A1(net77298), .A2(\REGFILE/reg_out[16][28] ), .ZN(n7012)
         );
  NAND2_X1 U6547 ( .A1(\REGFILE/reg_out[16][1] ), .A2(net77300), .ZN(n8201) );
  NAND2_X1 U6679 ( .A1(net77300), .A2(\REGFILE/reg_out[0][27] ), .ZN(n7076) );
  NAND2_X1 U6756 ( .A1(\REGFILE/reg_out[0][1] ), .A2(net77300), .ZN(n8221) );
  NAND2_X1 U6833 ( .A1(\REGFILE/reg_out[8][0] ), .A2(net77300), .ZN(n8255) );
  NAND2_X1 U6834 ( .A1(\REGFILE/reg_out[24][1] ), .A2(net77300), .ZN(n8191) );
  NAND2_X1 U6895 ( .A1(\REGFILE/reg_out[8][1] ), .A2(net77300), .ZN(n8211) );
  NAND4_X2 U6947 ( .A1(net75417), .A2(net75416), .A3(net75415), .A4(net75414), 
        .ZN(net73849) );
  NAND4_X2 U6962 ( .A1(n6927), .A2(n6928), .A3(n6926), .A4(n6925), .ZN(n8401)
         );
  INV_X16 U6984 ( .A(\PCLOGIC/imm26_32 [11]), .ZN(n5574) );
  OAI22_X2 U7135 ( .A1(n9640), .A2(n6130), .B1(n6053), .B2(n6169), .ZN(
        \REGFILE/REGISTER_FILE_32[24].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U7213 ( .A1(n9639), .A2(n6104), .B1(n6054), .B2(n6102), .ZN(
        \REGFILE/REGISTER_FILE_32[14].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI22_X2 U7363 ( .A1(n6193), .A2(n9638), .B1(n6054), .B2(n6195), .ZN(
        \REGFILE/REGISTER_FILE_32[11].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  OAI211_X2 U7428 ( .C1(n9967), .C2(net76646), .A(net70740), .B(n9966), .ZN(
        n9968) );
  NOR2_X2 U7492 ( .A1(n4815), .A2(n5571), .ZN(n4898) );
  NAND2_X1 U7494 ( .A1(n4890), .A2(\REGFILE/reg_out[8][12] ), .ZN(n9174) );
  NAND2_X1 U7495 ( .A1(\REGFILE/reg_out[8][12] ), .A2(net77308), .ZN(n7729) );
  INV_X32 U7626 ( .A(\PCLOGIC/imm26_32 [8]), .ZN(net73879) );
  AOI22_X2 U8002 ( .A1(\REGFILE/reg_out[1][30] ), .A2(net77514), .B1(
        \REGFILE/reg_out[0][30] ), .B2(net77298), .ZN(n6938) );
  INV_X4 U8019 ( .A(n5842), .ZN(n10953) );
  NAND2_X2 U8072 ( .A1(net77346), .A2(\REGFILE/reg_out[18][14] ), .ZN(n7632)
         );
  INV_X4 U8082 ( .A(net76260), .ZN(net75481) );
  INV_X8 U8092 ( .A(n6050), .ZN(n6048) );
  INV_X8 U8106 ( .A(n6050), .ZN(n6049) );
  INV_X8 U8116 ( .A(n6050), .ZN(n4801) );
  OAI211_X4 U8126 ( .C1(n9519), .C2(net76646), .A(net70740), .B(n9518), .ZN(
        n9520) );
  OAI22_X2 U8136 ( .A1(n5195), .A2(n6113), .B1(n6054), .B2(n6157), .ZN(
        \REGFILE/REGISTER_FILE_32[16].REGISTER32/REG_32BIT[5].REGISTER1/STORE_DATA/N3 ) );
  INV_X8 U8151 ( .A(dmem_addr_out[5]), .ZN(n9636) );
  OAI21_X2 U8161 ( .B1(net70509), .B2(n6072), .A(n10051), .ZN(
        \REGFILE/REGISTER_FILE_32[31].REGISTER32/REG_32BIT[3].REGISTER1/STORE_DATA/N3 ) );
  AOI21_X2 U8171 ( .B1(net73878), .B2(net81974), .A(net73997), .ZN(n8374) );
  OAI21_X2 U8181 ( .B1(net77114), .B2(n10534), .A(n10120), .ZN(
        \REGFILE/REGISTER_FILE_32[30].REGISTER32/REG_32BIT[2].REGISTER1/STORE_DATA/N3 ) );
  BUF_X4 U8196 ( .A(n10924), .Z(n5762) );
  MUX2_X2 U8574 ( .A(multOut[8]), .B(n9506), .S(net73585), .Z(n9515) );
  NAND2_X4 U8581 ( .A1(multOut[7]), .A2(net92392), .ZN(n9698) );
  NAND4_X4 U8996 ( .A1(n9630), .A2(n9631), .A3(n9632), .A4(n9629), .ZN(
        dmem_addr_out[5]) );
  NAND2_X4 U9003 ( .A1(multOut[5]), .A2(net92392), .ZN(n9630) );
  NAND2_X1 U9011 ( .A1(n4886), .A2(\REGFILE/reg_out[7][0] ), .ZN(n10632) );
  NAND2_X1 U9019 ( .A1(n4890), .A2(\REGFILE/reg_out[8][0] ), .ZN(n10635) );
  NAND2_X1 U9027 ( .A1(n4883), .A2(\REGFILE/reg_out[23][0] ), .ZN(n10589) );
  NAND2_X1 U9044 ( .A1(n4887), .A2(\REGFILE/reg_out[9][0] ), .ZN(n10638) );
  NAND2_X1 U9334 ( .A1(n4879), .A2(\REGFILE/reg_out[2][0] ), .ZN(n10612) );
  NAND2_X1 U9577 ( .A1(\REGFILE/reg_out[20][0] ), .A2(n4868), .ZN(n10580) );
  NAND2_X1 U10179 ( .A1(n4889), .A2(\REGFILE/reg_out[6][0] ), .ZN(n10629) );
  NAND2_X1 U10194 ( .A1(net76488), .A2(\REGFILE/reg_out[31][0] ), .ZN(n10618)
         );
  NAND2_X1 U10574 ( .A1(n6100), .A2(\REGFILE/reg_out[13][0] ), .ZN(n10558) );
  INV_X16 U10580 ( .A(net76508), .ZN(net76502) );
  NAND2_X1 U10694 ( .A1(n4888), .A2(\REGFILE/reg_out[22][1] ), .ZN(n10194) );
  NAND2_X1 U10710 ( .A1(\REGFILE/reg_out[3][12] ), .A2(n4871), .ZN(n9164) );
  NAND2_X1 U10711 ( .A1(\REGFILE/reg_out[3][12] ), .A2(net77416), .ZN(n7742)
         );
  AOI22_X4 U10714 ( .A1(\REGFILE/reg_out[14][16] ), .A2(net77780), .B1(n5611), 
        .B2(n5664), .ZN(n6569) );
  AOI22_X4 U10715 ( .A1(\REGFILE/reg_out[14][18] ), .A2(net77780), .B1(
        \REGFILE/reg_out[13][18] ), .B2(n6009), .ZN(n6537) );
  AOI22_X4 U10718 ( .A1(\REGFILE/reg_out[0][18] ), .A2(net120684), .B1(
        \REGFILE/reg_out[10][18] ), .B2(net83203), .ZN(n6534) );
  INV_X8 U10719 ( .A(\PCLOGIC/imm26_32 [11]), .ZN(net81974) );
  INV_X32 U10721 ( .A(\PCLOGIC/imm26_32 [11]), .ZN(net82618) );
  INV_X16 U10730 ( .A(\PCLOGIC/imm26_32 [11]), .ZN(n4820) );
  INV_X2 U10731 ( .A(net77328), .ZN(net77324) );
  INV_X4 U10733 ( .A(net77328), .ZN(net77320) );
  NAND2_X1 U10767 ( .A1(net82613), .A2(n5836), .ZN(n5942) );
  AOI21_X4 U10800 ( .B1(dmem_write_out[16]), .B2(net73509), .A(n5933), .ZN(
        n11001) );
  INV_X8 U11140 ( .A(n11001), .ZN(n10917) );
  INV_X8 U11326 ( .A(net78056), .ZN(net73509) );
endmodule

