
module single_cycle ( clk, reset, instructionAddr_out, instruction, 
        dmem_addr_out, dmem_write_out, dmem_read_in, dmem_writeEnable_out, 
        dmem_dsize );
  output [0:31] instructionAddr_out;
  input [0:31] instruction;
  output [0:31] dmem_addr_out;
  output [0:31] dmem_write_out;
  input [0:31] dmem_read_in;
  output [0:1] dmem_dsize;
  input clk, reset;
  output dmem_writeEnable_out;
  wire   n10944, REGFILE_reg_out_31__31_, REGFILE_reg_out_31__30_,
         REGFILE_reg_out_31__29_, REGFILE_reg_out_31__28_,
         REGFILE_reg_out_31__27_, REGFILE_reg_out_31__26_,
         REGFILE_reg_out_31__25_, REGFILE_reg_out_31__24_,
         REGFILE_reg_out_31__23_, REGFILE_reg_out_31__22_,
         REGFILE_reg_out_31__21_, REGFILE_reg_out_31__20_,
         REGFILE_reg_out_31__19_, REGFILE_reg_out_31__18_,
         REGFILE_reg_out_31__17_, REGFILE_reg_out_31__16_,
         REGFILE_reg_out_31__15_, REGFILE_reg_out_31__14_,
         REGFILE_reg_out_31__13_, REGFILE_reg_out_31__12_,
         REGFILE_reg_out_31__11_, REGFILE_reg_out_31__10_,
         REGFILE_reg_out_31__9_, REGFILE_reg_out_31__8_,
         REGFILE_reg_out_31__7_, REGFILE_reg_out_31__6_,
         REGFILE_reg_out_31__5_, REGFILE_reg_out_31__4_,
         REGFILE_reg_out_31__3_, REGFILE_reg_out_31__2_,
         REGFILE_reg_out_31__1_, REGFILE_reg_out_31__0_,
         REGFILE_reg_out_30__31_, REGFILE_reg_out_30__30_,
         REGFILE_reg_out_30__29_, REGFILE_reg_out_30__28_,
         REGFILE_reg_out_30__27_, REGFILE_reg_out_30__26_,
         REGFILE_reg_out_30__25_, REGFILE_reg_out_30__24_,
         REGFILE_reg_out_30__23_, REGFILE_reg_out_30__22_,
         REGFILE_reg_out_30__21_, REGFILE_reg_out_30__20_,
         REGFILE_reg_out_30__19_, REGFILE_reg_out_30__18_,
         REGFILE_reg_out_30__17_, REGFILE_reg_out_30__16_,
         REGFILE_reg_out_30__15_, REGFILE_reg_out_30__14_,
         REGFILE_reg_out_30__13_, REGFILE_reg_out_30__12_,
         REGFILE_reg_out_30__11_, REGFILE_reg_out_30__10_,
         REGFILE_reg_out_30__9_, REGFILE_reg_out_30__8_,
         REGFILE_reg_out_30__7_, REGFILE_reg_out_30__6_,
         REGFILE_reg_out_30__5_, REGFILE_reg_out_30__4_,
         REGFILE_reg_out_30__3_, REGFILE_reg_out_30__2_,
         REGFILE_reg_out_30__1_, REGFILE_reg_out_30__0_,
         REGFILE_reg_out_29__31_, REGFILE_reg_out_29__30_,
         REGFILE_reg_out_29__29_, REGFILE_reg_out_29__28_,
         REGFILE_reg_out_29__27_, REGFILE_reg_out_29__26_,
         REGFILE_reg_out_29__25_, REGFILE_reg_out_29__24_,
         REGFILE_reg_out_29__23_, REGFILE_reg_out_29__22_,
         REGFILE_reg_out_29__21_, REGFILE_reg_out_29__20_,
         REGFILE_reg_out_29__19_, REGFILE_reg_out_29__18_,
         REGFILE_reg_out_29__17_, REGFILE_reg_out_29__16_,
         REGFILE_reg_out_29__15_, REGFILE_reg_out_29__14_,
         REGFILE_reg_out_29__13_, REGFILE_reg_out_29__12_,
         REGFILE_reg_out_29__11_, REGFILE_reg_out_29__10_,
         REGFILE_reg_out_29__9_, REGFILE_reg_out_29__8_,
         REGFILE_reg_out_29__7_, REGFILE_reg_out_29__6_,
         REGFILE_reg_out_29__5_, REGFILE_reg_out_29__4_,
         REGFILE_reg_out_29__3_, REGFILE_reg_out_29__2_,
         REGFILE_reg_out_29__1_, REGFILE_reg_out_29__0_,
         REGFILE_reg_out_28__31_, REGFILE_reg_out_28__30_,
         REGFILE_reg_out_28__29_, REGFILE_reg_out_28__28_,
         REGFILE_reg_out_28__27_, REGFILE_reg_out_28__26_,
         REGFILE_reg_out_28__25_, REGFILE_reg_out_28__24_,
         REGFILE_reg_out_28__23_, REGFILE_reg_out_28__22_,
         REGFILE_reg_out_28__21_, REGFILE_reg_out_28__20_,
         REGFILE_reg_out_28__19_, REGFILE_reg_out_28__18_,
         REGFILE_reg_out_28__17_, REGFILE_reg_out_28__16_,
         REGFILE_reg_out_28__15_, REGFILE_reg_out_28__14_,
         REGFILE_reg_out_28__13_, REGFILE_reg_out_28__12_,
         REGFILE_reg_out_28__11_, REGFILE_reg_out_28__10_,
         REGFILE_reg_out_28__9_, REGFILE_reg_out_28__8_,
         REGFILE_reg_out_28__7_, REGFILE_reg_out_28__6_,
         REGFILE_reg_out_28__5_, REGFILE_reg_out_28__4_,
         REGFILE_reg_out_28__3_, REGFILE_reg_out_28__2_,
         REGFILE_reg_out_28__1_, REGFILE_reg_out_28__0_,
         REGFILE_reg_out_27__31_, REGFILE_reg_out_27__30_,
         REGFILE_reg_out_27__29_, REGFILE_reg_out_27__28_,
         REGFILE_reg_out_27__27_, REGFILE_reg_out_27__26_,
         REGFILE_reg_out_27__25_, REGFILE_reg_out_27__24_,
         REGFILE_reg_out_27__23_, REGFILE_reg_out_27__22_,
         REGFILE_reg_out_27__21_, REGFILE_reg_out_27__20_,
         REGFILE_reg_out_27__19_, REGFILE_reg_out_27__18_,
         REGFILE_reg_out_27__17_, REGFILE_reg_out_27__16_,
         REGFILE_reg_out_27__15_, REGFILE_reg_out_27__14_,
         REGFILE_reg_out_27__13_, REGFILE_reg_out_27__12_,
         REGFILE_reg_out_27__11_, REGFILE_reg_out_27__10_,
         REGFILE_reg_out_27__9_, REGFILE_reg_out_27__8_,
         REGFILE_reg_out_27__7_, REGFILE_reg_out_27__6_,
         REGFILE_reg_out_27__5_, REGFILE_reg_out_27__4_,
         REGFILE_reg_out_27__3_, REGFILE_reg_out_27__2_,
         REGFILE_reg_out_27__1_, REGFILE_reg_out_27__0_,
         REGFILE_reg_out_26__31_, REGFILE_reg_out_26__30_,
         REGFILE_reg_out_26__29_, REGFILE_reg_out_26__28_,
         REGFILE_reg_out_26__27_, REGFILE_reg_out_26__26_,
         REGFILE_reg_out_26__25_, REGFILE_reg_out_26__24_,
         REGFILE_reg_out_26__23_, REGFILE_reg_out_26__22_,
         REGFILE_reg_out_26__21_, REGFILE_reg_out_26__20_,
         REGFILE_reg_out_26__19_, REGFILE_reg_out_26__18_,
         REGFILE_reg_out_26__17_, REGFILE_reg_out_26__16_,
         REGFILE_reg_out_26__15_, REGFILE_reg_out_26__14_,
         REGFILE_reg_out_26__13_, REGFILE_reg_out_26__12_,
         REGFILE_reg_out_26__11_, REGFILE_reg_out_26__10_,
         REGFILE_reg_out_26__9_, REGFILE_reg_out_26__8_,
         REGFILE_reg_out_26__7_, REGFILE_reg_out_26__6_,
         REGFILE_reg_out_26__5_, REGFILE_reg_out_26__4_,
         REGFILE_reg_out_26__3_, REGFILE_reg_out_26__2_,
         REGFILE_reg_out_26__1_, REGFILE_reg_out_26__0_,
         REGFILE_reg_out_25__31_, REGFILE_reg_out_25__30_,
         REGFILE_reg_out_25__29_, REGFILE_reg_out_25__28_,
         REGFILE_reg_out_25__27_, REGFILE_reg_out_25__26_,
         REGFILE_reg_out_25__25_, REGFILE_reg_out_25__24_,
         REGFILE_reg_out_25__23_, REGFILE_reg_out_25__22_,
         REGFILE_reg_out_25__21_, REGFILE_reg_out_25__20_,
         REGFILE_reg_out_25__19_, REGFILE_reg_out_25__18_,
         REGFILE_reg_out_25__17_, REGFILE_reg_out_25__16_,
         REGFILE_reg_out_25__15_, REGFILE_reg_out_25__14_,
         REGFILE_reg_out_25__13_, REGFILE_reg_out_25__12_,
         REGFILE_reg_out_25__11_, REGFILE_reg_out_25__10_,
         REGFILE_reg_out_25__9_, REGFILE_reg_out_25__8_,
         REGFILE_reg_out_25__7_, REGFILE_reg_out_25__5_,
         REGFILE_reg_out_25__4_, REGFILE_reg_out_25__3_,
         REGFILE_reg_out_25__2_, REGFILE_reg_out_25__1_,
         REGFILE_reg_out_25__0_, REGFILE_reg_out_24__31_,
         REGFILE_reg_out_24__30_, REGFILE_reg_out_24__29_,
         REGFILE_reg_out_24__28_, REGFILE_reg_out_24__27_,
         REGFILE_reg_out_24__26_, REGFILE_reg_out_24__25_,
         REGFILE_reg_out_24__24_, REGFILE_reg_out_24__23_,
         REGFILE_reg_out_24__22_, REGFILE_reg_out_24__21_,
         REGFILE_reg_out_24__20_, REGFILE_reg_out_24__19_,
         REGFILE_reg_out_24__18_, REGFILE_reg_out_24__17_,
         REGFILE_reg_out_24__16_, REGFILE_reg_out_24__15_,
         REGFILE_reg_out_24__14_, REGFILE_reg_out_24__13_,
         REGFILE_reg_out_24__12_, REGFILE_reg_out_24__11_,
         REGFILE_reg_out_24__10_, REGFILE_reg_out_24__9_,
         REGFILE_reg_out_24__8_, REGFILE_reg_out_24__7_,
         REGFILE_reg_out_24__6_, REGFILE_reg_out_24__5_,
         REGFILE_reg_out_24__4_, REGFILE_reg_out_24__3_,
         REGFILE_reg_out_24__2_, REGFILE_reg_out_24__1_,
         REGFILE_reg_out_24__0_, REGFILE_reg_out_23__31_,
         REGFILE_reg_out_23__30_, REGFILE_reg_out_23__29_,
         REGFILE_reg_out_23__28_, REGFILE_reg_out_23__27_,
         REGFILE_reg_out_23__26_, REGFILE_reg_out_23__25_,
         REGFILE_reg_out_23__24_, REGFILE_reg_out_23__23_,
         REGFILE_reg_out_23__22_, REGFILE_reg_out_23__21_,
         REGFILE_reg_out_23__20_, REGFILE_reg_out_23__19_,
         REGFILE_reg_out_23__18_, REGFILE_reg_out_23__17_,
         REGFILE_reg_out_23__16_, REGFILE_reg_out_23__15_,
         REGFILE_reg_out_23__14_, REGFILE_reg_out_23__13_,
         REGFILE_reg_out_23__12_, REGFILE_reg_out_23__11_,
         REGFILE_reg_out_23__10_, REGFILE_reg_out_23__9_,
         REGFILE_reg_out_23__8_, REGFILE_reg_out_23__7_,
         REGFILE_reg_out_23__6_, REGFILE_reg_out_23__5_,
         REGFILE_reg_out_23__4_, REGFILE_reg_out_23__3_,
         REGFILE_reg_out_23__2_, REGFILE_reg_out_23__1_,
         REGFILE_reg_out_23__0_, REGFILE_reg_out_22__31_,
         REGFILE_reg_out_22__30_, REGFILE_reg_out_22__29_,
         REGFILE_reg_out_22__28_, REGFILE_reg_out_22__27_,
         REGFILE_reg_out_22__26_, REGFILE_reg_out_22__25_,
         REGFILE_reg_out_22__24_, REGFILE_reg_out_22__23_,
         REGFILE_reg_out_22__22_, REGFILE_reg_out_22__21_,
         REGFILE_reg_out_22__20_, REGFILE_reg_out_22__19_,
         REGFILE_reg_out_22__18_, REGFILE_reg_out_22__17_,
         REGFILE_reg_out_22__16_, REGFILE_reg_out_22__15_,
         REGFILE_reg_out_22__14_, REGFILE_reg_out_22__13_,
         REGFILE_reg_out_22__12_, REGFILE_reg_out_22__11_,
         REGFILE_reg_out_22__10_, REGFILE_reg_out_22__9_,
         REGFILE_reg_out_22__8_, REGFILE_reg_out_22__7_,
         REGFILE_reg_out_22__6_, REGFILE_reg_out_22__5_,
         REGFILE_reg_out_22__4_, REGFILE_reg_out_22__3_,
         REGFILE_reg_out_22__2_, REGFILE_reg_out_22__1_,
         REGFILE_reg_out_22__0_, REGFILE_reg_out_21__31_,
         REGFILE_reg_out_21__30_, REGFILE_reg_out_21__29_,
         REGFILE_reg_out_21__28_, REGFILE_reg_out_21__27_,
         REGFILE_reg_out_21__26_, REGFILE_reg_out_21__25_,
         REGFILE_reg_out_21__24_, REGFILE_reg_out_21__23_,
         REGFILE_reg_out_21__22_, REGFILE_reg_out_21__21_,
         REGFILE_reg_out_21__20_, REGFILE_reg_out_21__19_,
         REGFILE_reg_out_21__18_, REGFILE_reg_out_21__17_,
         REGFILE_reg_out_21__16_, REGFILE_reg_out_21__15_,
         REGFILE_reg_out_21__14_, REGFILE_reg_out_21__13_,
         REGFILE_reg_out_21__12_, REGFILE_reg_out_21__11_,
         REGFILE_reg_out_21__10_, REGFILE_reg_out_21__9_,
         REGFILE_reg_out_21__8_, REGFILE_reg_out_21__7_,
         REGFILE_reg_out_21__6_, REGFILE_reg_out_21__5_,
         REGFILE_reg_out_21__4_, REGFILE_reg_out_21__3_,
         REGFILE_reg_out_21__2_, REGFILE_reg_out_21__1_,
         REGFILE_reg_out_21__0_, REGFILE_reg_out_20__31_,
         REGFILE_reg_out_20__30_, REGFILE_reg_out_20__29_,
         REGFILE_reg_out_20__28_, REGFILE_reg_out_20__27_,
         REGFILE_reg_out_20__26_, REGFILE_reg_out_20__25_,
         REGFILE_reg_out_20__24_, REGFILE_reg_out_20__23_,
         REGFILE_reg_out_20__22_, REGFILE_reg_out_20__21_,
         REGFILE_reg_out_20__20_, REGFILE_reg_out_20__19_,
         REGFILE_reg_out_20__18_, REGFILE_reg_out_20__17_,
         REGFILE_reg_out_20__16_, REGFILE_reg_out_20__15_,
         REGFILE_reg_out_20__14_, REGFILE_reg_out_20__13_,
         REGFILE_reg_out_20__12_, REGFILE_reg_out_20__11_,
         REGFILE_reg_out_20__10_, REGFILE_reg_out_20__9_,
         REGFILE_reg_out_20__8_, REGFILE_reg_out_20__7_,
         REGFILE_reg_out_20__6_, REGFILE_reg_out_20__5_,
         REGFILE_reg_out_20__4_, REGFILE_reg_out_20__3_,
         REGFILE_reg_out_20__2_, REGFILE_reg_out_20__1_,
         REGFILE_reg_out_20__0_, REGFILE_reg_out_19__31_,
         REGFILE_reg_out_19__30_, REGFILE_reg_out_19__29_,
         REGFILE_reg_out_19__28_, REGFILE_reg_out_19__27_,
         REGFILE_reg_out_19__26_, REGFILE_reg_out_19__25_,
         REGFILE_reg_out_19__24_, REGFILE_reg_out_19__23_,
         REGFILE_reg_out_19__22_, REGFILE_reg_out_19__21_,
         REGFILE_reg_out_19__20_, REGFILE_reg_out_19__19_,
         REGFILE_reg_out_19__18_, REGFILE_reg_out_19__17_,
         REGFILE_reg_out_19__16_, REGFILE_reg_out_19__15_,
         REGFILE_reg_out_19__14_, REGFILE_reg_out_19__13_,
         REGFILE_reg_out_19__12_, REGFILE_reg_out_19__11_,
         REGFILE_reg_out_19__10_, REGFILE_reg_out_19__9_,
         REGFILE_reg_out_19__8_, REGFILE_reg_out_19__7_,
         REGFILE_reg_out_19__6_, REGFILE_reg_out_19__5_,
         REGFILE_reg_out_19__4_, REGFILE_reg_out_19__3_,
         REGFILE_reg_out_19__2_, REGFILE_reg_out_19__1_,
         REGFILE_reg_out_19__0_, REGFILE_reg_out_18__31_,
         REGFILE_reg_out_18__30_, REGFILE_reg_out_18__29_,
         REGFILE_reg_out_18__28_, REGFILE_reg_out_18__27_,
         REGFILE_reg_out_18__26_, REGFILE_reg_out_18__25_,
         REGFILE_reg_out_18__24_, REGFILE_reg_out_18__23_,
         REGFILE_reg_out_18__22_, REGFILE_reg_out_18__21_,
         REGFILE_reg_out_18__20_, REGFILE_reg_out_18__19_,
         REGFILE_reg_out_18__18_, REGFILE_reg_out_18__17_,
         REGFILE_reg_out_18__16_, REGFILE_reg_out_18__15_,
         REGFILE_reg_out_18__14_, REGFILE_reg_out_18__13_,
         REGFILE_reg_out_18__12_, REGFILE_reg_out_18__11_,
         REGFILE_reg_out_18__10_, REGFILE_reg_out_18__9_,
         REGFILE_reg_out_18__8_, REGFILE_reg_out_18__7_,
         REGFILE_reg_out_18__6_, REGFILE_reg_out_18__5_,
         REGFILE_reg_out_18__4_, REGFILE_reg_out_18__3_,
         REGFILE_reg_out_18__2_, REGFILE_reg_out_18__1_,
         REGFILE_reg_out_18__0_, REGFILE_reg_out_17__31_,
         REGFILE_reg_out_17__30_, REGFILE_reg_out_17__29_,
         REGFILE_reg_out_17__28_, REGFILE_reg_out_17__27_,
         REGFILE_reg_out_17__26_, REGFILE_reg_out_17__25_,
         REGFILE_reg_out_17__24_, REGFILE_reg_out_17__23_,
         REGFILE_reg_out_17__22_, REGFILE_reg_out_17__21_,
         REGFILE_reg_out_17__20_, REGFILE_reg_out_17__19_,
         REGFILE_reg_out_17__18_, REGFILE_reg_out_17__17_,
         REGFILE_reg_out_17__16_, REGFILE_reg_out_17__15_,
         REGFILE_reg_out_17__14_, REGFILE_reg_out_17__13_,
         REGFILE_reg_out_17__12_, REGFILE_reg_out_17__11_,
         REGFILE_reg_out_17__10_, REGFILE_reg_out_17__9_,
         REGFILE_reg_out_17__8_, REGFILE_reg_out_17__7_,
         REGFILE_reg_out_17__6_, REGFILE_reg_out_17__5_,
         REGFILE_reg_out_17__4_, REGFILE_reg_out_17__3_,
         REGFILE_reg_out_17__2_, REGFILE_reg_out_17__1_,
         REGFILE_reg_out_17__0_, REGFILE_reg_out_16__31_,
         REGFILE_reg_out_16__30_, REGFILE_reg_out_16__29_,
         REGFILE_reg_out_16__28_, REGFILE_reg_out_16__27_,
         REGFILE_reg_out_16__26_, REGFILE_reg_out_16__25_,
         REGFILE_reg_out_16__24_, REGFILE_reg_out_16__23_,
         REGFILE_reg_out_16__22_, REGFILE_reg_out_16__21_,
         REGFILE_reg_out_16__20_, REGFILE_reg_out_16__19_,
         REGFILE_reg_out_16__18_, REGFILE_reg_out_16__17_,
         REGFILE_reg_out_16__16_, REGFILE_reg_out_16__15_,
         REGFILE_reg_out_16__14_, REGFILE_reg_out_16__13_,
         REGFILE_reg_out_16__12_, REGFILE_reg_out_16__11_,
         REGFILE_reg_out_16__10_, REGFILE_reg_out_16__9_,
         REGFILE_reg_out_16__8_, REGFILE_reg_out_16__7_,
         REGFILE_reg_out_16__6_, REGFILE_reg_out_16__5_,
         REGFILE_reg_out_16__4_, REGFILE_reg_out_16__3_,
         REGFILE_reg_out_16__2_, REGFILE_reg_out_16__1_,
         REGFILE_reg_out_16__0_, REGFILE_reg_out_15__31_,
         REGFILE_reg_out_15__30_, REGFILE_reg_out_15__29_,
         REGFILE_reg_out_15__28_, REGFILE_reg_out_15__27_,
         REGFILE_reg_out_15__26_, REGFILE_reg_out_15__25_,
         REGFILE_reg_out_15__24_, REGFILE_reg_out_15__23_,
         REGFILE_reg_out_15__22_, REGFILE_reg_out_15__21_,
         REGFILE_reg_out_15__20_, REGFILE_reg_out_15__19_,
         REGFILE_reg_out_15__18_, REGFILE_reg_out_15__17_,
         REGFILE_reg_out_15__16_, REGFILE_reg_out_15__15_,
         REGFILE_reg_out_15__14_, REGFILE_reg_out_15__13_,
         REGFILE_reg_out_15__12_, REGFILE_reg_out_15__11_,
         REGFILE_reg_out_15__10_, REGFILE_reg_out_15__9_,
         REGFILE_reg_out_15__8_, REGFILE_reg_out_15__7_,
         REGFILE_reg_out_15__6_, REGFILE_reg_out_15__5_,
         REGFILE_reg_out_15__4_, REGFILE_reg_out_15__3_,
         REGFILE_reg_out_15__2_, REGFILE_reg_out_15__1_,
         REGFILE_reg_out_15__0_, REGFILE_reg_out_14__31_,
         REGFILE_reg_out_14__30_, REGFILE_reg_out_14__29_,
         REGFILE_reg_out_14__28_, REGFILE_reg_out_14__27_,
         REGFILE_reg_out_14__26_, REGFILE_reg_out_14__25_,
         REGFILE_reg_out_14__24_, REGFILE_reg_out_14__23_,
         REGFILE_reg_out_14__22_, REGFILE_reg_out_14__21_,
         REGFILE_reg_out_14__20_, REGFILE_reg_out_14__19_,
         REGFILE_reg_out_14__18_, REGFILE_reg_out_14__17_,
         REGFILE_reg_out_14__16_, REGFILE_reg_out_14__15_,
         REGFILE_reg_out_14__14_, REGFILE_reg_out_14__13_,
         REGFILE_reg_out_14__12_, REGFILE_reg_out_14__11_,
         REGFILE_reg_out_14__10_, REGFILE_reg_out_14__9_,
         REGFILE_reg_out_14__8_, REGFILE_reg_out_14__7_,
         REGFILE_reg_out_14__6_, REGFILE_reg_out_14__5_,
         REGFILE_reg_out_14__4_, REGFILE_reg_out_14__3_,
         REGFILE_reg_out_14__2_, REGFILE_reg_out_14__1_,
         REGFILE_reg_out_14__0_, REGFILE_reg_out_13__31_,
         REGFILE_reg_out_13__30_, REGFILE_reg_out_13__29_,
         REGFILE_reg_out_13__28_, REGFILE_reg_out_13__27_,
         REGFILE_reg_out_13__26_, REGFILE_reg_out_13__25_,
         REGFILE_reg_out_13__24_, REGFILE_reg_out_13__23_,
         REGFILE_reg_out_13__22_, REGFILE_reg_out_13__21_,
         REGFILE_reg_out_13__20_, REGFILE_reg_out_13__19_,
         REGFILE_reg_out_13__18_, REGFILE_reg_out_13__17_,
         REGFILE_reg_out_13__16_, REGFILE_reg_out_13__15_,
         REGFILE_reg_out_13__14_, REGFILE_reg_out_13__13_,
         REGFILE_reg_out_13__12_, REGFILE_reg_out_13__11_,
         REGFILE_reg_out_13__10_, REGFILE_reg_out_13__9_,
         REGFILE_reg_out_13__8_, REGFILE_reg_out_13__7_,
         REGFILE_reg_out_13__6_, REGFILE_reg_out_13__5_,
         REGFILE_reg_out_13__4_, REGFILE_reg_out_13__3_,
         REGFILE_reg_out_13__2_, REGFILE_reg_out_13__1_,
         REGFILE_reg_out_13__0_, REGFILE_reg_out_12__31_,
         REGFILE_reg_out_12__30_, REGFILE_reg_out_12__29_,
         REGFILE_reg_out_12__28_, REGFILE_reg_out_12__27_,
         REGFILE_reg_out_12__26_, REGFILE_reg_out_12__25_,
         REGFILE_reg_out_12__24_, REGFILE_reg_out_12__23_,
         REGFILE_reg_out_12__22_, REGFILE_reg_out_12__21_,
         REGFILE_reg_out_12__20_, REGFILE_reg_out_12__19_,
         REGFILE_reg_out_12__18_, REGFILE_reg_out_12__17_,
         REGFILE_reg_out_12__16_, REGFILE_reg_out_12__15_,
         REGFILE_reg_out_12__13_, REGFILE_reg_out_12__12_,
         REGFILE_reg_out_12__11_, REGFILE_reg_out_12__10_,
         REGFILE_reg_out_12__9_, REGFILE_reg_out_12__8_,
         REGFILE_reg_out_12__7_, REGFILE_reg_out_12__6_,
         REGFILE_reg_out_12__5_, REGFILE_reg_out_12__4_,
         REGFILE_reg_out_12__3_, REGFILE_reg_out_12__2_,
         REGFILE_reg_out_12__1_, REGFILE_reg_out_12__0_,
         REGFILE_reg_out_11__31_, REGFILE_reg_out_11__30_,
         REGFILE_reg_out_11__29_, REGFILE_reg_out_11__28_,
         REGFILE_reg_out_11__27_, REGFILE_reg_out_11__26_,
         REGFILE_reg_out_11__25_, REGFILE_reg_out_11__24_,
         REGFILE_reg_out_11__23_, REGFILE_reg_out_11__22_,
         REGFILE_reg_out_11__21_, REGFILE_reg_out_11__20_,
         REGFILE_reg_out_11__19_, REGFILE_reg_out_11__18_,
         REGFILE_reg_out_11__17_, REGFILE_reg_out_11__16_,
         REGFILE_reg_out_11__15_, REGFILE_reg_out_11__14_,
         REGFILE_reg_out_11__13_, REGFILE_reg_out_11__12_,
         REGFILE_reg_out_11__11_, REGFILE_reg_out_11__10_,
         REGFILE_reg_out_11__9_, REGFILE_reg_out_11__8_,
         REGFILE_reg_out_11__7_, REGFILE_reg_out_11__6_,
         REGFILE_reg_out_11__5_, REGFILE_reg_out_11__4_,
         REGFILE_reg_out_11__3_, REGFILE_reg_out_11__2_,
         REGFILE_reg_out_11__1_, REGFILE_reg_out_11__0_,
         REGFILE_reg_out_10__31_, REGFILE_reg_out_10__30_,
         REGFILE_reg_out_10__29_, REGFILE_reg_out_10__28_,
         REGFILE_reg_out_10__27_, REGFILE_reg_out_10__26_,
         REGFILE_reg_out_10__25_, REGFILE_reg_out_10__24_,
         REGFILE_reg_out_10__23_, REGFILE_reg_out_10__22_,
         REGFILE_reg_out_10__21_, REGFILE_reg_out_10__20_,
         REGFILE_reg_out_10__19_, REGFILE_reg_out_10__18_,
         REGFILE_reg_out_10__17_, REGFILE_reg_out_10__16_,
         REGFILE_reg_out_10__15_, REGFILE_reg_out_10__14_,
         REGFILE_reg_out_10__13_, REGFILE_reg_out_10__12_,
         REGFILE_reg_out_10__11_, REGFILE_reg_out_10__10_,
         REGFILE_reg_out_10__9_, REGFILE_reg_out_10__8_,
         REGFILE_reg_out_10__7_, REGFILE_reg_out_10__5_,
         REGFILE_reg_out_10__4_, REGFILE_reg_out_10__3_,
         REGFILE_reg_out_10__2_, REGFILE_reg_out_10__1_,
         REGFILE_reg_out_10__0_, REGFILE_reg_out_9__31_,
         REGFILE_reg_out_9__30_, REGFILE_reg_out_9__29_,
         REGFILE_reg_out_9__28_, REGFILE_reg_out_9__27_,
         REGFILE_reg_out_9__26_, REGFILE_reg_out_9__25_,
         REGFILE_reg_out_9__24_, REGFILE_reg_out_9__23_,
         REGFILE_reg_out_9__22_, REGFILE_reg_out_9__21_,
         REGFILE_reg_out_9__20_, REGFILE_reg_out_9__19_,
         REGFILE_reg_out_9__18_, REGFILE_reg_out_9__17_,
         REGFILE_reg_out_9__16_, REGFILE_reg_out_9__15_,
         REGFILE_reg_out_9__14_, REGFILE_reg_out_9__13_,
         REGFILE_reg_out_9__12_, REGFILE_reg_out_9__11_,
         REGFILE_reg_out_9__10_, REGFILE_reg_out_9__9_, REGFILE_reg_out_9__8_,
         REGFILE_reg_out_9__7_, REGFILE_reg_out_9__6_, REGFILE_reg_out_9__5_,
         REGFILE_reg_out_9__4_, REGFILE_reg_out_9__3_, REGFILE_reg_out_9__2_,
         REGFILE_reg_out_9__1_, REGFILE_reg_out_9__0_, REGFILE_reg_out_8__31_,
         REGFILE_reg_out_8__30_, REGFILE_reg_out_8__29_,
         REGFILE_reg_out_8__28_, REGFILE_reg_out_8__27_,
         REGFILE_reg_out_8__26_, REGFILE_reg_out_8__25_,
         REGFILE_reg_out_8__24_, REGFILE_reg_out_8__23_,
         REGFILE_reg_out_8__22_, REGFILE_reg_out_8__21_,
         REGFILE_reg_out_8__20_, REGFILE_reg_out_8__19_,
         REGFILE_reg_out_8__18_, REGFILE_reg_out_8__17_,
         REGFILE_reg_out_8__16_, REGFILE_reg_out_8__15_,
         REGFILE_reg_out_8__14_, REGFILE_reg_out_8__13_,
         REGFILE_reg_out_8__12_, REGFILE_reg_out_8__11_,
         REGFILE_reg_out_8__10_, REGFILE_reg_out_8__9_, REGFILE_reg_out_8__8_,
         REGFILE_reg_out_8__7_, REGFILE_reg_out_8__6_, REGFILE_reg_out_8__5_,
         REGFILE_reg_out_8__4_, REGFILE_reg_out_8__3_, REGFILE_reg_out_8__2_,
         REGFILE_reg_out_8__1_, REGFILE_reg_out_8__0_, REGFILE_reg_out_7__31_,
         REGFILE_reg_out_7__30_, REGFILE_reg_out_7__29_,
         REGFILE_reg_out_7__28_, REGFILE_reg_out_7__27_,
         REGFILE_reg_out_7__26_, REGFILE_reg_out_7__25_,
         REGFILE_reg_out_7__24_, REGFILE_reg_out_7__23_,
         REGFILE_reg_out_7__22_, REGFILE_reg_out_7__21_,
         REGFILE_reg_out_7__20_, REGFILE_reg_out_7__19_,
         REGFILE_reg_out_7__18_, REGFILE_reg_out_7__17_,
         REGFILE_reg_out_7__16_, REGFILE_reg_out_7__15_,
         REGFILE_reg_out_7__14_, REGFILE_reg_out_7__13_,
         REGFILE_reg_out_7__12_, REGFILE_reg_out_7__11_,
         REGFILE_reg_out_7__10_, REGFILE_reg_out_7__9_, REGFILE_reg_out_7__8_,
         REGFILE_reg_out_7__7_, REGFILE_reg_out_7__6_, REGFILE_reg_out_7__5_,
         REGFILE_reg_out_7__4_, REGFILE_reg_out_7__3_, REGFILE_reg_out_7__2_,
         REGFILE_reg_out_7__1_, REGFILE_reg_out_7__0_, REGFILE_reg_out_6__31_,
         REGFILE_reg_out_6__30_, REGFILE_reg_out_6__29_,
         REGFILE_reg_out_6__28_, REGFILE_reg_out_6__27_,
         REGFILE_reg_out_6__26_, REGFILE_reg_out_6__25_,
         REGFILE_reg_out_6__24_, REGFILE_reg_out_6__23_,
         REGFILE_reg_out_6__22_, REGFILE_reg_out_6__21_,
         REGFILE_reg_out_6__20_, REGFILE_reg_out_6__19_,
         REGFILE_reg_out_6__18_, REGFILE_reg_out_6__17_,
         REGFILE_reg_out_6__16_, REGFILE_reg_out_6__15_,
         REGFILE_reg_out_6__14_, REGFILE_reg_out_6__13_,
         REGFILE_reg_out_6__12_, REGFILE_reg_out_6__11_,
         REGFILE_reg_out_6__10_, REGFILE_reg_out_6__9_, REGFILE_reg_out_6__8_,
         REGFILE_reg_out_6__7_, REGFILE_reg_out_6__6_, REGFILE_reg_out_6__5_,
         REGFILE_reg_out_6__4_, REGFILE_reg_out_6__3_, REGFILE_reg_out_6__2_,
         REGFILE_reg_out_6__1_, REGFILE_reg_out_6__0_, REGFILE_reg_out_5__31_,
         REGFILE_reg_out_5__30_, REGFILE_reg_out_5__29_,
         REGFILE_reg_out_5__28_, REGFILE_reg_out_5__27_,
         REGFILE_reg_out_5__26_, REGFILE_reg_out_5__25_,
         REGFILE_reg_out_5__24_, REGFILE_reg_out_5__23_,
         REGFILE_reg_out_5__22_, REGFILE_reg_out_5__21_,
         REGFILE_reg_out_5__20_, REGFILE_reg_out_5__19_,
         REGFILE_reg_out_5__18_, REGFILE_reg_out_5__17_,
         REGFILE_reg_out_5__16_, REGFILE_reg_out_5__15_,
         REGFILE_reg_out_5__14_, REGFILE_reg_out_5__13_,
         REGFILE_reg_out_5__12_, REGFILE_reg_out_5__11_,
         REGFILE_reg_out_5__10_, REGFILE_reg_out_5__9_, REGFILE_reg_out_5__8_,
         REGFILE_reg_out_5__7_, REGFILE_reg_out_5__6_, REGFILE_reg_out_5__5_,
         REGFILE_reg_out_5__4_, REGFILE_reg_out_5__3_, REGFILE_reg_out_5__2_,
         REGFILE_reg_out_5__1_, REGFILE_reg_out_5__0_, REGFILE_reg_out_4__31_,
         REGFILE_reg_out_4__30_, REGFILE_reg_out_4__29_,
         REGFILE_reg_out_4__28_, REGFILE_reg_out_4__27_,
         REGFILE_reg_out_4__26_, REGFILE_reg_out_4__25_,
         REGFILE_reg_out_4__24_, REGFILE_reg_out_4__23_,
         REGFILE_reg_out_4__22_, REGFILE_reg_out_4__21_,
         REGFILE_reg_out_4__20_, REGFILE_reg_out_4__19_,
         REGFILE_reg_out_4__18_, REGFILE_reg_out_4__17_,
         REGFILE_reg_out_4__16_, REGFILE_reg_out_4__15_,
         REGFILE_reg_out_4__14_, REGFILE_reg_out_4__13_,
         REGFILE_reg_out_4__12_, REGFILE_reg_out_4__11_,
         REGFILE_reg_out_4__10_, REGFILE_reg_out_4__9_, REGFILE_reg_out_4__8_,
         REGFILE_reg_out_4__7_, REGFILE_reg_out_4__6_, REGFILE_reg_out_4__5_,
         REGFILE_reg_out_4__4_, REGFILE_reg_out_4__3_, REGFILE_reg_out_4__2_,
         REGFILE_reg_out_4__1_, REGFILE_reg_out_4__0_, REGFILE_reg_out_3__31_,
         REGFILE_reg_out_3__30_, REGFILE_reg_out_3__29_,
         REGFILE_reg_out_3__28_, REGFILE_reg_out_3__27_,
         REGFILE_reg_out_3__26_, REGFILE_reg_out_3__25_,
         REGFILE_reg_out_3__24_, REGFILE_reg_out_3__23_,
         REGFILE_reg_out_3__22_, REGFILE_reg_out_3__21_,
         REGFILE_reg_out_3__20_, REGFILE_reg_out_3__19_,
         REGFILE_reg_out_3__18_, REGFILE_reg_out_3__17_,
         REGFILE_reg_out_3__16_, REGFILE_reg_out_3__15_,
         REGFILE_reg_out_3__14_, REGFILE_reg_out_3__13_,
         REGFILE_reg_out_3__12_, REGFILE_reg_out_3__11_,
         REGFILE_reg_out_3__10_, REGFILE_reg_out_3__9_, REGFILE_reg_out_3__8_,
         REGFILE_reg_out_3__7_, REGFILE_reg_out_3__6_, REGFILE_reg_out_3__5_,
         REGFILE_reg_out_3__3_, REGFILE_reg_out_3__2_, REGFILE_reg_out_3__1_,
         REGFILE_reg_out_3__0_, REGFILE_reg_out_2__31_, REGFILE_reg_out_2__30_,
         REGFILE_reg_out_2__29_, REGFILE_reg_out_2__28_,
         REGFILE_reg_out_2__27_, REGFILE_reg_out_2__26_,
         REGFILE_reg_out_2__25_, REGFILE_reg_out_2__24_,
         REGFILE_reg_out_2__23_, REGFILE_reg_out_2__22_,
         REGFILE_reg_out_2__21_, REGFILE_reg_out_2__20_,
         REGFILE_reg_out_2__19_, REGFILE_reg_out_2__18_,
         REGFILE_reg_out_2__17_, REGFILE_reg_out_2__16_,
         REGFILE_reg_out_2__15_, REGFILE_reg_out_2__14_,
         REGFILE_reg_out_2__13_, REGFILE_reg_out_2__12_,
         REGFILE_reg_out_2__11_, REGFILE_reg_out_2__10_, REGFILE_reg_out_2__9_,
         REGFILE_reg_out_2__8_, REGFILE_reg_out_2__7_, REGFILE_reg_out_2__6_,
         REGFILE_reg_out_2__5_, REGFILE_reg_out_2__4_, REGFILE_reg_out_2__3_,
         REGFILE_reg_out_2__2_, REGFILE_reg_out_2__1_, REGFILE_reg_out_2__0_,
         REGFILE_reg_out_1__31_, REGFILE_reg_out_1__30_,
         REGFILE_reg_out_1__29_, REGFILE_reg_out_1__28_,
         REGFILE_reg_out_1__27_, REGFILE_reg_out_1__26_,
         REGFILE_reg_out_1__25_, REGFILE_reg_out_1__24_,
         REGFILE_reg_out_1__23_, REGFILE_reg_out_1__22_,
         REGFILE_reg_out_1__21_, REGFILE_reg_out_1__20_,
         REGFILE_reg_out_1__19_, REGFILE_reg_out_1__18_,
         REGFILE_reg_out_1__17_, REGFILE_reg_out_1__16_,
         REGFILE_reg_out_1__15_, REGFILE_reg_out_1__14_,
         REGFILE_reg_out_1__13_, REGFILE_reg_out_1__12_,
         REGFILE_reg_out_1__11_, REGFILE_reg_out_1__10_, REGFILE_reg_out_1__9_,
         REGFILE_reg_out_1__8_, REGFILE_reg_out_1__7_, REGFILE_reg_out_1__6_,
         REGFILE_reg_out_1__5_, REGFILE_reg_out_1__4_, REGFILE_reg_out_1__3_,
         REGFILE_reg_out_1__2_, REGFILE_reg_out_1__1_, REGFILE_reg_out_1__0_,
         REGFILE_reg_out_0__31_, REGFILE_reg_out_0__30_,
         REGFILE_reg_out_0__29_, REGFILE_reg_out_0__28_,
         REGFILE_reg_out_0__27_, REGFILE_reg_out_0__26_,
         REGFILE_reg_out_0__25_, REGFILE_reg_out_0__24_,
         REGFILE_reg_out_0__23_, REGFILE_reg_out_0__22_,
         REGFILE_reg_out_0__21_, REGFILE_reg_out_0__20_,
         REGFILE_reg_out_0__19_, REGFILE_reg_out_0__18_,
         REGFILE_reg_out_0__17_, REGFILE_reg_out_0__16_,
         REGFILE_reg_out_0__15_, REGFILE_reg_out_0__14_,
         REGFILE_reg_out_0__13_, REGFILE_reg_out_0__12_,
         REGFILE_reg_out_0__11_, REGFILE_reg_out_0__10_, REGFILE_reg_out_0__9_,
         REGFILE_reg_out_0__8_, REGFILE_reg_out_0__7_, REGFILE_reg_out_0__6_,
         REGFILE_reg_out_0__5_, REGFILE_reg_out_0__4_, REGFILE_reg_out_0__3_,
         REGFILE_reg_out_0__2_, REGFILE_reg_out_0__1_, REGFILE_reg_out_0__0_,
         PCLOGIC_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         PCLOGIC_PC_REG_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         WIRE_ALU_A_MUX2TO1_32BIT_1__MUX_N1,
         WIRE_ALU_A_MUX2TO1_32BIT_2__MUX_N1,
         WIRE_ALU_A_MUX2TO1_32BIT_3__MUX_N1,
         WIRE_ALU_A_MUX2TO1_32BIT_4__MUX_N1,
         WIRE_ALU_A_MUX2TO1_32BIT_5__MUX_N1,
         WIRE_ALU_A_MUX2TO1_32BIT_6__MUX_N1,
         WIRE_ALU_A_MUX2TO1_32BIT_7__MUX_N1,
         WIRE_ALU_A_MUX2TO1_32BIT_8__MUX_N1,
         WIRE_ALU_A_MUX2TO1_32BIT_9__MUX_N1,
         WIRE_ALU_A_MUX2TO1_32BIT_10__MUX_N1,
         WIRE_ALU_A_MUX2TO1_32BIT_11__MUX_N1,
         WIRE_ALU_A_MUX2TO1_32BIT_12__MUX_N1,
         WIRE_ALU_A_MUX2TO1_32BIT_13__MUX_N1,
         WIRE_ALU_A_MUX2TO1_32BIT_14__MUX_N1,
         WIRE_ALU_A_MUX2TO1_32BIT_15__MUX_N1, net36391, net36463, net36466,
         net36470, net36479, net36488, net70506, net70507, net70509, net70529,
         net70531, net70534, net70535, net70537, net70541, net70574, net70684,
         net70685, net70687, net70696, net70697, net70701, net70703, net70706,
         net70709, net70710, net70713, net70714, net70717, net70718, net70719,
         net70720, net70727, net70731, net70734, net70735, net70737, net70738,
         net70740, net70750, net70752, net70755, net70757, net70758, net70761,
         net70780, net70811, net70821, net70826, net70837, net70838, net70845,
         net70866, net70868, net70921, net71026, net71027, net71078, net71085,
         net71092, net71094, net71271, net71273, net71277, net71280, net71299,
         net71300, net71394, net71396, net71824, net71906, net71934, net71936,
         net72163, net72312, net72876, net72947, net72962, net73166, net73167,
         net73170, net73394, net73395, net73400, net73416, net73421, net73423,
         net73429, net73434, net73436, net73439, net73443, net73468, net73494,
         net73495, net73496, net73498, net73499, net73503, net73504, net73509,
         net73510, net73512, net73519, net73527, net73529, net73532, net73541,
         net73543, net73608, net73611, net73612, net73613, net73615, net73616,
         net73619, net73620, net73622, net73629, net73630, net73637, net73638,
         net73646, net73652, net73653, net73670, net73684, net73694, net73695,
         net73696, net73697, net73708, net73771, net73778, net73780, net73831,
         net73836, net73837, net73838, net73842, net73848, net73850, net73851,
         net73855, net73858, net73877, net73878, net73879, net73900, net73902,
         net73908, net73938, net73974, net73987, net73988, net73997, net74009,
         net74011, net74051, net74359, net74361, net74799, net74808, net75367,
         net75368, net75397, net75401, net75418, net75419, net75424, net75425,
         net75427, net75437, net75438, net75439, net75440, net75441, net75442,
         net75443, net75451, net75452, net75453, net75454, net75455, net75456,
         net75464, net75466, net75468, net75469, net75475, net75478, net75479,
         net75481, net75482, net75615, net75619, net75620, net75624, net75748,
         net75759, net75761, net75764, net75791, net75792, net75793, net75843,
         net75844, net75847, net75849, net75857, net75859, net75861, net75995,
         net76025, net76031, net76032, net76034, net76154, net76195, net76199,
         net76201, net76202, net76203, net76204, net76205, net76208, net76209,
         net76211, net76217, net76220, net76222, net76234, net76238, net76239,
         net76241, net76242, net76248, net76249, net76255, net76257, net76258,
         net76259, net76260, net76261, net76278, net76274, net76270, net76320,
         net76318, net76452, net76464, net76480, net76488, net76508, net76506,
         net76502, net76514, net76510, net76550, net76548, net76616, net76614,
         net76650, net76646, net76660, net76658, net76694, net76692, net76702,
         net76708, net76706, net76716, net76866, net76864, net76862, net77030,
         net77042, net77040, net77038, net77086, net77084, net77106, net77104,
         net77102, net77100, net77116, net77114, net77276, net77272, net77292,
         net77290, net77324, net77320, net77318, net77316, net77314, net77312,
         net77310, net77308, net77306, net77304, net77302, net77300, net77298,
         net77328, net77360, net77358, net77348, net77346, net77344, net77342,
         net77338, net77336, net77396, net77394, net77392, net77388, net77386,
         net77384, net77382, net77380, net77376, net77400, net77432, net77430,
         net77428, net77426, net77424, net77422, net77420, net77418, net77416,
         net77414, net77410, net77406, net77440, net77436, net77464, net77462,
         net77460, net77458, net77456, net77454, net77452, net77444, net77474,
         net77506, net77504, net77502, net77500, net77498, net77496, net77494,
         net77492, net77490, net77488, net77484, net77482, net77480, net77478,
         net77508, net77542, net77540, net77538, net77532, net77530, net77528,
         net77526, net77524, net77522, net77520, net77518, net77516, net77514,
         net77548, net77544, net77576, net77574, net77568, net77566, net77564,
         net77562, net77560, net77558, net77556, net77554, net77550, net77588,
         net77608, net77602, net77616, net77614, net77610, net77624, net77620,
         net77618, net77632, net77630, net77626, net77640, net77638, net77634,
         net77656, net77652, net77650, net77670, net77668, net77666, net77676,
         net77704, net77702, net77700, net77698, net77720, net77716, net77714,
         net77744, net77750, net77748, net77746, net77764, net77762, net77776,
         net77774, net77784, net77780, net77778, net77800, net77798, net77796,
         net77794, net77814, net77812, net77810, net77832, net77828, net77826,
         net77836, net77834, net77848, net77846, net77844, net77842, net77856,
         net77854, net77852, net77850, net77999, net78003, net78014, net78042,
         net78051, net78056, net78055, net78109, net78108, net78107, net78128,
         net78127, net78235, net80189, net80208, net80211, net80390, net80440,
         net80443, net81764, net81810, net82342, net82500, net82499, net82515,
         net82613, net82631, net82739, net83168, net83167, net83203, net83260,
         net84475, net84518, net84663, net84754, net84761, net85047, net85371,
         net86238, net86304, net86794, net86793, net87098, net87489, net87506,
         net87633, net88131, net88253, net89184, net90830, net90864, net91311,
         net91561, net91646, net92392, net92447, net93763, net105361,
         net105360, net105352, net105349, net87820, net85731, net76219,
         net75626, net75625, net75617, net72015, net87495, net76252, net76196,
         net76194, net75621, net75618, net75616, net83210, net82738, net81164,
         net80797, net76256, net76224, net76206, net75623, net120684,
         net121496, net123282, net123932, net124970, net77296, net82513,
         net78126, net77512, net77326, net75417, net75416, net75414, net74050,
         net73849, net123931, net76181, net75396, net75395, net74029, net78050,
         net77280, net73665, net70693, net36414, net105376, net105318,
         net87097, net78105, net75422, net75415, net70732, net70730, net70729,
         net70692, net70690, net70689, net70497, net78104, net75423, net73989,
         net89734, net88102, net87806, net82932, net77816, net76253, net75477,
         net148091, net148116, net148736, net148735, net83261, net72414,
         net91643, net76262, net73533, net77752, net76254, net76235, net75763,
         net75760, net75747, net75465, net73528, net122022, net73585, net92782,
         net81874, net81873, net70691, net70504, net70503, net70502, net73500,
         net71302, net71269, net71266, net73465, net73427, net71227, net71228,
         net75842, net81974, net76251, net76233, net75862, net73511, net83408,
         net82618, net82598, net81601, net77768, net76237, net76236, net76198,
         net75860, net75858, net75845, net75467, net148494, net123382,
         net92446, net87982, net87981, net84760, net84277, net82933, net80161,
         net76197, net75846, n10943, n4797, n4798, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4849, n4850, n4851, n4852, n4853, n4854, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5576, n5577, n5578,
         n5579, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5748, n5749, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5982, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10953, n11001, MULT_mult_6_n2378, MULT_mult_6_n2377,
         MULT_mult_6_n2376, MULT_mult_6_n2375, MULT_mult_6_n2374,
         MULT_mult_6_n2373, MULT_mult_6_n2372, MULT_mult_6_n2371,
         MULT_mult_6_n2370, MULT_mult_6_n2369, MULT_mult_6_n2368,
         MULT_mult_6_n2367, MULT_mult_6_n2366, MULT_mult_6_n2365,
         MULT_mult_6_n2364, MULT_mult_6_n2363, MULT_mult_6_n2362,
         MULT_mult_6_n2361, MULT_mult_6_n2360, MULT_mult_6_n2359,
         MULT_mult_6_n2358, MULT_mult_6_n2357, MULT_mult_6_n2356,
         MULT_mult_6_n2355, MULT_mult_6_n2354, MULT_mult_6_n2353,
         MULT_mult_6_n2352, MULT_mult_6_n2351, MULT_mult_6_n2350,
         MULT_mult_6_n2349, MULT_mult_6_n2348, MULT_mult_6_n2347,
         MULT_mult_6_n2346, MULT_mult_6_n2345, MULT_mult_6_n2344,
         MULT_mult_6_n2343, MULT_mult_6_n2342, MULT_mult_6_n2341,
         MULT_mult_6_n2340, MULT_mult_6_n2339, MULT_mult_6_n2338,
         MULT_mult_6_n2337, MULT_mult_6_n2336, MULT_mult_6_n2335,
         MULT_mult_6_n2334, MULT_mult_6_n2333, MULT_mult_6_n2332,
         MULT_mult_6_n2331, MULT_mult_6_n2330, MULT_mult_6_n2329,
         MULT_mult_6_n2328, MULT_mult_6_n2327, MULT_mult_6_n2326,
         MULT_mult_6_n2325, MULT_mult_6_n2324, MULT_mult_6_n2323,
         MULT_mult_6_n2322, MULT_mult_6_n2321, MULT_mult_6_n2320,
         MULT_mult_6_n2319, MULT_mult_6_n2318, MULT_mult_6_n2317,
         MULT_mult_6_n2316, MULT_mult_6_n2315, MULT_mult_6_n2314,
         MULT_mult_6_n2313, MULT_mult_6_n2312, MULT_mult_6_n2311,
         MULT_mult_6_n2310, MULT_mult_6_n2309, MULT_mult_6_n2308,
         MULT_mult_6_n2307, MULT_mult_6_n2306, MULT_mult_6_n2305,
         MULT_mult_6_n2304, MULT_mult_6_n2303, MULT_mult_6_n2302,
         MULT_mult_6_n2301, MULT_mult_6_n2300, MULT_mult_6_n2299,
         MULT_mult_6_n2298, MULT_mult_6_n2297, MULT_mult_6_n2296,
         MULT_mult_6_n2295, MULT_mult_6_n2294, MULT_mult_6_n2293,
         MULT_mult_6_n2292, MULT_mult_6_n2291, MULT_mult_6_n2290,
         MULT_mult_6_n2289, MULT_mult_6_n2288, MULT_mult_6_n2287,
         MULT_mult_6_n2286, MULT_mult_6_n2285, MULT_mult_6_n2284,
         MULT_mult_6_n2283, MULT_mult_6_n2282, MULT_mult_6_n2281,
         MULT_mult_6_n2280, MULT_mult_6_n2279, MULT_mult_6_n2278,
         MULT_mult_6_n2277, MULT_mult_6_n2276, MULT_mult_6_n2275,
         MULT_mult_6_n2274, MULT_mult_6_n2273, MULT_mult_6_n2272,
         MULT_mult_6_n2271, MULT_mult_6_n2270, MULT_mult_6_n2269,
         MULT_mult_6_n2268, MULT_mult_6_n2267, MULT_mult_6_n2266,
         MULT_mult_6_n2265, MULT_mult_6_n2264, MULT_mult_6_n2263,
         MULT_mult_6_n2262, MULT_mult_6_n2261, MULT_mult_6_n2260,
         MULT_mult_6_n2259, MULT_mult_6_n2258, MULT_mult_6_n2257,
         MULT_mult_6_n2256, MULT_mult_6_n2255, MULT_mult_6_n2254,
         MULT_mult_6_n2253, MULT_mult_6_n2252, MULT_mult_6_n2251,
         MULT_mult_6_n2250, MULT_mult_6_n2249, MULT_mult_6_n2248,
         MULT_mult_6_n2247, MULT_mult_6_n2246, MULT_mult_6_n2245,
         MULT_mult_6_n2244, MULT_mult_6_n2243, MULT_mult_6_n2242,
         MULT_mult_6_n2241, MULT_mult_6_n2240, MULT_mult_6_n2239,
         MULT_mult_6_n2238, MULT_mult_6_n2237, MULT_mult_6_n2236,
         MULT_mult_6_n2235, MULT_mult_6_n2234, MULT_mult_6_n2233,
         MULT_mult_6_n2232, MULT_mult_6_n2231, MULT_mult_6_n2230,
         MULT_mult_6_n2229, MULT_mult_6_n2228, MULT_mult_6_n2227,
         MULT_mult_6_n2226, MULT_mult_6_n2225, MULT_mult_6_n2224,
         MULT_mult_6_n2223, MULT_mult_6_n2222, MULT_mult_6_n2221,
         MULT_mult_6_n2220, MULT_mult_6_n2219, MULT_mult_6_n2218,
         MULT_mult_6_n2217, MULT_mult_6_n2216, MULT_mult_6_n2215,
         MULT_mult_6_n2214, MULT_mult_6_n2213, MULT_mult_6_n2212,
         MULT_mult_6_n2211, MULT_mult_6_n2210, MULT_mult_6_n2209,
         MULT_mult_6_n2208, MULT_mult_6_n2207, MULT_mult_6_n2206,
         MULT_mult_6_n2205, MULT_mult_6_n2204, MULT_mult_6_n2203,
         MULT_mult_6_n2202, MULT_mult_6_n2201, MULT_mult_6_n2200,
         MULT_mult_6_n2199, MULT_mult_6_n2198, MULT_mult_6_n2197,
         MULT_mult_6_n2196, MULT_mult_6_n2195, MULT_mult_6_n2194,
         MULT_mult_6_n2193, MULT_mult_6_n2192, MULT_mult_6_n2191,
         MULT_mult_6_n2190, MULT_mult_6_n2189, MULT_mult_6_n2188,
         MULT_mult_6_n2187, MULT_mult_6_n2186, MULT_mult_6_n2185,
         MULT_mult_6_n2184, MULT_mult_6_n2183, MULT_mult_6_n2182,
         MULT_mult_6_n2181, MULT_mult_6_n2180, MULT_mult_6_n2179,
         MULT_mult_6_n2178, MULT_mult_6_n2177, MULT_mult_6_n2176,
         MULT_mult_6_n2175, MULT_mult_6_n2174, MULT_mult_6_n2173,
         MULT_mult_6_n2172, MULT_mult_6_n2171, MULT_mult_6_n2170,
         MULT_mult_6_n2169, MULT_mult_6_n2168, MULT_mult_6_n2167,
         MULT_mult_6_n2166, MULT_mult_6_n2165, MULT_mult_6_n2164,
         MULT_mult_6_n2163, MULT_mult_6_n2162, MULT_mult_6_n2161,
         MULT_mult_6_n2160, MULT_mult_6_n2159, MULT_mult_6_n2158,
         MULT_mult_6_n2157, MULT_mult_6_n2156, MULT_mult_6_n2155,
         MULT_mult_6_n2154, MULT_mult_6_n2153, MULT_mult_6_n2152,
         MULT_mult_6_n2151, MULT_mult_6_n2150, MULT_mult_6_n2149,
         MULT_mult_6_n2148, MULT_mult_6_n2147, MULT_mult_6_n2146,
         MULT_mult_6_n2145, MULT_mult_6_n2144, MULT_mult_6_n2143,
         MULT_mult_6_n2142, MULT_mult_6_n2141, MULT_mult_6_n2140,
         MULT_mult_6_n2139, MULT_mult_6_n2138, MULT_mult_6_n2137,
         MULT_mult_6_n2136, MULT_mult_6_n2135, MULT_mult_6_n2134,
         MULT_mult_6_n2133, MULT_mult_6_n2132, MULT_mult_6_n2131,
         MULT_mult_6_n2130, MULT_mult_6_n2129, MULT_mult_6_n2128,
         MULT_mult_6_n2127, MULT_mult_6_n2126, MULT_mult_6_n2125,
         MULT_mult_6_n2124, MULT_mult_6_n2123, MULT_mult_6_n2122,
         MULT_mult_6_n2121, MULT_mult_6_n2120, MULT_mult_6_n2119,
         MULT_mult_6_n2118, MULT_mult_6_n2117, MULT_mult_6_n2116,
         MULT_mult_6_n2115, MULT_mult_6_n2114, MULT_mult_6_n2113,
         MULT_mult_6_n2112, MULT_mult_6_n2111, MULT_mult_6_n2110,
         MULT_mult_6_n2109, MULT_mult_6_n2108, MULT_mult_6_n2107,
         MULT_mult_6_n2106, MULT_mult_6_n2105, MULT_mult_6_n2104,
         MULT_mult_6_n2103, MULT_mult_6_n2102, MULT_mult_6_n2101,
         MULT_mult_6_n2100, MULT_mult_6_n2099, MULT_mult_6_n2098,
         MULT_mult_6_n2097, MULT_mult_6_n2096, MULT_mult_6_n2095,
         MULT_mult_6_n2094, MULT_mult_6_n2093, MULT_mult_6_n2092,
         MULT_mult_6_n2091, MULT_mult_6_n2090, MULT_mult_6_n2089,
         MULT_mult_6_n2088, MULT_mult_6_n2087, MULT_mult_6_n2086,
         MULT_mult_6_n2085, MULT_mult_6_n2084, MULT_mult_6_n2083,
         MULT_mult_6_n2082, MULT_mult_6_n2081, MULT_mult_6_n2080,
         MULT_mult_6_n2079, MULT_mult_6_n2078, MULT_mult_6_n2077,
         MULT_mult_6_n2076, MULT_mult_6_n2075, MULT_mult_6_n2074,
         MULT_mult_6_n2073, MULT_mult_6_n2072, MULT_mult_6_n2071,
         MULT_mult_6_n2070, MULT_mult_6_n2069, MULT_mult_6_n2068,
         MULT_mult_6_n2067, MULT_mult_6_n2066, MULT_mult_6_n2065,
         MULT_mult_6_n2064, MULT_mult_6_n2063, MULT_mult_6_n2062,
         MULT_mult_6_n2061, MULT_mult_6_n2060, MULT_mult_6_n2059,
         MULT_mult_6_n2058, MULT_mult_6_n2057, MULT_mult_6_n2056,
         MULT_mult_6_n2055, MULT_mult_6_n2054, MULT_mult_6_n2053,
         MULT_mult_6_n2052, MULT_mult_6_n2051, MULT_mult_6_n2050,
         MULT_mult_6_n2049, MULT_mult_6_n2048, MULT_mult_6_n2047,
         MULT_mult_6_n2046, MULT_mult_6_n2045, MULT_mult_6_n2044,
         MULT_mult_6_n2043, MULT_mult_6_n2042, MULT_mult_6_n2041,
         MULT_mult_6_n2040, MULT_mult_6_n2039, MULT_mult_6_n2038,
         MULT_mult_6_n2037, MULT_mult_6_n2036, MULT_mult_6_n2035,
         MULT_mult_6_n2034, MULT_mult_6_n2033, MULT_mult_6_n2032,
         MULT_mult_6_n2031, MULT_mult_6_n2030, MULT_mult_6_n2029,
         MULT_mult_6_n2028, MULT_mult_6_n2027, MULT_mult_6_n2026,
         MULT_mult_6_n2025, MULT_mult_6_n2024, MULT_mult_6_n2023,
         MULT_mult_6_n2022, MULT_mult_6_n2021, MULT_mult_6_n2020,
         MULT_mult_6_n2019, MULT_mult_6_n2018, MULT_mult_6_n2017,
         MULT_mult_6_n2016, MULT_mult_6_n2015, MULT_mult_6_n2014,
         MULT_mult_6_n2013, MULT_mult_6_n2012, MULT_mult_6_n2011,
         MULT_mult_6_n2010, MULT_mult_6_n2009, MULT_mult_6_n2008,
         MULT_mult_6_n2007, MULT_mult_6_n2006, MULT_mult_6_n2005,
         MULT_mult_6_n2004, MULT_mult_6_n2003, MULT_mult_6_n2002,
         MULT_mult_6_n2001, MULT_mult_6_n2000, MULT_mult_6_n1999,
         MULT_mult_6_n1998, MULT_mult_6_n1997, MULT_mult_6_n1996,
         MULT_mult_6_n1995, MULT_mult_6_n1994, MULT_mult_6_n1993,
         MULT_mult_6_n1992, MULT_mult_6_n1991, MULT_mult_6_n1990,
         MULT_mult_6_n1989, MULT_mult_6_n1988, MULT_mult_6_n1987,
         MULT_mult_6_n1986, MULT_mult_6_n1985, MULT_mult_6_n1984,
         MULT_mult_6_n1983, MULT_mult_6_n1982, MULT_mult_6_n1981,
         MULT_mult_6_n1980, MULT_mult_6_n1979, MULT_mult_6_n1978,
         MULT_mult_6_n1977, MULT_mult_6_n1976, MULT_mult_6_n1975,
         MULT_mult_6_n1974, MULT_mult_6_n1973, MULT_mult_6_n1972,
         MULT_mult_6_n1971, MULT_mult_6_n1970, MULT_mult_6_n1969,
         MULT_mult_6_n1968, MULT_mult_6_n1967, MULT_mult_6_n1966,
         MULT_mult_6_n1965, MULT_mult_6_n1964, MULT_mult_6_n1963,
         MULT_mult_6_n1962, MULT_mult_6_n1961, MULT_mult_6_n1960,
         MULT_mult_6_n1959, MULT_mult_6_n1958, MULT_mult_6_n1957,
         MULT_mult_6_n1956, MULT_mult_6_n1955, MULT_mult_6_n1954,
         MULT_mult_6_n1953, MULT_mult_6_n1952, MULT_mult_6_n1951,
         MULT_mult_6_n1950, MULT_mult_6_n1949, MULT_mult_6_n1948,
         MULT_mult_6_n1947, MULT_mult_6_n1946, MULT_mult_6_n1945,
         MULT_mult_6_n1944, MULT_mult_6_n1943, MULT_mult_6_n1942,
         MULT_mult_6_n1941, MULT_mult_6_n1940, MULT_mult_6_n1939,
         MULT_mult_6_n1938, MULT_mult_6_n1937, MULT_mult_6_n1936,
         MULT_mult_6_n1935, MULT_mult_6_n1934, MULT_mult_6_n1933,
         MULT_mult_6_n1932, MULT_mult_6_n1931, MULT_mult_6_n1930,
         MULT_mult_6_n1929, MULT_mult_6_n1928, MULT_mult_6_n1927,
         MULT_mult_6_n1926, MULT_mult_6_n1925, MULT_mult_6_n1924,
         MULT_mult_6_n1923, MULT_mult_6_n1922, MULT_mult_6_n1921,
         MULT_mult_6_n1920, MULT_mult_6_n1919, MULT_mult_6_n1918,
         MULT_mult_6_n1917, MULT_mult_6_n1916, MULT_mult_6_n1915,
         MULT_mult_6_n1914, MULT_mult_6_n1913, MULT_mult_6_n1912,
         MULT_mult_6_n1911, MULT_mult_6_n1910, MULT_mult_6_n1909,
         MULT_mult_6_n1908, MULT_mult_6_n1907, MULT_mult_6_n1906,
         MULT_mult_6_n1905, MULT_mult_6_n1904, MULT_mult_6_n1903,
         MULT_mult_6_n1902, MULT_mult_6_n1901, MULT_mult_6_n1900,
         MULT_mult_6_n1899, MULT_mult_6_n1898, MULT_mult_6_n1897,
         MULT_mult_6_n1896, MULT_mult_6_n1895, MULT_mult_6_n1894,
         MULT_mult_6_n1893, MULT_mult_6_n1892, MULT_mult_6_n1891,
         MULT_mult_6_n1890, MULT_mult_6_n1889, MULT_mult_6_n1888,
         MULT_mult_6_n1887, MULT_mult_6_n1886, MULT_mult_6_n1885,
         MULT_mult_6_n1884, MULT_mult_6_n1883, MULT_mult_6_n1882,
         MULT_mult_6_n1881, MULT_mult_6_n1880, MULT_mult_6_n1879,
         MULT_mult_6_n1878, MULT_mult_6_n1877, MULT_mult_6_n1876,
         MULT_mult_6_n1875, MULT_mult_6_n1874, MULT_mult_6_n1873,
         MULT_mult_6_n1872, MULT_mult_6_n1871, MULT_mult_6_n1870,
         MULT_mult_6_n1869, MULT_mult_6_n1868, MULT_mult_6_n1867,
         MULT_mult_6_n1866, MULT_mult_6_n1865, MULT_mult_6_n1864,
         MULT_mult_6_n1863, MULT_mult_6_n1862, MULT_mult_6_n1861,
         MULT_mult_6_n1860, MULT_mult_6_n1859, MULT_mult_6_n1858,
         MULT_mult_6_n1857, MULT_mult_6_n1856, MULT_mult_6_n1855,
         MULT_mult_6_n1854, MULT_mult_6_n1853, MULT_mult_6_n1852,
         MULT_mult_6_n1851, MULT_mult_6_n1850, MULT_mult_6_n1849,
         MULT_mult_6_n1848, MULT_mult_6_n1847, MULT_mult_6_n1846,
         MULT_mult_6_n1845, MULT_mult_6_n1844, MULT_mult_6_n1843,
         MULT_mult_6_n1842, MULT_mult_6_n1841, MULT_mult_6_n1840,
         MULT_mult_6_n1839, MULT_mult_6_n1838, MULT_mult_6_n1837,
         MULT_mult_6_n1836, MULT_mult_6_n1835, MULT_mult_6_n1834,
         MULT_mult_6_n1833, MULT_mult_6_n1832, MULT_mult_6_n1831,
         MULT_mult_6_n1830, MULT_mult_6_n1829, MULT_mult_6_n1828,
         MULT_mult_6_n1827, MULT_mult_6_n1826, MULT_mult_6_n1825,
         MULT_mult_6_n1824, MULT_mult_6_n1823, MULT_mult_6_n1822,
         MULT_mult_6_n1821, MULT_mult_6_n1820, MULT_mult_6_n1819,
         MULT_mult_6_n1818, MULT_mult_6_n1817, MULT_mult_6_n1816,
         MULT_mult_6_n1815, MULT_mult_6_n1814, MULT_mult_6_n1813,
         MULT_mult_6_n1812, MULT_mult_6_n1811, MULT_mult_6_n1810,
         MULT_mult_6_n1809, MULT_mult_6_n1808, MULT_mult_6_n1807,
         MULT_mult_6_n1806, MULT_mult_6_n1805, MULT_mult_6_n1804,
         MULT_mult_6_n1803, MULT_mult_6_n1802, MULT_mult_6_n1801,
         MULT_mult_6_n1800, MULT_mult_6_n1799, MULT_mult_6_n1798,
         MULT_mult_6_n1797, MULT_mult_6_n1796, MULT_mult_6_n1795,
         MULT_mult_6_n1794, MULT_mult_6_n1793, MULT_mult_6_n1792,
         MULT_mult_6_n1791, MULT_mult_6_n1790, MULT_mult_6_n1789,
         MULT_mult_6_n1788, MULT_mult_6_n1787, MULT_mult_6_n1786,
         MULT_mult_6_n1785, MULT_mult_6_n1784, MULT_mult_6_n1783,
         MULT_mult_6_n1782, MULT_mult_6_n1781, MULT_mult_6_n1780,
         MULT_mult_6_n1779, MULT_mult_6_n1778, MULT_mult_6_n1777,
         MULT_mult_6_n1776, MULT_mult_6_n1775, MULT_mult_6_n1774,
         MULT_mult_6_n1773, MULT_mult_6_n1772, MULT_mult_6_n1771,
         MULT_mult_6_n1770, MULT_mult_6_n1769, MULT_mult_6_n1768,
         MULT_mult_6_n1767, MULT_mult_6_n1766, MULT_mult_6_n1765,
         MULT_mult_6_n1764, MULT_mult_6_n1763, MULT_mult_6_n1762,
         MULT_mult_6_n1761, MULT_mult_6_n1760, MULT_mult_6_n1759,
         MULT_mult_6_n1758, MULT_mult_6_n1757, MULT_mult_6_n1756,
         MULT_mult_6_n1755, MULT_mult_6_n1754, MULT_mult_6_n1753,
         MULT_mult_6_n1752, MULT_mult_6_n1751, MULT_mult_6_n1750,
         MULT_mult_6_n1749, MULT_mult_6_n1748, MULT_mult_6_n1747,
         MULT_mult_6_n1746, MULT_mult_6_n1745, MULT_mult_6_n1744,
         MULT_mult_6_n1743, MULT_mult_6_n1742, MULT_mult_6_n1741,
         MULT_mult_6_n1740, MULT_mult_6_n1739, MULT_mult_6_n1738,
         MULT_mult_6_n1737, MULT_mult_6_n1736, MULT_mult_6_n1735,
         MULT_mult_6_n1734, MULT_mult_6_n1733, MULT_mult_6_n1732,
         MULT_mult_6_n1731, MULT_mult_6_n1730, MULT_mult_6_n1729,
         MULT_mult_6_n1728, MULT_mult_6_n1727, MULT_mult_6_n1726,
         MULT_mult_6_n1725, MULT_mult_6_n1724, MULT_mult_6_n1723,
         MULT_mult_6_n1722, MULT_mult_6_n1721, MULT_mult_6_n1720,
         MULT_mult_6_n1719, MULT_mult_6_n1718, MULT_mult_6_n1717,
         MULT_mult_6_n1716, MULT_mult_6_n1715, MULT_mult_6_n1714,
         MULT_mult_6_n1713, MULT_mult_6_n1712, MULT_mult_6_n1711,
         MULT_mult_6_n1710, MULT_mult_6_n1709, MULT_mult_6_n1708,
         MULT_mult_6_n1707, MULT_mult_6_n1706, MULT_mult_6_n1705,
         MULT_mult_6_n1704, MULT_mult_6_n1703, MULT_mult_6_n1702,
         MULT_mult_6_n1701, MULT_mult_6_n1700, MULT_mult_6_n1699,
         MULT_mult_6_n1698, MULT_mult_6_n1697, MULT_mult_6_n1696,
         MULT_mult_6_n1695, MULT_mult_6_n1694, MULT_mult_6_n1693,
         MULT_mult_6_n1692, MULT_mult_6_n1691, MULT_mult_6_n1690,
         MULT_mult_6_n1689, MULT_mult_6_n1688, MULT_mult_6_n1687,
         MULT_mult_6_n1686, MULT_mult_6_n1685, MULT_mult_6_n1684,
         MULT_mult_6_n1683, MULT_mult_6_n1682, MULT_mult_6_n1681,
         MULT_mult_6_n1680, MULT_mult_6_n1679, MULT_mult_6_n1678,
         MULT_mult_6_n1677, MULT_mult_6_n1676, MULT_mult_6_n1675,
         MULT_mult_6_n1674, MULT_mult_6_n1673, MULT_mult_6_n1672,
         MULT_mult_6_n1671, MULT_mult_6_n1670, MULT_mult_6_n1669,
         MULT_mult_6_n1668, MULT_mult_6_n1667, MULT_mult_6_n1666,
         MULT_mult_6_n1665, MULT_mult_6_n1664, MULT_mult_6_n1663,
         MULT_mult_6_n1662, MULT_mult_6_n1661, MULT_mult_6_n1660,
         MULT_mult_6_n1659, MULT_mult_6_n1658, MULT_mult_6_n1657,
         MULT_mult_6_n1656, MULT_mult_6_n1655, MULT_mult_6_n1654,
         MULT_mult_6_n1653, MULT_mult_6_n1652, MULT_mult_6_n1651,
         MULT_mult_6_n1650, MULT_mult_6_n1649, MULT_mult_6_n1648,
         MULT_mult_6_n1647, MULT_mult_6_n1646, MULT_mult_6_n1645,
         MULT_mult_6_n1644, MULT_mult_6_n1643, MULT_mult_6_n1642,
         MULT_mult_6_n1641, MULT_mult_6_n1640, MULT_mult_6_n1639,
         MULT_mult_6_n1638, MULT_mult_6_n1637, MULT_mult_6_n1636,
         MULT_mult_6_n1635, MULT_mult_6_n1634, MULT_mult_6_n1633,
         MULT_mult_6_n1632, MULT_mult_6_n1631, MULT_mult_6_n1630,
         MULT_mult_6_n1629, MULT_mult_6_n1628, MULT_mult_6_n1627,
         MULT_mult_6_n1626, MULT_mult_6_n1625, MULT_mult_6_n1624,
         MULT_mult_6_n1623, MULT_mult_6_n1622, MULT_mult_6_n1621,
         MULT_mult_6_n1620, MULT_mult_6_n1619, MULT_mult_6_n1618,
         MULT_mult_6_n1617, MULT_mult_6_n1616, MULT_mult_6_n1615,
         MULT_mult_6_n1614, MULT_mult_6_n1613, MULT_mult_6_n1612,
         MULT_mult_6_n1611, MULT_mult_6_n1610, MULT_mult_6_n1609,
         MULT_mult_6_n1608, MULT_mult_6_n1607, MULT_mult_6_n1606,
         MULT_mult_6_n1605, MULT_mult_6_n1604, MULT_mult_6_n1603,
         MULT_mult_6_n1602, MULT_mult_6_n1601, MULT_mult_6_n1600,
         MULT_mult_6_n1599, MULT_mult_6_n1598, MULT_mult_6_n1597,
         MULT_mult_6_n1596, MULT_mult_6_n1595, MULT_mult_6_n1594,
         MULT_mult_6_n1593, MULT_mult_6_n1592, MULT_mult_6_n1591,
         MULT_mult_6_n1590, MULT_mult_6_n1589, MULT_mult_6_n1588,
         MULT_mult_6_n1587, MULT_mult_6_n1586, MULT_mult_6_n1585,
         MULT_mult_6_n1584, MULT_mult_6_n1583, MULT_mult_6_n1582,
         MULT_mult_6_n1581, MULT_mult_6_n1580, MULT_mult_6_n1579,
         MULT_mult_6_n1578, MULT_mult_6_n1577, MULT_mult_6_n1576,
         MULT_mult_6_n1575, MULT_mult_6_n1574, MULT_mult_6_n1573,
         MULT_mult_6_n1572, MULT_mult_6_n1571, MULT_mult_6_n1570,
         MULT_mult_6_n1569, MULT_mult_6_n1568, MULT_mult_6_n1566,
         MULT_mult_6_n1565, MULT_mult_6_n1564, MULT_mult_6_n1563,
         MULT_mult_6_n1562, MULT_mult_6_n1561, MULT_mult_6_n1560,
         MULT_mult_6_n1559, MULT_mult_6_n1558, MULT_mult_6_n1557,
         MULT_mult_6_n1556, MULT_mult_6_n1555, MULT_mult_6_n1554,
         MULT_mult_6_n1553, MULT_mult_6_n1552, MULT_mult_6_n1551,
         MULT_mult_6_n1550, MULT_mult_6_n1549, MULT_mult_6_n1548,
         MULT_mult_6_n1547, MULT_mult_6_n1546, MULT_mult_6_n1545,
         MULT_mult_6_n1544, MULT_mult_6_n1543, MULT_mult_6_n1542,
         MULT_mult_6_n1541, MULT_mult_6_n1540, MULT_mult_6_n1539,
         MULT_mult_6_n1538, MULT_mult_6_n1537, MULT_mult_6_n1536,
         MULT_mult_6_n1535, MULT_mult_6_n1534, MULT_mult_6_n1533,
         MULT_mult_6_n1532, MULT_mult_6_n1531, MULT_mult_6_n1530,
         MULT_mult_6_n1529, MULT_mult_6_n1528, MULT_mult_6_n1527,
         MULT_mult_6_n1526, MULT_mult_6_n1525, MULT_mult_6_n1524,
         MULT_mult_6_n1523, MULT_mult_6_n1522, MULT_mult_6_n1521,
         MULT_mult_6_n1520, MULT_mult_6_n1519, MULT_mult_6_n1518,
         MULT_mult_6_n1517, MULT_mult_6_n1516, MULT_mult_6_n1515,
         MULT_mult_6_n1514, MULT_mult_6_n1513, MULT_mult_6_n1512,
         MULT_mult_6_n1511, MULT_mult_6_n1510, MULT_mult_6_n1509,
         MULT_mult_6_n1508, MULT_mult_6_n1507, MULT_mult_6_n1506,
         MULT_mult_6_n1505, MULT_mult_6_n1504, MULT_mult_6_n1503,
         MULT_mult_6_n1502, MULT_mult_6_n1501, MULT_mult_6_n1500,
         MULT_mult_6_n1499, MULT_mult_6_n1498, MULT_mult_6_n1497,
         MULT_mult_6_n1496, MULT_mult_6_n1495, MULT_mult_6_n1494,
         MULT_mult_6_n1493, MULT_mult_6_n1492, MULT_mult_6_n1491,
         MULT_mult_6_n1490, MULT_mult_6_n1489, MULT_mult_6_n1488,
         MULT_mult_6_n1487, MULT_mult_6_n1486, MULT_mult_6_n1485,
         MULT_mult_6_n1484, MULT_mult_6_n1483, MULT_mult_6_n1482,
         MULT_mult_6_n1481, MULT_mult_6_n1480, MULT_mult_6_n1479,
         MULT_mult_6_n1478, MULT_mult_6_n1477, MULT_mult_6_n1476,
         MULT_mult_6_n1475, MULT_mult_6_n1474, MULT_mult_6_n1473,
         MULT_mult_6_n1472, MULT_mult_6_n1471, MULT_mult_6_n1470,
         MULT_mult_6_n1469, MULT_mult_6_n1468, MULT_mult_6_n1467,
         MULT_mult_6_n1466, MULT_mult_6_n1465, MULT_mult_6_n1464,
         MULT_mult_6_n1463, MULT_mult_6_n1462, MULT_mult_6_n1461,
         MULT_mult_6_n1460, MULT_mult_6_n1459, MULT_mult_6_n1458,
         MULT_mult_6_n1457, MULT_mult_6_n1456, MULT_mult_6_n1455,
         MULT_mult_6_n1454, MULT_mult_6_n1453, MULT_mult_6_n1452,
         MULT_mult_6_n1451, MULT_mult_6_n1450, MULT_mult_6_n1449,
         MULT_mult_6_n1448, MULT_mult_6_n1447, MULT_mult_6_n1446,
         MULT_mult_6_n1445, MULT_mult_6_n1444, MULT_mult_6_n1443,
         MULT_mult_6_n1442, MULT_mult_6_n1441, MULT_mult_6_n1440,
         MULT_mult_6_n1439, MULT_mult_6_n1438, MULT_mult_6_n1437,
         MULT_mult_6_n1436, MULT_mult_6_n1435, MULT_mult_6_n1434,
         MULT_mult_6_n1433, MULT_mult_6_n1432, MULT_mult_6_n1431,
         MULT_mult_6_n1430, MULT_mult_6_n1429, MULT_mult_6_n1428,
         MULT_mult_6_n1427, MULT_mult_6_n1426, MULT_mult_6_n1425,
         MULT_mult_6_n1424, MULT_mult_6_n1423, MULT_mult_6_n1422,
         MULT_mult_6_n1421, MULT_mult_6_n1420, MULT_mult_6_n1419,
         MULT_mult_6_n1418, MULT_mult_6_n1417, MULT_mult_6_n1416,
         MULT_mult_6_n1415, MULT_mult_6_n1414, MULT_mult_6_n1413,
         MULT_mult_6_n1412, MULT_mult_6_n1411, MULT_mult_6_n1410,
         MULT_mult_6_n1409, MULT_mult_6_n1408, MULT_mult_6_n1407,
         MULT_mult_6_n1406, MULT_mult_6_n1405, MULT_mult_6_n1404,
         MULT_mult_6_n1403, MULT_mult_6_n1402, MULT_mult_6_n1401,
         MULT_mult_6_n1400, MULT_mult_6_n1399, MULT_mult_6_n1398,
         MULT_mult_6_n1397, MULT_mult_6_n1396, MULT_mult_6_n1395,
         MULT_mult_6_n1394, MULT_mult_6_n1393, MULT_mult_6_n1392,
         MULT_mult_6_n1391, MULT_mult_6_n1390, MULT_mult_6_n1389,
         MULT_mult_6_n1388, MULT_mult_6_n1387, MULT_mult_6_n1386,
         MULT_mult_6_n1385, MULT_mult_6_n1384, MULT_mult_6_n1383,
         MULT_mult_6_n1382, MULT_mult_6_n1381, MULT_mult_6_n1380,
         MULT_mult_6_n1379, MULT_mult_6_n1378, MULT_mult_6_n1377,
         MULT_mult_6_n1376, MULT_mult_6_n1375, MULT_mult_6_n1374,
         MULT_mult_6_n1373, MULT_mult_6_n1372, MULT_mult_6_n1371,
         MULT_mult_6_n1370, MULT_mult_6_n1369, MULT_mult_6_n1368,
         MULT_mult_6_n1367, MULT_mult_6_n1366, MULT_mult_6_n1365,
         MULT_mult_6_n1364, MULT_mult_6_n1363, MULT_mult_6_n1362,
         MULT_mult_6_n1361, MULT_mult_6_n1360, MULT_mult_6_n1359,
         MULT_mult_6_n1358, MULT_mult_6_n1357, MULT_mult_6_n1356,
         MULT_mult_6_n1355, MULT_mult_6_n1354, MULT_mult_6_n1353,
         MULT_mult_6_n1352, MULT_mult_6_n1351, MULT_mult_6_n1350,
         MULT_mult_6_n1349, MULT_mult_6_n1348, MULT_mult_6_n1347,
         MULT_mult_6_n1346, MULT_mult_6_n1345, MULT_mult_6_n1344,
         MULT_mult_6_n1343, MULT_mult_6_n1342, MULT_mult_6_n1341,
         MULT_mult_6_n1340, MULT_mult_6_n1339, MULT_mult_6_n1338,
         MULT_mult_6_n1337, MULT_mult_6_n1336, MULT_mult_6_n1335,
         MULT_mult_6_n1334, MULT_mult_6_n1333, MULT_mult_6_n1332,
         MULT_mult_6_n1331, MULT_mult_6_n1330, MULT_mult_6_n1329,
         MULT_mult_6_n1328, MULT_mult_6_n1327, MULT_mult_6_n1326,
         MULT_mult_6_n1325, MULT_mult_6_n1324, MULT_mult_6_n1323,
         MULT_mult_6_n1322, MULT_mult_6_n1321, MULT_mult_6_n1320,
         MULT_mult_6_n1319, MULT_mult_6_n1318, MULT_mult_6_n1317,
         MULT_mult_6_n1316, MULT_mult_6_n1315, MULT_mult_6_n1314,
         MULT_mult_6_n1313, MULT_mult_6_n1312, MULT_mult_6_n1311,
         MULT_mult_6_n1310, MULT_mult_6_n1309, MULT_mult_6_n1308,
         MULT_mult_6_n1307, MULT_mult_6_n1306, MULT_mult_6_n1305,
         MULT_mult_6_n1304, MULT_mult_6_n1303, MULT_mult_6_n1302,
         MULT_mult_6_n1301, MULT_mult_6_n1300, MULT_mult_6_n1299,
         MULT_mult_6_n1298, MULT_mult_6_n1297, MULT_mult_6_n1296,
         MULT_mult_6_n1295, MULT_mult_6_n1294, MULT_mult_6_n1293,
         MULT_mult_6_n1292, MULT_mult_6_n1291, MULT_mult_6_n1290,
         MULT_mult_6_n1289, MULT_mult_6_n1288, MULT_mult_6_n1287,
         MULT_mult_6_n1286, MULT_mult_6_n1285, MULT_mult_6_n1284,
         MULT_mult_6_n1283, MULT_mult_6_n1282, MULT_mult_6_n1281,
         MULT_mult_6_n1280, MULT_mult_6_n1279, MULT_mult_6_n1278,
         MULT_mult_6_n1277, MULT_mult_6_n1276, MULT_mult_6_n1275,
         MULT_mult_6_n1274, MULT_mult_6_n1273, MULT_mult_6_n1272,
         MULT_mult_6_n1271, MULT_mult_6_n1270, MULT_mult_6_n1269,
         MULT_mult_6_n1268, MULT_mult_6_n1267, MULT_mult_6_n1266,
         MULT_mult_6_n1265, MULT_mult_6_n1264, MULT_mult_6_n1263,
         MULT_mult_6_n1262, MULT_mult_6_n1261, MULT_mult_6_n1260,
         MULT_mult_6_n1259, MULT_mult_6_n1258, MULT_mult_6_n1257,
         MULT_mult_6_n1256, MULT_mult_6_n1255, MULT_mult_6_n1254,
         MULT_mult_6_n1253, MULT_mult_6_n1252, MULT_mult_6_n1251,
         MULT_mult_6_n1250, MULT_mult_6_n1249, MULT_mult_6_n1248,
         MULT_mult_6_n1247, MULT_mult_6_n1246, MULT_mult_6_n1245,
         MULT_mult_6_n1244, MULT_mult_6_n1243, MULT_mult_6_n1242,
         MULT_mult_6_n1241, MULT_mult_6_n1240, MULT_mult_6_n1239,
         MULT_mult_6_n1238, MULT_mult_6_n1237, MULT_mult_6_n1236,
         MULT_mult_6_n1235, MULT_mult_6_n1234, MULT_mult_6_n1233,
         MULT_mult_6_n1232, MULT_mult_6_n1231, MULT_mult_6_n1230,
         MULT_mult_6_n1229, MULT_mult_6_n1228, MULT_mult_6_n1227,
         MULT_mult_6_n1226, MULT_mult_6_n1225, MULT_mult_6_n1224,
         MULT_mult_6_n1223, MULT_mult_6_n1222, MULT_mult_6_n1221,
         MULT_mult_6_n1220, MULT_mult_6_n1219, MULT_mult_6_n1218,
         MULT_mult_6_n1217, MULT_mult_6_n1216, MULT_mult_6_n1215,
         MULT_mult_6_n1214, MULT_mult_6_n1213, MULT_mult_6_n1212,
         MULT_mult_6_n1211, MULT_mult_6_n1210, MULT_mult_6_n1209,
         MULT_mult_6_n1208, MULT_mult_6_n1207, MULT_mult_6_n1206,
         MULT_mult_6_n1205, MULT_mult_6_n1204, MULT_mult_6_n1203,
         MULT_mult_6_n1202, MULT_mult_6_n1201, MULT_mult_6_n1200,
         MULT_mult_6_n1199, MULT_mult_6_n1198, MULT_mult_6_n1197,
         MULT_mult_6_n1196, MULT_mult_6_n1195, MULT_mult_6_n1194,
         MULT_mult_6_n1193, MULT_mult_6_n1192, MULT_mult_6_n1191,
         MULT_mult_6_n1190, MULT_mult_6_n1189, MULT_mult_6_n1188,
         MULT_mult_6_n1187, MULT_mult_6_n1186, MULT_mult_6_n1185,
         MULT_mult_6_n1184, MULT_mult_6_n1183, MULT_mult_6_n1182,
         MULT_mult_6_n1181, MULT_mult_6_n1180, MULT_mult_6_n1179,
         MULT_mult_6_n1178, MULT_mult_6_n1177, MULT_mult_6_n1176,
         MULT_mult_6_n1175, MULT_mult_6_n1174, MULT_mult_6_n1173,
         MULT_mult_6_n1172, MULT_mult_6_n1171, MULT_mult_6_n1170,
         MULT_mult_6_n1169, MULT_mult_6_n1168, MULT_mult_6_n1167,
         MULT_mult_6_n1166, MULT_mult_6_n1165, MULT_mult_6_n1164,
         MULT_mult_6_n1163, MULT_mult_6_n1162, MULT_mult_6_n1161,
         MULT_mult_6_n1160, MULT_mult_6_n1159, MULT_mult_6_n1158,
         MULT_mult_6_n1157, MULT_mult_6_n1156, MULT_mult_6_n1155,
         MULT_mult_6_n1154, MULT_mult_6_n1153, MULT_mult_6_n1152,
         MULT_mult_6_n1151, MULT_mult_6_n1150, MULT_mult_6_n1149,
         MULT_mult_6_n1148, MULT_mult_6_n1147, MULT_mult_6_n1146,
         MULT_mult_6_n1145, MULT_mult_6_n1144, MULT_mult_6_n1143,
         MULT_mult_6_n1142, MULT_mult_6_n1141, MULT_mult_6_n1140,
         MULT_mult_6_n1139, MULT_mult_6_n1138, MULT_mult_6_n1137,
         MULT_mult_6_n1136, MULT_mult_6_n1135, MULT_mult_6_n1134,
         MULT_mult_6_n1133, MULT_mult_6_n1132, MULT_mult_6_n1131,
         MULT_mult_6_n1130, MULT_mult_6_n1129, MULT_mult_6_n1128,
         MULT_mult_6_n1127, MULT_mult_6_n1126, MULT_mult_6_n1125,
         MULT_mult_6_n1124, MULT_mult_6_n1123, MULT_mult_6_n1122,
         MULT_mult_6_n1121, MULT_mult_6_n1120, MULT_mult_6_n1119,
         MULT_mult_6_n1118, MULT_mult_6_n1117, MULT_mult_6_n1116,
         MULT_mult_6_n1115, MULT_mult_6_n1114, MULT_mult_6_n1113,
         MULT_mult_6_n1112, MULT_mult_6_n1111, MULT_mult_6_n1110,
         MULT_mult_6_n1109, MULT_mult_6_n1108, MULT_mult_6_n1107,
         MULT_mult_6_n1106, MULT_mult_6_n1105, MULT_mult_6_n1104,
         MULT_mult_6_n1103, MULT_mult_6_n1102, MULT_mult_6_n1101,
         MULT_mult_6_n1100, MULT_mult_6_n1099, MULT_mult_6_n1098,
         MULT_mult_6_n1097, MULT_mult_6_n1096, MULT_mult_6_n1095,
         MULT_mult_6_n1094, MULT_mult_6_n1093, MULT_mult_6_n1092,
         MULT_mult_6_n1091, MULT_mult_6_n1090, MULT_mult_6_n1089,
         MULT_mult_6_n1088, MULT_mult_6_n1087, MULT_mult_6_n1086,
         MULT_mult_6_n1085, MULT_mult_6_n1084, MULT_mult_6_n1083,
         MULT_mult_6_n1082, MULT_mult_6_n1081, MULT_mult_6_n1080,
         MULT_mult_6_n1079, MULT_mult_6_n1078, MULT_mult_6_n1077,
         MULT_mult_6_n1074, MULT_mult_6_n1073, MULT_mult_6_n1072,
         MULT_mult_6_n1071, MULT_mult_6_n1070, MULT_mult_6_n1069,
         MULT_mult_6_n1068, MULT_mult_6_n1067, MULT_mult_6_n1066,
         MULT_mult_6_n1065, MULT_mult_6_n1064, MULT_mult_6_n1063,
         MULT_mult_6_n1062, MULT_mult_6_n1061, MULT_mult_6_n1060,
         MULT_mult_6_n1059, MULT_mult_6_n1058, MULT_mult_6_n1057,
         MULT_mult_6_n1056, MULT_mult_6_n1055, MULT_mult_6_n1054,
         MULT_mult_6_n1053, MULT_mult_6_n1052, MULT_mult_6_n1051,
         MULT_mult_6_n1050, MULT_mult_6_n1049, MULT_mult_6_n1048,
         MULT_mult_6_n1047, MULT_mult_6_n1046, MULT_mult_6_n1045,
         MULT_mult_6_n1044, MULT_mult_6_n1043, MULT_mult_6_n1042,
         MULT_mult_6_n1041, MULT_mult_6_n1040, MULT_mult_6_n1039,
         MULT_mult_6_n1038, MULT_mult_6_n1037, MULT_mult_6_n1036,
         MULT_mult_6_n1035, MULT_mult_6_n1034, MULT_mult_6_n1033,
         MULT_mult_6_n1032, MULT_mult_6_n1031, MULT_mult_6_n1030,
         MULT_mult_6_n1029, MULT_mult_6_n1028, MULT_mult_6_n1027,
         MULT_mult_6_n1025, MULT_mult_6_n1024, MULT_mult_6_n1023,
         MULT_mult_6_n1022, MULT_mult_6_n1021, MULT_mult_6_n1020,
         MULT_mult_6_n1019, MULT_mult_6_n1018, MULT_mult_6_n1017,
         MULT_mult_6_n1016, MULT_mult_6_n1015, MULT_mult_6_n1014,
         MULT_mult_6_n1013, MULT_mult_6_n1012, MULT_mult_6_n1011,
         MULT_mult_6_n1010, MULT_mult_6_n1009, MULT_mult_6_n1008,
         MULT_mult_6_n1007, MULT_mult_6_n1006, MULT_mult_6_n1005,
         MULT_mult_6_n1004, MULT_mult_6_n1003, MULT_mult_6_n1002,
         MULT_mult_6_n1001, MULT_mult_6_n1000, MULT_mult_6_n999,
         MULT_mult_6_n998, MULT_mult_6_n997, MULT_mult_6_n996,
         MULT_mult_6_n995, MULT_mult_6_n994, MULT_mult_6_n993,
         MULT_mult_6_n992, MULT_mult_6_n991, MULT_mult_6_n990,
         MULT_mult_6_n989, MULT_mult_6_n988, MULT_mult_6_n987,
         MULT_mult_6_n986, MULT_mult_6_n985, MULT_mult_6_n984,
         MULT_mult_6_n983, MULT_mult_6_n982, MULT_mult_6_n981,
         MULT_mult_6_n980, MULT_mult_6_n979, MULT_mult_6_n978,
         MULT_mult_6_n977, MULT_mult_6_n976, MULT_mult_6_n975,
         MULT_mult_6_n974, MULT_mult_6_n973, MULT_mult_6_n972,
         MULT_mult_6_n971, MULT_mult_6_n970, MULT_mult_6_n969,
         MULT_mult_6_n968, MULT_mult_6_n967, MULT_mult_6_n966,
         MULT_mult_6_n965, MULT_mult_6_n964, MULT_mult_6_n963,
         MULT_mult_6_n962, MULT_mult_6_n961, MULT_mult_6_n960,
         MULT_mult_6_n959, MULT_mult_6_n958, MULT_mult_6_n957,
         MULT_mult_6_n956, MULT_mult_6_n955, MULT_mult_6_n954,
         MULT_mult_6_n953, MULT_mult_6_n952, MULT_mult_6_n951,
         MULT_mult_6_n950, MULT_mult_6_n949, MULT_mult_6_n948,
         MULT_mult_6_n947, MULT_mult_6_n946, MULT_mult_6_n945,
         MULT_mult_6_n944, MULT_mult_6_n943, MULT_mult_6_n942,
         MULT_mult_6_n941, MULT_mult_6_n940, MULT_mult_6_n939,
         MULT_mult_6_n938, MULT_mult_6_n937, MULT_mult_6_n936,
         MULT_mult_6_n935, MULT_mult_6_n934, MULT_mult_6_n933,
         MULT_mult_6_n932, MULT_mult_6_n931, MULT_mult_6_n930,
         MULT_mult_6_n929, MULT_mult_6_n928, MULT_mult_6_n927,
         MULT_mult_6_n926, MULT_mult_6_n925, MULT_mult_6_n924,
         MULT_mult_6_n923, MULT_mult_6_n922, MULT_mult_6_n921,
         MULT_mult_6_n920, MULT_mult_6_n919, MULT_mult_6_n918,
         MULT_mult_6_n917, MULT_mult_6_n916, MULT_mult_6_n915,
         MULT_mult_6_n914, MULT_mult_6_n913, MULT_mult_6_n912,
         MULT_mult_6_n911, MULT_mult_6_n910, MULT_mult_6_n909,
         MULT_mult_6_n908, MULT_mult_6_n907, MULT_mult_6_n906,
         MULT_mult_6_n905, MULT_mult_6_n904, MULT_mult_6_n903,
         MULT_mult_6_n902, MULT_mult_6_n901, MULT_mult_6_n900,
         MULT_mult_6_n899, MULT_mult_6_n898, MULT_mult_6_n897,
         MULT_mult_6_n896, MULT_mult_6_n895, MULT_mult_6_n894,
         MULT_mult_6_n893, MULT_mult_6_n892, MULT_mult_6_n891,
         MULT_mult_6_n890, MULT_mult_6_n889, MULT_mult_6_n888,
         MULT_mult_6_n887, MULT_mult_6_n886, MULT_mult_6_n885,
         MULT_mult_6_n884, MULT_mult_6_n883, MULT_mult_6_n882,
         MULT_mult_6_n881, MULT_mult_6_n880, MULT_mult_6_n879,
         MULT_mult_6_n878, MULT_mult_6_n877, MULT_mult_6_n876,
         MULT_mult_6_n875, MULT_mult_6_n874, MULT_mult_6_n873,
         MULT_mult_6_n872, MULT_mult_6_n871, MULT_mult_6_n870,
         MULT_mult_6_n869, MULT_mult_6_n868, MULT_mult_6_n867,
         MULT_mult_6_n866, MULT_mult_6_n865, MULT_mult_6_n864,
         MULT_mult_6_n863, MULT_mult_6_n862, MULT_mult_6_n861,
         MULT_mult_6_n860, MULT_mult_6_n859, MULT_mult_6_n858,
         MULT_mult_6_n857, MULT_mult_6_n856, MULT_mult_6_n855,
         MULT_mult_6_n854, MULT_mult_6_n853, MULT_mult_6_n852,
         MULT_mult_6_n851, MULT_mult_6_n850, MULT_mult_6_n849,
         MULT_mult_6_n848, MULT_mult_6_n847, MULT_mult_6_n846,
         MULT_mult_6_n845, MULT_mult_6_n844, MULT_mult_6_n843,
         MULT_mult_6_n842, MULT_mult_6_n841, MULT_mult_6_n840,
         MULT_mult_6_n839, MULT_mult_6_n838, MULT_mult_6_n837,
         MULT_mult_6_n836, MULT_mult_6_n835, MULT_mult_6_n834,
         MULT_mult_6_n833, MULT_mult_6_n832, MULT_mult_6_n831,
         MULT_mult_6_n830, MULT_mult_6_n829, MULT_mult_6_n828,
         MULT_mult_6_n827, MULT_mult_6_n826, MULT_mult_6_n825,
         MULT_mult_6_n824, MULT_mult_6_n823, MULT_mult_6_n822,
         MULT_mult_6_n821, MULT_mult_6_n820, MULT_mult_6_n819,
         MULT_mult_6_n818, MULT_mult_6_n817, MULT_mult_6_n816,
         MULT_mult_6_n815, MULT_mult_6_n814, MULT_mult_6_n813,
         MULT_mult_6_n812, MULT_mult_6_n811, MULT_mult_6_n810,
         MULT_mult_6_n809, MULT_mult_6_n808, MULT_mult_6_n807,
         MULT_mult_6_n806, MULT_mult_6_n805, MULT_mult_6_n804,
         MULT_mult_6_n803, MULT_mult_6_n802, MULT_mult_6_n801,
         MULT_mult_6_n800, MULT_mult_6_n799, MULT_mult_6_n798,
         MULT_mult_6_n797, MULT_mult_6_n796, MULT_mult_6_n795,
         MULT_mult_6_n794, MULT_mult_6_n793, MULT_mult_6_n792,
         MULT_mult_6_n791, MULT_mult_6_n790, MULT_mult_6_n789,
         MULT_mult_6_n788, MULT_mult_6_n787, MULT_mult_6_n786,
         MULT_mult_6_n785, MULT_mult_6_n784, MULT_mult_6_n783,
         MULT_mult_6_n782, MULT_mult_6_n781, MULT_mult_6_n780,
         MULT_mult_6_n779, MULT_mult_6_n778, MULT_mult_6_n777,
         MULT_mult_6_n776, MULT_mult_6_n775, MULT_mult_6_n774,
         MULT_mult_6_n773, MULT_mult_6_n772, MULT_mult_6_n771,
         MULT_mult_6_n770, MULT_mult_6_n769, MULT_mult_6_n768,
         MULT_mult_6_n767, MULT_mult_6_n766, MULT_mult_6_n765,
         MULT_mult_6_n764, MULT_mult_6_n763, MULT_mult_6_n762,
         MULT_mult_6_n761, MULT_mult_6_n760, MULT_mult_6_n759,
         MULT_mult_6_n758, MULT_mult_6_n757, MULT_mult_6_n756,
         MULT_mult_6_n755, MULT_mult_6_n754, MULT_mult_6_n753,
         MULT_mult_6_n752, MULT_mult_6_n751, MULT_mult_6_n750,
         MULT_mult_6_n749, MULT_mult_6_n748, MULT_mult_6_n747,
         MULT_mult_6_n746, MULT_mult_6_n745, MULT_mult_6_n744,
         MULT_mult_6_n743, MULT_mult_6_n742, MULT_mult_6_n741,
         MULT_mult_6_n740, MULT_mult_6_n739, MULT_mult_6_n738,
         MULT_mult_6_n737, MULT_mult_6_n736, MULT_mult_6_n735,
         MULT_mult_6_n734, MULT_mult_6_n733, MULT_mult_6_n732,
         MULT_mult_6_n731, MULT_mult_6_n730, MULT_mult_6_n729,
         MULT_mult_6_n728, MULT_mult_6_n727, MULT_mult_6_n726,
         MULT_mult_6_n725, MULT_mult_6_n724, MULT_mult_6_n723,
         MULT_mult_6_n722, MULT_mult_6_n721, MULT_mult_6_n720,
         MULT_mult_6_n719, MULT_mult_6_n718, MULT_mult_6_n717,
         MULT_mult_6_n716, MULT_mult_6_n715, MULT_mult_6_n714,
         MULT_mult_6_n713, MULT_mult_6_n712, MULT_mult_6_n711,
         MULT_mult_6_n710, MULT_mult_6_n709, MULT_mult_6_n708,
         MULT_mult_6_n707, MULT_mult_6_n706, MULT_mult_6_n705,
         MULT_mult_6_n704, MULT_mult_6_n703, MULT_mult_6_n702,
         MULT_mult_6_n701, MULT_mult_6_n700, MULT_mult_6_n699,
         MULT_mult_6_n698, MULT_mult_6_n697, MULT_mult_6_n696,
         MULT_mult_6_n695, MULT_mult_6_n694, MULT_mult_6_n693,
         MULT_mult_6_n692, MULT_mult_6_n691, MULT_mult_6_n690,
         MULT_mult_6_n689, MULT_mult_6_n688, MULT_mult_6_n687,
         MULT_mult_6_n686, MULT_mult_6_n685, MULT_mult_6_n684,
         MULT_mult_6_n683, MULT_mult_6_n682, MULT_mult_6_n681,
         MULT_mult_6_n680, MULT_mult_6_n679, MULT_mult_6_n678,
         MULT_mult_6_n677, MULT_mult_6_n676, MULT_mult_6_n675,
         MULT_mult_6_n674, MULT_mult_6_n673, MULT_mult_6_n672,
         MULT_mult_6_n671, MULT_mult_6_n670, MULT_mult_6_n669,
         MULT_mult_6_n668, MULT_mult_6_n667, MULT_mult_6_n666,
         MULT_mult_6_n665, MULT_mult_6_n664, MULT_mult_6_n663,
         MULT_mult_6_n662, MULT_mult_6_n661, MULT_mult_6_n660,
         MULT_mult_6_n659, MULT_mult_6_n658, MULT_mult_6_n657,
         MULT_mult_6_n656, MULT_mult_6_n655, MULT_mult_6_n654,
         MULT_mult_6_n653, MULT_mult_6_n652, MULT_mult_6_n651,
         MULT_mult_6_n649, MULT_mult_6_n648, MULT_mult_6_n647,
         MULT_mult_6_n646, MULT_mult_6_n645, MULT_mult_6_n644,
         MULT_mult_6_n643, MULT_mult_6_n642, MULT_mult_6_n641,
         MULT_mult_6_n640, MULT_mult_6_n639, MULT_mult_6_n638,
         MULT_mult_6_n637, MULT_mult_6_n636, MULT_mult_6_n635,
         MULT_mult_6_n634, MULT_mult_6_n633, MULT_mult_6_n632,
         MULT_mult_6_n631, MULT_mult_6_n630, MULT_mult_6_n629,
         MULT_mult_6_n628, MULT_mult_6_n627, MULT_mult_6_n626,
         MULT_mult_6_n625, MULT_mult_6_n624, MULT_mult_6_n623,
         MULT_mult_6_n622, MULT_mult_6_n621, MULT_mult_6_n620,
         MULT_mult_6_n619, MULT_mult_6_n618, MULT_mult_6_n617,
         MULT_mult_6_n616, MULT_mult_6_n615, MULT_mult_6_n614,
         MULT_mult_6_n613, MULT_mult_6_n612, MULT_mult_6_n611,
         MULT_mult_6_n610, MULT_mult_6_n609, MULT_mult_6_n608,
         MULT_mult_6_n607, MULT_mult_6_n606, MULT_mult_6_n605,
         MULT_mult_6_n604, MULT_mult_6_n603, MULT_mult_6_n602,
         MULT_mult_6_n601, MULT_mult_6_n600, MULT_mult_6_n599,
         MULT_mult_6_n598, MULT_mult_6_n597, MULT_mult_6_n596,
         MULT_mult_6_n595, MULT_mult_6_n594, MULT_mult_6_n593,
         MULT_mult_6_n592, MULT_mult_6_n591, MULT_mult_6_n590,
         MULT_mult_6_n589, MULT_mult_6_n588, MULT_mult_6_n587,
         MULT_mult_6_n586, MULT_mult_6_n585, MULT_mult_6_n584,
         MULT_mult_6_n583, MULT_mult_6_n582, MULT_mult_6_n581,
         MULT_mult_6_n580, MULT_mult_6_n579, MULT_mult_6_n578,
         MULT_mult_6_n577, MULT_mult_6_n576, MULT_mult_6_n575,
         MULT_mult_6_n574, MULT_mult_6_n573, MULT_mult_6_n572,
         MULT_mult_6_n571, MULT_mult_6_n570, MULT_mult_6_n569,
         MULT_mult_6_n568, MULT_mult_6_n567, MULT_mult_6_n566,
         MULT_mult_6_n565, MULT_mult_6_n564, MULT_mult_6_n563,
         MULT_mult_6_n562, MULT_mult_6_n561, MULT_mult_6_n560,
         MULT_mult_6_n559, MULT_mult_6_n558, MULT_mult_6_n557,
         MULT_mult_6_n556, MULT_mult_6_n555, MULT_mult_6_n554,
         MULT_mult_6_n553, MULT_mult_6_n552, MULT_mult_6_n551,
         MULT_mult_6_n550, MULT_mult_6_n549, MULT_mult_6_n548,
         MULT_mult_6_n547, MULT_mult_6_n546, MULT_mult_6_n545,
         MULT_mult_6_n544, MULT_mult_6_n543, MULT_mult_6_n542,
         MULT_mult_6_n541, MULT_mult_6_n540, MULT_mult_6_n539,
         MULT_mult_6_n538, MULT_mult_6_n537, MULT_mult_6_n536,
         MULT_mult_6_n535, MULT_mult_6_n534, MULT_mult_6_n533,
         MULT_mult_6_n532, MULT_mult_6_n531, MULT_mult_6_n530,
         MULT_mult_6_n529, MULT_mult_6_n528, MULT_mult_6_n527,
         MULT_mult_6_n526, MULT_mult_6_n525, MULT_mult_6_n524,
         MULT_mult_6_n523, MULT_mult_6_n522, MULT_mult_6_n521,
         MULT_mult_6_n520, MULT_mult_6_n519, MULT_mult_6_n518,
         MULT_mult_6_n517, MULT_mult_6_n516, MULT_mult_6_n515,
         MULT_mult_6_n514, MULT_mult_6_n513, MULT_mult_6_n512,
         MULT_mult_6_n511, MULT_mult_6_n510, MULT_mult_6_n509,
         MULT_mult_6_n508, MULT_mult_6_n507, MULT_mult_6_n506,
         MULT_mult_6_n505, MULT_mult_6_n504, MULT_mult_6_n503,
         MULT_mult_6_n502, MULT_mult_6_n501, MULT_mult_6_n500,
         MULT_mult_6_n499, MULT_mult_6_n498, MULT_mult_6_n497,
         MULT_mult_6_n496, MULT_mult_6_n495, MULT_mult_6_n494,
         MULT_mult_6_n493, MULT_mult_6_n492, MULT_mult_6_n491,
         MULT_mult_6_n490, MULT_mult_6_n489, MULT_mult_6_n488,
         MULT_mult_6_n487, MULT_mult_6_n486, MULT_mult_6_n485,
         MULT_mult_6_n484, MULT_mult_6_n483, MULT_mult_6_n482,
         MULT_mult_6_n481, MULT_mult_6_n480, MULT_mult_6_n479,
         MULT_mult_6_n478, MULT_mult_6_n477, MULT_mult_6_n476,
         MULT_mult_6_n475, MULT_mult_6_n474, MULT_mult_6_n473,
         MULT_mult_6_n472, MULT_mult_6_n471, MULT_mult_6_n470,
         MULT_mult_6_n469, MULT_mult_6_n468, MULT_mult_6_n467,
         MULT_mult_6_n466, MULT_mult_6_n465, MULT_mult_6_n464,
         MULT_mult_6_n463, MULT_mult_6_n462, MULT_mult_6_n461,
         MULT_mult_6_n460, MULT_mult_6_n459, MULT_mult_6_n458,
         MULT_mult_6_n457, MULT_mult_6_n456, MULT_mult_6_n455,
         MULT_mult_6_n454, MULT_mult_6_n453, MULT_mult_6_n452,
         MULT_mult_6_n451, MULT_mult_6_n450, MULT_mult_6_n449,
         MULT_mult_6_n448, MULT_mult_6_n447, MULT_mult_6_n446,
         MULT_mult_6_n445, MULT_mult_6_n444, MULT_mult_6_n443,
         MULT_mult_6_n442, MULT_mult_6_n441, MULT_mult_6_n440,
         MULT_mult_6_n439, MULT_mult_6_n438, MULT_mult_6_n437,
         MULT_mult_6_n436, MULT_mult_6_n435, MULT_mult_6_n434,
         MULT_mult_6_n433, MULT_mult_6_n432, MULT_mult_6_n431,
         MULT_mult_6_n430, MULT_mult_6_n429, MULT_mult_6_n428,
         MULT_mult_6_n427, MULT_mult_6_n426, MULT_mult_6_n425,
         MULT_mult_6_n424, MULT_mult_6_n423, MULT_mult_6_n422,
         MULT_mult_6_n421, MULT_mult_6_n420, MULT_mult_6_n419,
         MULT_mult_6_n418, MULT_mult_6_n417, MULT_mult_6_n416,
         MULT_mult_6_n415, MULT_mult_6_n414, MULT_mult_6_n413,
         MULT_mult_6_n412, MULT_mult_6_n411, MULT_mult_6_n410,
         MULT_mult_6_n409, MULT_mult_6_n408, MULT_mult_6_n407,
         MULT_mult_6_n406, MULT_mult_6_n405, MULT_mult_6_n404,
         MULT_mult_6_n403, MULT_mult_6_n402, MULT_mult_6_n401,
         MULT_mult_6_n400, MULT_mult_6_n399, MULT_mult_6_n398,
         MULT_mult_6_n397, MULT_mult_6_n396, MULT_mult_6_n395,
         MULT_mult_6_n394, MULT_mult_6_n393, MULT_mult_6_n392,
         MULT_mult_6_n391, MULT_mult_6_n390, MULT_mult_6_n389,
         MULT_mult_6_n388, MULT_mult_6_n387, MULT_mult_6_n386,
         MULT_mult_6_n385, MULT_mult_6_n384, MULT_mult_6_n383,
         MULT_mult_6_n382, MULT_mult_6_n381, MULT_mult_6_n380,
         MULT_mult_6_n379, MULT_mult_6_n378, MULT_mult_6_n377,
         MULT_mult_6_n376, MULT_mult_6_n375, MULT_mult_6_n374,
         MULT_mult_6_n373, MULT_mult_6_n372, MULT_mult_6_n371,
         MULT_mult_6_n370, MULT_mult_6_n369, MULT_mult_6_n368,
         MULT_mult_6_n367, MULT_mult_6_n366, MULT_mult_6_n365,
         MULT_mult_6_n364, MULT_mult_6_n363, MULT_mult_6_n362,
         MULT_mult_6_n361, MULT_mult_6_n360, MULT_mult_6_n359,
         MULT_mult_6_n357, MULT_mult_6_n356, MULT_mult_6_n355,
         MULT_mult_6_n354, MULT_mult_6_n353, MULT_mult_6_n352,
         MULT_mult_6_n351, MULT_mult_6_n350, MULT_mult_6_n349,
         MULT_mult_6_n348, MULT_mult_6_n347, MULT_mult_6_n346,
         MULT_mult_6_n345, MULT_mult_6_n344, MULT_mult_6_n343,
         MULT_mult_6_n342, MULT_mult_6_n341, MULT_mult_6_n340,
         MULT_mult_6_n339, MULT_mult_6_n338, MULT_mult_6_n337,
         MULT_mult_6_n336, MULT_mult_6_n335, MULT_mult_6_n334,
         MULT_mult_6_n333, MULT_mult_6_n332, MULT_mult_6_n331,
         MULT_mult_6_n330, MULT_mult_6_n329, MULT_mult_6_n328,
         MULT_mult_6_n327, MULT_mult_6_n326, MULT_mult_6_n325,
         MULT_mult_6_n324, MULT_mult_6_n323, MULT_mult_6_n322,
         MULT_mult_6_n321, MULT_mult_6_n320, MULT_mult_6_n319,
         MULT_mult_6_n318, MULT_mult_6_n317, MULT_mult_6_n316,
         MULT_mult_6_n315, MULT_mult_6_n314, MULT_mult_6_n313,
         MULT_mult_6_n312, MULT_mult_6_n311, MULT_mult_6_n310,
         MULT_mult_6_n309, MULT_mult_6_n308, MULT_mult_6_n307,
         MULT_mult_6_n306, MULT_mult_6_n305, MULT_mult_6_n304,
         MULT_mult_6_n303, MULT_mult_6_n302, MULT_mult_6_n301,
         MULT_mult_6_n300, MULT_mult_6_n299, MULT_mult_6_n298,
         MULT_mult_6_n297, MULT_mult_6_n296, MULT_mult_6_n295,
         MULT_mult_6_n294, MULT_mult_6_n293, MULT_mult_6_n292,
         MULT_mult_6_n291, MULT_mult_6_n290, MULT_mult_6_n289,
         MULT_mult_6_n288, MULT_mult_6_n287, MULT_mult_6_n286,
         MULT_mult_6_n285, MULT_mult_6_n284, MULT_mult_6_n283,
         MULT_mult_6_n282, MULT_mult_6_n281, MULT_mult_6_n280,
         MULT_mult_6_n279, MULT_mult_6_n278, MULT_mult_6_n277,
         MULT_mult_6_n276, MULT_mult_6_n275, MULT_mult_6_n274,
         MULT_mult_6_n273, MULT_mult_6_n272, MULT_mult_6_n271,
         MULT_mult_6_n270, MULT_mult_6_n269, MULT_mult_6_n268,
         MULT_mult_6_n267, MULT_mult_6_n266, MULT_mult_6_n265,
         MULT_mult_6_n264, MULT_mult_6_n263, MULT_mult_6_n262,
         MULT_mult_6_n261, MULT_mult_6_n260, MULT_mult_6_n259,
         MULT_mult_6_n258, MULT_mult_6_n257, MULT_mult_6_n256,
         MULT_mult_6_n255, MULT_mult_6_n254, MULT_mult_6_n253,
         MULT_mult_6_n252, MULT_mult_6_n251, MULT_mult_6_n250,
         MULT_mult_6_n249, MULT_mult_6_n248, MULT_mult_6_n247,
         MULT_mult_6_n246, MULT_mult_6_n245, MULT_mult_6_n244,
         MULT_mult_6_n243, MULT_mult_6_n242, MULT_mult_6_n241,
         MULT_mult_6_n240, MULT_mult_6_n239, MULT_mult_6_n238,
         MULT_mult_6_n237, MULT_mult_6_n236, MULT_mult_6_n235,
         MULT_mult_6_n234, MULT_mult_6_n233, MULT_mult_6_n232,
         MULT_mult_6_n231, MULT_mult_6_n230, MULT_mult_6_n229,
         MULT_mult_6_n228, MULT_mult_6_n227, MULT_mult_6_n226,
         MULT_mult_6_n225, MULT_mult_6_n224, MULT_mult_6_n223,
         MULT_mult_6_n222, MULT_mult_6_n221, MULT_mult_6_n220,
         MULT_mult_6_n219, MULT_mult_6_n218, MULT_mult_6_n217,
         MULT_mult_6_n216, MULT_mult_6_n215, MULT_mult_6_n214,
         MULT_mult_6_n213, MULT_mult_6_n212, MULT_mult_6_n211,
         MULT_mult_6_n210, MULT_mult_6_n209, MULT_mult_6_n208,
         MULT_mult_6_n207, MULT_mult_6_n206, MULT_mult_6_n204,
         MULT_mult_6_n203, MULT_mult_6_n202, MULT_mult_6_n201,
         MULT_mult_6_n200, MULT_mult_6_n199, MULT_mult_6_n198,
         MULT_mult_6_n197, MULT_mult_6_n196, MULT_mult_6_n195,
         MULT_mult_6_n194, MULT_mult_6_n193, MULT_mult_6_n192,
         MULT_mult_6_n191, MULT_mult_6_n190, MULT_mult_6_n189,
         MULT_mult_6_n188, MULT_mult_6_n187, MULT_mult_6_n186,
         MULT_mult_6_n185, MULT_mult_6_n184, MULT_mult_6_n183,
         MULT_mult_6_n182, MULT_mult_6_n181, MULT_mult_6_n180,
         MULT_mult_6_n179, MULT_mult_6_n178, MULT_mult_6_n177,
         MULT_mult_6_n176, MULT_mult_6_n175, MULT_mult_6_n174,
         MULT_mult_6_n173, MULT_mult_6_n172, MULT_mult_6_n171,
         MULT_mult_6_n170, MULT_mult_6_n169, MULT_mult_6_n168,
         MULT_mult_6_n167, MULT_mult_6_n166, MULT_mult_6_n165,
         MULT_mult_6_n164, MULT_mult_6_n163, MULT_mult_6_n162,
         MULT_mult_6_n161, MULT_mult_6_n160, MULT_mult_6_n159,
         MULT_mult_6_n158, MULT_mult_6_n157, MULT_mult_6_n156,
         MULT_mult_6_n155, MULT_mult_6_n154, MULT_mult_6_n153,
         MULT_mult_6_n152, MULT_mult_6_n151, MULT_mult_6_n150,
         MULT_mult_6_n149, MULT_mult_6_n148, MULT_mult_6_n147,
         MULT_mult_6_n146, MULT_mult_6_n145, MULT_mult_6_n144,
         MULT_mult_6_n143, MULT_mult_6_n142, MULT_mult_6_n141,
         MULT_mult_6_n140, MULT_mult_6_n139, MULT_mult_6_n138,
         MULT_mult_6_n137, MULT_mult_6_n136, MULT_mult_6_n135,
         MULT_mult_6_n134, MULT_mult_6_n133, MULT_mult_6_n132,
         MULT_mult_6_n131, MULT_mult_6_n130, MULT_mult_6_n129,
         MULT_mult_6_n128, MULT_mult_6_n127, MULT_mult_6_n126,
         MULT_mult_6_n125, MULT_mult_6_n124, MULT_mult_6_n123,
         MULT_mult_6_n122, MULT_mult_6_n120, MULT_mult_6_n119,
         MULT_mult_6_n118, MULT_mult_6_n117, MULT_mult_6_n116,
         MULT_mult_6_n115, MULT_mult_6_n114, MULT_mult_6_n113,
         MULT_mult_6_n112, MULT_mult_6_n111, MULT_mult_6_n110,
         MULT_mult_6_n109, MULT_mult_6_n108, MULT_mult_6_n107,
         MULT_mult_6_n106, MULT_mult_6_n105, MULT_mult_6_n104,
         MULT_mult_6_n103, MULT_mult_6_n102, MULT_mult_6_n101,
         MULT_mult_6_n100, MULT_mult_6_n99, MULT_mult_6_n98, MULT_mult_6_n97,
         MULT_mult_6_n96, MULT_mult_6_n95, MULT_mult_6_n94, MULT_mult_6_n93,
         MULT_mult_6_n92, MULT_mult_6_n91, MULT_mult_6_n90, MULT_mult_6_n89,
         MULT_mult_6_n88, MULT_mult_6_n87, MULT_mult_6_n86, MULT_mult_6_n85,
         MULT_mult_6_n84, MULT_mult_6_n83, MULT_mult_6_n82, MULT_mult_6_n81,
         MULT_mult_6_n80, MULT_mult_6_n79, MULT_mult_6_n78, MULT_mult_6_n77,
         MULT_mult_6_n76, MULT_mult_6_n75, MULT_mult_6_n74, MULT_mult_6_n73,
         MULT_mult_6_n72, MULT_mult_6_n71, MULT_mult_6_n70, MULT_mult_6_n69,
         MULT_mult_6_n68, MULT_mult_6_n67, MULT_mult_6_n66, MULT_mult_6_n65,
         MULT_mult_6_n64, MULT_mult_6_n63, MULT_mult_6_n62, MULT_mult_6_n61,
         MULT_mult_6_n60, MULT_mult_6_n59, MULT_mult_6_n58, MULT_mult_6_n57,
         MULT_mult_6_n56, MULT_mult_6_n55, MULT_mult_6_n54, MULT_mult_6_n53,
         MULT_mult_6_n52, MULT_mult_6_n51, MULT_mult_6_n50, MULT_mult_6_n49,
         MULT_mult_6_n48, MULT_mult_6_n47, MULT_mult_6_n46, MULT_mult_6_n45,
         MULT_mult_6_n44, MULT_mult_6_n43, MULT_mult_6_n42, MULT_mult_6_n41,
         MULT_mult_6_n40, MULT_mult_6_n39, MULT_mult_6_n38, MULT_mult_6_n37,
         MULT_mult_6_n36, MULT_mult_6_n35, MULT_mult_6_n34, MULT_mult_6_n33,
         MULT_mult_6_n32, MULT_mult_6_n31, MULT_mult_6_n30, MULT_mult_6_n29,
         MULT_mult_6_n28, MULT_mult_6_n27, MULT_mult_6_n26, MULT_mult_6_n25,
         MULT_mult_6_n24, MULT_mult_6_n23, MULT_mult_6_n22, MULT_mult_6_n21,
         MULT_mult_6_n20, MULT_mult_6_n19, MULT_mult_6_n18, MULT_mult_6_n17,
         MULT_mult_6_n16, MULT_mult_6_n15, MULT_mult_6_n14, MULT_mult_6_n13,
         MULT_mult_6_n12, MULT_mult_6_n11, MULT_mult_6_n10, MULT_mult_6_n9,
         MULT_mult_6_n8, MULT_mult_6_n7, MULT_mult_6_n6, MULT_mult_6_n5,
         MULT_mult_6_n4, MULT_mult_6_n3, MULT_mult_6_SUMB_6__12_,
         MULT_mult_6_net81209, MULT_mult_6_net83045, MULT_mult_6_net87460,
         MULT_mult_6_net87461, MULT_mult_6_net87462, MULT_mult_6_net88105,
         MULT_mult_6_net88106, MULT_mult_6_net88107, MULT_mult_6_net89021,
         MULT_mult_6__UDW__112699_net78589, MULT_mult_6_CARRYB_1__14_,
         MULT_mult_6_SUMB_1__15_, MULT_mult_6_SUMB_3__13_,
         MULT_mult_6_ab_0__16_, MULT_mult_6_net70466, MULT_mult_6_net81416,
         MULT_mult_6_net81694, MULT_mult_6_net84270, MULT_mult_6_net85493,
         MULT_mult_6_net88010, MULT_mult_6_net89227, MULT_mult_6_CARRYB_6__11_,
         MULT_mult_6_SUMB_5__12_, MULT_mult_6_ab_7__11_, MULT_mult_6_net84652,
         MULT_mult_6_CARRYB_4__11_, MULT_mult_6_CARRYB_5__11_,
         MULT_mult_6_SUMB_4__12_, MULT_mult_6_ab_5__11_, MULT_mult_6_net124527,
         MULT_mult_6_net82762, MULT_mult_6_net82763, MULT_mult_6_net88084,
         MULT_mult_6_net88085, MULT_mult_6__UDW__112699_net78591,
         MULT_mult_6_CARRYB_1__13_, MULT_mult_6_CARRYB_2__13_,
         MULT_mult_6_SUMB_1__14_, MULT_mult_6_ab_0__14_, MULT_mult_6_ab_2__13_,
         MULT_mult_6_net120391, MULT_mult_6_net120392, MULT_mult_6_net124833,
         MULT_mult_6_net70462, MULT_mult_6_SUMB_7__11_,
         MULT_mult_6_CARRYB_9__10_, MULT_mult_6_ab_10__10_,
         MULT_mult_6_net81001, MULT_mult_6_net81256, MULT_mult_6_net81643,
         MULT_mult_6_net83061, MULT_mult_6_net83062, MULT_mult_6_net87456,
         MULT_mult_6_net87457, MULT_mult_6_net87458, MULT_mult_6_net87459,
         MULT_mult_6_net91298, MULT_mult_6_CARRYB_12__8_,
         MULT_mult_6_SUMB_11__9_, MULT_mult_6_ab_13__8_, MULT_mult_6_net70450,
         MULT_mult_6_net77922, MULT_mult_6_net80505, MULT_mult_6_net80506,
         MULT_mult_6_net80507, MULT_mult_6_net81115, MULT_mult_6_net81116,
         MULT_mult_6_net88104, MULT_mult_6_CARRYB_8__10_,
         MULT_mult_6_SUMB_8__11_, MULT_mult_6_ab_9__10_, MULT_mult_6_net81215,
         MULT_mult_6_net81216, MULT_mult_6_CARRYB_11__8_,
         MULT_mult_6_ab_12__8_, MULT_mult_6_net121445, MULT_mult_6_net121446,
         MULT_mult_6_net121447, MULT_mult_6_net89537, MULT_mult_6_ab_6__11_,
         MULT_mult_6_net86151, MULT_mult_6_ab_1__14_, MULT_mult_6_net70493,
         MULT_mult_6_net77984, MULT_mult_6_net84070, MULT_mult_6_net84071,
         MULT_mult_6_net91259, MULT_mult_6_SUMB_10__10_,
         MULT_mult_6_SUMB_9__11_, MULT_mult_6_net83042, MULT_mult_6_net84069,
         MULT_mult_6_net84072, MULT_mult_6_CARRYB_10__9_, MULT_mult_6_net84267,
         MULT_mult_6_net84268, MULT_mult_6_net90735, MULT_mult_6_net93304,
         MULT_mult_6_net93305, MULT_mult_6_net93306, MULT_mult_6_net93307,
         MULT_mult_6_ab_11__9_, MULT_mult_6_net84654, MULT_mult_6_net84656,
         MULT_mult_6_net91419, MULT_mult_6_ab_0__15_, MULT_mult_6_ab_1__13_,
         MULT_mult_6_ab_3__13_, MULT_mult_6_CARRYB_7__10_,
         MULT_mult_6_CARRYB_13__8_, MULT_mult_6_SUMB_12__9_,
         MULT_mult_6_net122062, MULT_mult_6_net89168, MULT_mult_6_ab_8__10_,
         MULT_mult_6_ab_1__15_, MULT_mult_6_net87396, MULT_mult_6_ab_28__1_,
         MULT_mult_6_net79883, MULT_mult_6_net79884, MULT_mult_6_net79885,
         MULT_mult_6_net85287, MULT_mult_6_net86792, MULT_mult_6_net87798,
         MULT_mult_6_net92330, MULT_mult_6_net92331, MULT_mult_6_ab_5__14_,
         MULT_mult_6_net119908, MULT_mult_6_net119927, MULT_mult_6_net119948,
         MULT_mult_6_net148836, MULT_mult_6_net148837, MULT_mult_6_net148838,
         MULT_mult_6_net83918, MULT_mult_6_CARRYB_14__8_,
         MULT_mult_6_SUMB_14__8_, MULT_mult_6_SUMB_14__9_,
         MULT_mult_6_SUMB_15__8_, MULT_mult_6_net81666, MULT_mult_6_net81667,
         MULT_mult_6_net81668, MULT_mult_6_net83273, MULT_mult_6_net86536,
         MULT_mult_6_net86537, MULT_mult_6_net88904, MULT_mult_6_SUMB_21__5_,
         MULT_mult_6_net147924, MULT_mult_6_net147925, MULT_mult_6_net147926,
         MULT_mult_6_net149133, MULT_mult_6_net80862, MULT_mult_6_net83705,
         MULT_mult_6_net123365, MULT_mult_6_net80986, MULT_mult_6_net81867,
         MULT_mult_6_net83623, MULT_mult_6_net83624, MULT_mult_6_net83625,
         MULT_mult_6_net89460, MULT_mult_6_SUMB_16__7_, MULT_mult_6_net80906,
         MULT_mult_6_net82288, MULT_mult_6_net82289, MULT_mult_6_net85372,
         MULT_mult_6_CARRYB_22__5_, MULT_mult_6_SUMB_21__6_,
         MULT_mult_6_SUMB_22__5_, MULT_mult_6_SUMB_23__4_,
         MULT_mult_6_ab_22__5_, MULT_mult_6_net120364, MULT_mult_6_net120366,
         MULT_mult_6_net83101, MULT_mult_6_net84666, MULT_mult_6_net84667,
         MULT_mult_6_net84668, MULT_mult_6_net85109, MULT_mult_6_net86109,
         MULT_mult_6_net88648, MULT_mult_6_net89455, MULT_mult_6_net119909,
         MULT_mult_6_net119910, MULT_mult_6_net119955, MULT_mult_6_net119960,
         MULT_mult_6_net119974, MULT_mult_6_net123266, MULT_mult_6_net123267,
         MULT_mult_6_net123268, MULT_mult_6_net123269,
         MULT_mult_6_CARRYB_15__7_, MULT_mult_6_ab_16__7_,
         MULT_mult_6_net70448, MULT_mult_6_net77916, MULT_mult_6_net80536,
         MULT_mult_6_net80537, MULT_mult_6_net80538, MULT_mult_6_net86374,
         MULT_mult_6_net86375, MULT_mult_6_SUMB_13__9_, MULT_mult_6_ab_14__8_,
         MULT_mult_6_net148828, MULT_mult_6_net148829, MULT_mult_6_net87363,
         MULT_mult_6_net89652, MULT_mult_6_net119928, MULT_mult_6_net119951,
         MULT_mult_6_net123752, MULT_mult_6_net82152,
         MULT_mult_6_CARRYB_7__12_, MULT_mult_6_CARRYB_8__12_,
         MULT_mult_6_SUMB_7__13_, MULT_mult_6_ab_8__12_, MULT_mult_6_net70458,
         MULT_mult_6_net80847, MULT_mult_6_net80848, MULT_mult_6_CARRYB_21__3_,
         MULT_mult_6_CARRYB_22__3_, MULT_mult_6_CARRYB_24__2_,
         MULT_mult_6_SUMB_22__4_, MULT_mult_6_ab_23__3_, MULT_mult_6_net86519,
         MULT_mult_6_net86520, MULT_mult_6_net88665, MULT_mult_6_net92568,
         MULT_mult_6_net92569, MULT_mult_6_CARRYB_10__11_,
         MULT_mult_6_SUMB_11__11_, MULT_mult_6_net81165, MULT_mult_6_net84874,
         MULT_mult_6_net85537, MULT_mult_6_net85539, MULT_mult_6_net87043,
         MULT_mult_6_net88302, MULT_mult_6_net88303, MULT_mult_6_net89167,
         MULT_mult_6_net89369, MULT_mult_6_net89447, MULT_mult_6_net89840,
         MULT_mult_6_net92550, MULT_mult_6_net92551, MULT_mult_6_net92552,
         MULT_mult_6_net92553, MULT_mult_6_CARRYB_12__9_,
         MULT_mult_6_SUMB_12__10_, MULT_mult_6_net81182, MULT_mult_6_net82292,
         MULT_mult_6_net82294, MULT_mult_6_net82295, MULT_mult_6_net83848,
         MULT_mult_6_net86142, MULT_mult_6_net86144, MULT_mult_6_net86145,
         MULT_mult_6_net92622, MULT_mult_6_CARRYB_17__6_,
         MULT_mult_6_SUMB_17__6_, MULT_mult_6_SUMB_18__6_,
         MULT_mult_6_net120625, MULT_mult_6_net124589, MULT_mult_6_net81264,
         MULT_mult_6_net82403, MULT_mult_6_net82404, MULT_mult_6_net82748,
         MULT_mult_6_net85610, MULT_mult_6_net85611, MULT_mult_6_net86806,
         MULT_mult_6_net88878, MULT_mult_6_net90576, MULT_mult_6_net91377,
         MULT_mult_6_CARRYB_27__0_, MULT_mult_6_SUMB_27__1_,
         MULT_mult_6_net80771, MULT_mult_6_net80773,
         MULT_mult_6_CARRYB_11__10_, MULT_mult_6_ab_12__10_,
         MULT_mult_6_net121898, MULT_mult_6_net83880, MULT_mult_6_net83881,
         MULT_mult_6_net83882, MULT_mult_6_net84873, MULT_mult_6_net80564,
         MULT_mult_6_CARRYB_28__0_, MULT_mult_6_net70436, MULT_mult_6_net77864,
         MULT_mult_6_net82838, MULT_mult_6_net83876, MULT_mult_6_net87364,
         MULT_mult_6_net87365, MULT_mult_6_net87366, MULT_mult_6_net87367,
         MULT_mult_6_net91003, MULT_mult_6_SUMB_8__13_, MULT_mult_6_net81373,
         MULT_mult_6_net81374, MULT_mult_6_net81375, MULT_mult_6_net82837,
         MULT_mult_6_net84669, MULT_mult_6_net84670, MULT_mult_6_net84671,
         MULT_mult_6_net84672, MULT_mult_6_net84867, MULT_mult_6_net84868,
         MULT_mult_6_net84870, MULT_mult_6_net85459, MULT_mult_6_net85460,
         MULT_mult_6_net85461, MULT_mult_6_net88841, MULT_mult_6_net89149,
         MULT_mult_6_CARRYB_20__5_, MULT_mult_6_SUMB_19__6_,
         MULT_mult_6_ab_20__5_, MULT_mult_6_net120626, MULT_mult_6_net70444,
         MULT_mult_6_net77904, MULT_mult_6_net82405, MULT_mult_6_ab_19__6_,
         MULT_mult_6_net124627, MULT_mult_6_net81268, MULT_mult_6_net81270,
         MULT_mult_6_net81947, MULT_mult_6_net82009, MULT_mult_6_net90810,
         MULT_mult_6_net93914, MULT_mult_6_SUMB_10__11_, MULT_mult_6_ab_1__17_,
         MULT_mult_6_net82286, MULT_mult_6_net85688, MULT_mult_6_net86959,
         MULT_mult_6_net87050, MULT_mult_6_ab_9__12_, MULT_mult_6_ab_17__6_,
         MULT_mult_6_SUMB_25__2_, MULT_mult_6_net92790,
         MULT_mult_6_CARRYB_16__6_, MULT_mult_6_SUMB_17__7_,
         MULT_mult_6_net80540, MULT_mult_6_net80541, MULT_mult_6_net81269,
         MULT_mult_6_CARRYB_25__1_, MULT_mult_6_SUMB_24__2_,
         MULT_mult_6_net83975, MULT_mult_6_net83976, MULT_mult_6_net83977,
         MULT_mult_6_CARRYB_5__14_, MULT_mult_6_CARRYB_6__14_,
         MULT_mult_6_SUMB_6__14_, MULT_mult_6_net88660, MULT_mult_6_net90348,
         MULT_mult_6_net90897, MULT_mult_6__UDW__112684_net78549,
         MULT_mult_6_net77988, MULT_mult_6_net81630, MULT_mult_6_SUMB_4__16_,
         MULT_mult_6_SUMB_5__15_, MULT_mult_6_ab_6__14_, MULT_mult_6_net82297,
         MULT_mult_6_net84446, MULT_mult_6_net84856, MULT_mult_6_ab_21__5_,
         MULT_mult_6_ab_30__0_, MULT_mult_6_net36614, MULT_mult_6_net83536,
         MULT_mult_6_CARRYB_4__14_, MULT_mult_6_net84945, MULT_mult_6_net84946,
         MULT_mult_6_ab_27__1_, MULT_mult_6_SUMB_28__2_, MULT_mult_6_ab_29__1_,
         MULT_mult_6_net81158, MULT_mult_6_net86055, MULT_mult_6_net92337,
         MULT_mult_6__UDW__112689_net78561, MULT_mult_6_CARRYB_1__16_,
         MULT_mult_6_ab_0__17_, MULT_mult_6_net119899, MULT_mult_6_net119901,
         MULT_mult_6_net119952, MULT_mult_6_SUMB_1__18_, MULT_mult_6_net84327,
         MULT_mult_6_ab_24__3_, MULT_mult_6_net124949,
         MULT_mult_6_CARRYB_20__3_, MULT_mult_6_ab_22__3_,
         MULT_mult_6_net80509, MULT_mult_6_net80511, MULT_mult_6_SUMB_20__6_,
         MULT_mult_6_SUMB_17__8_, MULT_mult_6_SUMB_18__7_,
         MULT_mult_6_net83776, MULT_mult_6_net84374, MULT_mult_6_net88856,
         MULT_mult_6_net149916, MULT_mult_6_net149917, MULT_mult_6_net149611,
         MULT_mult_6_net149605, MULT_mult_6_net149580, MULT_mult_6_net149530,
         MULT_mult_6_net149526, MULT_mult_6_net149004, MULT_mult_6_net148754,
         MULT_mult_6_net148582, MULT_mult_6_net148302, MULT_mult_6_net148230,
         MULT_mult_6_net148233, MULT_mult_6_net148235, MULT_mult_6_net148179,
         MULT_mult_6_net148051, MULT_mult_6_net148053, MULT_mult_6_net148015,
         MULT_mult_6_net147998, MULT_mult_6_net147999, MULT_mult_6_net147920,
         MULT_mult_6_net147922, MULT_mult_6_net147928, MULT_mult_6_net147929,
         MULT_mult_6_net147930, MULT_mult_6_net147936, MULT_mult_6_net147938,
         MULT_mult_6_net147939, MULT_mult_6_net147940, MULT_mult_6_net147421,
         MULT_mult_6_net147444, MULT_mult_6_net147451,
         MULT_mult_6__UDW__112734_net78687, MULT_mult_6_CARRYB_1__7_,
         MULT_mult_6_CARRYB_2__7_, MULT_mult_6_CARRYB_3__5_,
         MULT_mult_6_CARRYB_4__5_, MULT_mult_6_SUMB_1__8_,
         MULT_mult_6_SUMB_2__7_, MULT_mult_6_SUMB_3__6_, MULT_mult_6_ab_2__7_,
         MULT_mult_6_net77976, MULT_mult_6_net84928, MULT_mult_6_net84929,
         MULT_mult_6_net87961, MULT_mult_6_net87962, MULT_mult_6_CARRYB_11__1_,
         MULT_mult_6_CARRYB_12__1_, MULT_mult_6_CARRYB_13__1_,
         MULT_mult_6_SUMB_11__2_, MULT_mult_6_SUMB_12__1_,
         MULT_mult_6_SUMB_12__2_, MULT_mult_6_ab_12__1_, MULT_mult_6_ab_13__1_,
         MULT_mult_6_net122130, MULT_mult_6_net85032, MULT_mult_6_net86129,
         MULT_mult_6_net86131, MULT_mult_6_CARRYB_16__1_,
         MULT_mult_6_CARRYB_17__1_, MULT_mult_6_CARRYB_18__1_,
         MULT_mult_6_SUMB_15__2_, MULT_mult_6_SUMB_16__1_,
         MULT_mult_6_SUMB_17__2_, MULT_mult_6_ab_16__1_,
         MULT_mult_6_CARRYB_22__1_, MULT_mult_6_CARRYB_23__1_,
         MULT_mult_6_SUMB_22__2_, MULT_mult_6_ab_23__1_, MULT_mult_6_net82541,
         MULT_mult_6_net82542, MULT_mult_6_net82543, MULT_mult_6_CARRYB_19__1_,
         MULT_mult_6_SUMB_18__2_, MULT_mult_6_ab_19__1_, MULT_mult_6_net81095,
         MULT_mult_6_net81097, MULT_mult_6_net93676, MULT_mult_6_CARRYB_2__6_,
         MULT_mult_6_SUMB_1__7_, MULT_mult_6_ab_0__7_, MULT_mult_6_ab_2__6_,
         MULT_mult_6_CARRYB_13__2_, MULT_mult_6_CARRYB_14__1_,
         MULT_mult_6_CARRYB_15__1_, MULT_mult_6_SUMB_13__3_,
         MULT_mult_6_SUMB_14__2_, MULT_mult_6_SUMB_15__1_,
         MULT_mult_6_ab_14__2_, MULT_mult_6_ab_15__1_, MULT_mult_6_net86134,
         MULT_mult_6_net86135, MULT_mult_6_CARRYB_6__4_,
         MULT_mult_6_CARRYB_7__4_, MULT_mult_6_CARRYB_8__4_,
         MULT_mult_6_SUMB_6__5_, MULT_mult_6_SUMB_7__4_,
         MULT_mult_6_SUMB_7__5_, MULT_mult_6_SUMB_8__4_, MULT_mult_6_ab_8__4_,
         MULT_mult_6_net88200, MULT_mult_6_SUMB_10__3_, MULT_mult_6_ab_11__2_,
         MULT_mult_6_SUMB_23__2_, MULT_mult_6_SUMB_24__1_,
         MULT_mult_6_ab_24__1_, MULT_mult_6_net122156, MULT_mult_6_net85902,
         MULT_mult_6_net85903, MULT_mult_6_net88776, MULT_mult_6_ab_5__5_,
         MULT_mult_6_net89958, MULT_mult_6_ab_1__8_, MULT_mult_6_CARRYB_7__3_,
         MULT_mult_6_CARRYB_8__3_, MULT_mult_6_SUMB_8__3_,
         MULT_mult_6_ab_7__4_, MULT_mult_6_net88198, MULT_mult_6_net88199,
         MULT_mult_6_SUMB_4__6_, MULT_mult_6_SUMB_5__5_, MULT_mult_6_net125691,
         MULT_mult_6_ab_0__8_, MULT_mult_6_ab_1__7_, MULT_mult_6_net124610,
         MULT_mult_6_CARRYB_28__1_, MULT_mult_6_net79880, MULT_mult_6_net79881,
         MULT_mult_6_net79882, MULT_mult_6_net85094, MULT_mult_6_net89103,
         MULT_mult_6_net89104, MULT_mult_6_net89110, MULT_mult_6_net123291,
         MULT_mult_6_net123293, MULT_mult_6_net87391, MULT_mult_6_net87949,
         MULT_mult_6_net87950, MULT_mult_6_net88699, MULT_mult_6_net90022,
         MULT_mult_6_net90818, MULT_mult_6_net93279, MULT_mult_6_net93683,
         MULT_mult_6_net81042, MULT_mult_6_net81552, MULT_mult_6_net81553,
         MULT_mult_6_net81555, MULT_mult_6_net87681, MULT_mult_6_CARRYB_23__4_,
         MULT_mult_6_ab_24__4_, MULT_mult_6_net124635, MULT_mult_6_net84000,
         MULT_mult_6_net84001, MULT_mult_6_net120647, MULT_mult_6_net120648,
         MULT_mult_6_net82158, MULT_mult_6_net84059, MULT_mult_6_net87934,
         MULT_mult_6_net87935, MULT_mult_6_net87936, MULT_mult_6_net87937,
         MULT_mult_6_net81559, MULT_mult_6_net81560, MULT_mult_6_net84349,
         MULT_mult_6_net88906, MULT_mult_6_SUMB_13__11_, MULT_mult_6_net120649,
         MULT_mult_6_net93277, MULT_mult_6_CARRYB_12__10_,
         MULT_mult_6_CARRYB_13__10_, MULT_mult_6_CARRYB_14__10_,
         MULT_mult_6_ab_14__10_, MULT_mult_6_net82160, MULT_mult_6_net82161,
         MULT_mult_6_net82162, MULT_mult_6_SUMB_25__3_, MULT_mult_6_net121449,
         MULT_mult_6_net121450, MULT_mult_6_net121451, MULT_mult_6_net121452,
         MULT_mult_6_net121770, MULT_mult_6_net123363, MULT_mult_6_net80927,
         MULT_mult_6_net83054, MULT_mult_6_net83055, MULT_mult_6_net83057,
         MULT_mult_6_net81372, MULT_mult_6_net87066, MULT_mult_6_net88880,
         MULT_mult_6_net88881, MULT_mult_6_net88943, MULT_mult_6_net89356,
         MULT_mult_6_net93800, MULT_mult_6_CARRYB_3__16_,
         MULT_mult_6_SUMB_3__17_, MULT_mult_6_ab_4__16_, MULT_mult_6_net119953,
         MULT_mult_6_net119976, MULT_mult_6_net80833, MULT_mult_6_net80834,
         MULT_mult_6_net84445, MULT_mult_6_net86162, MULT_mult_6_net80667,
         MULT_mult_6_net80668, MULT_mult_6_net85096, MULT_mult_6_CARRYB_16__9_,
         MULT_mult_6_ab_17__9_, MULT_mult_6_net120655, MULT_mult_6_net120656,
         MULT_mult_6_net120657, MULT_mult_6_net121214, MULT_mult_6_net79980,
         MULT_mult_6_net79981, MULT_mult_6_net81992, MULT_mult_6_net84208,
         MULT_mult_6_net79907, MULT_mult_6_net79908, MULT_mult_6_net80021,
         MULT_mult_6_SUMB_24__4_, MULT_mult_6_ab_25__3_, MULT_mult_6_net81006,
         MULT_mult_6_net81007, MULT_mult_6_net82544, MULT_mult_6_net86022,
         MULT_mult_6_net86023, MULT_mult_6_net86024, MULT_mult_6_net87938,
         MULT_mult_6_net87939, MULT_mult_6_net87940, MULT_mult_6_net87941,
         MULT_mult_6_net88123, MULT_mult_6_CARRYB_10__12_,
         MULT_mult_6_CARRYB_9__12_, MULT_mult_6_SUMB_9__13_,
         MULT_mult_6_ab_10__12_, MULT_mult_6_net80351, MULT_mult_6_net80352,
         MULT_mult_6_net80353, MULT_mult_6_net84819, MULT_mult_6_net84820,
         MULT_mult_6_net84822, MULT_mult_6_net85399, MULT_mult_6_net89065,
         MULT_mult_6_net89982, MULT_mult_6_net90996, MULT_mult_6_net89109,
         MULT_mult_6_CARRYB_24__3_, MULT_mult_6_net84678, MULT_mult_6_net84679,
         MULT_mult_6_net84680, MULT_mult_6_CARRYB_11__11_,
         MULT_mult_6_CARRYB_12__11_, MULT_mult_6_SUMB_11__12_,
         MULT_mult_6_ab_13__11_, MULT_mult_6_net82021, MULT_mult_6_net82022,
         MULT_mult_6_net84824, MULT_mult_6_net89670, MULT_mult_6_net90262,
         MULT_mult_6_net90604, MULT_mult_6_CARRYB_26__2_, MULT_mult_6_net80261,
         MULT_mult_6_net80262, MULT_mult_6_net80263, MULT_mult_6_net80987,
         MULT_mult_6_net80988, MULT_mult_6_net80989, MULT_mult_6_net80472,
         MULT_mult_6_net80473, MULT_mult_6_net80474, MULT_mult_6_net89453,
         MULT_mult_6_ab_27__2_, MULT_mult_6_net80686, MULT_mult_6_net93918,
         MULT_mult_6_CARRYB_21__5_, MULT_mult_6_net79989, MULT_mult_6_net79990,
         MULT_mult_6_net79991, MULT_mult_6_net80290, MULT_mult_6_net84213,
         MULT_mult_6_ab_12__11_, MULT_mult_6_net81087, MULT_mult_6_net81166,
         MULT_mult_6_net81167, MULT_mult_6_net81168, MULT_mult_6_net83631,
         MULT_mult_6_net87490, MULT_mult_6_CARRYB_17__8_,
         MULT_mult_6_SUMB_17__9_, MULT_mult_6_ab_18__8_, MULT_mult_6_net85807,
         MULT_mult_6_net85808, MULT_mult_6_net87945, MULT_mult_6_net93410,
         MULT_mult_6_CARRYB_15__10_, MULT_mult_6_SUMB_14__11_,
         MULT_mult_6_SUMB_15__11_, MULT_mult_6_ab_16__10_,
         MULT_mult_6_net125934, MULT_mult_6_net82559, MULT_mult_6_net82560,
         MULT_mult_6_net82561, MULT_mult_6_net86801, MULT_mult_6_net87688,
         MULT_mult_6_net87944, MULT_mult_6_ab_23__4_, MULT_mult_6_SUMB_15__10_,
         MULT_mult_6_ab_16__9_, MULT_mult_6_net86799, MULT_mult_6_net82030,
         MULT_mult_6_SUMB_23__5_, MULT_mult_6_net79909, MULT_mult_6_net84434,
         MULT_mult_6_net89008, MULT_mult_6_net93813, MULT_mult_6_ab_2__16_,
         MULT_mult_6_ab_11__12_, MULT_mult_6_net80250, MULT_mult_6_net80251,
         MULT_mult_6_net83628, MULT_mult_6_net83629, MULT_mult_6_net83630,
         MULT_mult_6_net120511, MULT_mult_6_net124908, MULT_mult_6_net88079,
         MULT_mult_6_ab_5__15_, MULT_mult_6_net88700,
         MULT_mult_6_CARRYB_8__13_, MULT_mult_6_net81371, MULT_mult_6_net87065,
         MULT_mult_6_net87067, MULT_mult_6_net87068, MULT_mult_6_net124392,
         MULT_mult_6_net87797, MULT_mult_6_ab_15__10_, MULT_mult_6_SUMB_18__9_,
         MULT_mult_6_CARRYB_15__9_, MULT_mult_6_SUMB_14__10_,
         MULT_mult_6_net82263, MULT_mult_6_net87942, MULT_mult_6_net93756,
         MULT_mult_6_SUMB_10__13_, MULT_mult_6_ab_9__13_, MULT_mult_6_net80346,
         MULT_mult_6_net83438, MULT_mult_6_SUMB_8__14_, MULT_mult_6_net84447,
         MULT_mult_6_SUMB_26__3_, MULT_mult_6_net83030, MULT_mult_6_net86884,
         MULT_mult_6_CARRYB_29__1_, MULT_mult_6_net81157, MULT_mult_6_net87654,
         MULT_mult_6_net87655, MULT_mult_6_net92317, MULT_mult_6_net92318,
         MULT_mult_6_net92325, MULT_mult_6_net93672, MULT_mult_6_net88668,
         MULT_mult_6_net90817, MULT_mult_6_net125375, MULT_mult_6_net125062,
         MULT_mult_6_net124874, MULT_mult_6_net124757, MULT_mult_6_net124723,
         MULT_mult_6_net124618, MULT_mult_6_net124563, MULT_mult_6_net124434,
         MULT_mult_6_net124367, MULT_mult_6_net124104, MULT_mult_6_net123897,
         MULT_mult_6_net123898, MULT_mult_6_net123899, MULT_mult_6_net123842,
         MULT_mult_6_net123843, MULT_mult_6_net123591, MULT_mult_6_net123592,
         MULT_mult_6_net123509, MULT_mult_6_net123427, MULT_mult_6_net123428,
         MULT_mult_6_net123429, MULT_mult_6_net123430, MULT_mult_6_net123303,
         MULT_mult_6_net123142, MULT_mult_6_net123143, MULT_mult_6_net123019,
         MULT_mult_6_net123028, MULT_mult_6_net123055, MULT_mult_6_net123062,
         MULT_mult_6_net123072, MULT_mult_6_net123000,
         MULT_mult_6_CARRYB_7__17_, MULT_mult_6_net80366, MULT_mult_6_net80657,
         MULT_mult_6_net80658, MULT_mult_6_net80660, MULT_mult_6_CARRYB_19__9_,
         MULT_mult_6_SUMB_19__10_, MULT_mult_6_SUMB_20__9_,
         MULT_mult_6_ab_20__9_, MULT_mult_6_net81953, MULT_mult_6_net81954,
         MULT_mult_6_net82255, MULT_mult_6_net82396, MULT_mult_6_net86403,
         MULT_mult_6_net86404, MULT_mult_6_net87009, MULT_mult_6_net87134,
         MULT_mult_6_net90802, MULT_mult_6_net122087, MULT_mult_6_net121926,
         MULT_mult_6_net121859, MULT_mult_6_net121814, MULT_mult_6_net121785,
         MULT_mult_6_net121606, MULT_mult_6_net121607, MULT_mult_6_net121523,
         MULT_mult_6_net121453, MULT_mult_6_net121454, MULT_mult_6_net121455,
         MULT_mult_6_net121380, MULT_mult_6_net121285, MULT_mult_6_net121150,
         MULT_mult_6_net120922, MULT_mult_6_net120651, MULT_mult_6_net120652,
         MULT_mult_6_net120653, MULT_mult_6_net120627, MULT_mult_6_net120628,
         MULT_mult_6_net120585, MULT_mult_6_net120586, MULT_mult_6_net120513,
         MULT_mult_6_net120514, MULT_mult_6_net120515, MULT_mult_6_net120517,
         MULT_mult_6_net120518, MULT_mult_6_net120519, MULT_mult_6_net120501,
         MULT_mult_6_net120463, MULT_mult_6_net120464, MULT_mult_6_net120466,
         MULT_mult_6_net120467, MULT_mult_6_net120468, MULT_mult_6_net120359,
         MULT_mult_6_net120174, MULT_mult_6_net119979, MULT_mult_6_net119982,
         MULT_mult_6_net119920, MULT_mult_6_net119921, MULT_mult_6_net119949,
         MULT_mult_6_net119855, MULT_mult_6_net119817,
         MULT_mult_6_CARRYB_26__1_, MULT_mult_6_SUMB_26__2_,
         MULT_mult_6_net81070, MULT_mult_6_net93791, MULT_mult_6_net93792,
         MULT_mult_6_SUMB_20__5_, MULT_mult_6_net83202,
         MULT_mult_6_SUMB_15__7_, MULT_mult_6_net83755, MULT_mult_6_ab_25__2_,
         MULT_mult_6_net80257, MULT_mult_6_SUMB_10__17_, MULT_mult_6_net80517,
         MULT_mult_6_net81394, MULT_mult_6_net86407, MULT_mult_6_net86409,
         MULT_mult_6_net88225, MULT_mult_6_net88226, MULT_mult_6_CARRYB_4__22_,
         MULT_mult_6_ab_5__22_, MULT_mult_6_net81284, MULT_mult_6_net81285,
         MULT_mult_6_net84311, MULT_mult_6_net84312, MULT_mult_6_net84313,
         MULT_mult_6_CARRYB_14__13_, MULT_mult_6_SUMB_14__14_,
         MULT_mult_6_net80484, MULT_mult_6_net80485, MULT_mult_6_net85119,
         MULT_mult_6_net93107, MULT_mult_6_net79868, MULT_mult_6_net86696,
         MULT_mult_6_net88916, MULT_mult_6_CARRYB_12__14_,
         MULT_mult_6_net82657, MULT_mult_6_net82658, MULT_mult_6_net88756,
         MULT_mult_6_net80794, MULT_mult_6_net80825, MULT_mult_6_CARRYB_3__22_,
         MULT_mult_6_SUMB_3__23_, MULT_mult_6_ab_4__22_, MULT_mult_6_net87855,
         MULT_mult_6_net90671, MULT_mult_6_SUMB_11__16_,
         MULT_mult_6_CARRYB_25__5_, MULT_mult_6_SUMB_24__6_,
         MULT_mult_6_ab_25__5_, MULT_mult_6_net79867, MULT_mult_6_SUMB_2__24_,
         MULT_mult_6_CARRYB_21__7_, MULT_mult_6_SUMB_21__8_,
         MULT_mult_6_net80268, MULT_mult_6_net81113, MULT_mult_6_net90801,
         MULT_mult_6_net82043, MULT_mult_6_net82044, MULT_mult_6_net82124,
         MULT_mult_6_net83044, MULT_mult_6_net83575, MULT_mult_6_net83576,
         MULT_mult_6_net88004, MULT_mult_6_CARRYB_26__4_,
         MULT_mult_6_SUMB_26__5_, MULT_mult_6_ab_26__5_, MULT_mult_6_ab_27__4_,
         MULT_mult_6_ab_31__0_, MULT_mult_6_net82807, MULT_mult_6_net84979,
         MULT_mult_6_net86937, MULT_mult_6_net92319, MULT_mult_6_net92320,
         MULT_mult_6_net92321, MULT_mult_6_net92323, MULT_mult_6_net84978,
         MULT_mult_6_CARRYB_24__6_, MULT_mult_6_ab_24__7_,
         MULT_mult_6_net79864, MULT_mult_6_net79865, MULT_mult_6_net81946,
         MULT_mult_6_CARRYB_2__23_, MULT_mult_6_ab_3__23_,
         MULT_mult_6_net70480, MULT_mult_6_net84357,
         MULT_mult_6_CARRYB_16__12_, MULT_mult_6_CARRYB_17__12_,
         MULT_mult_6_SUMB_15__14_, MULT_mult_6_SUMB_16__13_,
         MULT_mult_6_SUMB_17__12_, MULT_mult_6_ab_17__12_,
         MULT_mult_6_net81290, MULT_mult_6_net90103, MULT_mult_6_net90525,
         MULT_mult_6_CARRYB_13__14_, MULT_mult_6_ab_14__14_,
         MULT_mult_6_ab_1__24_, MULT_mult_6_SUMB_4__23_,
         MULT_mult_6_SUMB_5__22_, MULT_mult_6_SUMB_23__7_,
         MULT_mult_6_net79863, MULT_mult_6_net80110, MULT_mult_6_net83115,
         MULT_mult_6_net83116, MULT_mult_6_net89094,
         MULT_mult_6_CARRYB_11__15_, MULT_mult_6_ab_12__15_,
         MULT_mult_6_CARRYB_15__13_, MULT_mult_6_ab_15__13_,
         MULT_mult_6_CARRYB_22__7_, MULT_mult_6_ab_22__7_,
         MULT_mult_6_net80267, MULT_mult_6_net89461, MULT_mult_6_ab_13__14_,
         MULT_mult_6_SUMB_22__8_, MULT_mult_6_net88961,
         MULT_mult_6_CARRYB_20__8_, MULT_mult_6_SUMB_19__9_,
         MULT_mult_6_ab_21__8_, MULT_mult_6_CARRYB_9__17_,
         MULT_mult_6_SUMB_9__18_, MULT_mult_6_ab_10__17_, MULT_mult_6_net79950,
         MULT_mult_6_net80801, MULT_mult_6_net80802, MULT_mult_6_net80803,
         MULT_mult_6_ab_1__23_, MULT_mult_6_ab_2__23_,
         MULT_mult_6_CARRYB_7__19_, MULT_mult_6_SUMB_7__20_,
         MULT_mult_6_SUMB_8__19_, MULT_mult_6_ab_8__19_, MULT_mult_6_net81340,
         MULT_mult_6_net86231, MULT_mult_6_CARRYB_17__11_,
         MULT_mult_6_SUMB_18__11_, MULT_mult_6_ab_18__11_,
         MULT_mult_6_net88647, MULT_mult_6_net89353, MULT_mult_6_ab_16__13_,
         MULT_mult_6_ab_23__7_, MULT_mult_6_SUMB_13__15_, MULT_mult_6_net93674,
         MULT_mult_6_CARRYB_7__18_, MULT_mult_6_CARRYB_8__18_,
         MULT_mult_6_ab_9__18_, MULT_mult_6_net80302, MULT_mult_6_net80303,
         MULT_mult_6_ab_0__25_, MULT_mult_6_CARRYB_18__10_,
         MULT_mult_6_ab_19__10_, MULT_mult_6__UDW__112644_net78437,
         MULT_mult_6_SUMB_1__25_, MULT_mult_6_ab_0__26_, MULT_mult_6_ab_2__24_,
         MULT_mult_6_net84883, MULT_mult_6_CARRYB_5__21_,
         MULT_mult_6_CARRYB_6__20_, MULT_mult_6_CARRYB_6__21_,
         MULT_mult_6_SUMB_6__21_, MULT_mult_6_ab_6__21_, MULT_mult_6_net93880,
         MULT_mult_6_net93878, MULT_mult_6_net93840, MULT_mult_6_net93747,
         MULT_mult_6_net93713, MULT_mult_6_net93308, MULT_mult_6_net93309,
         MULT_mult_6_net93243, MULT_mult_6_net93203, MULT_mult_6_net92884,
         MULT_mult_6_net92862, MULT_mult_6_net92863, MULT_mult_6_net92716,
         MULT_mult_6_net92717, MULT_mult_6_net92718, MULT_mult_6_net92724,
         MULT_mult_6_net92542, MULT_mult_6_net92405, MULT_mult_6_net92378,
         MULT_mult_6_net92311, MULT_mult_6_net92314, MULT_mult_6_net92322,
         MULT_mult_6_net92341, MULT_mult_6_SUMB_25__1_, MULT_mult_6_net91660,
         MULT_mult_6_net91301, MULT_mult_6_net91243, MULT_mult_6_net91118,
         MULT_mult_6_net91088, MULT_mult_6_net91001, MULT_mult_6_net90731,
         MULT_mult_6_net90702, MULT_mult_6_net90687, MULT_mult_6_net90433,
         MULT_mult_6_net90347, MULT_mult_6_net90174, MULT_mult_6_net89997,
         MULT_mult_6_net89876, MULT_mult_6_net89819, MULT_mult_6_net89467,
         MULT_mult_6_net89402, MULT_mult_6_net89289, MULT_mult_6_net89255,
         MULT_mult_6_net89026, MULT_mult_6_net88934, MULT_mult_6_net88928,
         MULT_mult_6_net88887, MULT_mult_6_net88867, MULT_mult_6_net88868,
         MULT_mult_6_net88859, MULT_mult_6_net88860, MULT_mult_6_net88800,
         MULT_mult_6_net88712, MULT_mult_6_net88703, MULT_mult_6_net88704,
         MULT_mult_6_net88702, MULT_mult_6_net88692, MULT_mult_6_net88655,
         MULT_mult_6_net88656, MULT_mult_6_net88638, MULT_mult_6_net88525,
         MULT_mult_6_net88455, MULT_mult_6_net88449, MULT_mult_6_net88444,
         MULT_mult_6_net88407, MULT_mult_6_net88408, MULT_mult_6_net88410,
         MULT_mult_6_net88344, MULT_mult_6_net88295, MULT_mult_6_net88296,
         MULT_mult_6_net88297, MULT_mult_6_net88206, MULT_mult_6_net88207,
         MULT_mult_6_net88208, MULT_mult_6_net88209, MULT_mult_6_net88210,
         MULT_mult_6_net88211, MULT_mult_6_net88177, MULT_mult_6_net88166,
         MULT_mult_6_net88165, MULT_mult_6_net88156, MULT_mult_6_net88157,
         MULT_mult_6_net88086, MULT_mult_6_net87874, MULT_mult_6_net87682,
         MULT_mult_6_net87683, MULT_mult_6_net87619, MULT_mult_6_net87573,
         MULT_mult_6_net87464, MULT_mult_6_net87465, MULT_mult_6_net87411,
         MULT_mult_6_net87308, MULT_mult_6_net87309, MULT_mult_6_net87310,
         MULT_mult_6_net87133, MULT_mult_6_net87136, MULT_mult_6_net87064,
         MULT_mult_6_net87045, MULT_mult_6_net87003, MULT_mult_6_net87004,
         MULT_mult_6_net87005, MULT_mult_6_net87010, MULT_mult_6_net87011,
         MULT_mult_6_net87012, MULT_mult_6_net86893, MULT_mult_6_net86894,
         MULT_mult_6_net86895, MULT_mult_6_net86896, MULT_mult_6_net86864,
         MULT_mult_6_net86844, MULT_mult_6_net86697, MULT_mult_6_net86698,
         MULT_mult_6_net86699, MULT_mult_6_net86702, MULT_mult_6_net86703,
         MULT_mult_6_net86704, MULT_mult_6_net86661, MULT_mult_6_net86662,
         MULT_mult_6_net86649, MULT_mult_6_net86651, MULT_mult_6_net86652,
         MULT_mult_6_net86653, MULT_mult_6_net86654, MULT_mult_6_net86656,
         MULT_mult_6_net86629, MULT_mult_6_net86630, MULT_mult_6_net86601,
         MULT_mult_6_net86565, MULT_mult_6_net86557, MULT_mult_6_net86464,
         MULT_mult_6_net86440, MULT_mult_6_net86427, MULT_mult_6_net86412,
         MULT_mult_6_net86413, MULT_mult_6_net86414, MULT_mult_6_net86385,
         MULT_mult_6_net86170, MULT_mult_6_net86171, MULT_mult_6_net86172,
         MULT_mult_6_net86158, MULT_mult_6_net86159, MULT_mult_6_net86101,
         MULT_mult_6_net86054, MULT_mult_6_net85979, MULT_mult_6_net85734,
         MULT_mult_6_net85732, MULT_mult_6_net85716, MULT_mult_6_net85602,
         MULT_mult_6_net85603, MULT_mult_6_net85540, MULT_mult_6_net85543,
         MULT_mult_6_net85455, MULT_mult_6_net85456, MULT_mult_6_net85457,
         MULT_mult_6_net85465, MULT_mult_6_net85469, MULT_mult_6_net85373,
         MULT_mult_6_net85325, MULT_mult_6_net85251, MULT_mult_6_net85254,
         MULT_mult_6_net85212, MULT_mult_6_net85043, MULT_mult_6_net85044,
         MULT_mult_6_net85035, MULT_mult_6_net85036, MULT_mult_6_net85017,
         MULT_mult_6_net84998, MULT_mult_6_net84999, MULT_mult_6_net85000,
         MULT_mult_6_net84947, MULT_mult_6_net84948, MULT_mult_6_net84924,
         MULT_mult_6_net84925, MULT_mult_6_net84926, MULT_mult_6_net84902,
         MULT_mult_6_net84891, MULT_mult_6_net84817, MULT_mult_6_net84818,
         MULT_mult_6_net84825, MULT_mult_6_net84826, MULT_mult_6_net84746,
         MULT_mult_6_net84706, MULT_mult_6_net84707, MULT_mult_6_net84708,
         MULT_mult_6_net84710, MULT_mult_6_net84711, MULT_mult_6_net84712,
         MULT_mult_6_net84698, MULT_mult_6_net84657, MULT_mult_6_net84481,
         MULT_mult_6_net84358, MULT_mult_6_net84348, MULT_mult_6_net84297,
         MULT_mult_6_net84298, MULT_mult_6_net84299, MULT_mult_6_net84300,
         MULT_mult_6_net84301, MULT_mult_6_net84302, MULT_mult_6_net84303,
         MULT_mult_6_net84304, MULT_mult_6_net84305, MULT_mult_6_net84308,
         MULT_mult_6_net84309, MULT_mult_6_net84209, MULT_mult_6_net84211,
         MULT_mult_6_net84212, MULT_mult_6_net84163, MULT_mult_6_net84116,
         MULT_mult_6_net84118, MULT_mult_6_net84007, MULT_mult_6_net83919,
         MULT_mult_6_net83866, MULT_mult_6_net83850, MULT_mult_6_net83796,
         MULT_mult_6_net83797, MULT_mult_6_net83784, MULT_mult_6_net83736,
         MULT_mult_6_net83535, MULT_mult_6_net83445, MULT_mult_6_net83357,
         MULT_mult_6_net83358, MULT_mult_6_net83351, MULT_mult_6_net83296,
         MULT_mult_6_net83263, MULT_mult_6_net83172, MULT_mult_6_net83174,
         MULT_mult_6_net83175, MULT_mult_6_net83151, MULT_mult_6_net83134,
         MULT_mult_6_net83120, MULT_mult_6_net83121, MULT_mult_6_net82890,
         MULT_mult_6_net82848, MULT_mult_6_net82849, MULT_mult_6_net82850,
         MULT_mult_6_net82834, MULT_mult_6_net82757, MULT_mult_6_net82759,
         MULT_mult_6_net82760, MULT_mult_6_net82723, MULT_mult_6_net82678,
         MULT_mult_6_net82664, MULT_mult_6_net82665, MULT_mult_6_net82666,
         MULT_mult_6_net82667, MULT_mult_6_net82668, MULT_mult_6_net82669,
         MULT_mult_6_net82641, MULT_mult_6_net82601, MULT_mult_6_net82550,
         MULT_mult_6_net82551, MULT_mult_6_net82556, MULT_mult_6_net82557,
         MULT_mult_6_net82558, MULT_mult_6_net82548, MULT_mult_6_net82532,
         MULT_mult_6_net82534, MULT_mult_6_net82407, MULT_mult_6_net82408,
         MULT_mult_6_net82247, MULT_mult_6_net82238, MULT_mult_6_net82239,
         MULT_mult_6_net82159, MULT_mult_6_net82154, MULT_mult_6_net82149,
         MULT_mult_6_net82099, MULT_mult_6_net82101, MULT_mult_6_net82089,
         MULT_mult_6_net82045, MULT_mult_6_net82046, MULT_mult_6_net82024,
         MULT_mult_6_net82027, MULT_mult_6_net82028, MULT_mult_6_net82029,
         MULT_mult_6_net82031, MULT_mult_6_net81995, MULT_mult_6_net81983,
         MULT_mult_6_net81958, MULT_mult_6_net81955, MULT_mult_6_net81956,
         MULT_mult_6_net81945, MULT_mult_6_net81815, MULT_mult_6_net81782,
         MULT_mult_6_net81779, MULT_mult_6_net81780, MULT_mult_6_net81781,
         MULT_mult_6_net81756, MULT_mult_6_net81713, MULT_mult_6_net81714,
         MULT_mult_6_net81673, MULT_mult_6_net81663, MULT_mult_6_net81615,
         MULT_mult_6_net81616, MULT_mult_6_net81617, MULT_mult_6_net81586,
         MULT_mult_6_net81581, MULT_mult_6_net81548, MULT_mult_6_net81513,
         MULT_mult_6_net81514, MULT_mult_6_net81515, MULT_mult_6_net81530,
         MULT_mult_6_net81531, MULT_mult_6_net81533, MULT_mult_6_net81535,
         MULT_mult_6_net81493, MULT_mult_6_net81491, MULT_mult_6_net81431,
         MULT_mult_6_net81424, MULT_mult_6_net81365, MULT_mult_6_net81367,
         MULT_mult_6_net81354, MULT_mult_6_net81258, MULT_mult_6_net81259,
         MULT_mult_6_net81260, MULT_mult_6_net81261, MULT_mult_6_net81262,
         MULT_mult_6_net81265, MULT_mult_6_net81266, MULT_mult_6_net81267,
         MULT_mult_6_net81211, MULT_mult_6_net81212, MULT_mult_6_net81213,
         MULT_mult_6_net81204, MULT_mult_6_net81205, MULT_mult_6_net81206,
         MULT_mult_6_net81169, MULT_mult_6_net81178, MULT_mult_6_net81179,
         MULT_mult_6_net81180, MULT_mult_6_net81110, MULT_mult_6_net81111,
         MULT_mult_6_net81112, MULT_mult_6_net81080, MULT_mult_6_net81052,
         MULT_mult_6_net81053, MULT_mult_6_net81056, MULT_mult_6_net81057,
         MULT_mult_6_net81058, MULT_mult_6_net81059, MULT_mult_6_net81060,
         MULT_mult_6_net81065, MULT_mult_6_net81066, MULT_mult_6_net81067,
         MULT_mult_6_net81068, MULT_mult_6_net81069, MULT_mult_6_net81033,
         MULT_mult_6_net81034, MULT_mult_6_net81035, MULT_mult_6_net81036,
         MULT_mult_6_net81037, MULT_mult_6_net81038, MULT_mult_6_net80990,
         MULT_mult_6_net80991, MULT_mult_6_net80992, MULT_mult_6_net80993,
         MULT_mult_6_net80983, MULT_mult_6_net80940, MULT_mult_6_net80941,
         MULT_mult_6_net80942, MULT_mult_6_net80956, MULT_mult_6_net80957,
         MULT_mult_6_net80958, MULT_mult_6_net80920, MULT_mult_6_net80921,
         MULT_mult_6_net80922, MULT_mult_6_net80924, MULT_mult_6_net80925,
         MULT_mult_6_net80926, MULT_mult_6_net80879, MULT_mult_6_net80880,
         MULT_mult_6_net80835, MULT_mult_6_net80836, MULT_mult_6_net80838,
         MULT_mult_6_net80839, MULT_mult_6_net80840, MULT_mult_6_net80844,
         MULT_mult_6_net80845, MULT_mult_6_net80850, MULT_mult_6_net80852,
         MULT_mult_6_net80805, MULT_mult_6_net80806, MULT_mult_6_net80812,
         MULT_mult_6_net80813, MULT_mult_6_net80814, MULT_mult_6_net80816,
         MULT_mult_6_net80817, MULT_mult_6_net80818, MULT_mult_6_net80791,
         MULT_mult_6_net80792, MULT_mult_6_net80793, MULT_mult_6_net80795,
         MULT_mult_6_net80796, MULT_mult_6_net80767, MULT_mult_6_net80768,
         MULT_mult_6_net80769, MULT_mult_6_net80727, MULT_mult_6_net80694,
         MULT_mult_6_net80671, MULT_mult_6_net80672, MULT_mult_6_net80673,
         MULT_mult_6_net80674, MULT_mult_6_net80675, MULT_mult_6_net80676,
         MULT_mult_6_net80643, MULT_mult_6_net80561, MULT_mult_6_net80562,
         MULT_mult_6_net80563, MULT_mult_6_net80565, MULT_mult_6_net80566,
         MULT_mult_6_net80518, MULT_mult_6_net80519, MULT_mult_6_net80520,
         MULT_mult_6_net80521, MULT_mult_6_net80522, MULT_mult_6_net80523,
         MULT_mult_6_net80510, MULT_mult_6_net80478, MULT_mult_6_net80479,
         MULT_mult_6_net80480, MULT_mult_6_net80449, MULT_mult_6_net80451,
         MULT_mult_6_net80409, MULT_mult_6_net80392, MULT_mult_6_net80348,
         MULT_mult_6_net80349, MULT_mult_6_net80350, MULT_mult_6_net80355,
         MULT_mult_6_net80356, MULT_mult_6_net80264, MULT_mult_6_net80273,
         MULT_mult_6_net80274, MULT_mult_6_net80275, MULT_mult_6_net80246,
         MULT_mult_6_net80247, MULT_mult_6_net80248, MULT_mult_6_net80254,
         MULT_mult_6_net80255, MULT_mult_6_net80258, MULT_mult_6_net79992,
         MULT_mult_6_net79993, MULT_mult_6_net79968, MULT_mult_6_net79969,
         MULT_mult_6_net79970, MULT_mult_6_net79951, MULT_mult_6_net79952,
         MULT_mult_6_net79953, MULT_mult_6_net79955, MULT_mult_6_net79956,
         MULT_mult_6_net79957, MULT_mult_6_net79959, MULT_mult_6_net79960,
         MULT_mult_6_net79961, MULT_mult_6_net79935, MULT_mult_6_net79936,
         MULT_mult_6_net79937, MULT_mult_6_net79939, MULT_mult_6_net79891,
         MULT_mult_6_net79892, MULT_mult_6_net79893, MULT_mult_6_net79904,
         MULT_mult_6_net79905, MULT_mult_6_net79906,
         MULT_mult_6__UDW__112739_net78703, MULT_mult_6__UDW__112704_net78605,
         MULT_mult_6__UDW__112694_net78575, MULT_mult_6__UDW__112684_net78547,
         MULT_mult_6__UDW__112679_net78533, MULT_mult_6_net77970,
         MULT_mult_6_net77964, MULT_mult_6_net77966, MULT_mult_6_net77956,
         MULT_mult_6_net77946, MULT_mult_6_net77948, MULT_mult_6_net77938,
         MULT_mult_6_net77940, MULT_mult_6_net77930, MULT_mult_6_net77932,
         MULT_mult_6_net77924, MULT_mult_6_net77926, MULT_mult_6_net77920,
         MULT_mult_6_net77912, MULT_mult_6_net77914, MULT_mult_6_net77906,
         MULT_mult_6_net77908, MULT_mult_6_net77898, MULT_mult_6_net77900,
         MULT_mult_6_net77892, MULT_mult_6_net77882, MULT_mult_6_net77886,
         MULT_mult_6_net77878, MULT_mult_6_net77866, MULT_mult_6_net77868,
         MULT_mult_6_net77858, MULT_mult_6_net77860, MULT_mult_6_net70492,
         MULT_mult_6_net70491, MULT_mult_6_net70486, MULT_mult_6_net70482,
         MULT_mult_6_net70478, MULT_mult_6_net70477, MULT_mult_6_net70476,
         MULT_mult_6_net70475, MULT_mult_6_net70474, MULT_mult_6_net70473,
         MULT_mult_6_net70472, MULT_mult_6_net70471, MULT_mult_6_net70470,
         MULT_mult_6_net70469, MULT_mult_6_net70467, MULT_mult_6_net70465,
         MULT_mult_6_net70463, MULT_mult_6_net70461, MULT_mult_6_net70460,
         MULT_mult_6_net70459, MULT_mult_6_net70457, MULT_mult_6_net70456,
         MULT_mult_6_net70455, MULT_mult_6_net70454, MULT_mult_6_net70453,
         MULT_mult_6_net70452, MULT_mult_6_net70451, MULT_mult_6_net70449,
         MULT_mult_6_net70447, MULT_mult_6_net70445, MULT_mult_6_net70443,
         MULT_mult_6_net70441, MULT_mult_6_net70435, MULT_mult_6_SUMB_16__2_,
         MULT_mult_6_SUMB_16__3_, MULT_mult_6_SUMB_16__4_,
         MULT_mult_6_SUMB_16__5_, MULT_mult_6_SUMB_16__6_,
         MULT_mult_6_SUMB_16__8_, MULT_mult_6_SUMB_16__9_,
         MULT_mult_6_SUMB_16__11_, MULT_mult_6_SUMB_16__12_,
         MULT_mult_6_SUMB_16__14_, MULT_mult_6_SUMB_17__1_,
         MULT_mult_6_SUMB_17__3_, MULT_mult_6_SUMB_17__4_,
         MULT_mult_6_SUMB_17__5_, MULT_mult_6_SUMB_17__10_,
         MULT_mult_6_SUMB_17__11_, MULT_mult_6_SUMB_17__13_,
         MULT_mult_6_SUMB_17__14_, MULT_mult_6_SUMB_18__1_,
         MULT_mult_6_SUMB_18__3_, MULT_mult_6_SUMB_18__4_,
         MULT_mult_6_SUMB_18__5_, MULT_mult_6_SUMB_18__8_,
         MULT_mult_6_SUMB_18__12_, MULT_mult_6_SUMB_19__1_,
         MULT_mult_6_SUMB_19__2_, MULT_mult_6_SUMB_19__3_,
         MULT_mult_6_SUMB_19__4_, MULT_mult_6_SUMB_19__5_,
         MULT_mult_6_SUMB_19__11_, MULT_mult_6_SUMB_20__1_,
         MULT_mult_6_SUMB_20__2_, MULT_mult_6_SUMB_20__3_,
         MULT_mult_6_SUMB_20__4_, MULT_mult_6_SUMB_20__8_,
         MULT_mult_6_SUMB_20__10_, MULT_mult_6_SUMB_20__11_,
         MULT_mult_6_SUMB_21__1_, MULT_mult_6_SUMB_21__2_,
         MULT_mult_6_SUMB_21__3_, MULT_mult_6_SUMB_21__4_,
         MULT_mult_6_SUMB_21__7_, MULT_mult_6_SUMB_21__9_,
         MULT_mult_6_SUMB_21__10_, MULT_mult_6_SUMB_22__1_,
         MULT_mult_6_SUMB_22__3_, MULT_mult_6_SUMB_22__7_,
         MULT_mult_6_SUMB_22__9_, MULT_mult_6_SUMB_23__1_,
         MULT_mult_6_SUMB_23__6_, MULT_mult_6_SUMB_23__8_,
         MULT_mult_6_SUMB_24__5_, MULT_mult_6_SUMB_25__4_,
         MULT_mult_6_SUMB_25__5_, MULT_mult_6_SUMB_26__1_,
         MULT_mult_6_SUMB_26__4_, MULT_mult_6_CARRYB_16__0_,
         MULT_mult_6_CARRYB_16__2_, MULT_mult_6_CARRYB_16__3_,
         MULT_mult_6_CARRYB_16__5_, MULT_mult_6_CARRYB_16__7_,
         MULT_mult_6_CARRYB_16__8_, MULT_mult_6_CARRYB_16__11_,
         MULT_mult_6_CARRYB_16__13_, MULT_mult_6_CARRYB_16__14_,
         MULT_mult_6_CARRYB_17__0_, MULT_mult_6_CARRYB_17__2_,
         MULT_mult_6_CARRYB_17__3_, MULT_mult_6_CARRYB_17__4_,
         MULT_mult_6_CARRYB_17__5_, MULT_mult_6_CARRYB_17__9_,
         MULT_mult_6_CARRYB_17__10_, MULT_mult_6_CARRYB_17__13_,
         MULT_mult_6_CARRYB_18__0_, MULT_mult_6_CARRYB_18__2_,
         MULT_mult_6_CARRYB_18__3_, MULT_mult_6_CARRYB_18__4_,
         MULT_mult_6_CARRYB_18__5_, MULT_mult_6_CARRYB_18__7_,
         MULT_mult_6_CARRYB_18__8_, MULT_mult_6_CARRYB_18__9_,
         MULT_mult_6_CARRYB_18__11_, MULT_mult_6_CARRYB_18__12_,
         MULT_mult_6_CARRYB_19__0_, MULT_mult_6_CARRYB_19__2_,
         MULT_mult_6_CARRYB_19__3_, MULT_mult_6_CARRYB_19__4_,
         MULT_mult_6_CARRYB_19__6_, MULT_mult_6_CARRYB_19__7_,
         MULT_mult_6_CARRYB_19__8_, MULT_mult_6_CARRYB_19__10_,
         MULT_mult_6_CARRYB_19__11_, MULT_mult_6_CARRYB_20__0_,
         MULT_mult_6_CARRYB_20__1_, MULT_mult_6_CARRYB_20__2_,
         MULT_mult_6_CARRYB_20__4_, MULT_mult_6_CARRYB_20__6_,
         MULT_mult_6_CARRYB_20__7_, MULT_mult_6_CARRYB_20__9_,
         MULT_mult_6_CARRYB_20__10_, MULT_mult_6_CARRYB_21__0_,
         MULT_mult_6_CARRYB_21__1_, MULT_mult_6_CARRYB_21__2_,
         MULT_mult_6_CARRYB_21__4_, MULT_mult_6_CARRYB_21__6_,
         MULT_mult_6_CARRYB_21__8_, MULT_mult_6_CARRYB_21__9_,
         MULT_mult_6_CARRYB_22__0_, MULT_mult_6_CARRYB_22__2_,
         MULT_mult_6_CARRYB_22__4_, MULT_mult_6_CARRYB_22__6_,
         MULT_mult_6_CARRYB_22__8_, MULT_mult_6_CARRYB_23__0_,
         MULT_mult_6_CARRYB_23__2_, MULT_mult_6_CARRYB_23__5_,
         MULT_mult_6_CARRYB_23__6_, MULT_mult_6_CARRYB_23__7_,
         MULT_mult_6_CARRYB_24__0_, MULT_mult_6_CARRYB_24__1_,
         MULT_mult_6_CARRYB_24__4_, MULT_mult_6_CARRYB_24__5_,
         MULT_mult_6_CARRYB_25__0_, MULT_mult_6_CARRYB_25__2_,
         MULT_mult_6_CARRYB_25__3_, MULT_mult_6_CARRYB_25__4_,
         MULT_mult_6_CARRYB_26__0_, MULT_mult_6_CARRYB_26__3_,
         MULT_mult_6_CARRYB_27__1_, MULT_mult_6_CARRYB_27__2_,
         MULT_mult_6_SUMB_1__2_, MULT_mult_6_SUMB_1__3_,
         MULT_mult_6_SUMB_1__4_, MULT_mult_6_SUMB_1__5_,
         MULT_mult_6_SUMB_1__6_, MULT_mult_6_SUMB_1__9_,
         MULT_mult_6_SUMB_1__10_, MULT_mult_6_SUMB_1__11_,
         MULT_mult_6_SUMB_1__12_, MULT_mult_6_SUMB_1__13_,
         MULT_mult_6_SUMB_1__16_, MULT_mult_6_SUMB_1__19_,
         MULT_mult_6_SUMB_1__20_, MULT_mult_6_SUMB_1__21_,
         MULT_mult_6_SUMB_1__23_, MULT_mult_6_SUMB_1__26_,
         MULT_mult_6_SUMB_1__27_, MULT_mult_6_SUMB_1__28_,
         MULT_mult_6_SUMB_1__29_, MULT_mult_6_SUMB_2__1_,
         MULT_mult_6_SUMB_2__2_, MULT_mult_6_SUMB_2__3_,
         MULT_mult_6_SUMB_2__4_, MULT_mult_6_SUMB_2__5_,
         MULT_mult_6_SUMB_2__6_, MULT_mult_6_SUMB_2__8_,
         MULT_mult_6_SUMB_2__9_, MULT_mult_6_SUMB_2__10_,
         MULT_mult_6_SUMB_2__11_, MULT_mult_6_SUMB_2__12_,
         MULT_mult_6_SUMB_2__13_, MULT_mult_6_SUMB_2__14_,
         MULT_mult_6_SUMB_2__15_, MULT_mult_6_SUMB_2__18_,
         MULT_mult_6_SUMB_2__19_, MULT_mult_6_SUMB_2__20_,
         MULT_mult_6_SUMB_2__21_, MULT_mult_6_SUMB_2__22_,
         MULT_mult_6_SUMB_2__23_, MULT_mult_6_SUMB_2__25_,
         MULT_mult_6_SUMB_2__26_, MULT_mult_6_SUMB_2__27_,
         MULT_mult_6_SUMB_2__28_, MULT_mult_6_SUMB_2__29_,
         MULT_mult_6_SUMB_3__1_, MULT_mult_6_SUMB_3__2_,
         MULT_mult_6_SUMB_3__3_, MULT_mult_6_SUMB_3__4_,
         MULT_mult_6_SUMB_3__5_, MULT_mult_6_SUMB_3__7_,
         MULT_mult_6_SUMB_3__8_, MULT_mult_6_SUMB_3__9_,
         MULT_mult_6_SUMB_3__10_, MULT_mult_6_SUMB_3__11_,
         MULT_mult_6_SUMB_3__12_, MULT_mult_6_SUMB_3__14_,
         MULT_mult_6_SUMB_3__15_, MULT_mult_6_SUMB_3__18_,
         MULT_mult_6_SUMB_3__19_, MULT_mult_6_SUMB_3__20_,
         MULT_mult_6_SUMB_3__21_, MULT_mult_6_SUMB_3__22_,
         MULT_mult_6_SUMB_3__24_, MULT_mult_6_SUMB_3__25_,
         MULT_mult_6_SUMB_3__26_, MULT_mult_6_SUMB_3__27_,
         MULT_mult_6_SUMB_3__28_, MULT_mult_6_SUMB_4__1_,
         MULT_mult_6_SUMB_4__2_, MULT_mult_6_SUMB_4__3_,
         MULT_mult_6_SUMB_4__4_, MULT_mult_6_SUMB_4__5_,
         MULT_mult_6_SUMB_4__7_, MULT_mult_6_SUMB_4__8_,
         MULT_mult_6_SUMB_4__9_, MULT_mult_6_SUMB_4__10_,
         MULT_mult_6_SUMB_4__11_, MULT_mult_6_SUMB_4__13_,
         MULT_mult_6_SUMB_4__14_, MULT_mult_6_SUMB_4__17_,
         MULT_mult_6_SUMB_4__18_, MULT_mult_6_SUMB_4__19_,
         MULT_mult_6_SUMB_4__20_, MULT_mult_6_SUMB_4__21_,
         MULT_mult_6_SUMB_4__22_, MULT_mult_6_SUMB_4__24_,
         MULT_mult_6_SUMB_4__26_, MULT_mult_6_SUMB_4__27_,
         MULT_mult_6_SUMB_5__1_, MULT_mult_6_SUMB_5__2_,
         MULT_mult_6_SUMB_5__3_, MULT_mult_6_SUMB_5__4_,
         MULT_mult_6_SUMB_5__6_, MULT_mult_6_SUMB_5__7_,
         MULT_mult_6_SUMB_5__8_, MULT_mult_6_SUMB_5__9_,
         MULT_mult_6_SUMB_5__10_, MULT_mult_6_SUMB_5__11_,
         MULT_mult_6_SUMB_5__13_, MULT_mult_6_SUMB_5__14_,
         MULT_mult_6_SUMB_5__16_, MULT_mult_6_SUMB_5__17_,
         MULT_mult_6_SUMB_5__18_, MULT_mult_6_SUMB_5__19_,
         MULT_mult_6_SUMB_5__20_, MULT_mult_6_SUMB_5__21_,
         MULT_mult_6_SUMB_5__23_, MULT_mult_6_SUMB_5__24_,
         MULT_mult_6_SUMB_5__25_, MULT_mult_6_SUMB_5__26_,
         MULT_mult_6_SUMB_6__1_, MULT_mult_6_SUMB_6__2_,
         MULT_mult_6_SUMB_6__3_, MULT_mult_6_SUMB_6__4_,
         MULT_mult_6_SUMB_6__6_, MULT_mult_6_SUMB_6__7_,
         MULT_mult_6_SUMB_6__8_, MULT_mult_6_SUMB_6__9_,
         MULT_mult_6_SUMB_6__10_, MULT_mult_6_SUMB_6__11_,
         MULT_mult_6_SUMB_6__13_, MULT_mult_6_SUMB_6__15_,
         MULT_mult_6_SUMB_6__16_, MULT_mult_6_SUMB_6__17_,
         MULT_mult_6_SUMB_6__19_, MULT_mult_6_SUMB_6__20_,
         MULT_mult_6_SUMB_6__22_, MULT_mult_6_SUMB_6__23_,
         MULT_mult_6_SUMB_6__24_, MULT_mult_6_SUMB_6__25_,
         MULT_mult_6_SUMB_7__1_, MULT_mult_6_SUMB_7__2_,
         MULT_mult_6_SUMB_7__3_, MULT_mult_6_SUMB_7__7_,
         MULT_mult_6_SUMB_7__8_, MULT_mult_6_SUMB_7__9_,
         MULT_mult_6_SUMB_7__10_, MULT_mult_6_SUMB_7__12_,
         MULT_mult_6_SUMB_7__14_, MULT_mult_6_SUMB_7__15_,
         MULT_mult_6_SUMB_7__16_, MULT_mult_6_SUMB_7__17_,
         MULT_mult_6_SUMB_7__19_, MULT_mult_6_SUMB_7__21_,
         MULT_mult_6_SUMB_7__22_, MULT_mult_6_SUMB_7__23_,
         MULT_mult_6_SUMB_7__24_, MULT_mult_6_SUMB_8__1_,
         MULT_mult_6_SUMB_8__2_, MULT_mult_6_SUMB_8__5_,
         MULT_mult_6_SUMB_8__6_, MULT_mult_6_SUMB_8__7_,
         MULT_mult_6_SUMB_8__8_, MULT_mult_6_SUMB_8__9_,
         MULT_mult_6_SUMB_8__10_, MULT_mult_6_SUMB_8__15_,
         MULT_mult_6_SUMB_8__16_, MULT_mult_6_SUMB_8__20_,
         MULT_mult_6_SUMB_8__21_, MULT_mult_6_SUMB_8__22_,
         MULT_mult_6_SUMB_8__23_, MULT_mult_6_SUMB_9__1_,
         MULT_mult_6_SUMB_9__2_, MULT_mult_6_SUMB_9__4_,
         MULT_mult_6_SUMB_9__5_, MULT_mult_6_SUMB_9__6_,
         MULT_mult_6_SUMB_9__7_, MULT_mult_6_SUMB_9__8_,
         MULT_mult_6_SUMB_9__9_, MULT_mult_6_SUMB_9__10_,
         MULT_mult_6_SUMB_9__12_, MULT_mult_6_SUMB_9__14_,
         MULT_mult_6_SUMB_9__15_, MULT_mult_6_SUMB_9__16_,
         MULT_mult_6_SUMB_9__19_, MULT_mult_6_SUMB_9__20_,
         MULT_mult_6_SUMB_9__21_, MULT_mult_6_SUMB_9__22_,
         MULT_mult_6_SUMB_10__1_, MULT_mult_6_SUMB_10__2_,
         MULT_mult_6_SUMB_10__4_, MULT_mult_6_SUMB_10__5_,
         MULT_mult_6_SUMB_10__6_, MULT_mult_6_SUMB_10__7_,
         MULT_mult_6_SUMB_10__8_, MULT_mult_6_SUMB_10__9_,
         MULT_mult_6_SUMB_10__12_, MULT_mult_6_SUMB_10__14_,
         MULT_mult_6_SUMB_10__15_, MULT_mult_6_SUMB_10__16_,
         MULT_mult_6_SUMB_10__18_, MULT_mult_6_SUMB_10__19_,
         MULT_mult_6_SUMB_10__20_, MULT_mult_6_SUMB_10__21_,
         MULT_mult_6_SUMB_11__1_, MULT_mult_6_SUMB_11__3_,
         MULT_mult_6_SUMB_11__4_, MULT_mult_6_SUMB_11__5_,
         MULT_mult_6_SUMB_11__6_, MULT_mult_6_SUMB_11__7_,
         MULT_mult_6_SUMB_11__8_, MULT_mult_6_SUMB_11__10_,
         MULT_mult_6_SUMB_11__13_, MULT_mult_6_SUMB_11__14_,
         MULT_mult_6_SUMB_11__15_, MULT_mult_6_SUMB_11__17_,
         MULT_mult_6_SUMB_11__18_, MULT_mult_6_SUMB_11__19_,
         MULT_mult_6_SUMB_11__20_, MULT_mult_6_SUMB_12__3_,
         MULT_mult_6_SUMB_12__4_, MULT_mult_6_SUMB_12__5_,
         MULT_mult_6_SUMB_12__6_, MULT_mult_6_SUMB_12__7_,
         MULT_mult_6_SUMB_12__8_, MULT_mult_6_SUMB_12__11_,
         MULT_mult_6_SUMB_12__12_, MULT_mult_6_SUMB_12__13_,
         MULT_mult_6_SUMB_12__14_, MULT_mult_6_SUMB_12__15_,
         MULT_mult_6_SUMB_12__16_, MULT_mult_6_SUMB_12__17_,
         MULT_mult_6_SUMB_12__18_, MULT_mult_6_SUMB_12__19_,
         MULT_mult_6_SUMB_13__1_, MULT_mult_6_SUMB_13__2_,
         MULT_mult_6_SUMB_13__4_, MULT_mult_6_SUMB_13__5_,
         MULT_mult_6_SUMB_13__6_, MULT_mult_6_SUMB_13__7_,
         MULT_mult_6_SUMB_13__8_, MULT_mult_6_SUMB_13__10_,
         MULT_mult_6_SUMB_13__12_, MULT_mult_6_SUMB_13__13_,
         MULT_mult_6_SUMB_13__14_, MULT_mult_6_SUMB_13__16_,
         MULT_mult_6_SUMB_13__17_, MULT_mult_6_SUMB_13__18_,
         MULT_mult_6_SUMB_14__1_, MULT_mult_6_SUMB_14__3_,
         MULT_mult_6_SUMB_14__4_, MULT_mult_6_SUMB_14__5_,
         MULT_mult_6_SUMB_14__6_, MULT_mult_6_SUMB_14__7_,
         MULT_mult_6_SUMB_14__12_, MULT_mult_6_SUMB_14__13_,
         MULT_mult_6_SUMB_14__15_, MULT_mult_6_SUMB_14__16_,
         MULT_mult_6_SUMB_14__17_, MULT_mult_6_SUMB_15__3_,
         MULT_mult_6_SUMB_15__4_, MULT_mult_6_SUMB_15__5_,
         MULT_mult_6_SUMB_15__6_, MULT_mult_6_SUMB_15__9_,
         MULT_mult_6_SUMB_15__12_, MULT_mult_6_SUMB_15__13_,
         MULT_mult_6_SUMB_15__15_, MULT_mult_6_CARRYB_1__0_,
         MULT_mult_6_CARRYB_1__2_, MULT_mult_6_CARRYB_1__3_,
         MULT_mult_6_CARRYB_1__4_, MULT_mult_6_CARRYB_1__5_,
         MULT_mult_6_CARRYB_1__9_, MULT_mult_6_CARRYB_1__10_,
         MULT_mult_6_CARRYB_1__11_, MULT_mult_6_CARRYB_1__12_,
         MULT_mult_6_CARRYB_1__15_, MULT_mult_6_CARRYB_1__18_,
         MULT_mult_6_CARRYB_1__19_, MULT_mult_6_CARRYB_1__20_,
         MULT_mult_6_CARRYB_1__21_, MULT_mult_6_CARRYB_1__22_,
         MULT_mult_6_CARRYB_1__26_, MULT_mult_6_CARRYB_2__0_,
         MULT_mult_6_CARRYB_2__1_, MULT_mult_6_CARRYB_2__2_,
         MULT_mult_6_CARRYB_2__3_, MULT_mult_6_CARRYB_2__4_,
         MULT_mult_6_CARRYB_2__5_, MULT_mult_6_CARRYB_2__8_,
         MULT_mult_6_CARRYB_2__9_, MULT_mult_6_CARRYB_2__10_,
         MULT_mult_6_CARRYB_2__11_, MULT_mult_6_CARRYB_2__14_,
         MULT_mult_6_CARRYB_2__15_, MULT_mult_6_CARRYB_2__17_,
         MULT_mult_6_CARRYB_2__18_, MULT_mult_6_CARRYB_2__19_,
         MULT_mult_6_CARRYB_2__20_, MULT_mult_6_CARRYB_2__21_,
         MULT_mult_6_CARRYB_2__22_, MULT_mult_6_CARRYB_2__24_,
         MULT_mult_6_CARRYB_2__25_, MULT_mult_6_CARRYB_2__26_,
         MULT_mult_6_CARRYB_2__27_, MULT_mult_6_CARRYB_2__28_,
         MULT_mult_6_CARRYB_3__0_, MULT_mult_6_CARRYB_3__1_,
         MULT_mult_6_CARRYB_3__2_, MULT_mult_6_CARRYB_3__3_,
         MULT_mult_6_CARRYB_3__4_, MULT_mult_6_CARRYB_3__6_,
         MULT_mult_6_CARRYB_3__7_, MULT_mult_6_CARRYB_3__8_,
         MULT_mult_6_CARRYB_3__9_, MULT_mult_6_CARRYB_3__10_,
         MULT_mult_6_CARRYB_3__11_, MULT_mult_6_CARRYB_3__13_,
         MULT_mult_6_CARRYB_3__14_, MULT_mult_6_CARRYB_3__17_,
         MULT_mult_6_CARRYB_3__18_, MULT_mult_6_CARRYB_3__19_,
         MULT_mult_6_CARRYB_3__20_, MULT_mult_6_CARRYB_3__21_,
         MULT_mult_6_CARRYB_3__23_, MULT_mult_6_CARRYB_3__24_,
         MULT_mult_6_CARRYB_3__25_, MULT_mult_6_CARRYB_3__26_,
         MULT_mult_6_CARRYB_3__27_, MULT_mult_6_CARRYB_4__0_,
         MULT_mult_6_CARRYB_4__1_, MULT_mult_6_CARRYB_4__2_,
         MULT_mult_6_CARRYB_4__3_, MULT_mult_6_CARRYB_4__4_,
         MULT_mult_6_CARRYB_4__6_, MULT_mult_6_CARRYB_4__7_,
         MULT_mult_6_CARRYB_4__8_, MULT_mult_6_CARRYB_4__9_,
         MULT_mult_6_CARRYB_4__10_, MULT_mult_6_CARRYB_4__12_,
         MULT_mult_6_CARRYB_4__13_, MULT_mult_6_CARRYB_4__16_,
         MULT_mult_6_CARRYB_4__17_, MULT_mult_6_CARRYB_4__18_,
         MULT_mult_6_CARRYB_4__19_, MULT_mult_6_CARRYB_4__20_,
         MULT_mult_6_CARRYB_4__21_, MULT_mult_6_CARRYB_4__23_,
         MULT_mult_6_CARRYB_4__24_, MULT_mult_6_CARRYB_4__25_,
         MULT_mult_6_CARRYB_4__26_, MULT_mult_6_CARRYB_5__0_,
         MULT_mult_6_CARRYB_5__1_, MULT_mult_6_CARRYB_5__2_,
         MULT_mult_6_CARRYB_5__3_, MULT_mult_6_CARRYB_5__4_,
         MULT_mult_6_CARRYB_5__5_, MULT_mult_6_CARRYB_5__6_,
         MULT_mult_6_CARRYB_5__7_, MULT_mult_6_CARRYB_5__8_,
         MULT_mult_6_CARRYB_5__9_, MULT_mult_6_CARRYB_5__10_,
         MULT_mult_6_CARRYB_5__12_, MULT_mult_6_CARRYB_5__13_,
         MULT_mult_6_CARRYB_5__15_, MULT_mult_6_CARRYB_5__16_,
         MULT_mult_6_CARRYB_5__17_, MULT_mult_6_CARRYB_5__18_,
         MULT_mult_6_CARRYB_5__19_, MULT_mult_6_CARRYB_5__20_,
         MULT_mult_6_CARRYB_5__22_, MULT_mult_6_CARRYB_5__23_,
         MULT_mult_6_CARRYB_5__24_, MULT_mult_6_CARRYB_5__25_,
         MULT_mult_6_CARRYB_6__0_, MULT_mult_6_CARRYB_6__1_,
         MULT_mult_6_CARRYB_6__2_, MULT_mult_6_CARRYB_6__3_,
         MULT_mult_6_CARRYB_6__5_, MULT_mult_6_CARRYB_6__6_,
         MULT_mult_6_CARRYB_6__7_, MULT_mult_6_CARRYB_6__9_,
         MULT_mult_6_CARRYB_6__10_, MULT_mult_6_CARRYB_6__12_,
         MULT_mult_6_CARRYB_6__13_, MULT_mult_6_CARRYB_6__15_,
         MULT_mult_6_CARRYB_6__16_, MULT_mult_6_CARRYB_6__17_,
         MULT_mult_6_CARRYB_6__18_, MULT_mult_6_CARRYB_6__19_,
         MULT_mult_6_CARRYB_6__22_, MULT_mult_6_CARRYB_6__23_,
         MULT_mult_6_CARRYB_6__24_, MULT_mult_6_CARRYB_7__0_,
         MULT_mult_6_CARRYB_7__1_, MULT_mult_6_CARRYB_7__2_,
         MULT_mult_6_CARRYB_7__5_, MULT_mult_6_CARRYB_7__6_,
         MULT_mult_6_CARRYB_7__7_, MULT_mult_6_CARRYB_7__8_,
         MULT_mult_6_CARRYB_7__9_, MULT_mult_6_CARRYB_7__11_,
         MULT_mult_6_CARRYB_7__13_, MULT_mult_6_CARRYB_7__14_,
         MULT_mult_6_CARRYB_7__15_, MULT_mult_6_CARRYB_7__16_,
         MULT_mult_6_CARRYB_7__20_, MULT_mult_6_CARRYB_7__21_,
         MULT_mult_6_CARRYB_7__22_, MULT_mult_6_CARRYB_7__23_,
         MULT_mult_6_CARRYB_8__0_, MULT_mult_6_CARRYB_8__1_,
         MULT_mult_6_CARRYB_8__2_, MULT_mult_6_CARRYB_8__5_,
         MULT_mult_6_CARRYB_8__6_, MULT_mult_6_CARRYB_8__7_,
         MULT_mult_6_CARRYB_8__8_, MULT_mult_6_CARRYB_8__9_,
         MULT_mult_6_CARRYB_8__11_, MULT_mult_6_CARRYB_8__14_,
         MULT_mult_6_CARRYB_8__15_, MULT_mult_6_CARRYB_8__16_,
         MULT_mult_6_CARRYB_8__19_, MULT_mult_6_CARRYB_8__20_,
         MULT_mult_6_CARRYB_8__21_, MULT_mult_6_CARRYB_8__22_,
         MULT_mult_6_CARRYB_9__0_, MULT_mult_6_CARRYB_9__1_,
         MULT_mult_6_CARRYB_9__3_, MULT_mult_6_CARRYB_9__4_,
         MULT_mult_6_CARRYB_9__5_, MULT_mult_6_CARRYB_9__6_,
         MULT_mult_6_CARRYB_9__7_, MULT_mult_6_CARRYB_9__8_,
         MULT_mult_6_CARRYB_9__9_, MULT_mult_6_CARRYB_9__11_,
         MULT_mult_6_CARRYB_9__13_, MULT_mult_6_CARRYB_9__14_,
         MULT_mult_6_CARRYB_9__15_, MULT_mult_6_CARRYB_9__16_,
         MULT_mult_6_CARRYB_9__18_, MULT_mult_6_CARRYB_9__19_,
         MULT_mult_6_CARRYB_9__20_, MULT_mult_6_CARRYB_9__21_,
         MULT_mult_6_CARRYB_10__0_, MULT_mult_6_CARRYB_10__1_,
         MULT_mult_6_CARRYB_10__3_, MULT_mult_6_CARRYB_10__4_,
         MULT_mult_6_CARRYB_10__5_, MULT_mult_6_CARRYB_10__6_,
         MULT_mult_6_CARRYB_10__7_, MULT_mult_6_CARRYB_10__8_,
         MULT_mult_6_CARRYB_10__10_, MULT_mult_6_CARRYB_10__13_,
         MULT_mult_6_CARRYB_10__14_, MULT_mult_6_CARRYB_10__15_,
         MULT_mult_6_CARRYB_10__16_, MULT_mult_6_CARRYB_10__17_,
         MULT_mult_6_CARRYB_10__18_, MULT_mult_6_CARRYB_10__19_,
         MULT_mult_6_CARRYB_10__20_, MULT_mult_6_CARRYB_11__0_,
         MULT_mult_6_CARRYB_11__2_, MULT_mult_6_CARRYB_11__3_,
         MULT_mult_6_CARRYB_11__4_, MULT_mult_6_CARRYB_11__5_,
         MULT_mult_6_CARRYB_11__6_, MULT_mult_6_CARRYB_11__7_,
         MULT_mult_6_CARRYB_11__9_, MULT_mult_6_CARRYB_11__12_,
         MULT_mult_6_CARRYB_11__13_, MULT_mult_6_CARRYB_11__14_,
         MULT_mult_6_CARRYB_11__16_, MULT_mult_6_CARRYB_11__17_,
         MULT_mult_6_CARRYB_11__18_, MULT_mult_6_CARRYB_11__19_,
         MULT_mult_6_CARRYB_12__0_, MULT_mult_6_CARRYB_12__2_,
         MULT_mult_6_CARRYB_12__3_, MULT_mult_6_CARRYB_12__4_,
         MULT_mult_6_CARRYB_12__5_, MULT_mult_6_CARRYB_12__6_,
         MULT_mult_6_CARRYB_12__7_, MULT_mult_6_CARRYB_12__12_,
         MULT_mult_6_CARRYB_12__13_, MULT_mult_6_CARRYB_12__15_,
         MULT_mult_6_CARRYB_12__16_, MULT_mult_6_CARRYB_12__17_,
         MULT_mult_6_CARRYB_12__18_, MULT_mult_6_CARRYB_13__0_,
         MULT_mult_6_CARRYB_13__3_, MULT_mult_6_CARRYB_13__4_,
         MULT_mult_6_CARRYB_13__5_, MULT_mult_6_CARRYB_13__6_,
         MULT_mult_6_CARRYB_13__7_, MULT_mult_6_CARRYB_13__11_,
         MULT_mult_6_CARRYB_13__12_, MULT_mult_6_CARRYB_13__13_,
         MULT_mult_6_CARRYB_13__15_, MULT_mult_6_CARRYB_13__16_,
         MULT_mult_6_CARRYB_13__17_, MULT_mult_6_CARRYB_14__0_,
         MULT_mult_6_CARRYB_14__2_, MULT_mult_6_CARRYB_14__3_,
         MULT_mult_6_CARRYB_14__4_, MULT_mult_6_CARRYB_14__5_,
         MULT_mult_6_CARRYB_14__6_, MULT_mult_6_CARRYB_14__7_,
         MULT_mult_6_CARRYB_14__9_, MULT_mult_6_CARRYB_14__11_,
         MULT_mult_6_CARRYB_14__12_, MULT_mult_6_CARRYB_14__14_,
         MULT_mult_6_CARRYB_14__15_, MULT_mult_6_CARRYB_14__16_,
         MULT_mult_6_CARRYB_15__0_, MULT_mult_6_CARRYB_15__2_,
         MULT_mult_6_CARRYB_15__3_, MULT_mult_6_CARRYB_15__5_,
         MULT_mult_6_CARRYB_15__6_, MULT_mult_6_CARRYB_15__8_,
         MULT_mult_6_CARRYB_15__11_, MULT_mult_6_CARRYB_15__12_,
         MULT_mult_6_CARRYB_15__14_, MULT_mult_6_CARRYB_15__15_,
         MULT_mult_6_ab_0__1_, MULT_mult_6_ab_0__2_, MULT_mult_6_ab_0__3_,
         MULT_mult_6_ab_0__5_, MULT_mult_6_ab_0__6_, MULT_mult_6_ab_0__9_,
         MULT_mult_6_ab_0__11_, MULT_mult_6_ab_0__12_, MULT_mult_6_ab_0__13_,
         MULT_mult_6_ab_0__20_, MULT_mult_6_ab_0__21_, MULT_mult_6_ab_0__22_,
         MULT_mult_6_ab_0__23_, MULT_mult_6_ab_0__24_, MULT_mult_6_ab_0__27_,
         MULT_mult_6_ab_0__28_, MULT_mult_6_ab_0__29_, MULT_mult_6_ab_0__30_,
         MULT_mult_6_ab_0__31_, MULT_mult_6_ab_1__0_, MULT_mult_6_ab_1__1_,
         MULT_mult_6_ab_1__2_, MULT_mult_6_ab_1__3_, MULT_mult_6_ab_1__4_,
         MULT_mult_6_ab_1__5_, MULT_mult_6_ab_1__6_, MULT_mult_6_ab_1__9_,
         MULT_mult_6_ab_1__10_, MULT_mult_6_ab_1__11_, MULT_mult_6_ab_1__18_,
         MULT_mult_6_ab_1__19_, MULT_mult_6_ab_1__20_, MULT_mult_6_ab_1__21_,
         MULT_mult_6_ab_1__25_, MULT_mult_6_ab_1__26_, MULT_mult_6_ab_1__27_,
         MULT_mult_6_ab_1__28_, MULT_mult_6_ab_1__29_, MULT_mult_6_ab_1__30_,
         MULT_mult_6_ab_2__0_, MULT_mult_6_ab_2__1_, MULT_mult_6_ab_2__2_,
         MULT_mult_6_ab_2__3_, MULT_mult_6_ab_2__4_, MULT_mult_6_ab_2__5_,
         MULT_mult_6_ab_2__8_, MULT_mult_6_ab_2__9_, MULT_mult_6_ab_2__10_,
         MULT_mult_6_ab_2__11_, MULT_mult_6_ab_2__12_, MULT_mult_6_ab_2__14_,
         MULT_mult_6_ab_2__15_, MULT_mult_6_ab_2__17_, MULT_mult_6_ab_2__18_,
         MULT_mult_6_ab_2__19_, MULT_mult_6_ab_2__20_, MULT_mult_6_ab_2__21_,
         MULT_mult_6_ab_2__22_, MULT_mult_6_ab_2__25_, MULT_mult_6_ab_2__26_,
         MULT_mult_6_ab_2__27_, MULT_mult_6_ab_2__28_, MULT_mult_6_ab_2__29_,
         MULT_mult_6_ab_3__0_, MULT_mult_6_ab_3__1_, MULT_mult_6_ab_3__2_,
         MULT_mult_6_ab_3__3_, MULT_mult_6_ab_3__4_, MULT_mult_6_ab_3__5_,
         MULT_mult_6_ab_3__6_, MULT_mult_6_ab_3__7_, MULT_mult_6_ab_3__8_,
         MULT_mult_6_ab_3__9_, MULT_mult_6_ab_3__10_, MULT_mult_6_ab_3__11_,
         MULT_mult_6_ab_3__12_, MULT_mult_6_ab_3__14_, MULT_mult_6_ab_3__17_,
         MULT_mult_6_ab_3__18_, MULT_mult_6_ab_3__19_, MULT_mult_6_ab_3__20_,
         MULT_mult_6_ab_3__21_, MULT_mult_6_ab_3__22_, MULT_mult_6_ab_3__24_,
         MULT_mult_6_ab_3__25_, MULT_mult_6_ab_3__26_, MULT_mult_6_ab_3__27_,
         MULT_mult_6_ab_3__28_, MULT_mult_6_ab_4__0_, MULT_mult_6_ab_4__1_,
         MULT_mult_6_ab_4__2_, MULT_mult_6_ab_4__3_, MULT_mult_6_ab_4__4_,
         MULT_mult_6_ab_4__5_, MULT_mult_6_ab_4__6_, MULT_mult_6_ab_4__7_,
         MULT_mult_6_ab_4__8_, MULT_mult_6_ab_4__9_, MULT_mult_6_ab_4__10_,
         MULT_mult_6_ab_4__11_, MULT_mult_6_ab_4__12_, MULT_mult_6_ab_4__13_,
         MULT_mult_6_ab_4__14_, MULT_mult_6_ab_4__17_, MULT_mult_6_ab_4__18_,
         MULT_mult_6_ab_4__19_, MULT_mult_6_ab_4__20_, MULT_mult_6_ab_4__21_,
         MULT_mult_6_ab_4__23_, MULT_mult_6_ab_4__24_, MULT_mult_6_ab_4__25_,
         MULT_mult_6_ab_4__26_, MULT_mult_6_ab_4__27_, MULT_mult_6_ab_5__0_,
         MULT_mult_6_ab_5__1_, MULT_mult_6_ab_5__2_, MULT_mult_6_ab_5__3_,
         MULT_mult_6_ab_5__4_, MULT_mult_6_ab_5__6_, MULT_mult_6_ab_5__7_,
         MULT_mult_6_ab_5__8_, MULT_mult_6_ab_5__9_, MULT_mult_6_ab_5__10_,
         MULT_mult_6_ab_5__12_, MULT_mult_6_ab_5__13_, MULT_mult_6_ab_5__16_,
         MULT_mult_6_ab_5__17_, MULT_mult_6_ab_5__18_, MULT_mult_6_ab_5__19_,
         MULT_mult_6_ab_5__20_, MULT_mult_6_ab_5__21_, MULT_mult_6_ab_5__23_,
         MULT_mult_6_ab_5__24_, MULT_mult_6_ab_5__25_, MULT_mult_6_ab_5__26_,
         MULT_mult_6_ab_6__0_, MULT_mult_6_ab_6__1_, MULT_mult_6_ab_6__2_,
         MULT_mult_6_ab_6__3_, MULT_mult_6_ab_6__4_, MULT_mult_6_ab_6__5_,
         MULT_mult_6_ab_6__6_, MULT_mult_6_ab_6__7_, MULT_mult_6_ab_6__8_,
         MULT_mult_6_ab_6__9_, MULT_mult_6_ab_6__10_, MULT_mult_6_ab_6__12_,
         MULT_mult_6_ab_6__13_, MULT_mult_6_ab_6__15_, MULT_mult_6_ab_6__16_,
         MULT_mult_6_ab_6__17_, MULT_mult_6_ab_6__18_, MULT_mult_6_ab_6__19_,
         MULT_mult_6_ab_6__20_, MULT_mult_6_ab_6__22_, MULT_mult_6_ab_6__23_,
         MULT_mult_6_ab_6__24_, MULT_mult_6_ab_6__25_, MULT_mult_6_ab_7__0_,
         MULT_mult_6_ab_7__1_, MULT_mult_6_ab_7__2_, MULT_mult_6_ab_7__3_,
         MULT_mult_6_ab_7__5_, MULT_mult_6_ab_7__6_, MULT_mult_6_ab_7__7_,
         MULT_mult_6_ab_7__8_, MULT_mult_6_ab_7__9_, MULT_mult_6_ab_7__10_,
         MULT_mult_6_ab_7__12_, MULT_mult_6_ab_7__13_, MULT_mult_6_ab_7__14_,
         MULT_mult_6_ab_7__15_, MULT_mult_6_ab_7__16_, MULT_mult_6_ab_7__17_,
         MULT_mult_6_ab_7__18_, MULT_mult_6_ab_7__19_, MULT_mult_6_ab_7__20_,
         MULT_mult_6_ab_7__21_, MULT_mult_6_ab_7__22_, MULT_mult_6_ab_7__23_,
         MULT_mult_6_ab_7__24_, MULT_mult_6_ab_8__0_, MULT_mult_6_ab_8__1_,
         MULT_mult_6_ab_8__2_, MULT_mult_6_ab_8__3_, MULT_mult_6_ab_8__5_,
         MULT_mult_6_ab_8__6_, MULT_mult_6_ab_8__7_, MULT_mult_6_ab_8__8_,
         MULT_mult_6_ab_8__9_, MULT_mult_6_ab_8__11_, MULT_mult_6_ab_8__13_,
         MULT_mult_6_ab_8__14_, MULT_mult_6_ab_8__15_, MULT_mult_6_ab_8__16_,
         MULT_mult_6_ab_8__18_, MULT_mult_6_ab_8__20_, MULT_mult_6_ab_8__21_,
         MULT_mult_6_ab_8__22_, MULT_mult_6_ab_8__23_, MULT_mult_6_ab_9__0_,
         MULT_mult_6_ab_9__1_, MULT_mult_6_ab_9__2_, MULT_mult_6_ab_9__3_,
         MULT_mult_6_ab_9__4_, MULT_mult_6_ab_9__5_, MULT_mult_6_ab_9__6_,
         MULT_mult_6_ab_9__7_, MULT_mult_6_ab_9__8_, MULT_mult_6_ab_9__9_,
         MULT_mult_6_ab_9__11_, MULT_mult_6_ab_9__14_, MULT_mult_6_ab_9__15_,
         MULT_mult_6_ab_9__16_, MULT_mult_6_ab_9__19_, MULT_mult_6_ab_9__20_,
         MULT_mult_6_ab_9__21_, MULT_mult_6_ab_9__22_, MULT_mult_6_ab_10__0_,
         MULT_mult_6_ab_10__1_, MULT_mult_6_ab_10__3_, MULT_mult_6_ab_10__4_,
         MULT_mult_6_ab_10__5_, MULT_mult_6_ab_10__6_, MULT_mult_6_ab_10__7_,
         MULT_mult_6_ab_10__8_, MULT_mult_6_ab_10__9_, MULT_mult_6_ab_10__11_,
         MULT_mult_6_ab_10__13_, MULT_mult_6_ab_10__14_,
         MULT_mult_6_ab_10__15_, MULT_mult_6_ab_10__16_,
         MULT_mult_6_ab_10__18_, MULT_mult_6_ab_10__19_,
         MULT_mult_6_ab_10__20_, MULT_mult_6_ab_10__21_, MULT_mult_6_ab_11__0_,
         MULT_mult_6_ab_11__1_, MULT_mult_6_ab_11__3_, MULT_mult_6_ab_11__4_,
         MULT_mult_6_ab_11__5_, MULT_mult_6_ab_11__6_, MULT_mult_6_ab_11__7_,
         MULT_mult_6_ab_11__8_, MULT_mult_6_ab_11__10_, MULT_mult_6_ab_11__11_,
         MULT_mult_6_ab_11__13_, MULT_mult_6_ab_11__14_,
         MULT_mult_6_ab_11__15_, MULT_mult_6_ab_11__16_,
         MULT_mult_6_ab_11__17_, MULT_mult_6_ab_11__18_,
         MULT_mult_6_ab_11__19_, MULT_mult_6_ab_11__20_, MULT_mult_6_ab_12__0_,
         MULT_mult_6_ab_12__2_, MULT_mult_6_ab_12__3_, MULT_mult_6_ab_12__4_,
         MULT_mult_6_ab_12__5_, MULT_mult_6_ab_12__6_, MULT_mult_6_ab_12__7_,
         MULT_mult_6_ab_12__9_, MULT_mult_6_ab_12__12_, MULT_mult_6_ab_12__13_,
         MULT_mult_6_ab_12__14_, MULT_mult_6_ab_12__16_,
         MULT_mult_6_ab_12__17_, MULT_mult_6_ab_12__18_,
         MULT_mult_6_ab_12__19_, MULT_mult_6_ab_13__0_, MULT_mult_6_ab_13__2_,
         MULT_mult_6_ab_13__3_, MULT_mult_6_ab_13__4_, MULT_mult_6_ab_13__5_,
         MULT_mult_6_ab_13__6_, MULT_mult_6_ab_13__7_, MULT_mult_6_ab_13__9_,
         MULT_mult_6_ab_13__10_, MULT_mult_6_ab_13__12_,
         MULT_mult_6_ab_13__13_, MULT_mult_6_ab_13__15_,
         MULT_mult_6_ab_13__16_, MULT_mult_6_ab_13__17_,
         MULT_mult_6_ab_13__18_, MULT_mult_6_ab_14__0_, MULT_mult_6_ab_14__1_,
         MULT_mult_6_ab_14__3_, MULT_mult_6_ab_14__4_, MULT_mult_6_ab_14__5_,
         MULT_mult_6_ab_14__6_, MULT_mult_6_ab_14__7_, MULT_mult_6_ab_14__9_,
         MULT_mult_6_ab_14__11_, MULT_mult_6_ab_14__12_,
         MULT_mult_6_ab_14__13_, MULT_mult_6_ab_14__15_,
         MULT_mult_6_ab_14__16_, MULT_mult_6_ab_15__0_, MULT_mult_6_ab_15__2_,
         MULT_mult_6_ab_15__3_, MULT_mult_6_ab_15__4_, MULT_mult_6_ab_15__5_,
         MULT_mult_6_ab_15__6_, MULT_mult_6_ab_15__7_, MULT_mult_6_ab_15__8_,
         MULT_mult_6_ab_15__9_, MULT_mult_6_ab_15__11_, MULT_mult_6_ab_15__12_,
         MULT_mult_6_ab_15__14_, MULT_mult_6_ab_15__15_,
         MULT_mult_6_ab_15__16_, MULT_mult_6_ab_16__0_, MULT_mult_6_ab_16__2_,
         MULT_mult_6_ab_16__3_, MULT_mult_6_ab_16__4_, MULT_mult_6_ab_16__5_,
         MULT_mult_6_ab_16__6_, MULT_mult_6_ab_16__8_, MULT_mult_6_ab_16__11_,
         MULT_mult_6_ab_16__12_, MULT_mult_6_ab_16__14_,
         MULT_mult_6_ab_16__15_, MULT_mult_6_ab_17__0_, MULT_mult_6_ab_17__1_,
         MULT_mult_6_ab_17__2_, MULT_mult_6_ab_17__3_, MULT_mult_6_ab_17__4_,
         MULT_mult_6_ab_17__5_, MULT_mult_6_ab_17__7_, MULT_mult_6_ab_17__8_,
         MULT_mult_6_ab_17__10_, MULT_mult_6_ab_17__11_,
         MULT_mult_6_ab_17__13_, MULT_mult_6_ab_18__0_, MULT_mult_6_ab_18__1_,
         MULT_mult_6_ab_18__2_, MULT_mult_6_ab_18__3_, MULT_mult_6_ab_18__4_,
         MULT_mult_6_ab_18__5_, MULT_mult_6_ab_18__6_, MULT_mult_6_ab_18__7_,
         MULT_mult_6_ab_18__9_, MULT_mult_6_ab_18__10_, MULT_mult_6_ab_18__12_,
         MULT_mult_6_ab_18__13_, MULT_mult_6_ab_19__0_, MULT_mult_6_ab_19__2_,
         MULT_mult_6_ab_19__3_, MULT_mult_6_ab_19__4_, MULT_mult_6_ab_19__5_,
         MULT_mult_6_ab_19__7_, MULT_mult_6_ab_19__8_, MULT_mult_6_ab_19__9_,
         MULT_mult_6_ab_19__11_, MULT_mult_6_ab_19__12_, MULT_mult_6_ab_20__0_,
         MULT_mult_6_ab_20__1_, MULT_mult_6_ab_20__2_, MULT_mult_6_ab_20__3_,
         MULT_mult_6_ab_20__4_, MULT_mult_6_ab_20__6_, MULT_mult_6_ab_20__7_,
         MULT_mult_6_ab_20__8_, MULT_mult_6_ab_20__10_, MULT_mult_6_ab_21__0_,
         MULT_mult_6_ab_21__1_, MULT_mult_6_ab_21__2_, MULT_mult_6_ab_21__3_,
         MULT_mult_6_ab_21__4_, MULT_mult_6_ab_21__6_, MULT_mult_6_ab_21__7_,
         MULT_mult_6_ab_21__9_, MULT_mult_6_ab_21__10_, MULT_mult_6_ab_22__0_,
         MULT_mult_6_ab_22__1_, MULT_mult_6_ab_22__2_, MULT_mult_6_ab_22__4_,
         MULT_mult_6_ab_22__6_, MULT_mult_6_ab_22__8_, MULT_mult_6_ab_23__0_,
         MULT_mult_6_ab_23__2_, MULT_mult_6_ab_23__5_, MULT_mult_6_ab_23__6_,
         MULT_mult_6_ab_23__8_, MULT_mult_6_ab_24__0_, MULT_mult_6_ab_24__2_,
         MULT_mult_6_ab_24__5_, MULT_mult_6_ab_24__6_, MULT_mult_6_ab_25__0_,
         MULT_mult_6_ab_25__1_, MULT_mult_6_ab_25__4_, MULT_mult_6_ab_26__0_,
         MULT_mult_6_ab_26__1_, MULT_mult_6_ab_26__2_, MULT_mult_6_ab_26__3_,
         MULT_mult_6_ab_26__4_, MULT_mult_6_ab_27__0_, MULT_mult_6_ab_27__3_,
         MULT_mult_6_ab_28__2_;
  wire   [16:31] aluA;
  wire   [0:31] multOut;

  OAI22_X2 U181 ( .A1(n6223), .A2(n6219), .B1(n10936), .B2(n6217), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U183 ( .A1(n6222), .A2(n6219), .B1(n4940), .B2(n6217), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U184 ( .A1(n6221), .A2(n6219), .B1(n4950), .B2(n6217), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U216 ( .A1(n6223), .A2(net76318), .B1(n4938), .B2(n6215), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U218 ( .A1(n6222), .A2(net76318), .B1(n4957), .B2(n6215), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U219 ( .A1(n6221), .A2(net76318), .B1(n4952), .B2(n6215), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U386 ( .A1(n6223), .A2(n6213), .B1(n10937), .B2(n6176), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U388 ( .A1(n6222), .A2(n6213), .B1(n10934), .B2(n6176), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U389 ( .A1(n6221), .A2(n6214), .B1(n5543), .B2(n6176), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U421 ( .A1(n6223), .A2(n6211), .B1(n10938), .B2(n6209), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U423 ( .A1(n6222), .A2(n6211), .B1(n4937), .B2(n6209), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U424 ( .A1(n6221), .A2(n6211), .B1(n4958), .B2(n6209), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U660 ( .A1(n6223), .A2(n6207), .B1(n10939), .B2(n6205), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U662 ( .A1(n6222), .A2(n6207), .B1(n10935), .B2(n6205), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U663 ( .A1(n6221), .A2(n6207), .B1(n4951), .B2(n6205), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U729 ( .A1(n6223), .A2(n6203), .B1(n5898), .B2(n6202), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U731 ( .A1(n6222), .A2(n6203), .B1(n5397), .B2(n6202), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U732 ( .A1(n6221), .A2(n6203), .B1(n5433), .B2(n6202), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U969 ( .A1(n6223), .A2(n6198), .B1(n10940), .B2(n6196), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U971 ( .A1(n6222), .A2(n6198), .B1(n4956), .B2(n6197), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U972 ( .A1(n6221), .A2(n6198), .B1(n4961), .B2(n6196), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1005 ( .A1(n6223), .A2(n6194), .B1(n10941), .B2(n6192), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1007 ( .A1(n6222), .A2(n6194), .B1(n4959), .B2(n6192), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1008 ( .A1(n6221), .A2(n6194), .B1(n4960), .B2(n6192), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__31_), .QN(n5948) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[31]) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__31_), .QN(n5792) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__31_), .QN(n5891) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__31_), .QN(net78127) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__31_), .QN(net78128) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__31_), .QN(net80211) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__31_), .QN(net80440) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__31_), .QN(net82515) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__31_), .QN(n5949) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__31_), .QN(net80208) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__31_), .QN(net78108) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__31_), .QN(net78109) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__31_), .QN(n6002) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__31_), .QN(n6003) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__31_), .QN(n5823) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__31_), .QN(n5999) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__31_), .QN(n5717) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__31_), .QN(n4939) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__31_), .QN(n5765) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__31_), .QN(net82499) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__31_), .QN(n5026) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__31_), .QN(n5790) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__31_), .QN(n4917) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__31_), .QN(n5778) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__31_), .QN(n5788) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__31_), .QN(n5895) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__31_), .QN(n5811) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__31_), .QN(n5893) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__31_), .QN(n5824) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__31_), .QN(n5827) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__31_), .QN(net78235) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__15_), .QN(n4935) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__15_), .QN(n4927) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__15_), .QN(n4945) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__15_), .QN(n4948) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__15_), .QN(n5396) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__15_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__15_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__15_), .QN(n5917) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__15_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__15_), .QN(n10950) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__15_), .QN(n4944) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__15_), .QN(n5784) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__15_), .QN(n5251) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__15_), .QN(n4934) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__15_), .QN(n4919) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__15_), .QN(n4943) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__15_), .QN(n5431) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__15_), .QN(n5122) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__15_), .QN(n4942) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__15_), .QN(n5866) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__15_), .QN(n4941) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__15_), .QN(n5714) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__15_), .QN(n5856) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__15_), .QN(n5121) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__15_), .QN(n5852) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__15_), .QN(n5250) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__14_), .QN(n4933) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__14_), .QN(n4918) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__14_), .QN(n4932) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__14_), .QN(n4926) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__14_), .QN(n5395) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__14_), .QN(n4981) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__14_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__14_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__14_), .QN(n5838) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__14_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__14_), .QN(n4831) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__14_), .QN(n5839) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__14_), .QN(n4936) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__14_), .QN(n5879) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__14_), .QN(n5662) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__14_), .QN(n4931) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__14_), .QN(n5837) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__14_), .QN(n4930) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__14_), .QN(n5841) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__14_), .QN(n5394) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__14_), .QN(n5842) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__14_), .QN(n4929) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__14_), .QN(n5819) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__14_), .QN(n5883) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__14_), .QN(n4928) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__14_), .QN(n5843) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__14_), .QN(n5844) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__10_), .QN(n5249) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__10_), .QN(n5350) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__10_), .QN(n5248) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__10_), .QN(n5349) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__10_), .QN(n5083) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__10_), .QN(n5120) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__10_), .QN(n5114) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__10_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__10_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__10_), .QN(n5773) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__10_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__10_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__10_), .QN(n5877) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__10_), .QN(n5247) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__10_), .QN(n5025) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__10_), .QN(n5110) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__10_), .QN(n5109) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__10_), .QN(n5082) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__10_), .QN(n5246) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__10_), .QN(n5430) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__10_), .QN(n4979) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__10_), .QN(n5393) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__10_), .QN(n5774) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__10_), .QN(n5108) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__10_), .QN(n5245) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__10_), .QN(n5614) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__10_), .QN(n5107) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__10_), .QN(n5024) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__10_), .QN(n5775) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__10_), .QN(n5119) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__10_), .QN(n5875) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__10_), .QN(n5106) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__2_), .QN(n4987) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__2_), .QN(n5244) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__2_), .QN(n5243) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__2_), .QN(n5242) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__2_), .QN(n4986) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__2_), .QN(n5392) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__2_), .QN(n5241) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__20_), .QN(n5240) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__20_), .QN(n5346) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__20_), .QN(n5239) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__20_), .QN(n5345) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__20_), .QN(n5344) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__20_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__20_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__20_), .QN(n5023) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__20_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__20_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__20_), .QN(n5681) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__20_), .QN(n5238) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__20_), .QN(n5661) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__20_), .QN(n5237) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__20_), .QN(n5236) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__20_), .QN(n5343) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__20_), .QN(n5235) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__20_), .QN(n5342) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__20_), .QN(n5391) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__20_), .QN(n5341) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__20_), .QN(n5234) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__20_), .QN(n5105) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__20_), .QN(n5081) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__20_), .QN(n5233) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__20_), .QN(n5340) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__20_), .QN(n5682) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__20_), .QN(n5390) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__20_), .QN(n5821) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__20_), .QN(n5232) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__3_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__3_), .QN(n5429) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__3_), .QN(n5428) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__3_), .QN(n5389) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__19_), .QN(n5227) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__19_), .QN(n5337) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__19_), .QN(n5226) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__19_), .QN(n5336) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__19_), .QN(n5335) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__19_), .QN(n5388) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__19_), .QN(n5426) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__19_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__19_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__19_), .QN(n5651) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__19_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__19_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__19_), .QN(n5225) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__19_), .QN(n4973) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__19_), .QN(n5104) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__19_), .QN(n5224) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__19_), .QN(n5334) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__19_), .QN(n5223) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__19_), .QN(n5425) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__19_), .QN(n5080) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__19_), .QN(n5118) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__19_), .QN(n5333) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__19_), .QN(n5222) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__19_), .QN(n5221) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__19_), .QN(n4978) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__19_), .QN(n5220) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__19_), .QN(n5332) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__19_), .QN(n5387) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__19_), .QN(n5219) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__4_), .QN(n5218) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__4_), .QN(n5386) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__4_), .QN(n5217) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__4_), .QN(n5216) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__4_), .QN(n5215) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__11_), .QN(n5873) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__11_), .QN(n5858) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__11_), .QN(n5881) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__11_), .QN(n5908) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__11_), .QN(n5871) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__11_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__29_), .QN(n5987) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__29_), .QN(n5125) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__29_), .QN(n4940) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__29_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__29_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__29_), .QN(n5989) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__29_), .QN(n5985) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__29_), .QN(n4937) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__29_), .QN(n5214) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__29_), .QN(n4974) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__29_), .QN(n5123) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__29_), .QN(net87633) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__29_), .QN(n5988) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__29_), .QN(n4977) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__29_), .QN(n5397) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__29_), .QN(n5126) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__29_), .QN(n5213) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__29_), .QN(n5914) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__29_), .QN(n5991) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__29_), .QN(n5328) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__26_), .QN(n5422) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__26_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__26_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__26_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__26_), .QN(n5421) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__26_), .QN(n5212) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__26_), .QN(n5327) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__26_), .QN(n5211) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__26_), .QN(n5210) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__26_), .QN(n5326) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__26_), .QN(n5209) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__26_), .QN(n5420) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__26_), .QN(n5325) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__26_), .QN(n5385) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__26_), .QN(n5208) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__26_), .QN(n5324) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__26_), .QN(n5207) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__26_), .QN(n5323) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__7_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__6_), .QN(n5206) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__6_), .QN(n5322) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__6_), .QN(n5205) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__6_), .QN(n5321) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__6_), .QN(n5320) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__6_), .QN(n5384) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__6_), .QN(n5419) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__6_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__6_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__6_), .QN(n5319) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__6_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__6_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__6_), .QN(n5113) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__6_), .QN(n5103) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__6_), .QN(n5204) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__6_), .QN(n5203) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__6_), .QN(n5318) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__6_), .QN(n5202) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__6_), .QN(n5418) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__6_), .QN(n5317) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__6_), .QN(n5383) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__6_), .QN(n5316) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__6_), .QN(n5201) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__6_), .QN(n5200) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__6_), .QN(n5315) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__6_), .QN(n5417) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__6_), .QN(n5382) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__6_), .QN(n5437) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__5_), .QN(n5199) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__5_), .QN(n5314) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__5_), .QN(n4985) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__5_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__5_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__5_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__5_), .QN(n5416) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__5_), .QN(n5313) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__5_), .QN(n5198) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__5_), .QN(n5197) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__5_), .QN(n5381) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__5_), .QN(n5196) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__5_), .QN(n5195) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__5_), .QN(n5309) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__5_), .QN(n5308) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__21_), .QN(n5194) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__21_), .QN(n5307) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__21_), .QN(n5193) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__21_), .QN(n5306) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__21_), .QN(n5305) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__21_), .QN(n5414) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__21_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__21_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__21_), .QN(n5304) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__21_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__21_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__21_), .QN(n5192) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__21_), .QN(n5191) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__21_), .QN(n5190) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__21_), .QN(n5303) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__21_), .QN(n5189) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__21_), .QN(n5302) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__21_), .QN(n5380) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__21_), .QN(n5301) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__21_), .QN(n5188) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__21_), .QN(n5187) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__21_), .QN(n5300) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__21_), .QN(n5186) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__21_), .QN(n5299) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__21_), .QN(n5810) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__21_), .QN(n5379) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__21_), .QN(n5808) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__21_), .QN(n5185) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[21]), .QN(n5085) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__8_), .QN(n5102) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__8_), .QN(n4972) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__8_), .QN(n5101) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__8_), .QN(n5079) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__8_), .QN(n5686) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__8_), .QN(n5378) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__8_), .QN(n5028) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__8_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__8_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__8_), .QN(n5911) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__8_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__8_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__8_), .QN(n5978) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__8_), .QN(n5184) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__8_), .QN(n5183) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__8_), .QN(n5182) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__8_), .QN(n5298) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__8_), .QN(n5181) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__8_), .QN(n5413) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__8_), .QN(n5297) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__8_), .QN(n5377) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__8_), .QN(n5296) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__8_), .QN(n5180) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__8_), .QN(n5179) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__8_), .QN(n5910) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__8_), .QN(n5178) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__8_), .QN(n5295) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__8_), .QN(n5950) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__8_), .QN(n5376) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__8_), .QN(n5977) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__8_), .QN(n5127) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__13_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__13_), .QN(n5715) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__13_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__13_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__13_), .QN(n5816) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__13_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__13_), .QN(n5801) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__13_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__13_), .QN(n5835) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__13_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__13_), .QN(n5767) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__13_), .QN(n5937) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__13_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__13_), .QN(n5939) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__13_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__13_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__13_), .QN(n5799) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__13_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__13_), .QN(n5719) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__13_), .QN(n4850) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__13_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__13_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__13_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__13_), .QN(n4845) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__13_), .QN(net83260) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__13_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__13_), .QN(n5803) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__13_), .QN(net84518) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__13_), .QN(n5813) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__13_) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[13]) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[10]) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__9_), .QN(n5177) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__9_), .QN(n5294) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__9_), .QN(n5176) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__9_), .QN(n5293) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__9_), .QN(n5292) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__9_), .QN(n5375) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__9_), .QN(n5112) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__9_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__9_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__9_), .QN(n5022) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__9_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__9_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__9_), .QN(n5412) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__9_), .QN(n5175) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__9_), .QN(n5021) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__9_), .QN(n5100) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__9_), .QN(n5174) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__9_), .QN(n5291) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__9_), .QN(n5173) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__9_), .QN(n5411) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__9_), .QN(n5290) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__9_), .QN(n5374) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__9_), .QN(n5289) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__9_), .QN(n5172) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__9_), .QN(n5171) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__9_), .QN(n4976) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__9_), .QN(n5170) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__9_), .QN(n5288) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__9_), .QN(n5653) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__9_), .QN(n5373) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__9_), .QN(n5616) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__9_), .QN(n5169) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__23_), .QN(n5168) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__23_), .QN(n5287) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__23_), .QN(n5286) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__23_), .QN(n5372) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__23_), .QN(n5410) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__23_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__23_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__23_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__23_), .QN(n5409) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__23_), .QN(n5167) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__23_), .QN(n5166) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__23_), .QN(n5285) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__23_), .QN(n5165) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__23_), .QN(n5408) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__23_), .QN(n5284) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__23_), .QN(n5371) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__23_), .QN(n5164) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__23_), .QN(n5283) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__23_), .QN(n5163) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__23_), .QN(n5282) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[23]), .QN(n5086) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[20]) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[19]), .QN(n5063) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__16_), .QN(n5667) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__16_), .QN(n4859) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__16_), .QN(n5755) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__16_), .QN(n5676) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__16_), .QN(n5786) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__16_), .QN(n5612) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__16_), .QN(n5665) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__16_), .QN(n5610) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__16_), .QN(n5617) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__16_), .QN(n5771) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__16_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__12_), .QN(n5862) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__12_), .QN(n5860) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__12_), .QN(n5864) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__12_), .QN(n4825) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__12_), .QN(n5673) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__12_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__17_), .QN(n5099) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__17_), .QN(n5078) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__17_), .QN(n5098) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__17_), .QN(n5077) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__17_), .QN(n5076) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__17_), .QN(n5117) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__17_), .QN(n5111) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__17_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__17_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__17_), .QN(n5020) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__17_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__17_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__17_), .QN(n5027) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__17_), .QN(n5097) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__17_), .QN(n5019) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__17_), .QN(n5096) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__17_), .QN(n5162) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__17_), .QN(n5281) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__17_), .QN(n5161) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__17_), .QN(n5407) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__17_), .QN(n5075) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__17_), .QN(n5116) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__17_), .QN(n5074) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__17_), .QN(n5095) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__17_), .QN(n5094) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__17_), .QN(n5018) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__17_), .QN(n5160) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__17_), .QN(n5280) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__17_), .QN(n5620) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__17_), .QN(n5370) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__17_), .QN(n5073) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__17_), .QN(n5093) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__25_), .QN(n5279) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__25_), .QN(n5369) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__25_), .QN(n5406) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__25_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__25_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__25_), .QN(n5405) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__25_), .QN(n5159) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__25_), .QN(n5278) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__25_), .QN(n5158) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__25_), .QN(n5157) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__25_), .QN(n5277) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__25_), .QN(n5156) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__25_), .QN(n5404) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__25_), .QN(n5155) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__25_), .QN(n5276) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__25_), .QN(n5154) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__25_), .QN(n5275) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__25_), .QN(n5274) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__25_), .QN(n5153) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[25]), .QN(n5087) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[22]) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__22_), .QN(n5152) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__22_), .QN(n5273) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__22_), .QN(n5151) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__22_), .QN(n5272) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__22_), .QN(n5271) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__22_), .QN(n5403) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__22_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__22_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__22_), .QN(n5270) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__22_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__22_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__22_), .QN(n5402) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__22_), .QN(n5150) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__22_), .QN(n5269) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__22_), .QN(n5149) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__22_), .QN(n5148) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__22_), .QN(n5268) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__22_), .QN(n5147) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__22_), .QN(n5267) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__22_), .QN(n5368) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__22_), .QN(n5266) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__22_), .QN(n5146) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__22_), .QN(n5092) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__22_), .QN(n5017) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__22_), .QN(n5145) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__22_), .QN(n5265) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__22_), .QN(n5621) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__22_), .QN(n5367) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__22_), .QN(n5144) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__27_), .QN(n5356) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__27_), .QN(n5362) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__27_), .QN(n5436) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__27_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__27_), .QN(n5361) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__27_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__27_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__27_), .QN(n5435) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__27_), .QN(n5355) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__27_), .QN(n5360) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__27_), .QN(n5354) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__27_), .QN(n5353) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__27_), .QN(n5352) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__27_), .QN(n5434) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__27_), .QN(n5359) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__27_), .QN(n5432) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__27_), .QN(n4949) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__18_), .QN(n5091) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__18_), .QN(n5072) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__18_), .QN(n5143) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__18_), .QN(n5264) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__18_), .QN(n5366) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__18_), .QN(n5685) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__18_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__18_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__18_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__18_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__18_), .QN(n5913) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__18_), .QN(n5142) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__18_), .QN(n5857) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__18_), .QN(n5141) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__18_), .QN(n5090) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__18_), .QN(n5071) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__18_), .QN(n5140) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__18_), .QN(n5401) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__18_), .QN(n5263) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__18_), .QN(n5365) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__18_), .QN(n5262) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__18_), .QN(n5139) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__18_), .QN(n5138) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__18_), .QN(n5878) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__18_), .QN(n5089) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__18_), .QN(n4925) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__18_), .QN(n4980) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__18_), .QN(n5115) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__18_), .QN(n5886) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__18_), .QN(n5088) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[18]) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[17]), .QN(n5084) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__28_), .QN(n5358) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__28_), .QN(n4950) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__28_), .QN(n4952) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__28_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__28_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__28_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__28_), .QN(n5351) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__28_), .QN(n5069) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__28_), .QN(n4951) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__28_), .QN(n5357) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__28_), .QN(n5433) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__30_), .QN(n5927) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__30_), .QN(n5961) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__30_), .QN(n5070) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__30_), .QN(n4938) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__30_), .QN(n5794) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__30_), .QN(n5925) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__30_), .QN(n5680) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__30_), .QN(n5833) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__30_), .QN(n5963) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__30_), .QN(n5920) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__30_), .QN(n5967) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__30_), .QN(n5924) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__30_), .QN(n5969) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__30_), .QN(n5934) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__30_), .QN(n5973) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__30_), .QN(n5922) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__30_), .QN(n5965) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__30_), .QN(n5124) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__30_), .QN(n5898) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__30_), .QN(n5971) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__30_), .QN(n5854) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__30_), .QN(n5929) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__30_), .QN(n5918) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__30_), .QN(n5992) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__30_), .QN(n5958) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__30_), .QN(n5994) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__30_), .QN(n5959) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__30_), .QN(n5996) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__30_), .QN(n4975) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[28]) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[26]) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__24_), .QN(n5137) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__24_), .QN(n5261) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__24_), .QN(n5136) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__24_), .QN(n5260) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__24_), .QN(n5259) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__24_), .QN(n5364) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__24_), .QN(n5400) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__24_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__24_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__24_), .QN(n5258) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__24_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__24_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__24_), .QN(n5399) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__24_), .QN(n5135) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__24_), .QN(n5257) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__24_), .QN(n5134) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__24_), .QN(n5133) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__24_), .QN(n5256) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__24_), .QN(n5132) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__24_), .QN(n5398) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__24_), .QN(n5255) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__24_), .QN(n5363) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__24_), .QN(n5254) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__24_), .QN(n5131) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__24_), .QN(n5130) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__24_), .QN(n4947) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__24_), .QN(n5129) );
  DFF_X2 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__24_), .QN(n4946) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__24_), .QN(n5253) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__24_), .QN(n5128) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[24]) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[16]) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[14]) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[9]) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[6]) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[5]) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[3]) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[1]) );
  DFF_X1 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__3_), .QN(n5956) );
  DFF_X1 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__11_), .QN(n5906) );
  DFF_X1 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__16_), .QN(n5903) );
  DFF_X1 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__1_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__8_), .QN(n5869) );
  DFF_X1 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__13_), .QN(n5849) );
  DFF_X1 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__14_), .QN(n5831) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5845) );
  DFF_X1 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__21_), .QN(n5807) );
  DFF_X1 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__14_), .QN(n5780) );
  DFF_X1 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__14_), .QN(n5776) );
  DFF_X1 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__4_), .QN(n5770) );
  DFF_X1 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__1_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__30_), .QN(n5671) );
  DFF_X1 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__5_), .QN(n5660) );
  DFF_X1 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__15_), .QN(n5656) );
  DFF_X1 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__13_), .QN(net148735) );
  DFF_X1 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__28_), .QN(n5569) );
  DFF_X1 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__28_), .QN(n5568) );
  DFF_X1 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__27_), .QN(n5567) );
  DFF_X1 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__27_), .QN(n5566) );
  DFF_X1 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__28_), .QN(n5565) );
  DFF_X1 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__24_), .QN(n5564) );
  DFF_X1 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__24_), .QN(n5563) );
  DFF_X1 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__27_), .QN(n5562) );
  DFF_X1 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__3_), .QN(n5559) );
  DFF_X1 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__26_), .QN(n5556) );
  DFF_X1 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__26_), .QN(n5555) );
  DFF_X1 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__5_), .QN(n5554) );
  DFF_X1 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__23_), .QN(n5553) );
  DFF_X1 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__25_), .QN(n5551) );
  DFF_X1 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__27_), .QN(n5550) );
  DFF_X1 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__27_), .QN(n5549) );
  DFF_X1 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__27_), .QN(n5548) );
  DFF_X1 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__28_), .QN(n5547) );
  DFF_X1 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__28_), .QN(n5546) );
  DFF_X1 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__28_), .QN(n5545) );
  DFF_X1 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__28_), .QN(n5544) );
  DFF_X1 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__28_), .QN(n5543) );
  DFF_X1 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__27_), .QN(n5542) );
  DFF_X1 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__3_), .QN(n5534) );
  DFF_X1 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__3_), .QN(n5533) );
  DFF_X1 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__3_), .QN(n5530) );
  DFF_X1 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__29_), .QN(n5523) );
  DFF_X1 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__29_), .QN(n5522) );
  DFF_X1 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__26_), .QN(n5521) );
  DFF_X1 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__26_), .QN(n5518) );
  DFF_X1 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__6_), .QN(n5517) );
  DFF_X1 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__5_), .QN(n5516) );
  DFF_X1 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__5_), .QN(n5515) );
  DFF_X1 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__23_), .QN(n5514) );
  DFF_X1 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__23_), .QN(n5513) );
  DFF_X1 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__25_), .QN(n5508) );
  DFF_X1 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__30_), .QN(n5507) );
  DFF_X1 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__20_), .QN(n5506) );
  DFF_X1 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__21_), .QN(n5505) );
  DFF_X1 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__22_), .QN(n5504) );
  DFF_X1 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__26_), .QN(n5503) );
  DFF_X1 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__23_), .QN(n5502) );
  DFF_X1 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__25_), .QN(n5501) );
  DFF_X1 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__20_), .QN(n5500) );
  DFF_X1 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__21_), .QN(n5499) );
  DFF_X1 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__22_), .QN(n5498) );
  DFF_X1 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__27_), .QN(n5497) );
  DFF_X1 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__27_), .QN(n5496) );
  DFF_X1 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__28_), .QN(n5495) );
  DFF_X1 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__28_), .QN(n5494) );
  DFF_X1 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__27_), .QN(n5493) );
  DFF_X1 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__28_), .QN(n5491) );
  DFF_X1 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__27_), .QN(n5490) );
  DFF_X1 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__27_), .QN(n5489) );
  DFF_X1 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__28_), .QN(n5488) );
  DFF_X1 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__28_), .QN(n5487) );
  DFF_X1 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__28_), .QN(n5486) );
  DFF_X1 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__28_), .QN(n5485) );
  DFF_X1 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__28_), .QN(n5484) );
  DFF_X1 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__3_), .QN(n5476) );
  DFF_X1 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__3_), .QN(n5475) );
  DFF_X1 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__3_), .QN(n5474) );
  DFF_X1 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__4_), .QN(n5468) );
  DFF_X1 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__4_), .QN(n5464) );
  DFF_X1 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__29_), .QN(n5463) );
  DFF_X1 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__29_), .QN(n5462) );
  DFF_X1 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__29_), .QN(n5461) );
  DFF_X1 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__29_), .QN(n5460) );
  DFF_X1 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__29_), .QN(n5459) );
  DFF_X1 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__29_), .QN(n5458) );
  DFF_X1 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__26_), .QN(n5457) );
  DFF_X1 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__26_), .QN(n5456) );
  DFF_X1 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__26_), .QN(n5455) );
  DFF_X1 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__26_), .QN(n5454) );
  DFF_X1 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__26_), .QN(n5453) );
  DFF_X1 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__26_), .QN(n5452) );
  DFF_X1 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__5_), .QN(n5451) );
  DFF_X1 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__23_), .QN(n5450) );
  DFF_X1 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__23_), .QN(n5449) );
  DFF_X1 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__23_), .QN(n5448) );
  DFF_X1 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__23_), .QN(n5447) );
  DFF_X1 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__23_), .QN(n5446) );
  DFF_X1 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__25_), .QN(n5445) );
  DFF_X1 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__25_), .QN(n5444) );
  DFF_X1 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__25_), .QN(n5443) );
  DFF_X1 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__25_), .QN(n5442) );
  DFF_X1 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__25_), .QN(n5441) );
  DFF_X1 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__30_), .QN(n5440) );
  DFF_X1 PCLOGIC_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[0]), .QN(n5439) );
  DFF_X1 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__5_), .QN(n5310) );
  DFF_X1 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__3_), .QN(n5231) );
  DFF_X1 PCLOGIC_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[7]), .QN(n5059) );
  DFF_X1 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__28_), .QN(n5047) );
  DFF_X1 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__3_), .QN(n5046) );
  DFF_X1 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__3_), .QN(n5045) );
  DFF_X1 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__5_), .QN(n5044) );
  DFF_X1 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__5_), .QN(n5043) );
  DFF_X1 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__15_), .QN(n5038) );
  DFF_X1 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__20_), .QN(n5037) );
  DFF_X1 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__19_), .QN(n5036) );
  DFF_X1 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__19_), .QN(n5035) );
  DFF_X1 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__21_), .QN(n5034) );
  DFF_X1 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__4_), .QN(n5033) );
  DFF_X1 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__28_), .QN(n5032) );
  DFF_X1 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__18_), .QN(n5030) );
  DFF_X1 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__14_), .QN(n5029) );
  DFF_X1 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__29_), .QN(n4988) );
  DFF_X1 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__5_), .QN(n4984) );
  DFF_X1 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__22_), .QN(n4983) );
  DFF_X1 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__6_), .QN(n4982) );
  DFF_X1 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__28_), .QN(n4961) );
  DFF_X1 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__28_), .QN(n4960) );
  DFF_X1 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__29_), .QN(n4959) );
  DFF_X1 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__28_), .QN(n4958) );
  DFF_X1 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__29_), .QN(n4957) );
  DFF_X1 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__29_), .QN(n4956) );
  DFF_X1 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__27_), .QN(n4955) );
  DFF_X1 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__15_), .QN(n4954) );
  DFF_X1 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__31_), .QN(n4953) );
  DFF_X1 PCLOGIC_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[4]), .QN(n4924) );
  DFF_X1 PCLOGIC_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[2]), .QN(n4923) );
  DFF_X1 PCLOGIC_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[8]), .QN(n4909) );
  DFF_X1 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__15_), .QN(n4902) );
  DFF_X1 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__1_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__15_), .QN(n5683) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__19_), .QN(n5031) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__15_), .QN(n4901) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__18_), .QN(n5785) );
  INV_X2 U4891 ( .A(net77744), .ZN(net81764) );
  INV_X2 U4893 ( .A(net88131), .ZN(n4797) );
  INV_X4 U4894 ( .A(net76242), .ZN(n5587) );
  INV_X4 U4895 ( .A(n5083), .ZN(n4798) );
  AOI22_X4 U4896 ( .A1(REGFILE_reg_out_16__12_), .A2(net77764), .B1(
        REGFILE_reg_out_15__12_), .B2(net75468), .ZN(n6650) );
  AOI22_X2 U4897 ( .A1(REGFILE_reg_out_19__8_), .A2(net77810), .B1(
        REGFILE_reg_out_1__8_), .B2(net75478), .ZN(n6733) );
  OAI21_X2 U4898 ( .B1(net76502), .B2(n10581), .A(n10580), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U4899 ( .B1(net76506), .B2(n10593), .A(n10592), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  INV_X1 U4902 ( .A(n10141), .ZN(dmem_addr_out[10]) );
  OAI211_X4 U4903 ( .C1(n10141), .C2(net76646), .A(net70740), .B(n10140), .ZN(
        n10142) );
  NAND4_X4 U4904 ( .A1(n9370), .A2(n9371), .A3(n9372), .A4(n9369), .ZN(
        dmem_addr_out[9]) );
  NAND2_X4 U4905 ( .A1(multOut[9]), .A2(net92392), .ZN(n9370) );
  OAI211_X4 U4906 ( .C1(n9377), .C2(net76646), .A(net70740), .B(n9376), .ZN(
        n9378) );
  INV_X8 U4907 ( .A(net77436), .ZN(net77430) );
  INV_X16 U4908 ( .A(net77436), .ZN(net77428) );
  INV_X8 U4909 ( .A(net77430), .ZN(net77416) );
  INV_X8 U4910 ( .A(net77430), .ZN(net77418) );
  INV_X8 U4911 ( .A(net77430), .ZN(net77420) );
  NAND4_X4 U4912 ( .A1(n6543), .A2(n6542), .A3(n6541), .A4(n6540), .ZN(n6549)
         );
  AOI22_X1 U4913 ( .A1(REGFILE_reg_out_14__28_), .A2(net77780), .B1(
        REGFILE_reg_out_13__28_), .B2(n5663), .ZN(n6304) );
  AOI22_X2 U4915 ( .A1(REGFILE_reg_out_14__17_), .A2(net77780), .B1(
        REGFILE_reg_out_13__17_), .B2(n5663), .ZN(net75859) );
  AOI22_X2 U4916 ( .A1(REGFILE_reg_out_14__13_), .A2(net77780), .B1(n5804), 
        .B2(n5664), .ZN(net75761) );
  INV_X16 U4918 ( .A(n9528), .ZN(n6050) );
  NAND4_X4 U4919 ( .A1(n9698), .A2(n9697), .A3(n9696), .A4(n9695), .ZN(
        dmem_addr_out[7]) );
  NAND2_X4 U4920 ( .A1(net76650), .A2(dmem_addr_out[7]), .ZN(n9702) );
  NAND3_X4 U4921 ( .A1(n9702), .A2(net70740), .A3(n9701), .ZN(n9703) );
  INV_X16 U4922 ( .A(n6058), .ZN(n4802) );
  INV_X16 U4923 ( .A(n6069), .ZN(n4803) );
  INV_X16 U4924 ( .A(n9974), .ZN(n6069) );
  AOI21_X4 U4925 ( .B1(multOut[2]), .B2(net92392), .A(n5749), .ZN(net71394) );
  MUX2_X2 U4926 ( .A(multOut[6]), .B(n9662), .S(net73585), .Z(n9668) );
  OAI211_X4 U4927 ( .C1(n9673), .C2(net76646), .A(net70740), .B(n9672), .ZN(
        n9674) );
  INV_X2 U4928 ( .A(n9673), .ZN(dmem_addr_out[6]) );
  OAI21_X2 U4931 ( .B1(n6214), .B2(n6072), .A(n10048), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U4932 ( .B1(n10534), .B2(n6072), .A(n10050), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U4933 ( .B1(n10532), .B2(n6072), .A(n10049), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  NAND2_X1 U4935 ( .A1(n6100), .A2(REGFILE_reg_out_13__1_), .ZN(n10176) );
  INV_X16 U4936 ( .A(net77752), .ZN(net77746) );
  INV_X4 U4937 ( .A(net77436), .ZN(net77432) );
  INV_X8 U4938 ( .A(net77432), .ZN(net77414) );
  INV_X16 U4939 ( .A(net77432), .ZN(net77410) );
  INV_X8 U4940 ( .A(n4830), .ZN(n4897) );
  OAI21_X2 U4941 ( .B1(dmem_write_out[1]), .B2(net75427), .A(n10945), .ZN(
        net70921) );
  INV_X2 U4942 ( .A(net70921), .ZN(net36466) );
  INV_X8 U4943 ( .A(net80161), .ZN(n5576) );
  AND2_X4 U4944 ( .A1(net76270), .A2(n10521), .ZN(n4804) );
  AND2_X4 U4945 ( .A1(net76270), .A2(n10519), .ZN(n4805) );
  AND2_X4 U4946 ( .A1(n4874), .A2(n8673), .ZN(n4806) );
  INV_X32 U4947 ( .A(instruction[11]), .ZN(net87820) );
  XOR2_X1 U4948 ( .A(n9057), .B(n10463), .Z(n4807) );
  XOR2_X1 U4949 ( .A(n5762), .B(net77040), .Z(n4808) );
  AND2_X2 U4950 ( .A1(n5712), .A2(net70696), .ZN(n4809) );
  NAND2_X4 U4951 ( .A1(n10303), .A2(net70697), .ZN(net70710) );
  NAND2_X4 U4952 ( .A1(n8985), .A2(net70697), .ZN(n9606) );
  NAND2_X4 U4953 ( .A1(n8861), .A2(net70697), .ZN(n9854) );
  NAND2_X1 U4954 ( .A1(n6005), .A2(net71026), .ZN(n10544) );
  INV_X8 U4955 ( .A(n10544), .ZN(n6082) );
  NAND2_X1 U4956 ( .A1(net71026), .A2(n10099), .ZN(net70718) );
  XOR2_X1 U4957 ( .A(n5783), .B(net77038), .Z(n4810) );
  AND2_X2 U4958 ( .A1(n10465), .A2(net78051), .ZN(n4811) );
  AND4_X4 U4959 ( .A1(n9805), .A2(n8717), .A3(n8716), .A4(n8715), .ZN(n4812)
         );
  INV_X16 U4960 ( .A(n8679), .ZN(n6022) );
  NAND2_X4 U4961 ( .A1(net76270), .A2(n8668), .ZN(n8679) );
  XOR2_X1 U4962 ( .A(n10110), .B(n10404), .Z(n4813) );
  INV_X16 U4963 ( .A(n9325), .ZN(n6039) );
  NAND2_X4 U4964 ( .A1(net76270), .A2(n9320), .ZN(n9325) );
  INV_X16 U4965 ( .A(n8961), .ZN(n6028) );
  NAND2_X4 U4966 ( .A1(net76270), .A2(n8956), .ZN(n8961) );
  INV_X16 U4967 ( .A(n9579), .ZN(n6052) );
  NAND2_X4 U4968 ( .A1(net76270), .A2(n9573), .ZN(n9579) );
  XOR2_X1 U4969 ( .A(n4856), .B(net77038), .Z(n4814) );
  INV_X8 U4970 ( .A(dmem_write_out[19]), .ZN(n6529) );
  NAND2_X4 U4971 ( .A1(net76270), .A2(n9425), .ZN(n9426) );
  AND2_X2 U4972 ( .A1(multOut[2]), .A2(net92392), .ZN(n4815) );
  NAND2_X4 U4973 ( .A1(net76270), .A2(n9867), .ZN(n9868) );
  INV_X8 U4974 ( .A(net70541), .ZN(net76514) );
  NAND2_X4 U4975 ( .A1(net76270), .A2(n9113), .ZN(n4816) );
  INV_X8 U4976 ( .A(net77464), .ZN(net77452) );
  AOI22_X1 U4977 ( .A1(REGFILE_reg_out_11__6_), .A2(net77746), .B1(
        REGFILE_reg_out_12__6_), .B2(net83168), .ZN(n6769) );
  AOI22_X2 U4978 ( .A1(REGFILE_reg_out_11__12_), .A2(net77748), .B1(n4826), 
        .B2(net83168), .ZN(n6649) );
  AOI22_X4 U4979 ( .A1(REGFILE_reg_out_9__10_), .A2(net77698), .B1(
        REGFILE_reg_out_8__10_), .B2(net75454), .ZN(n6700) );
  NAND2_X1 U4980 ( .A1(REGFILE_reg_out_3__10_), .A2(net77414), .ZN(n7830) );
  INV_X4 U4981 ( .A(n5775), .ZN(n4817) );
  NAND4_X2 U4982 ( .A1(net75623), .A2(net75624), .A3(net75625), .A4(net75626), 
        .ZN(net75617) );
  AOI22_X2 U4983 ( .A1(REGFILE_reg_out_19__26_), .A2(net77814), .B1(
        REGFILE_reg_out_1__26_), .B2(net82631), .ZN(n6345) );
  INV_X32 U4984 ( .A(net77816), .ZN(net77814) );
  INV_X8 U4985 ( .A(net77640), .ZN(net77634) );
  AOI22_X4 U4986 ( .A1(REGFILE_reg_out_29__16_), .A2(net77652), .B1(n5787), 
        .B2(n6911), .ZN(n6579) );
  AOI22_X4 U4987 ( .A1(REGFILE_reg_out_29__21_), .A2(net77652), .B1(
        REGFILE_reg_out_28__21_), .B2(n6911), .ZN(n6475) );
  AOI22_X4 U4988 ( .A1(REGFILE_reg_out_9__20_), .A2(net77700), .B1(
        REGFILE_reg_out_8__20_), .B2(n4829), .ZN(n6494) );
  AOI22_X2 U4989 ( .A1(REGFILE_reg_out_16__4_), .A2(net77764), .B1(
        REGFILE_reg_out_15__4_), .B2(n5579), .ZN(n6814) );
  AOI22_X2 U4990 ( .A1(REGFILE_reg_out_24__19_), .A2(net75437), .B1(
        REGFILE_reg_out_25__19_), .B2(net75438), .ZN(n6520) );
  AOI22_X2 U4991 ( .A1(REGFILE_reg_out_24__20_), .A2(net75437), .B1(n4836), 
        .B2(net75438), .ZN(n6496) );
  INV_X8 U4992 ( .A(net75438), .ZN(net77616) );
  AOI22_X2 U4993 ( .A1(REGFILE_reg_out_26__14_), .A2(net75439), .B1(n5840), 
        .B2(net89184), .ZN(n6623) );
  AOI22_X2 U4994 ( .A1(REGFILE_reg_out_16__18_), .A2(net75467), .B1(
        REGFILE_reg_out_15__18_), .B2(net75468), .ZN(n6536) );
  AOI22_X2 U4995 ( .A1(REGFILE_reg_out_16__16_), .A2(net87506), .B1(n5666), 
        .B2(net75468), .ZN(n6568) );
  INV_X16 U4996 ( .A(net75465), .ZN(net77752) );
  INV_X8 U4997 ( .A(net76235), .ZN(net75465) );
  INV_X32 U4998 ( .A(net77752), .ZN(net77748) );
  INV_X4 U4999 ( .A(n5913), .ZN(n4818) );
  INV_X32 U5000 ( .A(net76201), .ZN(net75439) );
  NOR2_X4 U5001 ( .A1(n6420), .A2(n6419), .ZN(n6431) );
  INV_X4 U5002 ( .A(net81601), .ZN(net83408) );
  NOR2_X4 U5003 ( .A1(n6805), .A2(n6804), .ZN(n6806) );
  INV_X16 U5004 ( .A(instruction[12]), .ZN(net73533) );
  NAND4_X4 U5005 ( .A1(n6561), .A2(n6560), .A3(n6559), .A4(n6558), .ZN(
        net75847) );
  AOI22_X4 U5006 ( .A1(REGFILE_reg_out_26__24_), .A2(net77618), .B1(
        REGFILE_reg_out_27__24_), .B2(net77630), .ZN(n6402) );
  AOI22_X2 U5007 ( .A1(REGFILE_reg_out_24__18_), .A2(net75437), .B1(n5684), 
        .B2(net75438), .ZN(n6544) );
  NAND2_X1 U5008 ( .A1(REGFILE_reg_out_13__15_), .A2(net77454), .ZN(n7593) );
  NAND2_X1 U5009 ( .A1(n6100), .A2(REGFILE_reg_out_13__12_), .ZN(n9122) );
  NAND2_X1 U5010 ( .A1(REGFILE_reg_out_13__12_), .A2(net77452), .ZN(n7725) );
  BUF_X32 U5011 ( .A(n6505), .Z(n4819) );
  INV_X16 U5012 ( .A(net84760), .ZN(net84761) );
  NAND4_X2 U5013 ( .A1(n6959), .A2(n6958), .A3(n6957), .A4(n6956), .ZN(n6965)
         );
  NAND2_X4 U5014 ( .A1(REGFILE_reg_out_1__29_), .A2(net77516), .ZN(n6956) );
  INV_X32 U5015 ( .A(instruction[15]), .ZN(net82739) );
  AOI22_X4 U5016 ( .A1(REGFILE_reg_out_0__17_), .A2(net82342), .B1(
        REGFILE_reg_out_10__17_), .B2(net83203), .ZN(net75862) );
  BUF_X16 U5017 ( .A(n10916), .Z(n4864) );
  AOI22_X2 U5018 ( .A1(REGFILE_reg_out_21__14_), .A2(net77844), .B1(
        REGFILE_reg_out_20__14_), .B2(net77852), .ZN(n6611) );
  NAND2_X4 U5019 ( .A1(n6526), .A2(n6527), .ZN(dmem_write_out[19]) );
  NAND3_X4 U5020 ( .A1(n4842), .A2(instruction[15]), .A3(instruction[13]), 
        .ZN(n4821) );
  NAND3_X2 U5021 ( .A1(n4842), .A2(instruction[15]), .A3(instruction[13]), 
        .ZN(net76261) );
  NAND2_X4 U5022 ( .A1(n5642), .A2(net77272), .ZN(n4822) );
  INV_X32 U5023 ( .A(n4822), .ZN(n4963) );
  NAND2_X4 U5024 ( .A1(net73533), .A2(instruction[11]), .ZN(n4823) );
  INV_X8 U5025 ( .A(net77768), .ZN(net77764) );
  INV_X8 U5026 ( .A(net77768), .ZN(net77762) );
  INV_X2 U5027 ( .A(n4917), .ZN(n4824) );
  INV_X2 U5028 ( .A(n4825), .ZN(n4826) );
  AOI22_X2 U5029 ( .A1(REGFILE_reg_out_26__10_), .A2(net75439), .B1(
        REGFILE_reg_out_27__10_), .B2(net89184), .ZN(n6703) );
  NOR2_X4 U5030 ( .A1(n6525), .A2(n6524), .ZN(n6526) );
  NAND2_X1 U5031 ( .A1(REGFILE_reg_out_28__18_), .A2(net77384), .ZN(n7449) );
  INV_X2 U5032 ( .A(n5026), .ZN(n4827) );
  NAND4_X2 U5033 ( .A1(n6625), .A2(n6624), .A3(n6623), .A4(n6622), .ZN(n6626)
         );
  AOI22_X2 U5034 ( .A1(REGFILE_reg_out_30__14_), .A2(net77638), .B1(net82613), 
        .B2(n4838), .ZN(n6624) );
  BUF_X32 U5035 ( .A(n10914), .Z(n4828) );
  INV_X16 U5037 ( .A(net76220), .ZN(n4829) );
  INV_X8 U5038 ( .A(net76220), .ZN(net75454) );
  NAND4_X4 U5039 ( .A1(n7041), .A2(n7040), .A3(n7039), .A4(n7038), .ZN(n8451)
         );
  NAND2_X2 U5040 ( .A1(n8451), .A2(net123282), .ZN(n5657) );
  INV_X32 U5041 ( .A(net77464), .ZN(net77456) );
  INV_X8 U5042 ( .A(net76251), .ZN(net76204) );
  NOR2_X4 U5044 ( .A1(n6515), .A2(n6514), .ZN(n6527) );
  AOI22_X2 U5045 ( .A1(n5921), .A2(net77406), .B1(n5968), .B2(n6014), .ZN(
        n6943) );
  AOI22_X4 U5046 ( .A1(REGFILE_reg_out_26__7_), .A2(net75439), .B1(
        REGFILE_reg_out_27__7_), .B2(net77626), .ZN(net75621) );
  NAND2_X4 U5047 ( .A1(REGFILE_reg_out_31__29_), .A2(net77498), .ZN(n6990) );
  AOI22_X4 U5048 ( .A1(REGFILE_reg_out_0__15_), .A2(net82342), .B1(n5853), 
        .B2(net83203), .ZN(n6588) );
  INV_X2 U5050 ( .A(n4831), .ZN(n4832) );
  INV_X1 U5051 ( .A(net73831), .ZN(n4833) );
  INV_X4 U5052 ( .A(n4833), .ZN(n4834) );
  NAND2_X1 U5053 ( .A1(n4884), .A2(REGFILE_reg_out_18__16_), .ZN(n9224) );
  INV_X4 U5054 ( .A(n5784), .ZN(n4835) );
  AOI22_X2 U5055 ( .A1(REGFILE_reg_out_24__15_), .A2(net75437), .B1(n4835), 
        .B2(net124970), .ZN(n6598) );
  NAND2_X2 U5056 ( .A1(n8411), .A2(net77272), .ZN(n6946) );
  INV_X16 U5057 ( .A(instruction[2]), .ZN(net74029) );
  INV_X16 U5058 ( .A(instruction[14]), .ZN(n4843) );
  AOI22_X2 U5059 ( .A1(REGFILE_reg_out_30__17_), .A2(net84761), .B1(
        REGFILE_reg_out_2__17_), .B2(net82613), .ZN(n5584) );
  AOI22_X2 U5061 ( .A1(REGFILE_reg_out_30__15_), .A2(net77638), .B1(n4837), 
        .B2(net82613), .ZN(n6600) );
  AOI22_X2 U5062 ( .A1(REGFILE_reg_out_30__12_), .A2(net84761), .B1(n5863), 
        .B2(net82613), .ZN(n6660) );
  AOI22_X2 U5063 ( .A1(REGFILE_reg_out_30__9_), .A2(net77634), .B1(
        REGFILE_reg_out_2__9_), .B2(net82613), .ZN(n6726) );
  AOI22_X2 U5064 ( .A1(REGFILE_reg_out_30__7_), .A2(net77634), .B1(
        REGFILE_reg_out_2__7_), .B2(net82613), .ZN(net75620) );
  AOI22_X2 U5065 ( .A1(REGFILE_reg_out_30__8_), .A2(net77634), .B1(n5912), 
        .B2(net75442), .ZN(n6748) );
  INV_X16 U5067 ( .A(net75418), .ZN(net77328) );
  INV_X16 U5068 ( .A(net74050), .ZN(net77512) );
  NOR2_X2 U5069 ( .A1(net87633), .A2(net77512), .ZN(net91561) );
  INV_X1 U5070 ( .A(net75464), .ZN(net77744) );
  AOI22_X2 U5071 ( .A1(REGFILE_reg_out_0__20_), .A2(net82342), .B1(
        REGFILE_reg_out_10__20_), .B2(net83203), .ZN(n6486) );
  INV_X4 U5072 ( .A(net77550), .ZN(net77576) );
  INV_X8 U5073 ( .A(net77576), .ZN(net77554) );
  INV_X4 U5074 ( .A(n5661), .ZN(n4836) );
  NAND2_X4 U5075 ( .A1(n6731), .A2(n6730), .ZN(dmem_write_out[9]) );
  INV_X4 U5076 ( .A(n5917), .ZN(n4837) );
  NAND2_X1 U5077 ( .A1(net77406), .A2(REGFILE_reg_out_19__27_), .ZN(n7059) );
  NAND2_X1 U5078 ( .A1(net77406), .A2(REGFILE_reg_out_27__28_), .ZN(n7005) );
  NAND2_X1 U5079 ( .A1(net77406), .A2(REGFILE_reg_out_19__28_), .ZN(n7015) );
  NAND2_X1 U5080 ( .A1(net77406), .A2(REGFILE_reg_out_3__28_), .ZN(n7035) );
  AOI22_X2 U5081 ( .A1(n4827), .A2(net77406), .B1(n5791), .B2(n6014), .ZN(
        n6922) );
  OAI21_X2 U5082 ( .B1(n7007), .B2(n7006), .A(n6011), .ZN(n7041) );
  INV_X4 U5084 ( .A(n5838), .ZN(n4838) );
  INV_X2 U5085 ( .A(n5683), .ZN(n4839) );
  INV_X16 U5086 ( .A(net77440), .ZN(net77436) );
  INV_X2 U5087 ( .A(net75437), .ZN(net77608) );
  AOI22_X4 U5088 ( .A1(REGFILE_reg_out_11__14_), .A2(net77748), .B1(n5846), 
        .B2(net83167), .ZN(n6613) );
  OAI21_X2 U5089 ( .B1(net76502), .B2(n10619), .A(n10618), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  AOI22_X4 U5090 ( .A1(REGFILE_reg_out_16__22_), .A2(net77764), .B1(
        REGFILE_reg_out_15__22_), .B2(n5579), .ZN(n6440) );
  NAND2_X1 U5091 ( .A1(REGFILE_reg_out_30__13_), .A2(net75441), .ZN(n5941) );
  AOI22_X1 U5092 ( .A1(REGFILE_reg_out_19__28_), .A2(net77814), .B1(
        REGFILE_reg_out_1__28_), .B2(net82631), .ZN(n6298) );
  AOI22_X1 U5093 ( .A1(REGFILE_reg_out_19__27_), .A2(net77814), .B1(
        REGFILE_reg_out_1__27_), .B2(net82631), .ZN(n6322) );
  AOI22_X2 U5095 ( .A1(REGFILE_reg_out_16__14_), .A2(net75467), .B1(n5884), 
        .B2(net75468), .ZN(n6614) );
  INV_X32 U5096 ( .A(net77624), .ZN(net77620) );
  INV_X16 U5097 ( .A(net75439), .ZN(net77624) );
  INV_X32 U5098 ( .A(instruction[14]), .ZN(n4840) );
  INV_X32 U5099 ( .A(instruction[14]), .ZN(n4841) );
  INV_X32 U5100 ( .A(instruction[14]), .ZN(n4842) );
  OAI21_X1 U5101 ( .B1(dmem_write_out[0]), .B2(net75427), .A(n10945), .ZN(
        net71027) );
  OAI21_X2 U5102 ( .B1(dmem_write_out[4]), .B2(net75427), .A(n10945), .ZN(
        n10400) );
  NAND2_X1 U5103 ( .A1(REGFILE_reg_out_6__29_), .A2(net77550), .ZN(n6963) );
  NAND2_X1 U5104 ( .A1(REGFILE_reg_out_22__29_), .A2(net77550), .ZN(n6981) );
  AOI22_X4 U5105 ( .A1(REGFILE_reg_out_14__15_), .A2(net77780), .B1(
        REGFILE_reg_out_13__15_), .B2(n5664), .ZN(n6591) );
  INV_X16 U5106 ( .A(n6074), .ZN(n6072) );
  INV_X16 U5107 ( .A(n6074), .ZN(n6073) );
  AOI22_X1 U5108 ( .A1(REGFILE_reg_out_26__26_), .A2(net77620), .B1(
        REGFILE_reg_out_27__26_), .B2(net89184), .ZN(n6359) );
  AOI22_X2 U5109 ( .A1(REGFILE_reg_out_26__11_), .A2(net75439), .B1(net89184), 
        .B2(n5859), .ZN(n6681) );
  INV_X16 U5110 ( .A(net77776), .ZN(n5579) );
  NAND3_X2 U5111 ( .A1(instruction[15]), .A2(instruction[14]), .A3(
        instruction[13]), .ZN(n4844) );
  INV_X8 U5112 ( .A(net75440), .ZN(net77632) );
  NAND3_X4 U5113 ( .A1(net87495), .A2(n4841), .A3(instruction[15]), .ZN(
        net76252) );
  INV_X8 U5114 ( .A(net76252), .ZN(net76196) );
  AOI22_X2 U5115 ( .A1(REGFILE_reg_out_24__5_), .A2(net75437), .B1(
        REGFILE_reg_out_25__5_), .B2(net77610), .ZN(n6800) );
  AOI22_X2 U5116 ( .A1(REGFILE_reg_out_24__29_), .A2(net77602), .B1(
        REGFILE_reg_out_25__29_), .B2(net77610), .ZN(n6287) );
  AOI22_X2 U5117 ( .A1(n5935), .A2(net77478), .B1(n5974), .B2(net77550), .ZN(
        n6937) );
  OAI21_X4 U5118 ( .B1(n6964), .B2(n6965), .A(net73838), .ZN(n6997) );
  NAND4_X4 U5119 ( .A1(n6963), .A2(n6962), .A3(n6961), .A4(n6960), .ZN(n6964)
         );
  NAND2_X1 U5120 ( .A1(n4805), .A2(REGFILE_reg_out_14__13_), .ZN(n9437) );
  NAND2_X1 U5121 ( .A1(REGFILE_reg_out_14__13_), .A2(net77560), .ZN(n7684) );
  INV_X2 U5122 ( .A(n4845), .ZN(n4846) );
  NAND2_X1 U5123 ( .A1(n4875), .A2(REGFILE_reg_out_24__13_), .ZN(n9459) );
  NAND2_X1 U5124 ( .A1(REGFILE_reg_out_24__13_), .A2(net77308), .ZN(n7665) );
  INV_X1 U5125 ( .A(n4819), .ZN(dmem_write_out[20]) );
  OR2_X4 U5126 ( .A1(n10040), .A2(n10039), .ZN(dmem_addr_out[3]) );
  OAI22_X2 U5127 ( .A1(n10038), .A2(net70691), .B1(n10037), .B2(n5752), .ZN(
        n10039) );
  INV_X32 U5128 ( .A(instruction[1]), .ZN(net73496) );
  INV_X4 U5129 ( .A(net77550), .ZN(net77574) );
  INV_X8 U5130 ( .A(net77574), .ZN(net77564) );
  INV_X8 U5131 ( .A(net77574), .ZN(net77562) );
  INV_X8 U5132 ( .A(net77574), .ZN(net77560) );
  INV_X8 U5133 ( .A(net77574), .ZN(net77568) );
  INV_X8 U5134 ( .A(net77576), .ZN(net77566) );
  INV_X8 U5135 ( .A(net77576), .ZN(net77556) );
  INV_X8 U5136 ( .A(net77576), .ZN(net77558) );
  NAND4_X4 U5137 ( .A1(n6630), .A2(n6631), .A3(n6633), .A4(n6632), .ZN(
        net75759) );
  AOI22_X2 U5138 ( .A1(REGFILE_reg_out_19__21_), .A2(net77812), .B1(
        REGFILE_reg_out_1__21_), .B2(net75478), .ZN(n6459) );
  INV_X4 U5139 ( .A(n5680), .ZN(n4849) );
  AOI22_X2 U5140 ( .A1(REGFILE_reg_out_3__30_), .A2(net77406), .B1(n4849), 
        .B2(n6014), .ZN(n6939) );
  AND2_X2 U5141 ( .A1(n5654), .A2(n5655), .ZN(n6941) );
  INV_X2 U5142 ( .A(n4850), .ZN(n4851) );
  NAND2_X2 U5143 ( .A1(n10207), .A2(n10206), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  INV_X8 U5144 ( .A(n9835), .ZN(n10915) );
  INV_X16 U5145 ( .A(n5697), .ZN(net75456) );
  AOI22_X2 U5146 ( .A1(REGFILE_reg_out_7__3_), .A2(net75455), .B1(
        REGFILE_reg_out_6__3_), .B2(net75456), .ZN(n6843) );
  OAI21_X1 U5147 ( .B1(n6553), .B2(net78056), .A(n6552), .ZN(n4852) );
  INV_X8 U5148 ( .A(dmem_write_out[18]), .ZN(n6553) );
  AOI22_X2 U5149 ( .A1(REGFILE_reg_out_24__14_), .A2(net75437), .B1(n5880), 
        .B2(net124970), .ZN(n6622) );
  INV_X4 U5150 ( .A(n5843), .ZN(n4853) );
  AOI22_X4 U5151 ( .A1(REGFILE_reg_out_11__13_), .A2(net77748), .B1(n5608), 
        .B2(net83167), .ZN(net75763) );
  INV_X4 U5152 ( .A(n5915), .ZN(n5916) );
  NOR2_X2 U5153 ( .A1(n6501), .A2(n6500), .ZN(n6502) );
  INV_X4 U5154 ( .A(n5856), .ZN(n4854) );
  NAND2_X2 U5155 ( .A1(net77100), .A2(n4990), .ZN(n10171) );
  NAND2_X2 U5156 ( .A1(net77104), .A2(n4806), .ZN(n10207) );
  NAND2_X2 U5157 ( .A1(n10203), .A2(n10202), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U5158 ( .A1(n10197), .A2(n10196), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U5159 ( .A1(n10205), .A2(n10204), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U5160 ( .A1(n10191), .A2(n10190), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U5161 ( .A1(n10185), .A2(n10184), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U5162 ( .A1(n10169), .A2(n10168), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U5163 ( .A1(n10219), .A2(n10218), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U5164 ( .A1(n10221), .A2(n10220), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U5165 ( .A1(n10187), .A2(n10186), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U5166 ( .A1(n10171), .A2(n10170), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  INV_X8 U5167 ( .A(n5578), .ZN(net77454) );
  INV_X16 U5169 ( .A(net75467), .ZN(net77768) );
  INV_X16 U5170 ( .A(net77768), .ZN(net87506) );
  INV_X8 U5172 ( .A(net123382), .ZN(net76198) );
  NAND2_X1 U5173 ( .A1(n6175), .A2(REGFILE_reg_out_28__15_), .ZN(n10299) );
  NAND2_X1 U5174 ( .A1(net77382), .A2(REGFILE_reg_out_28__15_), .ZN(n7579) );
  NAND2_X2 U5176 ( .A1(net73851), .A2(n4963), .ZN(net75396) );
  OAI22_X4 U5177 ( .A1(net82515), .A2(n5648), .B1(net80208), .B2(net85371), 
        .ZN(net82513) );
  AOI22_X4 U5178 ( .A1(REGFILE_reg_out_19__13_), .A2(net77812), .B1(n4851), 
        .B2(net75478), .ZN(n6631) );
  AOI22_X2 U5179 ( .A1(REGFILE_reg_out_16__17_), .A2(net75467), .B1(
        REGFILE_reg_out_15__17_), .B2(net75468), .ZN(net75860) );
  NAND2_X4 U5180 ( .A1(net76238), .A2(n5607), .ZN(net76253) );
  AOI22_X2 U5181 ( .A1(REGFILE_reg_out_0__10_), .A2(net120684), .B1(n5876), 
        .B2(net83203), .ZN(n6692) );
  INV_X8 U5182 ( .A(net76194), .ZN(net75438) );
  INV_X8 U5183 ( .A(net77616), .ZN(net77610) );
  AOI22_X2 U5184 ( .A1(REGFILE_reg_out_24__2_), .A2(net75437), .B1(
        REGFILE_reg_out_25__2_), .B2(net77610), .ZN(n6866) );
  NOR2_X2 U5186 ( .A1(n6339), .A2(n6340), .ZN(n6341) );
  INV_X8 U5187 ( .A(n6000), .ZN(n6010) );
  INV_X16 U5188 ( .A(n6010), .ZN(n5664) );
  NAND4_X4 U5189 ( .A1(n6969), .A2(n6968), .A3(n6967), .A4(n6966), .ZN(n6975)
         );
  OAI21_X2 U5190 ( .B1(n6982), .B2(n6983), .A(net77588), .ZN(n6995) );
  AOI22_X2 U5191 ( .A1(REGFILE_reg_out_16__5_), .A2(net87506), .B1(
        REGFILE_reg_out_15__5_), .B2(net77774), .ZN(n6792) );
  NOR2_X2 U5192 ( .A1(n6795), .A2(n6794), .ZN(n6807) );
  INV_X4 U5193 ( .A(n5845), .ZN(n5846) );
  INV_X4 U5194 ( .A(n5996), .ZN(n5997) );
  INV_X2 U5195 ( .A(n9306), .ZN(n4856) );
  AOI22_X4 U5196 ( .A1(REGFILE_reg_out_19__17_), .A2(net77812), .B1(
        REGFILE_reg_out_1__17_), .B2(net75478), .ZN(n6555) );
  AOI22_X2 U5197 ( .A1(REGFILE_reg_out_24__26_), .A2(net75437), .B1(
        REGFILE_reg_out_25__26_), .B2(net77614), .ZN(n6358) );
  INV_X32 U5198 ( .A(instruction[14]), .ZN(net86793) );
  INV_X1 U5199 ( .A(n6994), .ZN(n4857) );
  INV_X4 U5200 ( .A(n4857), .ZN(n4858) );
  INV_X8 U5201 ( .A(n10288), .ZN(n5851) );
  INV_X2 U5202 ( .A(n4859), .ZN(n4860) );
  AOI22_X4 U5203 ( .A1(n5919), .A2(net77474), .B1(n5995), .B2(net77400), .ZN(
        n6948) );
  INV_X4 U5204 ( .A(n5994), .ZN(n5995) );
  INV_X4 U5205 ( .A(n8408), .ZN(n6952) );
  NAND2_X4 U5206 ( .A1(n5607), .A2(net122022), .ZN(net76235) );
  INV_X16 U5207 ( .A(n5689), .ZN(n5696) );
  NOR2_X4 U5208 ( .A1(n9963), .A2(n9962), .ZN(n9967) );
  OR2_X1 U5209 ( .A1(n5991), .A2(net75424), .ZN(n6971) );
  INV_X16 U5210 ( .A(net75424), .ZN(net77550) );
  OAI21_X2 U5211 ( .B1(n10532), .B2(net77114), .A(n10119), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  NOR2_X4 U5212 ( .A1(n6363), .A2(n6362), .ZN(n6364) );
  OAI21_X2 U5213 ( .B1(net70509), .B2(net77116), .A(n5690), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  INV_X8 U5214 ( .A(net86304), .ZN(net77506) );
  NAND2_X4 U5215 ( .A1(multOut[3]), .A2(n4861), .ZN(n4862) );
  NAND2_X4 U5216 ( .A1(n10032), .A2(net73585), .ZN(n4863) );
  NAND2_X4 U5217 ( .A1(n4862), .A2(n4863), .ZN(n10040) );
  INV_X4 U5218 ( .A(net73585), .ZN(n4861) );
  AOI22_X2 U5219 ( .A1(REGFILE_reg_out_19__19_), .A2(net77812), .B1(
        REGFILE_reg_out_1__19_), .B2(net75478), .ZN(n6507) );
  AOI22_X4 U5220 ( .A1(REGFILE_reg_out_19__16_), .A2(net77812), .B1(
        REGFILE_reg_out_1__16_), .B2(net75478), .ZN(n6563) );
  INV_X8 U5221 ( .A(net75478), .ZN(n5624) );
  AOI22_X1 U5222 ( .A1(REGFILE_reg_out_16__0_), .A2(net87506), .B1(
        REGFILE_reg_out_15__0_), .B2(net77774), .ZN(n6903) );
  AOI22_X1 U5223 ( .A1(REGFILE_reg_out_16__2_), .A2(net75467), .B1(
        REGFILE_reg_out_15__2_), .B2(net77774), .ZN(n6858) );
  AOI22_X1 U5224 ( .A1(REGFILE_reg_out_16__27_), .A2(net75467), .B1(
        REGFILE_reg_out_15__27_), .B2(net77774), .ZN(n6327) );
  AOI22_X1 U5225 ( .A1(REGFILE_reg_out_16__29_), .A2(net77762), .B1(
        REGFILE_reg_out_15__29_), .B2(net77774), .ZN(n6279) );
  AOI22_X1 U5226 ( .A1(REGFILE_reg_out_16__26_), .A2(net87506), .B1(
        REGFILE_reg_out_15__26_), .B2(n5579), .ZN(n6350) );
  AOI22_X1 U5227 ( .A1(REGFILE_reg_out_16__3_), .A2(net77764), .B1(
        REGFILE_reg_out_15__3_), .B2(n5579), .ZN(n6836) );
  INV_X4 U5228 ( .A(net88131), .ZN(net122022) );
  AOI22_X2 U5229 ( .A1(REGFILE_reg_out_24__6_), .A2(net75437), .B1(n5764), 
        .B2(net124970), .ZN(n6778) );
  AOI22_X4 U5230 ( .A1(REGFILE_reg_out_19__24_), .A2(net77814), .B1(
        REGFILE_reg_out_1__24_), .B2(net82631), .ZN(n5622) );
  NAND4_X4 U5231 ( .A1(net76031), .A2(net76032), .A3(n5622), .A4(net76034), 
        .ZN(net76025) );
  NOR2_X4 U5232 ( .A1(instruction[2]), .A2(instruction[4]), .ZN(n4865) );
  INV_X32 U5233 ( .A(net77392), .ZN(net77386) );
  NAND2_X2 U5234 ( .A1(REGFILE_reg_out_5__29_), .A2(net77444), .ZN(n6960) );
  INV_X16 U5235 ( .A(n5588), .ZN(net83203) );
  AOI22_X2 U5236 ( .A1(REGFILE_reg_out_11__18_), .A2(net77748), .B1(
        REGFILE_reg_out_12__18_), .B2(net83167), .ZN(n6535) );
  CLKBUF_X3 U5237 ( .A(net77272), .Z(n4866) );
  INV_X16 U5238 ( .A(net77464), .ZN(net77444) );
  INV_X16 U5239 ( .A(net77464), .ZN(net77458) );
  INV_X8 U5240 ( .A(net77272), .ZN(net77276) );
  NAND2_X1 U5241 ( .A1(REGFILE_reg_out_25__26_), .A2(net77514), .ZN(n7088) );
  NAND2_X1 U5242 ( .A1(REGFILE_reg_out_17__26_), .A2(net77514), .ZN(n7098) );
  NAND2_X1 U5243 ( .A1(REGFILE_reg_out_9__26_), .A2(net77514), .ZN(n7108) );
  NAND2_X1 U5244 ( .A1(REGFILE_reg_out_1__26_), .A2(net77514), .ZN(n7118) );
  NAND2_X1 U5245 ( .A1(net77514), .A2(REGFILE_reg_out_17__27_), .ZN(n7054) );
  NAND2_X1 U5246 ( .A1(net77514), .A2(REGFILE_reg_out_25__28_), .ZN(n7000) );
  NAND2_X1 U5247 ( .A1(net77514), .A2(REGFILE_reg_out_17__28_), .ZN(n7010) );
  AOI22_X2 U5248 ( .A1(n4824), .A2(net77514), .B1(n5779), .B2(net77298), .ZN(
        n6921) );
  INV_X4 U5249 ( .A(net77514), .ZN(net86238) );
  AOI22_X2 U5250 ( .A1(n5818), .A2(net77514), .B1(n5970), .B2(net77298), .ZN(
        n6942) );
  AOI22_X2 U5251 ( .A1(n5855), .A2(net77514), .B1(n5930), .B2(net77298), .ZN(
        n6934) );
  AOI22_X2 U5252 ( .A1(n5928), .A2(net77514), .B1(n5962), .B2(net77298), .ZN(
        n6950) );
  NAND2_X2 U5253 ( .A1(REGFILE_reg_out_17__29_), .A2(net77514), .ZN(n6976) );
  INV_X4 U5254 ( .A(net77320), .ZN(net77314) );
  INV_X4 U5255 ( .A(net77320), .ZN(net77316) );
  AOI22_X2 U5256 ( .A1(REGFILE_reg_out_14__11_), .A2(net77780), .B1(
        REGFILE_reg_out_13__11_), .B2(n5664), .ZN(n6673) );
  AOI22_X2 U5257 ( .A1(REGFILE_reg_out_14__10_), .A2(net77778), .B1(
        REGFILE_reg_out_13__10_), .B2(n5664), .ZN(n6695) );
  NAND2_X4 U5258 ( .A1(n9968), .A2(net76270), .ZN(n9974) );
  AOI22_X2 U5259 ( .A1(REGFILE_reg_out_24__25_), .A2(net75437), .B1(
        REGFILE_reg_out_25__25_), .B2(net77610), .ZN(n6382) );
  NAND2_X1 U5260 ( .A1(net77474), .A2(REGFILE_reg_out_5__28_), .ZN(n7028) );
  AOI22_X2 U5261 ( .A1(n5834), .A2(net77474), .B1(n5964), .B2(net77400), .ZN(
        n6944) );
  NOR2_X4 U5262 ( .A1(n10040), .A2(n10039), .ZN(n10045) );
  OAI21_X2 U5263 ( .B1(n6993), .B2(n6992), .A(n8411), .ZN(n6994) );
  NAND4_X4 U5264 ( .A1(n6987), .A2(n6986), .A3(n6985), .A4(n6984), .ZN(n6993)
         );
  NOR2_X2 U5265 ( .A1(n6491), .A2(n6490), .ZN(n6503) );
  AOI22_X2 U5266 ( .A1(REGFILE_reg_out_24__10_), .A2(net75437), .B1(
        REGFILE_reg_out_25__10_), .B2(net75438), .ZN(n6702) );
  AOI22_X2 U5267 ( .A1(REGFILE_reg_out_24__9_), .A2(net75437), .B1(
        REGFILE_reg_out_25__9_), .B2(net124970), .ZN(n6724) );
  INV_X16 U5268 ( .A(net76237), .ZN(net75467) );
  NAND4_X4 U5269 ( .A1(n6557), .A2(n6556), .A3(n6555), .A4(n6554), .ZN(
        net75857) );
  AOI22_X4 U5270 ( .A1(REGFILE_reg_out_23__17_), .A2(net77828), .B1(
        REGFILE_reg_out_22__17_), .B2(net77836), .ZN(n6556) );
  INV_X32 U5271 ( .A(net77816), .ZN(net77812) );
  INV_X32 U5272 ( .A(instruction[15]), .ZN(net73511) );
  NAND2_X4 U5273 ( .A1(multOut[0]), .A2(net105376), .ZN(net105318) );
  INV_X16 U5274 ( .A(n5588), .ZN(net75464) );
  NAND4_X4 U5275 ( .A1(net75849), .A2(n5584), .A3(n5586), .A4(n5585), .ZN(
        n5583) );
  NAND2_X1 U5276 ( .A1(net75844), .A2(instruction[30]), .ZN(n5639) );
  INV_X8 U5277 ( .A(n5645), .ZN(net77440) );
  OAI21_X2 U5278 ( .B1(n10367), .B2(n10366), .A(n10365), .ZN(n10370) );
  INV_X8 U5279 ( .A(n5646), .ZN(n5645) );
  INV_X16 U5280 ( .A(net77394), .ZN(net77384) );
  INV_X16 U5281 ( .A(net77394), .ZN(net77380) );
  INV_X4 U5282 ( .A(n10944), .ZN(n6505) );
  NAND3_X1 U5283 ( .A1(n8564), .A2(instruction[5]), .A3(net73496), .ZN(n8542)
         );
  INV_X16 U5284 ( .A(n6920), .ZN(n6014) );
  INV_X16 U5285 ( .A(net85371), .ZN(net77336) );
  NOR3_X1 U5286 ( .A1(n8438), .A2(n8437), .A3(n8436), .ZN(n8439) );
  NOR2_X1 U5287 ( .A1(net70868), .A2(net71273), .ZN(n8614) );
  OAI21_X2 U5288 ( .B1(n9033), .B2(n9032), .A(n9031), .ZN(n9053) );
  OAI21_X2 U5289 ( .B1(n9833), .B2(n9356), .A(n9355), .ZN(n10131) );
  AOI21_X2 U5290 ( .B1(net73638), .B2(net73646), .A(n8568), .ZN(n8569) );
  INV_X4 U5292 ( .A(n10385), .ZN(n10912) );
  NOR3_X2 U5293 ( .A1(n8559), .A2(instruction[2]), .A3(instruction[0]), .ZN(
        n8553) );
  INV_X4 U5294 ( .A(dmem_write_out[22]), .ZN(n6457) );
  OAI21_X2 U5295 ( .B1(n8270), .B2(n8269), .A(net77290), .ZN(n8271) );
  INV_X16 U5296 ( .A(net77360), .ZN(net77338) );
  OAI21_X1 U5297 ( .B1(n7214), .B2(n7213), .A(net77588), .ZN(n7215) );
  OAI21_X2 U5298 ( .B1(n7139), .B2(n7138), .A(n6011), .ZN(n7173) );
  OAI21_X1 U5299 ( .B1(n7259), .B2(n7258), .A(net77588), .ZN(n7260) );
  OAI21_X1 U5300 ( .B1(n7349), .B2(n7348), .A(net77588), .ZN(n7350) );
  INV_X8 U5301 ( .A(net75479), .ZN(net77832) );
  INV_X4 U5302 ( .A(net76257), .ZN(net75479) );
  INV_X8 U5303 ( .A(net75469), .ZN(net77784) );
  INV_X4 U5304 ( .A(net76241), .ZN(net75469) );
  OAI21_X1 U5305 ( .B1(net36488), .B2(net70535), .A(net70838), .ZN(net70837)
         );
  NOR2_X1 U5306 ( .A1(net70868), .A2(n10404), .ZN(n8611) );
  NOR2_X2 U5307 ( .A1(n8624), .A2(n8623), .ZN(n8625) );
  NOR2_X1 U5308 ( .A1(net70868), .A2(n9954), .ZN(n8623) );
  OAI21_X2 U5309 ( .B1(n8818), .B2(n10054), .A(n8817), .ZN(n9993) );
  NOR2_X1 U5310 ( .A1(net70868), .A2(n10109), .ZN(n8620) );
  OAI21_X2 U5311 ( .B1(n9511), .B2(n9510), .A(n9509), .ZN(n9611) );
  OAI21_X2 U5312 ( .B1(n9581), .B2(net71273), .A(n9580), .ZN(n10091) );
  OAI21_X2 U5313 ( .B1(net70535), .B2(n9581), .A(n9580), .ZN(net70727) );
  OAI21_X2 U5314 ( .B1(n7125), .B2(n7124), .A(net77290), .ZN(n7126) );
  OAI21_X2 U5315 ( .B1(n7428), .B2(n7427), .A(n6019), .ZN(n7440) );
  NOR3_X1 U5316 ( .A1(n8418), .A2(n8417), .A3(n8416), .ZN(n8429) );
  NOR3_X1 U5317 ( .A1(n8425), .A2(n8424), .A3(n8423), .ZN(n8426) );
  NOR2_X1 U5318 ( .A1(n8422), .A2(n8421), .ZN(n8427) );
  NOR2_X1 U5319 ( .A1(n8431), .A2(n8430), .ZN(n8442) );
  NOR2_X1 U5320 ( .A1(n8433), .A2(n8432), .ZN(n8441) );
  NOR2_X1 U5321 ( .A1(n8435), .A2(n8434), .ZN(n8440) );
  NOR2_X1 U5322 ( .A1(n10494), .A2(net73541), .ZN(n8580) );
  AOI222_X1 U5323 ( .A1(n6083), .A2(n8976), .B1(n8728), .B2(n10466), .C1(
        n10465), .C2(net71026), .ZN(n9801) );
  AOI222_X1 U5324 ( .A1(n6083), .A2(n8928), .B1(n8891), .B2(n8759), .C1(n8758), 
        .C2(net71026), .ZN(n9804) );
  NAND3_X2 U5325 ( .A1(n8853), .A2(n8852), .A3(n8851), .ZN(n9011) );
  INV_X4 U5326 ( .A(n5065), .ZN(net78003) );
  OAI21_X2 U5327 ( .B1(net70731), .B2(net70732), .A(n5627), .ZN(net70730) );
  OAI21_X2 U5328 ( .B1(instructionAddr_out[28]), .B2(instructionAddr_out[29]), 
        .A(n8337), .ZN(n8331) );
  OAI21_X1 U5329 ( .B1(n7452), .B2(n7451), .A(n6012), .ZN(n7486) );
  OAI21_X1 U5330 ( .B1(n7462), .B2(n7461), .A(net77588), .ZN(n7485) );
  OAI21_X1 U5331 ( .B1(n7482), .B2(n7481), .A(net77292), .ZN(n7483) );
  OAI21_X1 U5332 ( .B1(n7680), .B2(n7679), .A(net77588), .ZN(n7703) );
  OAI21_X1 U5333 ( .B1(n7670), .B2(n7669), .A(n6012), .ZN(n7704) );
  OAI21_X1 U5334 ( .B1(n7700), .B2(n7699), .A(net77292), .ZN(n7701) );
  AOI21_X2 U5335 ( .B1(n9531), .B2(net77030), .A(n9517), .ZN(n9518) );
  AOI21_X2 U5336 ( .B1(n9634), .B2(net77030), .A(n9633), .ZN(n9635) );
  AOI21_X1 U5337 ( .B1(n9671), .B2(net77030), .A(n9670), .ZN(n9672) );
  AOI21_X1 U5338 ( .B1(n9965), .B2(net77030), .A(n9964), .ZN(n9966) );
  AOI21_X1 U5339 ( .B1(n10043), .B2(net77030), .A(n10042), .ZN(n10044) );
  AOI21_X1 U5340 ( .B1(net71396), .B2(net77030), .A(n5693), .ZN(n5692) );
  AOI21_X1 U5341 ( .B1(n10139), .B2(net77030), .A(n10138), .ZN(n10140) );
  NAND3_X2 U5342 ( .A1(dmem_read_in[0]), .A2(n4899), .A3(net73170), .ZN(
        net70740) );
  NOR2_X2 U5343 ( .A1(n8592), .A2(net70691), .ZN(n8780) );
  OAI21_X2 U5344 ( .B1(n4909), .B2(n8379), .A(n5059), .ZN(n8297) );
  NOR2_X1 U5345 ( .A1(n10430), .A2(n10429), .ZN(n10440) );
  INV_X8 U5346 ( .A(net77336), .ZN(net77358) );
  INV_X4 U5347 ( .A(dmem_write_out[21]), .ZN(n6481) );
  NAND4_X2 U5348 ( .A1(n6950), .A2(n6949), .A3(n6948), .A4(n6947), .ZN(n8408)
         );
  NAND3_X2 U5349 ( .A1(n6930), .A2(net75401), .A3(n6931), .ZN(n5915) );
  NOR3_X2 U5350 ( .A1(n10308), .A2(n10307), .A3(n10394), .ZN(n10455) );
  NAND3_X1 U5351 ( .A1(n8564), .A2(net73496), .A3(net73503), .ZN(n8551) );
  NAND3_X2 U5352 ( .A1(n8553), .A2(net73498), .A3(net73503), .ZN(n8554) );
  NOR2_X2 U5353 ( .A1(instruction[31]), .A2(n8563), .ZN(n8552) );
  NAND3_X2 U5354 ( .A1(net73684), .A2(instruction[28]), .A3(n5605), .ZN(
        net73695) );
  AOI21_X1 U5355 ( .B1(n8545), .B2(net73646), .A(n5252), .ZN(n8546) );
  NAND3_X1 U5356 ( .A1(n9066), .A2(n9093), .A3(n8850), .ZN(n9978) );
  OAI21_X2 U5357 ( .B1(n9683), .B2(n9614), .A(n9613), .ZN(n9663) );
  OAI21_X2 U5358 ( .B1(n7920), .B2(n7919), .A(net77290), .ZN(n7921) );
  OAI21_X2 U5359 ( .B1(n7962), .B2(n7961), .A(net77290), .ZN(n7963) );
  OAI21_X2 U5360 ( .B1(n8240), .B2(n8239), .A(n6011), .ZN(n8274) );
  OAI21_X2 U5361 ( .B1(n8260), .B2(n8259), .A(n6019), .ZN(n8272) );
  OAI21_X2 U5362 ( .B1(n8250), .B2(n8249), .A(net77588), .ZN(n8273) );
  OAI21_X2 U5363 ( .B1(n7876), .B2(n7875), .A(net77290), .ZN(n7877) );
  OAI21_X1 U5364 ( .B1(n7724), .B2(n7723), .A(net77588), .ZN(n7747) );
  OAI21_X1 U5365 ( .B1(n7714), .B2(n7713), .A(n6012), .ZN(n7748) );
  OAI21_X1 U5366 ( .B1(n7734), .B2(n7733), .A(n6019), .ZN(n7746) );
  OAI21_X1 U5367 ( .B1(n7184), .B2(n7183), .A(n6011), .ZN(n7218) );
  OAI21_X1 U5368 ( .B1(n7194), .B2(n7193), .A(net77290), .ZN(n7217) );
  OAI21_X1 U5369 ( .B1(n7204), .B2(n7203), .A(n6019), .ZN(n7216) );
  NAND4_X2 U5370 ( .A1(n6991), .A2(n6990), .A3(n6989), .A4(n6988), .ZN(n6992)
         );
  NAND4_X2 U5371 ( .A1(n6934), .A2(n6937), .A3(n6936), .A4(n6935), .ZN(
        net73831) );
  AOI22_X2 U5372 ( .A1(REGFILE_reg_out_5__30_), .A2(net77454), .B1(
        REGFILE_reg_out_4__30_), .B2(net77386), .ZN(n6940) );
  OAI21_X1 U5373 ( .B1(n7149), .B2(n7148), .A(net77290), .ZN(n7172) );
  OAI21_X1 U5374 ( .B1(n7159), .B2(n7158), .A(n6019), .ZN(n7171) );
  OAI21_X1 U5375 ( .B1(n7169), .B2(n7168), .A(net77588), .ZN(n7170) );
  NOR2_X2 U5376 ( .A1(net77999), .A2(n9373), .ZN(n8997) );
  NOR2_X2 U5377 ( .A1(net70811), .A2(n5597), .ZN(net72947) );
  AOI21_X1 U5378 ( .B1(n9000), .B2(net77030), .A(n8999), .ZN(n9001) );
  NOR2_X2 U5379 ( .A1(net76464), .A2(n8998), .ZN(n8999) );
  OAI21_X1 U5380 ( .B1(n7229), .B2(n7228), .A(n6012), .ZN(n7263) );
  OAI21_X1 U5381 ( .B1(n7239), .B2(n7238), .A(net77292), .ZN(n7262) );
  OAI21_X1 U5382 ( .B1(n7249), .B2(n7248), .A(n6019), .ZN(n7261) );
  OAI21_X1 U5383 ( .B1(n7822), .B2(n7821), .A(n6019), .ZN(n7834) );
  NOR2_X1 U5384 ( .A1(n8420), .A2(n8419), .ZN(n8428) );
  OAI21_X1 U5385 ( .B1(n7319), .B2(n7318), .A(n6012), .ZN(n7353) );
  OAI21_X1 U5386 ( .B1(n7329), .B2(n7328), .A(net77292), .ZN(n7352) );
  OAI21_X1 U5387 ( .B1(n7339), .B2(n7338), .A(n6019), .ZN(n7351) );
  OAI21_X2 U5388 ( .B1(n9393), .B2(n9062), .A(n9061), .ZN(n9353) );
  INV_X16 U5389 ( .A(net70718), .ZN(net77084) );
  NAND3_X2 U5390 ( .A1(n9584), .A2(n9583), .A3(n9582), .ZN(n9934) );
  AOI21_X2 U5391 ( .B1(n8728), .B2(n10013), .A(n5015), .ZN(n9582) );
  NOR2_X2 U5392 ( .A1(n10152), .A2(n9606), .ZN(n10105) );
  OAI21_X2 U5393 ( .B1(n8152), .B2(n8151), .A(n6011), .ZN(n8186) );
  OAI21_X2 U5394 ( .B1(n8162), .B2(n8161), .A(net77588), .ZN(n8185) );
  OAI21_X2 U5395 ( .B1(n8172), .B2(n8171), .A(n6019), .ZN(n8184) );
  OAI21_X2 U5396 ( .B1(n8064), .B2(n8063), .A(n6011), .ZN(n8098) );
  OAI21_X2 U5397 ( .B1(n8074), .B2(n8073), .A(net77588), .ZN(n8097) );
  OAI21_X2 U5398 ( .B1(n8084), .B2(n8083), .A(n6019), .ZN(n8096) );
  OAI21_X2 U5399 ( .B1(n8196), .B2(n8195), .A(n6011), .ZN(n8230) );
  OAI21_X2 U5400 ( .B1(n8216), .B2(n8215), .A(n6019), .ZN(n8228) );
  OAI21_X2 U5401 ( .B1(n8226), .B2(n8225), .A(net77290), .ZN(n8227) );
  OAI21_X2 U5402 ( .B1(n8108), .B2(n8107), .A(n6011), .ZN(n8142) );
  OAI21_X2 U5403 ( .B1(n8118), .B2(n8117), .A(net77588), .ZN(n8141) );
  OAI21_X1 U5404 ( .B1(n8128), .B2(n8127), .A(n6019), .ZN(n8140) );
  OAI21_X2 U5405 ( .B1(n8020), .B2(n8019), .A(n6011), .ZN(n8054) );
  OAI21_X1 U5406 ( .B1(n8030), .B2(n8029), .A(net77588), .ZN(n8053) );
  OAI21_X2 U5407 ( .B1(n8040), .B2(n8039), .A(n6019), .ZN(n8052) );
  OAI21_X2 U5408 ( .B1(n7976), .B2(n7975), .A(n6011), .ZN(n8010) );
  OAI21_X2 U5409 ( .B1(n7986), .B2(n7985), .A(net77588), .ZN(n8009) );
  OAI21_X2 U5410 ( .B1(n7996), .B2(n7995), .A(n6019), .ZN(n8008) );
  OAI21_X1 U5411 ( .B1(n7626), .B2(n7625), .A(n6012), .ZN(n7660) );
  OAI21_X1 U5412 ( .B1(n7636), .B2(n7635), .A(net77588), .ZN(n7659) );
  OAI21_X1 U5413 ( .B1(n7656), .B2(n7655), .A(net77292), .ZN(n7657) );
  OAI21_X1 U5414 ( .B1(n7582), .B2(n7581), .A(n6012), .ZN(n7616) );
  OAI21_X1 U5415 ( .B1(n7592), .B2(n7591), .A(net77588), .ZN(n7615) );
  OAI21_X1 U5416 ( .B1(n7612), .B2(n7611), .A(net77292), .ZN(n7613) );
  OAI21_X1 U5417 ( .B1(n7548), .B2(n7547), .A(net77588), .ZN(n7571) );
  OAI21_X1 U5418 ( .B1(n7558), .B2(n7557), .A(n6019), .ZN(n7570) );
  OAI21_X1 U5419 ( .B1(n7768), .B2(n7767), .A(net77588), .ZN(n7791) );
  OAI21_X1 U5420 ( .B1(n7758), .B2(n7757), .A(n6011), .ZN(n7792) );
  OAI21_X1 U5421 ( .B1(n7788), .B2(n7787), .A(net77290), .ZN(n7789) );
  NOR2_X2 U5422 ( .A1(n8661), .A2(n8660), .ZN(n8666) );
  OAI21_X2 U5423 ( .B1(n7095), .B2(n7094), .A(n6011), .ZN(n7129) );
  OAI21_X2 U5424 ( .B1(n7105), .B2(n7104), .A(net77588), .ZN(n7128) );
  OAI21_X2 U5425 ( .B1(n7115), .B2(n7114), .A(n6019), .ZN(n7127) );
  NAND4_X2 U5426 ( .A1(n7085), .A2(n7084), .A3(n7083), .A4(n7082), .ZN(n8450)
         );
  OAI21_X1 U5427 ( .B1(n7496), .B2(n7495), .A(n6012), .ZN(n7528) );
  OAI21_X1 U5428 ( .B1(n7506), .B2(n7505), .A(net77588), .ZN(n7527) );
  OAI21_X1 U5429 ( .B1(n7515), .B2(n7514), .A(n6019), .ZN(n7526) );
  NOR2_X2 U5430 ( .A1(n10000), .A2(n8949), .ZN(n8954) );
  OAI21_X2 U5431 ( .B1(n7274), .B2(n7273), .A(n6012), .ZN(n7308) );
  OAI21_X1 U5432 ( .B1(n7284), .B2(n7283), .A(net77292), .ZN(n7307) );
  OAI21_X1 U5433 ( .B1(n7294), .B2(n7293), .A(n6019), .ZN(n7306) );
  NOR2_X2 U5434 ( .A1(net77999), .A2(n5597), .ZN(net72876) );
  AOI21_X1 U5435 ( .B1(n9041), .B2(net77030), .A(n9040), .ZN(n9042) );
  NOR2_X2 U5436 ( .A1(net76464), .A2(n9039), .ZN(n9040) );
  AOI21_X2 U5437 ( .B1(dmem_read_in[0]), .B2(n4911), .A(n10000), .ZN(n9204) );
  AOI222_X2 U5438 ( .A1(net76650), .A2(dmem_addr_out[16]), .B1(
        dmem_read_in[16]), .B2(dmem_dsize[0]), .C1(n9203), .C2(net77030), .ZN(
        n9205) );
  OAI21_X2 U5439 ( .B1(n7408), .B2(n7407), .A(n6012), .ZN(n7442) );
  OAI21_X2 U5440 ( .B1(n7418), .B2(n7417), .A(net77588), .ZN(n7441) );
  OAI21_X2 U5441 ( .B1(n7438), .B2(n7437), .A(net77292), .ZN(n7439) );
  OAI21_X1 U5442 ( .B1(n7364), .B2(n7363), .A(n6012), .ZN(n7398) );
  OAI21_X1 U5443 ( .B1(n7374), .B2(n7373), .A(net77588), .ZN(n7397) );
  OAI21_X1 U5444 ( .B1(n7384), .B2(n7383), .A(n6019), .ZN(n7396) );
  NOR2_X2 U5445 ( .A1(n10000), .A2(n9313), .ZN(n9318) );
  AOI21_X2 U5446 ( .B1(n9375), .B2(net77030), .A(n9374), .ZN(n9376) );
  NOR2_X2 U5447 ( .A1(n10000), .A2(n9566), .ZN(n9571) );
  INV_X8 U5448 ( .A(n9800), .ZN(n6064) );
  NOR2_X2 U5449 ( .A1(n9788), .A2(net71906), .ZN(n9793) );
  INV_X16 U5450 ( .A(n10090), .ZN(n6077) );
  NOR2_X2 U5451 ( .A1(n10504), .A2(net76464), .ZN(n10293) );
  NAND3_X2 U5452 ( .A1(n4907), .A2(net73429), .A3(net73443), .ZN(n8677) );
  NAND4_X2 U5453 ( .A1(n6488), .A2(n6489), .A3(n6487), .A4(n6486), .ZN(n6490)
         );
  AOI22_X2 U5454 ( .A1(REGFILE_reg_out_7__8_), .A2(net77716), .B1(
        REGFILE_reg_out_6__8_), .B2(net75456), .ZN(n6745) );
  AOI22_X2 U5455 ( .A1(REGFILE_reg_out_26__6_), .A2(net77618), .B1(
        REGFILE_reg_out_27__6_), .B2(net77626), .ZN(n6779) );
  NOR3_X1 U5456 ( .A1(n8729), .A2(net71026), .A3(net78003), .ZN(n8730) );
  NOR2_X1 U5457 ( .A1(n4812), .A2(n9854), .ZN(n8718) );
  NOR3_X1 U5458 ( .A1(net78003), .A2(n10099), .A3(n10312), .ZN(n9806) );
  NOR2_X1 U5459 ( .A1(n10442), .A2(net78014), .ZN(n9811) );
  OAI21_X1 U5460 ( .B1(n9804), .B2(n10472), .A(n8764), .ZN(n8770) );
  NOR2_X1 U5461 ( .A1(n8601), .A2(net78014), .ZN(n8602) );
  NOR2_X1 U5462 ( .A1(n10336), .A2(net78014), .ZN(n9291) );
  NOR3_X1 U5463 ( .A1(n9306), .A2(n10334), .A3(net78003), .ZN(n9307) );
  NOR2_X1 U5464 ( .A1(n8921), .A2(net78014), .ZN(n8922) );
  NOR3_X1 U5465 ( .A1(n10338), .A2(n8967), .A3(net78003), .ZN(n8943) );
  NOR2_X1 U5466 ( .A1(n10343), .A2(net78014), .ZN(n9544) );
  NOR2_X1 U5467 ( .A1(n8833), .A2(net70710), .ZN(n8834) );
  AOI21_X2 U5468 ( .B1(n8863), .B2(n8862), .A(net72163), .ZN(n8864) );
  OAI21_X2 U5469 ( .B1(n8848), .B2(n9606), .A(n8847), .ZN(n8866) );
  OAI21_X2 U5470 ( .B1(n9414), .B2(n9854), .A(n9413), .ZN(n9415) );
  NOR2_X1 U5471 ( .A1(net70710), .A2(n9366), .ZN(n9367) );
  NOR2_X2 U5472 ( .A1(n9606), .A2(n9348), .ZN(n9350) );
  NOR2_X1 U5473 ( .A1(n10418), .A2(net78014), .ZN(n9349) );
  NOR2_X1 U5474 ( .A1(net70710), .A2(n9626), .ZN(n9627) );
  INV_X4 U5475 ( .A(net70691), .ZN(net71271) );
  NOR2_X2 U5476 ( .A1(n9606), .A2(n9605), .ZN(n9608) );
  NOR3_X1 U5477 ( .A1(net73630), .A2(n5605), .A3(net73532), .ZN(n5602) );
  NOR2_X1 U5478 ( .A1(n5604), .A2(net73629), .ZN(n5603) );
  NAND3_X2 U5479 ( .A1(net105361), .A2(n5637), .A3(n5636), .ZN(net105376) );
  AOI21_X2 U5480 ( .B1(n5710), .B2(net70701), .A(n4809), .ZN(net105361) );
  NOR2_X2 U5481 ( .A1(n10000), .A2(net73166), .ZN(n8875) );
  AOI21_X2 U5482 ( .B1(n8873), .B2(net77030), .A(n8872), .ZN(n8874) );
  NOR2_X2 U5483 ( .A1(n10000), .A2(n9999), .ZN(n10005) );
  AOI21_X1 U5484 ( .B1(n10003), .B2(net77030), .A(n10002), .ZN(n10004) );
  NOR2_X2 U5485 ( .A1(n5592), .A2(net70531), .ZN(net70529) );
  OAI21_X2 U5486 ( .B1(n8479), .B2(n8480), .A(n8395), .ZN(n8473) );
  OAI21_X2 U5487 ( .B1(n8493), .B2(n8494), .A(n8386), .ZN(n8487) );
  OAI21_X1 U5488 ( .B1(n4908), .B2(n8308), .A(n5060), .ZN(n8304) );
  OAI21_X2 U5489 ( .B1(n9107), .B2(n8372), .A(n8523), .ZN(n8373) );
  NOR2_X2 U5490 ( .A1(n8739), .A2(n8738), .ZN(n8740) );
  NOR2_X2 U5491 ( .A1(n8785), .A2(n8784), .ZN(n8790) );
  INV_X4 U5492 ( .A(n5002), .ZN(n6172) );
  OAI21_X2 U5493 ( .B1(n8502), .B2(n8503), .A(n8366), .ZN(n9388) );
  INV_X4 U5494 ( .A(n4992), .ZN(net76660) );
  INV_X4 U5495 ( .A(n4994), .ZN(n6158) );
  INV_X4 U5496 ( .A(n4999), .ZN(n6160) );
  INV_X4 U5497 ( .A(n5000), .ZN(n6162) );
  INV_X4 U5498 ( .A(n4997), .ZN(net76616) );
  INV_X4 U5499 ( .A(n4903), .ZN(n6208) );
  INV_X4 U5500 ( .A(n4904), .ZN(n6164) );
  INV_X4 U5501 ( .A(n4905), .ZN(n6166) );
  INV_X4 U5502 ( .A(n4906), .ZN(n6168) );
  INV_X4 U5503 ( .A(n4995), .ZN(n6170) );
  INV_X4 U5504 ( .A(n5003), .ZN(n6174) );
  INV_X4 U5505 ( .A(n5005), .ZN(net76550) );
  INV_X4 U5506 ( .A(n4996), .ZN(n6220) );
  INV_X4 U5507 ( .A(n5006), .ZN(n6183) );
  INV_X4 U5508 ( .A(n5007), .ZN(n6185) );
  INV_X4 U5509 ( .A(n4991), .ZN(n6187) );
  INV_X4 U5510 ( .A(n5008), .ZN(n6189) );
  INV_X4 U5511 ( .A(n4993), .ZN(n6199) );
  INV_X4 U5512 ( .A(n4998), .ZN(n6195) );
  INV_X4 U5513 ( .A(n5001), .ZN(n6204) );
  INV_X4 U5514 ( .A(n5004), .ZN(n6212) );
  INV_X4 U5515 ( .A(n5009), .ZN(net76320) );
  AOI21_X1 U5516 ( .B1(n9700), .B2(net77030), .A(n9699), .ZN(n9701) );
  NOR2_X2 U5517 ( .A1(n9819), .A2(n9818), .ZN(n9824) );
  INV_X4 U5518 ( .A(n4992), .ZN(net76658) );
  INV_X4 U5519 ( .A(n4990), .ZN(n6155) );
  INV_X4 U5520 ( .A(n4998), .ZN(n6194) );
  INV_X4 U5521 ( .A(n4993), .ZN(n6198) );
  INV_X4 U5522 ( .A(n4994), .ZN(n6157) );
  INV_X4 U5523 ( .A(n4999), .ZN(n6159) );
  INV_X4 U5524 ( .A(n5000), .ZN(n6161) );
  INV_X4 U5525 ( .A(n5001), .ZN(n6203) );
  INV_X4 U5526 ( .A(n4997), .ZN(net76614) );
  INV_X4 U5527 ( .A(n4903), .ZN(n6207) );
  INV_X4 U5528 ( .A(n4904), .ZN(n6163) );
  INV_X4 U5529 ( .A(n4905), .ZN(n6165) );
  INV_X4 U5530 ( .A(n4906), .ZN(n6167) );
  INV_X4 U5531 ( .A(n4995), .ZN(n6169) );
  INV_X4 U5532 ( .A(n5002), .ZN(n6171) );
  INV_X4 U5533 ( .A(n5003), .ZN(n6173) );
  INV_X4 U5534 ( .A(n5004), .ZN(n6211) );
  INV_X4 U5535 ( .A(n4806), .ZN(n6214) );
  INV_X4 U5536 ( .A(n5005), .ZN(net76548) );
  INV_X4 U5537 ( .A(n5009), .ZN(net76318) );
  INV_X4 U5538 ( .A(n4996), .ZN(n6219) );
  INV_X4 U5539 ( .A(n5006), .ZN(n6182) );
  INV_X4 U5540 ( .A(n5007), .ZN(n6184) );
  INV_X4 U5541 ( .A(n4991), .ZN(n6186) );
  INV_X4 U5542 ( .A(n5008), .ZN(n6188) );
  NAND2_X2 U5543 ( .A1(n6829), .A2(n6828), .ZN(dmem_write_out[4]) );
  NOR2_X1 U5544 ( .A1(n6005), .A2(n10312), .ZN(n10313) );
  NAND3_X2 U5545 ( .A1(net73509), .A2(instruction[26]), .A3(net73696), .ZN(
        net73620) );
  INV_X4 U5546 ( .A(net77336), .ZN(net77360) );
  NAND3_X2 U5547 ( .A1(n10440), .A2(n10439), .A3(n10438), .ZN(n10451) );
  NAND3_X2 U5548 ( .A1(n8637), .A2(n9499), .A3(n8627), .ZN(n8892) );
  NOR2_X1 U5549 ( .A1(n8655), .A2(n8565), .ZN(n8566) );
  NAND3_X2 U5550 ( .A1(n8576), .A2(net73498), .A3(net73503), .ZN(n8535) );
  OAI21_X1 U5551 ( .B1(n7744), .B2(n7743), .A(net77292), .ZN(n7745) );
  NAND4_X2 U5552 ( .A1(n7011), .A2(n7010), .A3(n7009), .A4(n7008), .ZN(n7017)
         );
  NOR2_X1 U5553 ( .A1(instruction[2]), .A2(net73499), .ZN(net73504) );
  NAND4_X2 U5554 ( .A1(net75859), .A2(net75861), .A3(net75862), .A4(net75860), 
        .ZN(net75858) );
  OAI21_X1 U5555 ( .B1(net70868), .B2(n10247), .A(n9076), .ZN(n8708) );
  NOR2_X1 U5556 ( .A1(net70866), .A2(n9656), .ZN(n8709) );
  NAND3_X2 U5557 ( .A1(n9343), .A2(n8724), .A3(n8723), .ZN(n8978) );
  OAI21_X2 U5558 ( .B1(n6005), .B2(n8936), .A(n8935), .ZN(n9302) );
  NAND3_X1 U5559 ( .A1(n9070), .A2(n9069), .A3(n9068), .ZN(n9838) );
  NAND3_X1 U5560 ( .A1(n9341), .A2(n9340), .A3(n9339), .ZN(n9839) );
  OAI21_X2 U5561 ( .B1(n8576), .B2(net73637), .A(instruction[5]), .ZN(n8577)
         );
  OAI21_X2 U5562 ( .B1(net73638), .B2(net73616), .A(instruction[31]), .ZN(
        n8578) );
  OAI21_X2 U5563 ( .B1(n9959), .B2(n9958), .A(n9957), .ZN(n10035) );
  NOR2_X1 U5564 ( .A1(n10093), .A2(n9606), .ZN(n10029) );
  NOR2_X2 U5565 ( .A1(n9941), .A2(n9940), .ZN(n9942) );
  OAI21_X2 U5566 ( .B1(n8182), .B2(n8181), .A(net77290), .ZN(n8183) );
  OAI21_X1 U5567 ( .B1(n8094), .B2(n8093), .A(net77290), .ZN(n8095) );
  OAI21_X2 U5568 ( .B1(n8206), .B2(n8205), .A(net77588), .ZN(n8229) );
  OAI21_X2 U5569 ( .B1(n8138), .B2(n8137), .A(net77290), .ZN(n8139) );
  OAI21_X2 U5570 ( .B1(n8050), .B2(n8049), .A(net77290), .ZN(n8051) );
  OAI21_X2 U5571 ( .B1(n8006), .B2(n8005), .A(net77290), .ZN(n8007) );
  OAI21_X1 U5572 ( .B1(n7646), .B2(n7645), .A(n6019), .ZN(n7658) );
  OAI21_X1 U5573 ( .B1(n7602), .B2(n7601), .A(n6019), .ZN(n7614) );
  OAI21_X1 U5574 ( .B1(n7568), .B2(n7567), .A(net77292), .ZN(n7569) );
  OAI21_X1 U5575 ( .B1(n7778), .B2(n7777), .A(n6019), .ZN(n7790) );
  NOR2_X2 U5576 ( .A1(net77999), .A2(n9516), .ZN(n8661) );
  NOR2_X2 U5577 ( .A1(net70811), .A2(n10540), .ZN(n8660) );
  AOI21_X2 U5578 ( .B1(n8664), .B2(net77030), .A(n8663), .ZN(n8665) );
  NOR2_X2 U5579 ( .A1(net76464), .A2(n8662), .ZN(n8663) );
  OAI21_X1 U5580 ( .B1(n7524), .B2(n7523), .A(net77292), .ZN(n7525) );
  OAI21_X1 U5581 ( .B1(n7472), .B2(n7471), .A(n6019), .ZN(n7484) );
  NOR2_X2 U5582 ( .A1(net77999), .A2(n9669), .ZN(n8949) );
  AOI21_X2 U5583 ( .B1(n8964), .B2(net77030), .A(n8952), .ZN(n8953) );
  NOR2_X2 U5584 ( .A1(net76464), .A2(n8951), .ZN(n8952) );
  OAI21_X1 U5585 ( .B1(n7304), .B2(n7303), .A(net77588), .ZN(n7305) );
  NOR2_X2 U5586 ( .A1(net76464), .A2(n9108), .ZN(n9109) );
  OAI21_X1 U5587 ( .B1(n7394), .B2(n7393), .A(net77292), .ZN(n7395) );
  NOR2_X2 U5588 ( .A1(net77999), .A2(n10505), .ZN(n9313) );
  AOI21_X1 U5589 ( .B1(n9316), .B2(net77030), .A(n9315), .ZN(n9317) );
  NOR2_X2 U5590 ( .A1(net76464), .A2(n9314), .ZN(n9315) );
  NOR2_X2 U5591 ( .A1(net76464), .A2(n9373), .ZN(n9374) );
  OAI21_X1 U5592 ( .B1(n7690), .B2(n7689), .A(n6019), .ZN(n7702) );
  AOI21_X2 U5593 ( .B1(n9422), .B2(net77030), .A(n9421), .ZN(n9423) );
  NOR2_X2 U5594 ( .A1(net76464), .A2(n9816), .ZN(n9421) );
  NOR2_X2 U5595 ( .A1(net76464), .A2(n9516), .ZN(n9517) );
  NOR2_X2 U5596 ( .A1(net77999), .A2(n9817), .ZN(n9566) );
  AOI21_X1 U5597 ( .B1(n9569), .B2(net77030), .A(n9568), .ZN(n9570) );
  NOR2_X2 U5598 ( .A1(net76464), .A2(n9567), .ZN(n9568) );
  NOR2_X2 U5599 ( .A1(net76464), .A2(n9817), .ZN(n9633) );
  NOR2_X2 U5600 ( .A1(net76464), .A2(n9669), .ZN(n9670) );
  NOR2_X2 U5601 ( .A1(net77999), .A2(n10137), .ZN(n9788) );
  NOR2_X2 U5602 ( .A1(net70811), .A2(n5694), .ZN(net71906) );
  AOI21_X1 U5603 ( .B1(n9791), .B2(net77030), .A(n9790), .ZN(n9792) );
  NOR2_X2 U5604 ( .A1(net76464), .A2(n9789), .ZN(n9790) );
  AOI21_X1 U5605 ( .B1(n9864), .B2(net77030), .A(n9863), .ZN(n9865) );
  NOR2_X2 U5606 ( .A1(net76464), .A2(n9862), .ZN(n9863) );
  NOR2_X2 U5607 ( .A1(net76464), .A2(n10083), .ZN(n9964) );
  NOR2_X2 U5608 ( .A1(net76464), .A2(n10041), .ZN(n10042) );
  NOR2_X2 U5609 ( .A1(net76464), .A2(n5694), .ZN(n5693) );
  NOR2_X2 U5610 ( .A1(net76464), .A2(n10137), .ZN(n10138) );
  NOR2_X1 U5611 ( .A1(n10484), .A2(net77040), .ZN(n10458) );
  AOI21_X2 U5612 ( .B1(n10495), .B2(n10494), .A(n10493), .ZN(n10496) );
  NOR2_X1 U5613 ( .A1(n10494), .A2(net77040), .ZN(n10492) );
  AOI21_X1 U5614 ( .B1(n10484), .B2(net77042), .A(n10494), .ZN(n10488) );
  NOR2_X2 U5615 ( .A1(n8575), .A2(n8581), .ZN(n8556) );
  NAND3_X2 U5616 ( .A1(n8619), .A2(n8618), .A3(n8617), .ZN(n9294) );
  NAND3_X2 U5617 ( .A1(n9981), .A2(n9980), .A3(n9979), .ZN(n10057) );
  NAND3_X2 U5618 ( .A1(n9551), .A2(n9550), .A3(n9549), .ZN(n10059) );
  AOI21_X1 U5619 ( .B1(net71085), .B2(n9182), .A(n9023), .ZN(n9024) );
  AOI21_X1 U5620 ( .B1(net71085), .B2(n10282), .A(n5058), .ZN(n10283) );
  AOI21_X2 U5621 ( .B1(net71085), .B2(n10248), .A(n5057), .ZN(n10249) );
  NAND3_X1 U5622 ( .A1(n9067), .A2(n9066), .A3(n10462), .ZN(n10239) );
  OAI21_X2 U5623 ( .B1(n9094), .B2(n10327), .A(n9017), .ZN(n10238) );
  OAI21_X2 U5624 ( .B1(n9094), .B2(net72312), .A(n9082), .ZN(n9395) );
  AOI21_X1 U5625 ( .B1(net71085), .B2(n10126), .A(n5056), .ZN(n10127) );
  AOI21_X2 U5626 ( .B1(net71085), .B2(n9685), .A(n5051), .ZN(n9503) );
  NAND3_X1 U5627 ( .A1(n9361), .A2(n9360), .A3(n9359), .ZN(n9945) );
  NAND3_X1 U5628 ( .A1(n9078), .A2(n9077), .A3(n9076), .ZN(n9500) );
  NAND3_X2 U5629 ( .A1(n9588), .A2(n9587), .A3(n9586), .ZN(n9655) );
  AOI21_X1 U5630 ( .B1(net77084), .B2(n9585), .A(n5015), .ZN(n9586) );
  AOI21_X1 U5631 ( .B1(net71085), .B2(n10016), .A(n5055), .ZN(n9950) );
  INV_X8 U5632 ( .A(net78003), .ZN(net71078) );
  NOR2_X1 U5633 ( .A1(net70709), .A2(n9606), .ZN(net71280) );
  AOI222_X1 U5634 ( .A1(n6083), .A2(n10103), .B1(n10102), .B2(n10541), .C1(
        net70713), .C2(net71026), .ZN(n10152) );
  OAI21_X1 U5635 ( .B1(net71299), .B2(net70718), .A(net71300), .ZN(n10151) );
  AOI21_X2 U5636 ( .B1(n5638), .B2(net70727), .A(net76452), .ZN(net70693) );
  OAI21_X1 U5637 ( .B1(net71027), .B2(net105349), .A(net72163), .ZN(n5712) );
  OAI21_X2 U5638 ( .B1(n7890), .B2(n7889), .A(n6011), .ZN(n7924) );
  OAI21_X1 U5639 ( .B1(n7900), .B2(n7899), .A(net77588), .ZN(n7923) );
  OAI21_X1 U5640 ( .B1(n7910), .B2(n7909), .A(n6019), .ZN(n7922) );
  NOR2_X2 U5641 ( .A1(net76464), .A2(n8871), .ZN(n8872) );
  NOR2_X2 U5642 ( .A1(net77999), .A2(n5694), .ZN(net73166) );
  NOR2_X2 U5643 ( .A1(net76464), .A2(n10001), .ZN(n10002) );
  NOR2_X2 U5644 ( .A1(net77999), .A2(n10041), .ZN(n9999) );
  OAI21_X2 U5645 ( .B1(n7934), .B2(n7933), .A(n6011), .ZN(n7966) );
  OAI21_X2 U5646 ( .B1(n7944), .B2(n7943), .A(net77588), .ZN(n7965) );
  OAI21_X2 U5647 ( .B1(n7954), .B2(n7953), .A(n6019), .ZN(n7964) );
  OAI21_X2 U5648 ( .B1(net76464), .B2(n5597), .A(net70740), .ZN(n5596) );
  AOI21_X1 U5649 ( .B1(net73878), .B2(n8295), .A(net73997), .ZN(n8385) );
  INV_X4 U5650 ( .A(net70531), .ZN(net73858) );
  OAI21_X2 U5651 ( .B1(n7846), .B2(n7845), .A(n6011), .ZN(n7880) );
  OAI21_X1 U5652 ( .B1(n7856), .B2(n7855), .A(net77588), .ZN(n7879) );
  OAI21_X1 U5653 ( .B1(n7866), .B2(n7865), .A(n6019), .ZN(n7878) );
  NAND4_X2 U5654 ( .A1(n6996), .A2(n6995), .A3(n6997), .A4(n6994), .ZN(n5936)
         );
  NOR2_X2 U5655 ( .A1(net76464), .A2(n8737), .ZN(n8738) );
  NOR2_X2 U5656 ( .A1(n5014), .A2(net70738), .ZN(n8739) );
  NOR2_X2 U5657 ( .A1(net77999), .A2(n9108), .ZN(n8785) );
  NOR2_X2 U5658 ( .A1(net70811), .A2(n10083), .ZN(n8784) );
  AOI21_X1 U5659 ( .B1(n8788), .B2(net77030), .A(n8787), .ZN(n8789) );
  NOR2_X2 U5660 ( .A1(net76464), .A2(n8786), .ZN(n8787) );
  AOI21_X1 U5661 ( .B1(n8908), .B2(net77030), .A(n8907), .ZN(n8909) );
  NOR2_X2 U5662 ( .A1(net76464), .A2(n8906), .ZN(n8907) );
  NOR2_X2 U5663 ( .A1(n8905), .A2(n8904), .ZN(n8910) );
  NOR2_X2 U5664 ( .A1(net70811), .A2(n10041), .ZN(n8904) );
  NOR2_X2 U5665 ( .A1(net77999), .A2(n9862), .ZN(n8905) );
  INV_X8 U5666 ( .A(n9009), .ZN(n6031) );
  NOR2_X2 U5667 ( .A1(n8997), .A2(net72947), .ZN(n9002) );
  OAI21_X2 U5668 ( .B1(n7802), .B2(n7801), .A(n6011), .ZN(n7836) );
  OAI21_X1 U5669 ( .B1(n7812), .B2(n7811), .A(net77588), .ZN(n7835) );
  OAI21_X2 U5670 ( .B1(n7832), .B2(n7831), .A(net77290), .ZN(n7833) );
  OAI21_X1 U5671 ( .B1(net73519), .B2(n8461), .A(net73780), .ZN(n8463) );
  NOR2_X2 U5672 ( .A1(n10505), .A2(net76464), .ZN(n9699) );
  NOR2_X2 U5673 ( .A1(net77999), .A2(n9816), .ZN(n9819) );
  NOR2_X2 U5674 ( .A1(net70811), .A2(n9817), .ZN(n9818) );
  NOR2_X2 U5675 ( .A1(n9822), .A2(n9821), .ZN(n9823) );
  NOR2_X1 U5676 ( .A1(instructionAddr_out[29]), .A2(net70738), .ZN(n9822) );
  NOR2_X2 U5677 ( .A1(net76464), .A2(n9820), .ZN(n9821) );
  OAI21_X1 U5678 ( .B1(net73496), .B2(net73780), .A(reset), .ZN(n10650) );
  NOR2_X2 U5679 ( .A1(net76646), .A2(n10503), .ZN(n10508) );
  NOR2_X2 U5680 ( .A1(net77999), .A2(n10504), .ZN(n10507) );
  NOR2_X2 U5681 ( .A1(net70811), .A2(n10505), .ZN(n10506) );
  NOR2_X1 U5682 ( .A1(net73503), .A2(net73499), .ZN(n8658) );
  NOR2_X1 U5683 ( .A1(net73498), .A2(net73499), .ZN(n8659) );
  NAND3_X1 U5684 ( .A1(n8655), .A2(net73170), .A3(n8654), .ZN(net70506) );
  NOR2_X2 U5685 ( .A1(instruction[1]), .A2(n8653), .ZN(n8654) );
  NAND4_X2 U5686 ( .A1(n6575), .A2(n6574), .A3(n6572), .A4(n6573), .ZN(n6581)
         );
  AOI22_X2 U5687 ( .A1(REGFILE_reg_out_19__15_), .A2(net77812), .B1(
        REGFILE_reg_out_1__15_), .B2(net75478), .ZN(n6585) );
  NAND3_X2 U5688 ( .A1(n10107), .A2(n5042), .A3(n10106), .ZN(n10108) );
  AOI21_X1 U5689 ( .B1(n10261), .B2(net77030), .A(n10260), .ZN(n10262) );
  NOR2_X2 U5690 ( .A1(net76464), .A2(n10259), .ZN(n10260) );
  NOR2_X2 U5691 ( .A1(n10000), .A2(net72876), .ZN(n9043) );
  INV_X4 U5692 ( .A(n4878), .ZN(n6132) );
  INV_X4 U5693 ( .A(n4867), .ZN(n6088) );
  INV_X4 U5694 ( .A(n4990), .ZN(n6156) );
  INV_X4 U5695 ( .A(n6093), .ZN(n6091) );
  INV_X4 U5696 ( .A(n6100), .ZN(n6097) );
  INV_X4 U5697 ( .A(n4804), .ZN(n6108) );
  INV_X4 U5698 ( .A(n4891), .ZN(n6112) );
  INV_X4 U5699 ( .A(n4892), .ZN(n6115) );
  INV_X4 U5700 ( .A(n4884), .ZN(n6118) );
  INV_X4 U5701 ( .A(n4877), .ZN(net76862) );
  INV_X4 U5702 ( .A(n4882), .ZN(n6121) );
  INV_X4 U5703 ( .A(n4888), .ZN(n6124) );
  INV_X4 U5704 ( .A(n4883), .ZN(n6127) );
  INV_X4 U5705 ( .A(n4875), .ZN(n6129) );
  INV_X4 U5706 ( .A(n4893), .ZN(n6136) );
  INV_X4 U5707 ( .A(n4879), .ZN(n6139) );
  INV_X4 U5708 ( .A(n4885), .ZN(n6144) );
  INV_X4 U5709 ( .A(n4889), .ZN(net76706) );
  INV_X4 U5710 ( .A(n4886), .ZN(net76692) );
  INV_X4 U5711 ( .A(n4890), .ZN(n6150) );
  INV_X4 U5712 ( .A(n4887), .ZN(n6153) );
  INV_X4 U5713 ( .A(n4876), .ZN(n6200) );
  INV_X4 U5714 ( .A(n4876), .ZN(n6202) );
  INV_X4 U5715 ( .A(n4867), .ZN(n6089) );
  INV_X4 U5716 ( .A(n6093), .ZN(n6092) );
  INV_X4 U5717 ( .A(n6100), .ZN(n6098) );
  INV_X4 U5718 ( .A(n4804), .ZN(n6109) );
  INV_X4 U5719 ( .A(n4891), .ZN(n6113) );
  INV_X4 U5720 ( .A(n4892), .ZN(n6116) );
  INV_X4 U5721 ( .A(n4884), .ZN(n6119) );
  INV_X4 U5722 ( .A(n4877), .ZN(net76864) );
  INV_X4 U5723 ( .A(n4882), .ZN(n6122) );
  INV_X4 U5724 ( .A(n4888), .ZN(n6125) );
  INV_X4 U5725 ( .A(n4883), .ZN(n6128) );
  INV_X4 U5726 ( .A(n4875), .ZN(n6130) );
  INV_X4 U5727 ( .A(n4878), .ZN(n6133) );
  INV_X4 U5728 ( .A(n4893), .ZN(n6137) );
  INV_X4 U5729 ( .A(n4879), .ZN(n6140) );
  INV_X4 U5730 ( .A(n4885), .ZN(n6145) );
  INV_X4 U5731 ( .A(n4889), .ZN(net76708) );
  INV_X4 U5732 ( .A(n4886), .ZN(net76694) );
  INV_X4 U5733 ( .A(n4890), .ZN(n6151) );
  INV_X4 U5734 ( .A(n4887), .ZN(n6154) );
  AOI21_X1 U5735 ( .B1(n10294), .B2(net77030), .A(n10293), .ZN(n10295) );
  INV_X4 U5736 ( .A(n4867), .ZN(n6090) );
  INV_X4 U5737 ( .A(n6100), .ZN(n6099) );
  INV_X4 U5738 ( .A(n6096), .ZN(n6094) );
  INV_X4 U5739 ( .A(n4804), .ZN(n6110) );
  INV_X4 U5740 ( .A(n6107), .ZN(n6105) );
  INV_X4 U5741 ( .A(n4876), .ZN(n6201) );
  INV_X4 U5742 ( .A(n4877), .ZN(net76866) );
  INV_X4 U5743 ( .A(n4875), .ZN(n6131) );
  INV_X4 U5744 ( .A(n4878), .ZN(n6134) );
  INV_X4 U5745 ( .A(n4879), .ZN(n6141) );
  INV_X4 U5746 ( .A(n6148), .ZN(n6146) );
  NOR2_X2 U5747 ( .A1(n6190), .A2(n10651), .ZN(n10652) );
  NOR2_X2 U5748 ( .A1(instruction[31]), .A2(n10650), .ZN(n10651) );
  NAND2_X2 U5749 ( .A1(n6408), .A2(n6407), .ZN(dmem_write_out[24]) );
  NAND2_X2 U5750 ( .A1(n6454), .A2(n6455), .ZN(dmem_write_out[22]) );
  NAND2_X2 U5751 ( .A1(n6479), .A2(n6478), .ZN(dmem_write_out[21]) );
  NAND2_X2 U5752 ( .A1(n6503), .A2(n6502), .ZN(n10944) );
  NAND2_X2 U5753 ( .A1(n6753), .A2(n6752), .ZN(dmem_write_out[8]) );
  NAND2_X2 U5754 ( .A1(n6850), .A2(n6851), .ZN(dmem_write_out[3]) );
  NAND2_X2 U5755 ( .A1(n6895), .A2(n6894), .ZN(dmem_write_out[1]) );
  NAND3_X2 U5756 ( .A1(n8734), .A2(n8733), .A3(n8732), .ZN(n8735) );
  NAND3_X2 U5757 ( .A1(n9815), .A2(n9814), .A3(n9813), .ZN(dmem_addr_out[29])
         );
  AOI21_X2 U5758 ( .B1(net71271), .B2(n9812), .A(n9811), .ZN(n9813) );
  OAI21_X2 U5759 ( .B1(n8770), .B2(n8769), .A(net70697), .ZN(n8782) );
  OAI21_X1 U5760 ( .B1(n8900), .B2(n8899), .A(net70697), .ZN(n8902) );
  AOI21_X2 U5761 ( .B1(net71271), .B2(n8889), .A(n8888), .ZN(n8903) );
  OAI21_X1 U5762 ( .B1(n9773), .B2(n9772), .A(net70697), .ZN(n9786) );
  AOI21_X2 U5763 ( .B1(n9784), .B2(n9783), .A(n9782), .ZN(n9785) );
  AOI21_X2 U5764 ( .B1(net71271), .B2(n8603), .A(n8602), .ZN(n8649) );
  AOI21_X2 U5765 ( .B1(net71271), .B2(n9292), .A(n9291), .ZN(n9312) );
  AOI21_X2 U5766 ( .B1(net71271), .B2(n8923), .A(n8922), .ZN(n8948) );
  AOI21_X2 U5767 ( .B1(net71271), .B2(n9545), .A(n9544), .ZN(n9565) );
  AOI21_X2 U5768 ( .B1(net71271), .B2(n8835), .A(n8834), .ZN(n8869) );
  AOI21_X1 U5769 ( .B1(n10064), .B2(n9182), .A(n9181), .ZN(n9200) );
  NOR2_X2 U5770 ( .A1(n9198), .A2(n9197), .ZN(n9199) );
  AOI21_X1 U5771 ( .B1(n10064), .B2(n10248), .A(n5050), .ZN(n9418) );
  AOI21_X1 U5772 ( .B1(n10064), .B2(n9403), .A(n5049), .ZN(n9104) );
  AOI21_X1 U5773 ( .B1(n10064), .B2(n9837), .A(n5054), .ZN(n9859) );
  AOI21_X1 U5774 ( .B1(net70697), .B2(n9338), .A(n9337), .ZN(n9372) );
  AOI21_X2 U5775 ( .B1(net71271), .B2(n9368), .A(n9367), .ZN(n9369) );
  AOI21_X1 U5776 ( .B1(n10064), .B2(n9685), .A(n5053), .ZN(n9696) );
  AOI21_X2 U5777 ( .B1(net71271), .B2(n9628), .A(n9627), .ZN(n9629) );
  AOI21_X1 U5778 ( .B1(n10649), .B2(n10642), .A(n6190), .ZN(n10646) );
  NOR2_X2 U5779 ( .A1(net73855), .A2(n8462), .ZN(n8468) );
  NOR2_X2 U5780 ( .A1(n8474), .A2(n8473), .ZN(n8478) );
  NOR2_X2 U5781 ( .A1(n8488), .A2(n8487), .ZN(n8492) );
  NOR2_X2 U5782 ( .A1(n8522), .A2(n8521), .ZN(n8526) );
  NAND3_X2 U5783 ( .A1(n8705), .A2(n8704), .A3(n8703), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  NAND3_X1 U5784 ( .A1(n10649), .A2(n8702), .A3(n8701), .ZN(n8704) );
  OAI21_X2 U5785 ( .B1(n6223), .B2(n6138), .A(n8753), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5786 ( .B1(n6223), .B2(n10534), .A(n8754), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5787 ( .B1(n6221), .B2(n10532), .A(n8793), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5788 ( .B1(n6221), .B2(n6142), .A(n8794), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5789 ( .B1(n6221), .B2(net70509), .A(n8795), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5790 ( .B1(n6213), .B2(n6023), .A(n8878), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5791 ( .B1(n6138), .B2(n6023), .A(n8879), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5792 ( .B1(n6142), .B2(n6023), .A(n8880), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5793 ( .B1(net76480), .B2(n6023), .A(n8881), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5794 ( .B1(n6213), .B2(n6025), .A(n8913), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5795 ( .B1(n6138), .B2(n6025), .A(n8914), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5796 ( .B1(n6142), .B2(n6025), .A(n8915), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5797 ( .B1(net76480), .B2(n6025), .A(n8916), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  NAND3_X2 U5798 ( .A1(n8973), .A2(n8972), .A3(n8971), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5799 ( .B1(n6213), .B2(n6032), .A(n9046), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5800 ( .B1(n6138), .B2(n6032), .A(n9047), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5801 ( .B1(n6142), .B2(n6032), .A(n9048), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5802 ( .B1(net76480), .B2(n6032), .A(n9049), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  NOR2_X1 U5803 ( .A1(n4968), .A2(n9271), .ZN(n9276) );
  NAND3_X2 U5804 ( .A1(n9288), .A2(n9287), .A3(n9286), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  NAND3_X2 U5805 ( .A1(n9541), .A2(n9540), .A3(n9539), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5806 ( .B1(n6056), .B2(n6138), .A(n9678), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5807 ( .B1(n6142), .B2(n4802), .A(n9679), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5808 ( .B1(net76480), .B2(n6057), .A(n9680), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5809 ( .B1(n6222), .B2(n10532), .A(n9829), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5810 ( .B1(n6222), .B2(n10534), .A(n9830), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5811 ( .B1(n6222), .B2(net70509), .A(n9831), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5812 ( .B1(n6214), .B2(n6068), .A(n9969), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5813 ( .B1(n10532), .B2(n4803), .A(n9970), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5814 ( .B1(n10534), .B2(n4803), .A(n9971), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5815 ( .B1(net70509), .B2(n6068), .A(n9972), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5816 ( .B1(n6214), .B2(n6070), .A(n10008), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5817 ( .B1(n10532), .B2(n6070), .A(n10009), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5818 ( .B1(n10534), .B2(n6070), .A(n10010), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5819 ( .B1(net70509), .B2(n6070), .A(n10011), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5820 ( .B1(n6214), .B2(n6085), .A(n10271), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5821 ( .B1(n10532), .B2(n6085), .A(n10272), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5822 ( .B1(n10534), .B2(n6085), .A(n10273), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5823 ( .B1(net70509), .B2(n6085), .A(n10274), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5824 ( .B1(n6214), .B2(n6087), .A(n10299), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5825 ( .B1(n10532), .B2(n6087), .A(n10300), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5826 ( .B1(n10534), .B2(n6087), .A(n10301), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5827 ( .B1(net70509), .B2(n6087), .A(n10302), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5828 ( .B1(n6214), .B2(n6191), .A(n10530), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5829 ( .B1(n6191), .B2(n6138), .A(n10531), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U5830 ( .B1(n6191), .B2(n6142), .A(n10533), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  NOR2_X2 U5831 ( .A1(net76278), .A2(net76658), .ZN(n10546) );
  NOR2_X2 U5832 ( .A1(net76278), .A2(n6155), .ZN(n10549) );
  NOR2_X2 U5833 ( .A1(n6194), .A2(net76274), .ZN(n10552) );
  NOR2_X2 U5834 ( .A1(n6198), .A2(net76274), .ZN(n10555) );
  NAND3_X2 U5835 ( .A1(n6096), .A2(reset), .A3(net76510), .ZN(n10559) );
  NAND3_X2 U5836 ( .A1(n6101), .A2(reset), .A3(net76510), .ZN(n10561) );
  NAND3_X2 U5837 ( .A1(n6107), .A2(reset), .A3(net76510), .ZN(n10563) );
  NOR2_X2 U5838 ( .A1(net76278), .A2(n6157), .ZN(n10564) );
  NOR2_X2 U5839 ( .A1(net76278), .A2(n6159), .ZN(n10567) );
  NOR2_X2 U5840 ( .A1(net76278), .A2(n6161), .ZN(n10570) );
  NOR2_X2 U5841 ( .A1(n6203), .A2(net76274), .ZN(n10573) );
  NOR2_X2 U5842 ( .A1(net76278), .A2(net76614), .ZN(n10576) );
  NOR2_X2 U5843 ( .A1(n6207), .A2(net76274), .ZN(n10579) );
  NOR2_X2 U5844 ( .A1(net76278), .A2(n6163), .ZN(n10582) );
  NOR2_X2 U5845 ( .A1(net76278), .A2(n6165), .ZN(n10585) );
  NOR2_X2 U5846 ( .A1(net76278), .A2(n6167), .ZN(n10588) );
  NOR2_X2 U5847 ( .A1(net76278), .A2(n6169), .ZN(n10591) );
  NOR2_X2 U5848 ( .A1(net76278), .A2(n6171), .ZN(n10594) );
  NOR2_X2 U5849 ( .A1(net76278), .A2(n6173), .ZN(n10597) );
  NOR2_X2 U5850 ( .A1(n6211), .A2(net76274), .ZN(n10600) );
  NOR2_X2 U5851 ( .A1(n6214), .A2(net76274), .ZN(n10603) );
  NAND3_X2 U5852 ( .A1(n10607), .A2(reset), .A3(net76510), .ZN(n10610) );
  NOR2_X2 U5853 ( .A1(net76278), .A2(net76548), .ZN(n10611) );
  NAND3_X2 U5854 ( .A1(n10614), .A2(reset), .A3(net76510), .ZN(n10617) );
  NAND3_X2 U5855 ( .A1(net70574), .A2(reset), .A3(net76510), .ZN(n10619) );
  NOR2_X2 U5856 ( .A1(net76318), .A2(net76274), .ZN(n10620) );
  NOR2_X2 U5857 ( .A1(n6219), .A2(net76274), .ZN(n10623) );
  NOR2_X2 U5858 ( .A1(net76278), .A2(n6182), .ZN(n10626) );
  NAND3_X2 U5859 ( .A1(n6148), .A2(reset), .A3(net76510), .ZN(n10630) );
  NOR2_X2 U5860 ( .A1(net76278), .A2(n6184), .ZN(n10631) );
  NOR2_X2 U5861 ( .A1(net76278), .A2(n6186), .ZN(n10634) );
  NOR2_X2 U5862 ( .A1(net76278), .A2(n6188), .ZN(n10637) );
  OAI21_X2 U5863 ( .B1(n6191), .B2(net76480), .A(n10656), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  AND2_X4 U5864 ( .A1(reset), .A2(net76660), .ZN(n4867) );
  AND2_X4 U5865 ( .A1(net76270), .A2(n6208), .ZN(n4868) );
  AND2_X4 U5866 ( .A1(net76270), .A2(n6195), .ZN(n4869) );
  AND2_X4 U5867 ( .A1(net76270), .A2(n6220), .ZN(n4870) );
  AND2_X4 U5868 ( .A1(net76270), .A2(net76320), .ZN(n4871) );
  AND2_X4 U5869 ( .A1(net76270), .A2(n6212), .ZN(n4872) );
  AND2_X4 U5870 ( .A1(net76270), .A2(n6199), .ZN(n4873) );
  AND2_X4 U5871 ( .A1(n8669), .A2(n8672), .ZN(n4874) );
  INV_X4 U5872 ( .A(n10604), .ZN(n6176) );
  INV_X16 U5873 ( .A(n9765), .ZN(n6061) );
  INV_X4 U5874 ( .A(n10012), .ZN(n6071) );
  INV_X16 U5875 ( .A(n6071), .ZN(n6070) );
  AND2_X4 U5876 ( .A1(net76270), .A2(n6170), .ZN(n4875) );
  AND2_X4 U5877 ( .A1(net76270), .A2(n6204), .ZN(n4876) );
  AND2_X4 U5878 ( .A1(net76270), .A2(net76616), .ZN(n4877) );
  AND2_X4 U5879 ( .A1(net76270), .A2(n6172), .ZN(n4878) );
  AND2_X4 U5880 ( .A1(net76270), .A2(net76550), .ZN(n4879) );
  AND2_X4 U5881 ( .A1(n6005), .A2(net78051), .ZN(n4880) );
  INV_X4 U5882 ( .A(n6101), .ZN(n6102) );
  INV_X4 U5883 ( .A(n6148), .ZN(n6147) );
  AND2_X4 U5884 ( .A1(net75791), .A2(net73697), .ZN(n4881) );
  INV_X8 U5885 ( .A(n5642), .ZN(n5644) );
  INV_X8 U5886 ( .A(n8402), .ZN(n6020) );
  INV_X4 U5887 ( .A(n10276), .ZN(n6086) );
  INV_X16 U5888 ( .A(n6086), .ZN(n6085) );
  INV_X4 U5889 ( .A(net76274), .ZN(net76270) );
  AND2_X4 U5890 ( .A1(net76270), .A2(n6164), .ZN(n4882) );
  AND2_X4 U5891 ( .A1(net76270), .A2(n6168), .ZN(n4883) );
  AND2_X4 U5892 ( .A1(net76270), .A2(n6162), .ZN(n4884) );
  AND2_X4 U5893 ( .A1(net76270), .A2(n6183), .ZN(n4885) );
  AND2_X4 U5894 ( .A1(net76270), .A2(n6185), .ZN(n4886) );
  AND2_X4 U5895 ( .A1(net76270), .A2(n6189), .ZN(n4887) );
  AND2_X4 U5896 ( .A1(net76270), .A2(n6166), .ZN(n4888) );
  AND2_X4 U5897 ( .A1(net76270), .A2(n10535), .ZN(n4889) );
  AND2_X4 U5898 ( .A1(net76270), .A2(n6187), .ZN(n4890) );
  AND2_X4 U5899 ( .A1(net76270), .A2(n6158), .ZN(n4891) );
  AND2_X4 U5900 ( .A1(net76270), .A2(n6160), .ZN(n4892) );
  AND2_X4 U5901 ( .A1(net76270), .A2(n6174), .ZN(n4893) );
  NAND4_X2 U5902 ( .A1(n6941), .A2(n6938), .A3(n6940), .A4(n6939), .ZN(
        net73837) );
  INV_X4 U5903 ( .A(net76650), .ZN(net76646) );
  INV_X4 U5904 ( .A(net73877), .ZN(net73997) );
  AND3_X4 U5905 ( .A1(n4900), .A2(net73429), .A3(net73443), .ZN(n4894) );
  NOR2_X2 U5906 ( .A1(n8677), .A2(net73434), .ZN(net70574) );
  NOR2_X2 U5907 ( .A1(n8677), .A2(net73439), .ZN(n10607) );
  NOR2_X2 U5908 ( .A1(n8677), .A2(net73436), .ZN(n10614) );
  AND3_X4 U5909 ( .A1(net73427), .A2(n4900), .A3(net73429), .ZN(n4895) );
  INV_X4 U5910 ( .A(n4872), .ZN(n6210) );
  INV_X4 U5911 ( .A(n4869), .ZN(n6193) );
  INV_X4 U5912 ( .A(n4868), .ZN(n6206) );
  INV_X4 U5913 ( .A(n4871), .ZN(n6216) );
  INV_X4 U5914 ( .A(n4870), .ZN(n6218) );
  INV_X4 U5915 ( .A(n4880), .ZN(n6084) );
  INV_X4 U5916 ( .A(n6084), .ZN(n6083) );
  AND2_X4 U5917 ( .A1(n8766), .A2(n8765), .ZN(n4896) );
  INV_X4 U5918 ( .A(n10544), .ZN(n6081) );
  INV_X4 U5920 ( .A(n8882), .ZN(n6024) );
  INV_X16 U5921 ( .A(n6024), .ZN(n6023) );
  INV_X4 U5922 ( .A(n9268), .ZN(n6037) );
  INV_X8 U5923 ( .A(n6037), .ZN(n6036) );
  INV_X8 U5924 ( .A(n6037), .ZN(n6035) );
  INV_X16 U5925 ( .A(n4816), .ZN(n6034) );
  INV_X16 U5926 ( .A(n4816), .ZN(n6033) );
  INV_X16 U5927 ( .A(n9426), .ZN(n6047) );
  INV_X16 U5928 ( .A(n9426), .ZN(n6046) );
  INV_X16 U5929 ( .A(n9868), .ZN(n6066) );
  INV_X16 U5930 ( .A(n9868), .ZN(n6065) );
  NAND2_X1 U5931 ( .A1(n4966), .A2(net73495), .ZN(net70738) );
  INV_X4 U5932 ( .A(net70738), .ZN(net77030) );
  INV_X4 U5933 ( .A(net80189), .ZN(net73608) );
  AND2_X4 U5934 ( .A1(net73494), .A2(net70507), .ZN(n4899) );
  AND2_X4 U5935 ( .A1(n5589), .A2(n5066), .ZN(n4900) );
  INV_X4 U5936 ( .A(net70718), .ZN(net105360) );
  AND2_X4 U5937 ( .A1(n5010), .A2(n4874), .ZN(n4903) );
  AND2_X4 U5938 ( .A1(n5010), .A2(net73416), .ZN(n4904) );
  AND2_X4 U5939 ( .A1(n5010), .A2(net73423), .ZN(n4905) );
  AND2_X4 U5940 ( .A1(n5010), .A2(net73421), .ZN(n4906) );
  NAND2_X2 U5941 ( .A1(n8464), .A2(n8463), .ZN(n9533) );
  INV_X4 U5942 ( .A(n9533), .ZN(n10649) );
  AND2_X4 U5943 ( .A1(n5066), .A2(net73468), .ZN(n4907) );
  AND2_X2 U5944 ( .A1(net70821), .A2(n8580), .ZN(n4910) );
  NAND2_X1 U5945 ( .A1(net78051), .A2(n10099), .ZN(n10094) );
  AND2_X4 U5946 ( .A1(dmem_dsize[1]), .A2(n4899), .ZN(n4911) );
  AND2_X2 U5947 ( .A1(n8728), .A2(n6041), .ZN(n4912) );
  AND2_X4 U5948 ( .A1(n5068), .A2(net73443), .ZN(n4913) );
  AND2_X4 U5949 ( .A1(n5067), .A2(net73443), .ZN(n4914) );
  NAND2_X2 U5950 ( .A1(net73500), .A2(net70738), .ZN(n4915) );
  INV_X4 U5951 ( .A(n8917), .ZN(n6026) );
  INV_X16 U5952 ( .A(n6026), .ZN(n6025) );
  AND2_X4 U5953 ( .A1(net73427), .A2(n5068), .ZN(n4916) );
  INV_X4 U5954 ( .A(reset), .ZN(net76274) );
  AND2_X4 U5955 ( .A1(n5067), .A2(net73427), .ZN(n4920) );
  AND2_X4 U5956 ( .A1(n8301), .A2(net73877), .ZN(n4921) );
  NAND2_X2 U5957 ( .A1(n4910), .A2(net73585), .ZN(net70691) );
  AND2_X4 U5958 ( .A1(n8768), .A2(n8767), .ZN(n4922) );
  NOR2_X2 U5959 ( .A1(net70574), .A2(net76274), .ZN(n5688) );
  NOR2_X2 U5960 ( .A1(n10607), .A2(net76274), .ZN(n10608) );
  NAND3_X2 U5961 ( .A1(reset), .A2(instruction[1]), .A3(n5591), .ZN(n4962) );
  INV_X4 U5962 ( .A(n10517), .ZN(n6100) );
  INV_X2 U5963 ( .A(net77276), .ZN(net123282) );
  INV_X16 U5964 ( .A(net77784), .ZN(net77780) );
  INV_X16 U5965 ( .A(net77832), .ZN(net77828) );
  INV_X16 U5966 ( .A(net75468), .ZN(net77776) );
  INV_X8 U5967 ( .A(n8411), .ZN(n6013) );
  INV_X16 U5968 ( .A(n6013), .ZN(n6012) );
  INV_X8 U5969 ( .A(net73838), .ZN(net77296) );
  INV_X16 U5970 ( .A(net77296), .ZN(net77292) );
  INV_X16 U5971 ( .A(net75443), .ZN(net77656) );
  AND2_X4 U5972 ( .A1(net76270), .A2(n9045), .ZN(n4964) );
  AND2_X4 U5973 ( .A1(reset), .A2(n10297), .ZN(n4965) );
  AND3_X4 U5974 ( .A1(instruction[4]), .A2(net74029), .A3(net73499), .ZN(n4966) );
  AND3_X4 U5975 ( .A1(net73684), .A2(instruction[29]), .A3(net73619), .ZN(
        n4967) );
  XOR2_X2 U5976 ( .A(instruction[19]), .B(n10003), .Z(n4968) );
  AND4_X2 U5977 ( .A1(n5593), .A2(net71266), .A3(n5594), .A4(n5595), .ZN(n4970) );
  OR2_X2 U5978 ( .A1(instruction[28]), .A2(instruction[29]), .ZN(n4971) );
  INV_X8 U5979 ( .A(n5628), .ZN(net77042) );
  INV_X4 U5980 ( .A(n5797), .ZN(n5955) );
  INV_X4 U5981 ( .A(net77504), .ZN(net77484) );
  INV_X8 U5982 ( .A(net77504), .ZN(net77482) );
  AND2_X4 U5983 ( .A1(net73423), .A2(n4913), .ZN(n4990) );
  AND2_X4 U5984 ( .A1(n4874), .A2(n4913), .ZN(n4991) );
  AND2_X4 U5985 ( .A1(n4916), .A2(n4874), .ZN(n4992) );
  AND2_X4 U5986 ( .A1(n4894), .A2(n4874), .ZN(n4993) );
  AND2_X4 U5987 ( .A1(n4920), .A2(n4874), .ZN(n4994) );
  AND2_X4 U5988 ( .A1(n4914), .A2(n4874), .ZN(n4995) );
  AND2_X4 U5989 ( .A1(n4895), .A2(n4874), .ZN(n4996) );
  AND2_X4 U5990 ( .A1(n4916), .A2(net73416), .ZN(n4997) );
  AND2_X4 U5991 ( .A1(n4913), .A2(net73421), .ZN(n4998) );
  AND2_X4 U5992 ( .A1(n4920), .A2(net73416), .ZN(n4999) );
  AND2_X4 U5993 ( .A1(n4920), .A2(net73423), .ZN(n5000) );
  AND2_X4 U5994 ( .A1(n4920), .A2(net73421), .ZN(n5001) );
  AND2_X4 U5995 ( .A1(n4914), .A2(net73416), .ZN(n5002) );
  AND2_X4 U5996 ( .A1(n4914), .A2(net73423), .ZN(n5003) );
  AND2_X4 U5997 ( .A1(n4914), .A2(net73421), .ZN(n5004) );
  AND2_X4 U5998 ( .A1(n4916), .A2(net73423), .ZN(n5005) );
  AND2_X4 U5999 ( .A1(n4895), .A2(net73416), .ZN(n5006) );
  AND2_X4 U6000 ( .A1(n4895), .A2(net73421), .ZN(n5007) );
  AND2_X4 U6001 ( .A1(n4913), .A2(net73416), .ZN(n5008) );
  AND2_X4 U6002 ( .A1(n4916), .A2(net73421), .ZN(n5009) );
  INV_X4 U6003 ( .A(n5577), .ZN(n5944) );
  AND3_X4 U6004 ( .A1(net73427), .A2(n4907), .A3(net73429), .ZN(n5010) );
  NAND3_X2 U6005 ( .A1(n8539), .A2(instruction[1]), .A3(net73170), .ZN(n8565)
         );
  AND2_X4 U6006 ( .A1(net76270), .A2(n8742), .ZN(n5011) );
  AND2_X4 U6007 ( .A1(net76270), .A2(n8792), .ZN(n5012) );
  AND2_X4 U6008 ( .A1(net76270), .A2(n9826), .ZN(n5013) );
  INV_X4 U6009 ( .A(n10400), .ZN(n10909) );
  AND2_X2 U6010 ( .A1(n4880), .A2(net70696), .ZN(n5015) );
  INV_X4 U6011 ( .A(net85047), .ZN(net84663) );
  AND2_X2 U6012 ( .A1(net70701), .A2(n10416), .ZN(n5039) );
  AND2_X2 U6013 ( .A1(net70701), .A2(n10415), .ZN(n5040) );
  AND2_X2 U6014 ( .A1(net70701), .A2(n10414), .ZN(n5041) );
  OR2_X4 U6015 ( .A1(n10093), .A2(net70710), .ZN(n5042) );
  NAND2_X2 U6016 ( .A1(n8464), .A2(n8463), .ZN(n6008) );
  AND2_X2 U6017 ( .A1(net70701), .A2(n10373), .ZN(n5049) );
  AND2_X2 U6018 ( .A1(net70701), .A2(n9402), .ZN(n5050) );
  AND2_X2 U6019 ( .A1(net70701), .A2(n10387), .ZN(n5051) );
  AND2_X2 U6020 ( .A1(net70701), .A2(n10394), .ZN(n5052) );
  AND2_X2 U6021 ( .A1(net70701), .A2(n10307), .ZN(n5053) );
  AND2_X2 U6022 ( .A1(net70701), .A2(n9836), .ZN(n5054) );
  AND2_X2 U6023 ( .A1(net70701), .A2(n10402), .ZN(n5055) );
  AND2_X2 U6024 ( .A1(net70701), .A2(n10380), .ZN(n5056) );
  AND2_X2 U6025 ( .A1(net70701), .A2(n10366), .ZN(n5057) );
  AND2_X2 U6026 ( .A1(net70701), .A2(n10281), .ZN(n5058) );
  AND3_X4 U6027 ( .A1(n8981), .A2(n8980), .A3(n8979), .ZN(n5061) );
  AND3_X4 U6028 ( .A1(n10542), .A2(net80189), .A3(net71094), .ZN(n5062) );
  AND2_X4 U6029 ( .A1(net70706), .A2(net73541), .ZN(n5065) );
  AND3_X4 U6030 ( .A1(n5590), .A2(net70506), .A3(net73519), .ZN(n5066) );
  AND2_X4 U6031 ( .A1(net73465), .A2(n4907), .ZN(n5067) );
  AND2_X4 U6032 ( .A1(net73465), .A2(n4900), .ZN(n5068) );
  AND2_X2 U6033 ( .A1(n8553), .A2(n8536), .ZN(n5252) );
  INV_X4 U6034 ( .A(n8527), .ZN(n6190) );
  INV_X4 U6035 ( .A(n4911), .ZN(net77999) );
  INV_X4 U6036 ( .A(n10608), .ZN(n6179) );
  INV_X4 U6037 ( .A(n6179), .ZN(n6178) );
  INV_X4 U6038 ( .A(n10615), .ZN(n6181) );
  NOR2_X2 U6039 ( .A1(n10614), .A2(net76274), .ZN(n10615) );
  INV_X4 U6040 ( .A(n6181), .ZN(n6180) );
  INV_X4 U6041 ( .A(n5688), .ZN(n5695) );
  INV_X4 U6042 ( .A(n5695), .ZN(net76488) );
  OR2_X4 U6043 ( .A1(n10152), .A2(net70710), .ZN(n5570) );
  INV_X1 U6044 ( .A(net148116), .ZN(dmem_write_out[17]) );
  INV_X4 U6045 ( .A(n9330), .ZN(n6042) );
  INV_X8 U6046 ( .A(n6042), .ZN(n6040) );
  INV_X8 U6047 ( .A(n6042), .ZN(n6041) );
  AND2_X2 U6048 ( .A1(n10108), .A2(net73585), .ZN(n5571) );
  INV_X1 U6049 ( .A(n5867), .ZN(n5868) );
  INV_X4 U6050 ( .A(net70507), .ZN(dmem_dsize[0]) );
  NAND3_X1 U6051 ( .A1(net73495), .A2(net73496), .A3(n8659), .ZN(net70507) );
  INV_X4 U6052 ( .A(dmem_dsize[0]), .ZN(net76464) );
  INV_X4 U6053 ( .A(net70718), .ZN(net77086) );
  OR2_X4 U6054 ( .A1(net76464), .A2(n10540), .ZN(n5572) );
  INV_X4 U6055 ( .A(n10535), .ZN(n6148) );
  INV_X4 U6056 ( .A(n10519), .ZN(n6101) );
  OR2_X4 U6057 ( .A1(net76464), .A2(n10078), .ZN(n5573) );
  INV_X8 U6058 ( .A(net78050), .ZN(net78051) );
  INV_X1 U6059 ( .A(net78051), .ZN(net72962) );
  INV_X4 U6060 ( .A(n6176), .ZN(n6175) );
  INV_X4 U6061 ( .A(n6176), .ZN(n6177) );
  INV_X4 U6062 ( .A(n10607), .ZN(n6138) );
  INV_X4 U6063 ( .A(n10614), .ZN(n6142) );
  INV_X4 U6064 ( .A(net70574), .ZN(net76480) );
  INV_X4 U6065 ( .A(n10516), .ZN(n6096) );
  INV_X4 U6066 ( .A(n6096), .ZN(n6095) );
  INV_X4 U6067 ( .A(n10521), .ZN(n6107) );
  INV_X4 U6068 ( .A(n6107), .ZN(n6106) );
  INV_X4 U6069 ( .A(n4869), .ZN(n6192) );
  INV_X4 U6070 ( .A(n4873), .ZN(n6196) );
  INV_X4 U6071 ( .A(n4873), .ZN(n6197) );
  INV_X4 U6072 ( .A(n4868), .ZN(n6205) );
  INV_X4 U6073 ( .A(n4872), .ZN(n6209) );
  INV_X4 U6074 ( .A(n4871), .ZN(n6215) );
  INV_X4 U6075 ( .A(n4870), .ZN(n6217) );
  INV_X4 U6076 ( .A(n10512), .ZN(n6093) );
  INV_X4 U6077 ( .A(n4805), .ZN(n6103) );
  INV_X4 U6078 ( .A(n4805), .ZN(n6104) );
  INV_X4 U6079 ( .A(n4891), .ZN(n6111) );
  INV_X4 U6080 ( .A(n4892), .ZN(n6114) );
  INV_X4 U6081 ( .A(n4884), .ZN(n6117) );
  INV_X4 U6082 ( .A(n4882), .ZN(n6120) );
  INV_X4 U6083 ( .A(n4888), .ZN(n6123) );
  INV_X4 U6084 ( .A(n4883), .ZN(n6126) );
  INV_X4 U6085 ( .A(n4893), .ZN(n6135) );
  INV_X4 U6086 ( .A(n4885), .ZN(n6143) );
  INV_X4 U6087 ( .A(n4889), .ZN(net76716) );
  INV_X4 U6088 ( .A(n4886), .ZN(net76702) );
  INV_X4 U6089 ( .A(n4890), .ZN(n6149) );
  INV_X4 U6090 ( .A(n4887), .ZN(n6152) );
  INV_X4 U6091 ( .A(n4806), .ZN(n6213) );
  INV_X4 U6092 ( .A(n4915), .ZN(net76650) );
  INV_X4 U6093 ( .A(reset), .ZN(net76278) );
  INV_X16 U6094 ( .A(n10149), .ZN(n6080) );
  NAND2_X4 U6095 ( .A1(n10142), .A2(reset), .ZN(n10149) );
  OAI21_X2 U6096 ( .B1(n6078), .B2(net70509), .A(n10148), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6097 ( .B1(n6078), .B2(n6142), .A(n10147), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6098 ( .B1(n6078), .B2(n6214), .A(n10145), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6099 ( .B1(n6078), .B2(n6138), .A(n10146), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6100 ( .B1(net76480), .B2(n6043), .A(n9382), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6101 ( .B1(n6138), .B2(n6043), .A(n9380), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6102 ( .B1(n6213), .B2(n6043), .A(n9379), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6103 ( .B1(n6142), .B2(n6043), .A(n9381), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X16 U6104 ( .A(n6080), .ZN(n6079) );
  INV_X16 U6105 ( .A(n6080), .ZN(n6078) );
  INV_X16 U6106 ( .A(n6045), .ZN(n6043) );
  NAND2_X4 U6107 ( .A1(n9378), .A2(net76270), .ZN(n9383) );
  INV_X16 U6108 ( .A(n6045), .ZN(n6044) );
  MUX2_X2 U6109 ( .A(multOut[10]), .B(n10130), .S(net73585), .Z(n10136) );
  INV_X16 U6110 ( .A(n9383), .ZN(n6045) );
  OAI21_X2 U6112 ( .B1(net76480), .B2(n4801), .A(n9526), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6113 ( .B1(n6142), .B2(n4801), .A(n9525), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6114 ( .B1(n6138), .B2(n6048), .A(n9523), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6115 ( .B1(n6213), .B2(n6048), .A(n9522), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6116 ( .A1(n5127), .A2(n6088), .B1(net76660), .B2(n6048), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  NAND2_X4 U6119 ( .A1(net76270), .A2(n9520), .ZN(n9528) );
  INV_X16 U6120 ( .A(n9704), .ZN(n9765) );
  NAND2_X4 U6121 ( .A1(net76270), .A2(n9703), .ZN(n9704) );
  OAI21_X2 U6122 ( .B1(n6213), .B2(n6056), .A(n9677), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  INV_X16 U6123 ( .A(n6058), .ZN(n6056) );
  NAND2_X4 U6124 ( .A1(n9674), .A2(net76270), .ZN(n9681) );
  INV_X16 U6125 ( .A(n6058), .ZN(n6057) );
  INV_X16 U6126 ( .A(n9681), .ZN(n6058) );
  OAI21_X2 U6127 ( .B1(n6053), .B2(net76480), .A(n9645), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6128 ( .B1(n6053), .B2(n6138), .A(n9643), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6129 ( .B1(n6053), .B2(n6213), .A(n9642), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6130 ( .B1(n6053), .B2(n6142), .A(n9644), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  INV_X16 U6131 ( .A(n6055), .ZN(n6054) );
  INV_X16 U6132 ( .A(n6055), .ZN(n6053) );
  NAND2_X1 U6133 ( .A1(n6178), .A2(REGFILE_reg_out_29__3_), .ZN(n10049) );
  INV_X16 U6134 ( .A(n9646), .ZN(n6055) );
  OAI21_X2 U6135 ( .B1(net76506), .B2(n10563), .A(n10562), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6136 ( .B1(net76506), .B2(n10596), .A(n10595), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6137 ( .B1(net76506), .B2(n10587), .A(n10586), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6138 ( .B1(net76506), .B2(n10584), .A(n10583), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6139 ( .B1(net76506), .B2(n10561), .A(n10560), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6140 ( .B1(net76506), .B2(n10559), .A(n10558), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6141 ( .B1(net76502), .B2(n10636), .A(n10635), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6142 ( .B1(net76502), .B2(n10630), .A(n10629), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6143 ( .B1(net76502), .B2(n10633), .A(n10632), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6144 ( .B1(net76502), .B2(n10639), .A(n10638), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6145 ( .B1(net76502), .B2(n10610), .A(n10609), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6146 ( .B1(net76506), .B2(n10617), .A(n10616), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6147 ( .B1(net76502), .B2(n10590), .A(n10589), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6148 ( .B1(net76506), .B2(n10578), .A(n10577), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6149 ( .B1(net76506), .B2(n10575), .A(n10574), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6150 ( .B1(net76502), .B2(n10628), .A(n10627), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  INV_X2 U6151 ( .A(n9519), .ZN(dmem_addr_out[8]) );
  OAI21_X2 U6152 ( .B1(net76506), .B2(n10572), .A(n10571), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6153 ( .B1(net76506), .B2(n10625), .A(n10624), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6154 ( .B1(net76506), .B2(n10566), .A(n10565), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6155 ( .B1(net76506), .B2(n10622), .A(n10621), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6156 ( .B1(net76506), .B2(n10557), .A(n10556), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6157 ( .B1(net76502), .B2(n10613), .A(n10612), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6158 ( .B1(net76506), .B2(n10554), .A(n10553), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6159 ( .B1(net76506), .B2(n10606), .A(n10605), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6160 ( .B1(net76506), .B2(n10602), .A(n10601), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6161 ( .B1(net76506), .B2(n10599), .A(n10598), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI21_X2 U6162 ( .B1(net76506), .B2(n10551), .A(n10550), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  NAND2_X1 U6163 ( .A1(n4892), .A2(REGFILE_reg_out_17__0_), .ZN(n10568) );
  OAI21_X2 U6164 ( .B1(net76502), .B2(n10569), .A(n10568), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  NAND2_X1 U6165 ( .A1(n4867), .A2(REGFILE_reg_out_0__0_), .ZN(n10547) );
  OAI21_X2 U6166 ( .B1(net76502), .B2(n10548), .A(n10547), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  NAND2_X1 U6167 ( .A1(REGFILE_reg_out_3__20_), .A2(net77422), .ZN(n7392) );
  INV_X8 U6168 ( .A(net77632), .ZN(net77630) );
  AOI22_X2 U6169 ( .A1(REGFILE_reg_out_26__19_), .A2(net75439), .B1(
        REGFILE_reg_out_27__19_), .B2(net89184), .ZN(n6521) );
  INV_X8 U6170 ( .A(net75441), .ZN(net84760) );
  OAI21_X2 U6171 ( .B1(n6214), .B2(net77116), .A(n10118), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  NAND2_X1 U6172 ( .A1(n5009), .A2(n10947), .ZN(n10217) );
  INV_X16 U6173 ( .A(n5582), .ZN(net77106) );
  NAND2_X4 U6174 ( .A1(instruction[11]), .A2(instruction[12]), .ZN(net80161)
         );
  AOI21_X4 U6175 ( .B1(net81874), .B2(n4970), .A(net76274), .ZN(n5582) );
  AOI22_X1 U6176 ( .A1(REGFILE_reg_out_16__6_), .A2(net77762), .B1(
        REGFILE_reg_out_15__6_), .B2(net75468), .ZN(n6770) );
  AOI22_X2 U6177 ( .A1(REGFILE_reg_out_16__10_), .A2(net75467), .B1(n5615), 
        .B2(net75468), .ZN(n6694) );
  AOI22_X2 U6178 ( .A1(n4846), .A2(net75467), .B1(net83261), .B2(net75468), 
        .ZN(n5606) );
  NAND2_X1 U6179 ( .A1(net92782), .A2(net81874), .ZN(dmem_addr_out[1]) );
  INV_X4 U6180 ( .A(net77300), .ZN(net93763) );
  NAND2_X1 U6181 ( .A1(REGFILE_reg_out_2__10_), .A2(net77342), .ZN(n7828) );
  BUF_X8 U6182 ( .A(n5943), .Z(n5577) );
  INV_X8 U6183 ( .A(net76194), .ZN(net124970) );
  AOI22_X4 U6184 ( .A1(REGFILE_reg_out_23__15_), .A2(net77828), .B1(
        REGFILE_reg_out_22__15_), .B2(net77836), .ZN(n6586) );
  INV_X4 U6185 ( .A(net77406), .ZN(n5648) );
  NAND3_X2 U6186 ( .A1(instruction[8]), .A2(net73989), .A3(instruction[10]), 
        .ZN(n5578) );
  INV_X8 U6187 ( .A(net77776), .ZN(net77774) );
  INV_X8 U6188 ( .A(net72414), .ZN(net36470) );
  AOI22_X4 U6189 ( .A1(REGFILE_reg_out_29__10_), .A2(net77650), .B1(
        REGFILE_reg_out_28__10_), .B2(n5751), .ZN(n6705) );
  AOI22_X2 U6190 ( .A1(REGFILE_reg_out_30__5_), .A2(net77634), .B1(
        REGFILE_reg_out_2__5_), .B2(net75442), .ZN(n6802) );
  AOI22_X1 U6191 ( .A1(REGFILE_reg_out_16__30_), .A2(net77764), .B1(
        REGFILE_reg_out_15__30_), .B2(n5579), .ZN(n6257) );
  AOI22_X2 U6192 ( .A1(REGFILE_reg_out_26__29_), .A2(net77620), .B1(
        REGFILE_reg_out_27__29_), .B2(net77630), .ZN(n6288) );
  AOI22_X2 U6193 ( .A1(REGFILE_reg_out_17__15_), .A2(net77796), .B1(
        REGFILE_reg_out_18__15_), .B2(n5890), .ZN(n6584) );
  AOI22_X2 U6194 ( .A1(REGFILE_reg_out_17__18_), .A2(net77796), .B1(
        REGFILE_reg_out_18__18_), .B2(n6896), .ZN(n6530) );
  INV_X4 U6195 ( .A(n10943), .ZN(net75842) );
  AOI22_X4 U6196 ( .A1(REGFILE_reg_out_7__13_), .A2(net77714), .B1(
        REGFILE_reg_out_6__13_), .B2(net75456), .ZN(n6637) );
  AOI22_X4 U6197 ( .A1(REGFILE_reg_out_17__10_), .A2(net77794), .B1(
        REGFILE_reg_out_18__10_), .B2(n6896), .ZN(n6688) );
  AOI22_X2 U6198 ( .A1(REGFILE_reg_out_19__29_), .A2(net77814), .B1(
        REGFILE_reg_out_1__29_), .B2(net82631), .ZN(n6274) );
  NOR2_X2 U6199 ( .A1(n4806), .A2(net76274), .ZN(n10604) );
  INV_X16 U6200 ( .A(n5624), .ZN(net82631) );
  AOI22_X4 U6201 ( .A1(REGFILE_reg_out_7__14_), .A2(net77714), .B1(
        REGFILE_reg_out_6__14_), .B2(net75456), .ZN(n6621) );
  AOI22_X4 U6202 ( .A1(REGFILE_reg_out_31__14_), .A2(net77668), .B1(
        REGFILE_reg_out_3__14_), .B2(net77676), .ZN(n6618) );
  AOI22_X4 U6203 ( .A1(REGFILE_reg_out_4__12_), .A2(n5678), .B1(
        REGFILE_reg_out_5__12_), .B2(net75452), .ZN(n6655) );
  NAND2_X4 U6204 ( .A1(n5631), .A2(net77400), .ZN(net78105) );
  BUF_X32 U6205 ( .A(aluA[31]), .Z(net80189) );
  NAND2_X2 U6206 ( .A1(net71227), .A2(net71228), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U6207 ( .A1(n4877), .A2(REGFILE_reg_out_1__1_), .ZN(net71228) );
  NAND2_X1 U6208 ( .A1(net77420), .A2(REGFILE_reg_out_27__18_), .ZN(n7450) );
  INV_X32 U6209 ( .A(instruction[15]), .ZN(net82738) );
  INV_X8 U6210 ( .A(net77508), .ZN(net77502) );
  INV_X4 U6211 ( .A(net77508), .ZN(net77504) );
  OAI211_X1 U6212 ( .C1(n4865), .C2(net73170), .A(net73496), .B(n8658), .ZN(
        n8870) );
  NAND4_X1 U6213 ( .A1(n4865), .A2(net73503), .A3(n6607), .A4(net73496), .ZN(
        net75793) );
  NAND2_X2 U6214 ( .A1(n4898), .A2(n5581), .ZN(dmem_addr_out[2]) );
  INV_X1 U6215 ( .A(n10115), .ZN(n5581) );
  NAND2_X4 U6216 ( .A1(net75845), .A2(net75846), .ZN(n10943) );
  NOR2_X4 U6217 ( .A1(net75847), .A2(n5583), .ZN(net75846) );
  AOI22_X4 U6218 ( .A1(REGFILE_reg_out_26__17_), .A2(net75439), .B1(
        REGFILE_reg_out_27__17_), .B2(net75440), .ZN(n5585) );
  INV_X8 U6219 ( .A(net76199), .ZN(net75440) );
  AOI22_X4 U6220 ( .A1(REGFILE_reg_out_24__17_), .A2(net75437), .B1(
        REGFILE_reg_out_25__17_), .B2(net75438), .ZN(n5586) );
  INV_X32 U6221 ( .A(net76197), .ZN(net75437) );
  NAND2_X4 U6222 ( .A1(net84277), .A2(n5576), .ZN(net76197) );
  INV_X8 U6223 ( .A(net87982), .ZN(net84277) );
  AND2_X4 U6224 ( .A1(net91646), .A2(net76204), .ZN(net120684) );
  NAND2_X4 U6225 ( .A1(net84277), .A2(net76204), .ZN(net76233) );
  NAND3_X4 U6226 ( .A1(net92446), .A2(net86794), .A3(net87981), .ZN(net87982)
         );
  INV_X32 U6227 ( .A(instruction[13]), .ZN(net87981) );
  MUX2_X2 U6228 ( .A(net87981), .B(net73529), .S(net73509), .Z(net73527) );
  INV_X32 U6229 ( .A(instruction[14]), .ZN(net82933) );
  NAND3_X4 U6230 ( .A1(net73511), .A2(n4843), .A3(net82598), .ZN(net76239) );
  NAND3_X4 U6231 ( .A1(net73511), .A2(net82933), .A3(net82598), .ZN(net123382)
         );
  AOI21_X1 U6232 ( .B1(net73878), .B2(net86794), .A(net73997), .ZN(net73900)
         );
  INV_X32 U6233 ( .A(instruction[15]), .ZN(net92446) );
  NAND3_X4 U6234 ( .A1(net89734), .A2(net92446), .A3(instruction[14]), .ZN(
        net90830) );
  NAND2_X4 U6235 ( .A1(net84754), .A2(n5576), .ZN(net76201) );
  INV_X16 U6236 ( .A(net76203), .ZN(net82613) );
  NOR2_X4 U6237 ( .A1(net75857), .A2(net75858), .ZN(net75845) );
  INV_X16 U6238 ( .A(net76236), .ZN(net75468) );
  NAND2_X4 U6239 ( .A1(net148494), .A2(net83408), .ZN(net76236) );
  NAND2_X2 U6240 ( .A1(net76206), .A2(net83408), .ZN(net76241) );
  NAND2_X2 U6241 ( .A1(net87806), .A2(n4797), .ZN(net76222) );
  NAND2_X4 U6242 ( .A1(net82618), .A2(instruction[12]), .ZN(net81601) );
  NAND2_X4 U6243 ( .A1(net87820), .A2(instruction[12]), .ZN(net88131) );
  INV_X8 U6244 ( .A(net76217), .ZN(net148494) );
  NAND2_X4 U6245 ( .A1(net148494), .A2(net76204), .ZN(net76224) );
  NAND2_X2 U6246 ( .A1(net91643), .A2(net148494), .ZN(net76257) );
  NAND2_X4 U6247 ( .A1(net91643), .A2(net76198), .ZN(net76237) );
  INV_X32 U6248 ( .A(instruction[13]), .ZN(net82598) );
  NAND3_X2 U6249 ( .A1(net82598), .A2(instruction[14]), .A3(instruction[15]), 
        .ZN(net85731) );
  AOI21_X1 U6250 ( .B1(net73878), .B2(net73511), .A(net73997), .ZN(net73902)
         );
  INV_X16 U6251 ( .A(net76233), .ZN(net82342) );
  NAND2_X4 U6252 ( .A1(net88253), .A2(net82618), .ZN(net76251) );
  NAND2_X4 U6253 ( .A1(net88253), .A2(n4820), .ZN(net81164) );
  INV_X32 U6254 ( .A(instruction[12]), .ZN(net88253) );
  NAND2_X2 U6255 ( .A1(REGFILE_reg_out_0__17_), .A2(net77312), .ZN(net74799)
         );
  NAND2_X2 U6256 ( .A1(REGFILE_reg_out_10__17_), .A2(net77348), .ZN(net74808)
         );
  NAND2_X4 U6257 ( .A1(n5587), .A2(net76202), .ZN(n5588) );
  NAND2_X4 U6258 ( .A1(net76208), .A2(n5587), .ZN(net76234) );
  OAI21_X4 U6259 ( .B1(net75842), .B2(net73697), .A(net75843), .ZN(net36463)
         );
  BUF_X32 U6260 ( .A(net75842), .Z(net148116) );
  INV_X4 U6261 ( .A(net73439), .ZN(net73416) );
  NAND2_X2 U6262 ( .A1(n5591), .A2(net70738), .ZN(n5590) );
  INV_X4 U6263 ( .A(net73780), .ZN(n5591) );
  INV_X4 U6264 ( .A(net73468), .ZN(n5589) );
  NAND2_X2 U6265 ( .A1(net77104), .A2(n4997), .ZN(net71227) );
  INV_X4 U6266 ( .A(net73429), .ZN(net73465) );
  INV_X4 U6267 ( .A(net73443), .ZN(net73427) );
  INV_X16 U6268 ( .A(net77106), .ZN(net77102) );
  NAND2_X2 U6269 ( .A1(net71269), .A2(net76650), .ZN(n5595) );
  INV_X4 U6270 ( .A(net70502), .ZN(net71269) );
  NAND2_X2 U6271 ( .A1(n5592), .A2(net77030), .ZN(n5594) );
  INV_X4 U6272 ( .A(net73771), .ZN(n5592) );
  XNOR2_X2 U6273 ( .A(n5592), .B(net73858), .ZN(net73778) );
  INV_X4 U6274 ( .A(net70504), .ZN(net71266) );
  NOR2_X2 U6275 ( .A1(n5596), .A2(net71302), .ZN(n5593) );
  INV_X4 U6276 ( .A(net70503), .ZN(net71302) );
  INV_X4 U6277 ( .A(dmem_read_in[1]), .ZN(n5597) );
  OAI211_X2 U6278 ( .C1(net73495), .C2(net73498), .A(net73496), .B(net73504), 
        .ZN(net73500) );
  INV_X4 U6279 ( .A(net73500), .ZN(net73494) );
  NOR2_X2 U6280 ( .A1(n5601), .A2(n5598), .ZN(net92782) );
  NAND2_X1 U6281 ( .A1(net70502), .A2(net70503), .ZN(n5598) );
  AND2_X2 U6282 ( .A1(net70504), .A2(net73585), .ZN(n5601) );
  NAND2_X4 U6283 ( .A1(multOut[1]), .A2(net81873), .ZN(net81874) );
  INV_X4 U6284 ( .A(net73585), .ZN(net81873) );
  NAND2_X2 U6285 ( .A1(net71271), .A2(n5599), .ZN(net70502) );
  XNOR2_X2 U6286 ( .A(net70731), .B(net70735), .ZN(n5599) );
  NAND3_X1 U6287 ( .A1(net71078), .A2(WIRE_ALU_A_MUX2TO1_32BIT_1__MUX_N1), 
        .A3(net36466), .ZN(net70503) );
  INV_X4 U6288 ( .A(net71273), .ZN(WIRE_ALU_A_MUX2TO1_32BIT_1__MUX_N1) );
  NAND3_X2 U6289 ( .A1(net71277), .A2(n5570), .A3(n5600), .ZN(net70504) );
  NOR2_X4 U6290 ( .A1(net71280), .A2(n5039), .ZN(n5600) );
  NAND2_X2 U6291 ( .A1(n5602), .A2(n5603), .ZN(net73585) );
  XNOR2_X2 U6292 ( .A(instruction[27]), .B(instruction[28]), .ZN(n5604) );
  INV_X4 U6293 ( .A(instruction[29]), .ZN(n5605) );
  OAI22_X2 U6294 ( .A1(instructionAddr_out[29]), .A2(n5605), .B1(net73394), 
        .B2(net73938), .ZN(net73400) );
  INV_X16 U6295 ( .A(net73629), .ZN(net74011) );
  INV_X4 U6296 ( .A(net73630), .ZN(net73646) );
  OAI211_X4 U6297 ( .C1(net73532), .C2(net73622), .A(net75792), .B(net75793), 
        .ZN(net75791) );
  INV_X4 U6298 ( .A(net73532), .ZN(net73495) );
  NAND2_X4 U6299 ( .A1(net75748), .A2(net75747), .ZN(dmem_write_out[13]) );
  OAI21_X4 U6300 ( .B1(dmem_write_out[13]), .B2(net75427), .A(n10945), .ZN(
        net72414) );
  NOR2_X4 U6301 ( .A1(net75759), .A2(net75760), .ZN(net75747) );
  NAND4_X2 U6302 ( .A1(net75764), .A2(net75761), .A3(n5606), .A4(net75763), 
        .ZN(net75760) );
  INV_X8 U6303 ( .A(net76234), .ZN(net83167) );
  INV_X2 U6304 ( .A(net84518), .ZN(n5608) );
  INV_X8 U6305 ( .A(net77752), .ZN(net77750) );
  NAND2_X4 U6306 ( .A1(net122022), .A2(net91646), .ZN(net76220) );
  INV_X8 U6307 ( .A(net76254), .ZN(n5607) );
  NAND2_X4 U6308 ( .A1(net76195), .A2(n5607), .ZN(net76199) );
  NAND3_X4 U6309 ( .A1(net73528), .A2(instruction[14]), .A3(instruction[15]), 
        .ZN(net76254) );
  INV_X32 U6310 ( .A(instruction[13]), .ZN(net73528) );
  NAND2_X1 U6311 ( .A1(net73878), .A2(net73528), .ZN(net73974) );
  INV_X4 U6312 ( .A(net76262), .ZN(net91643) );
  NAND2_X4 U6313 ( .A1(net91643), .A2(net121496), .ZN(net76258) );
  NAND2_X4 U6314 ( .A1(net73533), .A2(instruction[11]), .ZN(net76262) );
  INV_X8 U6315 ( .A(n4823), .ZN(net76238) );
  INV_X16 U6316 ( .A(net75791), .ZN(net75427) );
  INV_X2 U6317 ( .A(net83260), .ZN(net83261) );
  INV_X16 U6318 ( .A(net75481), .ZN(net77848) );
  INV_X8 U6319 ( .A(net77848), .ZN(net77846) );
  INV_X16 U6320 ( .A(n5704), .ZN(n5609) );
  NAND2_X1 U6321 ( .A1(n4888), .A2(REGFILE_reg_out_22__16_), .ZN(n9234) );
  AOI22_X4 U6322 ( .A1(REGFILE_reg_out_17__16_), .A2(net77796), .B1(
        REGFILE_reg_out_18__16_), .B2(n5890), .ZN(n6562) );
  AOI22_X4 U6323 ( .A1(REGFILE_reg_out_4__16_), .A2(n5678), .B1(n5756), .B2(
        net75452), .ZN(n6573) );
  INV_X2 U6324 ( .A(n5610), .ZN(n5611) );
  NAND2_X4 U6325 ( .A1(net77460), .A2(REGFILE_reg_out_21__28_), .ZN(n7008) );
  INV_X2 U6326 ( .A(n5612), .ZN(n5613) );
  OAI21_X2 U6327 ( .B1(n7027), .B2(n7026), .A(n6019), .ZN(n7039) );
  INV_X16 U6328 ( .A(instruction[9]), .ZN(net87097) );
  AOI22_X4 U6329 ( .A1(REGFILE_reg_out_31__12_), .A2(net77668), .B1(
        REGFILE_reg_out_3__12_), .B2(net77676), .ZN(n6654) );
  AOI22_X4 U6330 ( .A1(REGFILE_reg_out_23__18_), .A2(net77828), .B1(
        REGFILE_reg_out_22__18_), .B2(net77836), .ZN(n6532) );
  NAND2_X1 U6331 ( .A1(n4889), .A2(REGFILE_reg_out_6__16_), .ZN(n9262) );
  INV_X2 U6332 ( .A(n5614), .ZN(n5615) );
  AOI22_X4 U6333 ( .A1(REGFILE_reg_out_31__10_), .A2(net77666), .B1(
        REGFILE_reg_out_3__10_), .B2(n5609), .ZN(n6698) );
  AOI22_X2 U6334 ( .A1(REGFILE_reg_out_24__8_), .A2(net75437), .B1(
        REGFILE_reg_out_25__8_), .B2(net75438), .ZN(n6746) );
  AOI22_X1 U6335 ( .A1(REGFILE_reg_out_24__4_), .A2(net75437), .B1(
        REGFILE_reg_out_25__4_), .B2(net75438), .ZN(n6822) );
  AOI22_X2 U6336 ( .A1(REGFILE_reg_out_19__10_), .A2(net77810), .B1(
        REGFILE_reg_out_1__10_), .B2(net75478), .ZN(n6689) );
  AOI22_X2 U6337 ( .A1(REGFILE_reg_out_24__22_), .A2(net75437), .B1(
        REGFILE_reg_out_25__22_), .B2(net124970), .ZN(n6448) );
  AOI22_X2 U6338 ( .A1(REGFILE_reg_out_0__9_), .A2(net82342), .B1(
        REGFILE_reg_out_10__9_), .B2(net75464), .ZN(n6714) );
  INV_X16 U6339 ( .A(net77720), .ZN(net77716) );
  INV_X2 U6340 ( .A(n5617), .ZN(n5618) );
  NAND2_X1 U6341 ( .A1(REGFILE_reg_out_20__0_), .A2(net77386), .ZN(n8247) );
  NAND2_X1 U6342 ( .A1(REGFILE_reg_out_20__1_), .A2(net77386), .ZN(n8203) );
  NAND2_X1 U6343 ( .A1(REGFILE_reg_out_28__19_), .A2(net77386), .ZN(n7405) );
  NAND2_X1 U6344 ( .A1(REGFILE_reg_out_28__20_), .A2(net77386), .ZN(n7361) );
  NAND2_X1 U6345 ( .A1(REGFILE_reg_out_20__20_), .A2(net77386), .ZN(n7371) );
  NAND2_X1 U6346 ( .A1(REGFILE_reg_out_12__20_), .A2(net77386), .ZN(n7381) );
  NAND2_X1 U6347 ( .A1(REGFILE_reg_out_4__20_), .A2(net77386), .ZN(n7391) );
  NAND2_X1 U6348 ( .A1(REGFILE_reg_out_28__21_), .A2(net77386), .ZN(n7312) );
  NAND2_X1 U6349 ( .A1(REGFILE_reg_out_4__21_), .A2(net77386), .ZN(n7322) );
  NAND2_X1 U6350 ( .A1(REGFILE_reg_out_12__21_), .A2(net77386), .ZN(n7332) );
  NAND2_X1 U6351 ( .A1(REGFILE_reg_out_20__21_), .A2(net77386), .ZN(n7342) );
  NAND2_X1 U6352 ( .A1(REGFILE_reg_out_4__22_), .A2(net77386), .ZN(n7277) );
  NAND2_X1 U6353 ( .A1(REGFILE_reg_out_12__22_), .A2(net77386), .ZN(n7287) );
  NAND2_X1 U6354 ( .A1(REGFILE_reg_out_20__22_), .A2(net77386), .ZN(n7297) );
  NAND2_X1 U6355 ( .A1(net77386), .A2(REGFILE_reg_out_28__27_), .ZN(n7048) );
  NAND2_X1 U6356 ( .A1(net77386), .A2(REGFILE_reg_out_12__27_), .ZN(n7068) );
  NAND2_X1 U6357 ( .A1(net77386), .A2(REGFILE_reg_out_4__27_), .ZN(n7078) );
  NAND2_X1 U6358 ( .A1(net77386), .A2(REGFILE_reg_out_12__28_), .ZN(n7024) );
  INV_X16 U6359 ( .A(net77320), .ZN(net77318) );
  INV_X16 U6360 ( .A(n5703), .ZN(net77668) );
  INV_X16 U6361 ( .A(n5703), .ZN(net77666) );
  INV_X16 U6362 ( .A(n5703), .ZN(net77670) );
  NAND2_X1 U6363 ( .A1(REGFILE_reg_out_5__18_), .A2(net77456), .ZN(n7473) );
  AOI22_X2 U6364 ( .A1(REGFILE_reg_out_4__18_), .A2(net75451), .B1(
        REGFILE_reg_out_5__18_), .B2(net75452), .ZN(n6541) );
  AOI22_X4 U6365 ( .A1(REGFILE_reg_out_9__16_), .A2(net77700), .B1(n5668), 
        .B2(net75454), .ZN(n6574) );
  INV_X8 U6366 ( .A(net76239), .ZN(net91646) );
  AOI22_X2 U6367 ( .A1(REGFILE_reg_out_9__13_), .A2(net77700), .B1(n5716), 
        .B2(net75454), .ZN(n6636) );
  AOI22_X4 U6368 ( .A1(REGFILE_reg_out_7__17_), .A2(net77714), .B1(
        REGFILE_reg_out_6__17_), .B2(net75456), .ZN(n6561) );
  INV_X4 U6369 ( .A(net148735), .ZN(net148736) );
  NAND2_X1 U6370 ( .A1(n4891), .A2(REGFILE_reg_out_16__13_), .ZN(n9441) );
  NAND2_X1 U6371 ( .A1(net77308), .A2(REGFILE_reg_out_16__13_), .ZN(n7675) );
  BUF_X32 U6372 ( .A(net73851), .Z(n5619) );
  OAI22_X1 U6373 ( .A1(net78235), .A2(n6090), .B1(n6191), .B2(net76658), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  NAND2_X1 U6374 ( .A1(REGFILE_reg_out_1__16_), .A2(net77526), .ZN(n7561) );
  INV_X32 U6375 ( .A(net77800), .ZN(net77796) );
  INV_X16 U6376 ( .A(n6224), .ZN(n6896) );
  AOI22_X4 U6377 ( .A1(REGFILE_reg_out_29__17_), .A2(net77652), .B1(
        REGFILE_reg_out_28__17_), .B2(n5751), .ZN(net75849) );
  AOI22_X4 U6378 ( .A1(REGFILE_reg_out_11__10_), .A2(net77746), .B1(n4817), 
        .B2(net75466), .ZN(n6693) );
  NOR2_X4 U6379 ( .A1(n6453), .A2(n6452), .ZN(n6454) );
  NAND2_X1 U6381 ( .A1(REGFILE_reg_out_28__12_), .A2(n6177), .ZN(n9154) );
  NAND2_X1 U6382 ( .A1(REGFILE_reg_out_28__12_), .A2(net77380), .ZN(n7711) );
  NAND4_X2 U6383 ( .A1(n6924), .A2(n6923), .A3(n6921), .A4(n6922), .ZN(
        net73851) );
  NAND2_X1 U6384 ( .A1(REGFILE_reg_out_18__16_), .A2(net77346), .ZN(n7544) );
  INV_X8 U6385 ( .A(net77704), .ZN(net77702) );
  INV_X16 U6386 ( .A(net77704), .ZN(net77698) );
  INV_X16 U6387 ( .A(net75453), .ZN(net77704) );
  NAND2_X1 U6388 ( .A1(net77550), .A2(REGFILE_reg_out_30__28_), .ZN(n7001) );
  NAND2_X1 U6389 ( .A1(net77550), .A2(REGFILE_reg_out_22__28_), .ZN(n7011) );
  NAND2_X1 U6390 ( .A1(net77550), .A2(REGFILE_reg_out_6__28_), .ZN(n7031) );
  INV_X16 U6391 ( .A(net77848), .ZN(net77844) );
  INV_X16 U6392 ( .A(net77848), .ZN(net77842) );
  AOI22_X2 U6393 ( .A1(REGFILE_reg_out_11__17_), .A2(net77748), .B1(
        REGFILE_reg_out_12__17_), .B2(net75466), .ZN(net75861) );
  INV_X4 U6394 ( .A(n10378), .ZN(n10914) );
  NAND2_X4 U6395 ( .A1(n6551), .A2(n6550), .ZN(dmem_write_out[18]) );
  AOI22_X1 U6396 ( .A1(REGFILE_reg_out_0__3_), .A2(net82342), .B1(
        REGFILE_reg_out_10__3_), .B2(net75464), .ZN(n6834) );
  NAND2_X1 U6397 ( .A1(REGFILE_reg_out_28__11_), .A2(n6175), .ZN(n9909) );
  NAND2_X1 U6398 ( .A1(REGFILE_reg_out_28__11_), .A2(net77380), .ZN(n7755) );
  AOI22_X2 U6399 ( .A1(REGFILE_reg_out_29__11_), .A2(net77652), .B1(
        REGFILE_reg_out_28__11_), .B2(n5751), .ZN(n6683) );
  AOI22_X4 U6400 ( .A1(REGFILE_reg_out_23__10_), .A2(net77826), .B1(
        REGFILE_reg_out_22__10_), .B2(net77834), .ZN(n6690) );
  NAND2_X1 U6401 ( .A1(REGFILE_reg_out_13__10_), .A2(net77456), .ZN(n7813) );
  NAND2_X1 U6402 ( .A1(REGFILE_reg_out_6__16_), .A2(net77562), .ZN(n7562) );
  NAND2_X1 U6403 ( .A1(REGFILE_reg_out_2__3_), .A2(net77338), .ZN(n8134) );
  AOI22_X2 U6404 ( .A1(REGFILE_reg_out_14__23_), .A2(net77778), .B1(
        REGFILE_reg_out_13__23_), .B2(n6009), .ZN(n6418) );
  AOI22_X2 U6405 ( .A1(REGFILE_reg_out_14__8_), .A2(net77778), .B1(
        REGFILE_reg_out_13__8_), .B2(n6009), .ZN(n6739) );
  AOI22_X2 U6406 ( .A1(REGFILE_reg_out_23__3_), .A2(net77826), .B1(
        REGFILE_reg_out_22__3_), .B2(net77834), .ZN(n6832) );
  NAND2_X1 U6407 ( .A1(REGFILE_reg_out_12__12_), .A2(n4873), .ZN(n9120) );
  NAND2_X1 U6408 ( .A1(net77380), .A2(REGFILE_reg_out_12__12_), .ZN(n7731) );
  NAND3_X4 U6409 ( .A1(net92447), .A2(net82932), .A3(instruction[13]), .ZN(
        net148091) );
  NAND2_X1 U6410 ( .A1(n4804), .A2(REGFILE_reg_out_15__12_), .ZN(n9126) );
  NAND2_X1 U6411 ( .A1(REGFILE_reg_out_15__12_), .A2(net77488), .ZN(n7726) );
  AOI22_X4 U6412 ( .A1(REGFILE_reg_out_11__16_), .A2(net77748), .B1(n5618), 
        .B2(net83168), .ZN(n6567) );
  INV_X16 U6413 ( .A(n5623), .ZN(net75478) );
  NAND2_X4 U6414 ( .A1(net76204), .A2(net87806), .ZN(n5623) );
  INV_X8 U6415 ( .A(net88102), .ZN(net87806) );
  NAND2_X4 U6416 ( .A1(net76238), .A2(net87806), .ZN(net76249) );
  NAND3_X4 U6417 ( .A1(net89734), .A2(n4840), .A3(instruction[15]), .ZN(
        net88102) );
  INV_X32 U6418 ( .A(instruction[14]), .ZN(net82932) );
  INV_X16 U6419 ( .A(instruction[13]), .ZN(net89734) );
  INV_X16 U6420 ( .A(net75477), .ZN(net77816) );
  INV_X16 U6421 ( .A(net77816), .ZN(net77810) );
  INV_X8 U6422 ( .A(net76253), .ZN(net75477) );
  OR2_X2 U6423 ( .A1(n5578), .A2(net80211), .ZN(net78104) );
  AND2_X4 U6424 ( .A1(net78104), .A2(net78105), .ZN(net75415) );
  NAND3_X4 U6425 ( .A1(instruction[8]), .A2(net73989), .A3(instruction[10]), 
        .ZN(net75423) );
  OAI22_X2 U6426 ( .A1(net78108), .A2(net77464), .B1(net78109), .B2(net75422), 
        .ZN(net78107) );
  INV_X16 U6427 ( .A(net75423), .ZN(net77474) );
  INV_X32 U6428 ( .A(instruction[9]), .ZN(net73989) );
  NAND2_X2 U6429 ( .A1(net105318), .A2(net70497), .ZN(dmem_addr_out[0]) );
  INV_X4 U6430 ( .A(net70689), .ZN(net70497) );
  NAND2_X2 U6431 ( .A1(net70685), .A2(net70497), .ZN(net70687) );
  OAI22_X2 U6432 ( .A1(net70690), .A2(net70691), .B1(net81873), .B2(net70692), 
        .ZN(net70689) );
  INV_X4 U6433 ( .A(net105376), .ZN(net70692) );
  AOI22_X2 U6434 ( .A1(net70692), .A2(net70684), .B1(net70685), .B2(n4915), 
        .ZN(net70541) );
  XNOR2_X2 U6435 ( .A(n5625), .B(n5626), .ZN(net70690) );
  INV_X4 U6436 ( .A(net70730), .ZN(n5626) );
  NAND2_X2 U6437 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_1__MUX_N1), .A2(net70734), 
        .ZN(n5627) );
  INV_X4 U6438 ( .A(net70735), .ZN(net70732) );
  XNOR2_X2 U6439 ( .A(net70729), .B(net71027), .ZN(n5625) );
  XNOR2_X2 U6440 ( .A(net77042), .B(net70535), .ZN(net70729) );
  NAND4_X2 U6441 ( .A1(net73611), .A2(net73612), .A3(net73613), .A4(n5629), 
        .ZN(n5628) );
  NOR3_X4 U6442 ( .A1(net73615), .A2(net73616), .A3(n5630), .ZN(n5629) );
  NOR3_X4 U6443 ( .A1(n4971), .A2(net73619), .A3(net73620), .ZN(n5630) );
  INV_X4 U6444 ( .A(instruction[30]), .ZN(net73619) );
  INV_X16 U6445 ( .A(net75422), .ZN(net77400) );
  INV_X2 U6446 ( .A(net80440), .ZN(n5631) );
  NAND3_X4 U6447 ( .A1(net73987), .A2(net87097), .A3(instruction[8]), .ZN(
        net75422) );
  NAND2_X2 U6448 ( .A1(net73878), .A2(net87097), .ZN(net73988) );
  INV_X32 U6449 ( .A(instruction[10]), .ZN(net73987) );
  NOR2_X4 U6450 ( .A1(multOut[0]), .A2(net70687), .ZN(net70537) );
  NOR2_X4 U6451 ( .A1(n5634), .A2(n5635), .ZN(n5636) );
  INV_X4 U6452 ( .A(net70693), .ZN(n5635) );
  INV_X4 U6453 ( .A(net73585), .ZN(net76452) );
  NOR2_X4 U6454 ( .A1(n9854), .A2(net70718), .ZN(n5638) );
  NOR2_X4 U6455 ( .A1(net70709), .A2(net70710), .ZN(n5634) );
  INV_X4 U6456 ( .A(n5632), .ZN(n5637) );
  AOI21_X4 U6457 ( .B1(net105352), .B2(n5633), .A(n9606), .ZN(n5632) );
  NAND2_X2 U6458 ( .A1(net70713), .A2(net78051), .ZN(n5633) );
  INV_X4 U6459 ( .A(net36414), .ZN(net78050) );
  OAI21_X2 U6460 ( .B1(net76154), .B2(net78056), .A(n5639), .ZN(net36414) );
  INV_X8 U6461 ( .A(n5640), .ZN(net75844) );
  NAND2_X2 U6462 ( .A1(net77272), .A2(net78055), .ZN(n5640) );
  INV_X32 U6463 ( .A(net77280), .ZN(net77272) );
  INV_X16 U6464 ( .A(net73665), .ZN(net77280) );
  NOR2_X4 U6465 ( .A1(net77280), .A2(net73908), .ZN(net75792) );
  NAND2_X4 U6466 ( .A1(net76181), .A2(n5641), .ZN(net73665) );
  NOR3_X4 U6467 ( .A1(net74029), .A2(instruction[1]), .A3(instruction[0]), 
        .ZN(n5641) );
  NAND3_X4 U6468 ( .A1(net75397), .A2(net75395), .A3(net75396), .ZN(aluA[31])
         );
  AOI22_X4 U6469 ( .A1(net77276), .A2(instruction[30]), .B1(net73831), .B2(
        n4963), .ZN(net75367) );
  NOR2_X4 U6470 ( .A1(n5643), .A2(net73503), .ZN(net76181) );
  NAND2_X4 U6471 ( .A1(instruction[3]), .A2(instruction[4]), .ZN(n5643) );
  INV_X32 U6472 ( .A(instruction[5]), .ZN(net73503) );
  INV_X32 U6473 ( .A(n5644), .ZN(net77588) );
  INV_X4 U6474 ( .A(net73836), .ZN(n5642) );
  AOI22_X4 U6475 ( .A1(net77276), .A2(instruction[31]), .B1(net73849), .B2(
        n4897), .ZN(net75395) );
  NAND2_X4 U6476 ( .A1(net73837), .A2(n4897), .ZN(net75368) );
  INV_X32 U6477 ( .A(net77296), .ZN(net77290) );
  BUF_X32 U6478 ( .A(net73849), .Z(net80390) );
  INV_X4 U6479 ( .A(net78126), .ZN(net75414) );
  OAI22_X2 U6480 ( .A1(net78127), .A2(net77512), .B1(net78128), .B2(net75424), 
        .ZN(net78126) );
  INV_X32 U6481 ( .A(net77512), .ZN(net77508) );
  INV_X8 U6482 ( .A(net75425), .ZN(net74050) );
  INV_X4 U6483 ( .A(net82513), .ZN(net75416) );
  INV_X32 U6484 ( .A(n5647), .ZN(net77406) );
  INV_X8 U6485 ( .A(n5645), .ZN(n5647) );
  NAND3_X4 U6486 ( .A1(instruction[10]), .A2(net123931), .A3(instruction[9]), 
        .ZN(n5646) );
  INV_X32 U6487 ( .A(instruction[8]), .ZN(net123931) );
  NAND3_X4 U6488 ( .A1(net123931), .A2(net73987), .A3(instruction[9]), .ZN(
        net85371) );
  AOI22_X4 U6489 ( .A1(net82500), .A2(net77514), .B1(net80443), .B2(net77298), 
        .ZN(net75417) );
  INV_X16 U6490 ( .A(net77326), .ZN(net77298) );
  INV_X16 U6491 ( .A(net77328), .ZN(net77326) );
  INV_X16 U6492 ( .A(net77326), .ZN(net77300) );
  NAND2_X2 U6494 ( .A1(net76238), .A2(net84754), .ZN(n6224) );
  NAND2_X1 U6495 ( .A1(net77562), .A2(REGFILE_reg_out_14__27_), .ZN(n7065) );
  NAND2_X1 U6496 ( .A1(REGFILE_reg_out_30__0_), .A2(net77550), .ZN(n8234) );
  NAND2_X1 U6497 ( .A1(REGFILE_reg_out_30__1_), .A2(net77554), .ZN(n8190) );
  NAND2_X1 U6498 ( .A1(REGFILE_reg_out_14__1_), .A2(net77554), .ZN(n8210) );
  NAND2_X1 U6499 ( .A1(net77550), .A2(REGFILE_reg_out_6__27_), .ZN(n7075) );
  NAND2_X1 U6500 ( .A1(net77550), .A2(REGFILE_reg_out_14__28_), .ZN(n7021) );
  NAND2_X1 U6501 ( .A1(REGFILE_reg_out_22__1_), .A2(net77550), .ZN(n8200) );
  NAND2_X1 U6502 ( .A1(REGFILE_reg_out_22__0_), .A2(net77550), .ZN(n8244) );
  NAND2_X1 U6503 ( .A1(REGFILE_reg_out_14__0_), .A2(net77550), .ZN(n8254) );
  NAND2_X1 U6504 ( .A1(REGFILE_reg_out_6__1_), .A2(net77554), .ZN(n8220) );
  NAND2_X1 U6505 ( .A1(net77550), .A2(REGFILE_reg_out_30__27_), .ZN(n7045) );
  NAND4_X2 U6506 ( .A1(n6973), .A2(n6972), .A3(n6971), .A4(n6970), .ZN(n6974)
         );
  AOI22_X2 U6507 ( .A1(n5789), .A2(net77478), .B1(n5896), .B2(net77550), .ZN(
        n6927) );
  AOI22_X2 U6508 ( .A1(REGFILE_reg_out_23__31_), .A2(net77478), .B1(n5718), 
        .B2(net77550), .ZN(n6924) );
  AOI22_X2 U6509 ( .A1(n5795), .A2(net77478), .B1(n5926), .B2(net77550), .ZN(
        n6945) );
  INV_X16 U6510 ( .A(net77428), .ZN(net77422) );
  INV_X16 U6511 ( .A(net77400), .ZN(net77392) );
  INV_X16 U6512 ( .A(net77394), .ZN(net77382) );
  NOR2_X2 U6513 ( .A1(n5988), .A2(net77392), .ZN(n5754) );
  INV_X16 U6514 ( .A(instruction[13]), .ZN(net87495) );
  INV_X32 U6515 ( .A(net77720), .ZN(net77714) );
  NOR2_X2 U6516 ( .A1(n6751), .A2(n6750), .ZN(n6752) );
  INV_X16 U6517 ( .A(net77430), .ZN(net77424) );
  NAND2_X4 U6518 ( .A1(net88253), .A2(net87820), .ZN(n5706) );
  AOI22_X2 U6519 ( .A1(REGFILE_reg_out_11__11_), .A2(net77748), .B1(n5872), 
        .B2(net83168), .ZN(n6671) );
  NAND2_X4 U6520 ( .A1(net84754), .A2(net76238), .ZN(n5649) );
  AOI22_X1 U6521 ( .A1(REGFILE_reg_out_0__4_), .A2(net82342), .B1(
        REGFILE_reg_out_10__4_), .B2(net75464), .ZN(n6812) );
  NAND4_X2 U6522 ( .A1(n6393), .A2(n6394), .A3(n6395), .A4(n6392), .ZN(n6396)
         );
  INV_X4 U6523 ( .A(net77616), .ZN(net77614) );
  OAI21_X1 U6524 ( .B1(n6529), .B2(net78055), .A(n6528), .ZN(n5650) );
  OAI21_X1 U6525 ( .B1(dmem_write_out[27]), .B2(net78056), .A(n6343), .ZN(
        n5652) );
  OAI21_X2 U6526 ( .B1(n10355), .B2(n10354), .A(n10353), .ZN(n10358) );
  AOI22_X4 U6527 ( .A1(REGFILE_reg_out_4__11_), .A2(n5679), .B1(
        REGFILE_reg_out_5__11_), .B2(net84475), .ZN(n6677) );
  NAND2_X1 U6528 ( .A1(REGFILE_reg_out_16__15_), .A2(net77310), .ZN(n7587) );
  AOI22_X2 U6529 ( .A1(REGFILE_reg_out_29__25_), .A2(net77650), .B1(
        REGFILE_reg_out_28__25_), .B2(n6911), .ZN(n6385) );
  AOI22_X1 U6530 ( .A1(REGFILE_reg_out_24__3_), .A2(net75437), .B1(
        REGFILE_reg_out_25__3_), .B2(net75438), .ZN(n6844) );
  OAI211_X4 U6531 ( .C1(n10045), .C2(net76646), .A(net70740), .B(n10044), .ZN(
        n10046) );
  AOI22_X2 U6532 ( .A1(REGFILE_reg_out_11__22_), .A2(net77750), .B1(
        REGFILE_reg_out_12__22_), .B2(net75466), .ZN(n6439) );
  AOI22_X1 U6533 ( .A1(REGFILE_reg_out_11__4_), .A2(net77746), .B1(
        REGFILE_reg_out_12__4_), .B2(net75466), .ZN(n6813) );
  AOI22_X1 U6534 ( .A1(REGFILE_reg_out_30__26_), .A2(net77638), .B1(
        REGFILE_reg_out_2__26_), .B2(net75442), .ZN(n6360) );
  AOI22_X1 U6535 ( .A1(REGFILE_reg_out_30__2_), .A2(net77634), .B1(
        REGFILE_reg_out_2__2_), .B2(net75442), .ZN(n6868) );
  INV_X32 U6536 ( .A(instruction[8]), .ZN(net123932) );
  AOI22_X4 U6538 ( .A1(REGFILE_reg_out_31__11_), .A2(net77668), .B1(
        REGFILE_reg_out_3__11_), .B2(net77676), .ZN(n6676) );
  NAND2_X1 U6539 ( .A1(REGFILE_reg_out_5__15_), .A2(net77454), .ZN(n7603) );
  AOI22_X2 U6540 ( .A1(REGFILE_reg_out_4__15_), .A2(net75451), .B1(
        REGFILE_reg_out_5__15_), .B2(net84475), .ZN(n6595) );
  NAND2_X1 U6541 ( .A1(net73878), .A2(net90864), .ZN(n8380) );
  NAND2_X2 U6542 ( .A1(REGFILE_reg_out_7__30_), .A2(net77478), .ZN(n5654) );
  NAND2_X2 U6543 ( .A1(REGFILE_reg_out_6__30_), .A2(net77550), .ZN(n5655) );
  INV_X16 U6544 ( .A(net77506), .ZN(net77478) );
  NAND2_X1 U6545 ( .A1(net77298), .A2(REGFILE_reg_out_24__28_), .ZN(n7002) );
  NAND2_X1 U6548 ( .A1(REGFILE_reg_out_27__17_), .A2(net77420), .ZN(n7494) );
  INV_X8 U6549 ( .A(net76256), .ZN(net76206) );
  AOI22_X1 U6550 ( .A1(REGFILE_reg_out_19__3_), .A2(net77810), .B1(
        REGFILE_reg_out_1__3_), .B2(net75478), .ZN(n6831) );
  AOI22_X1 U6551 ( .A1(REGFILE_reg_out_19__25_), .A2(net77814), .B1(
        REGFILE_reg_out_1__25_), .B2(net75478), .ZN(n6369) );
  INV_X16 U6552 ( .A(net77832), .ZN(net77826) );
  NAND2_X1 U6553 ( .A1(REGFILE_reg_out_29__0_), .A2(net77444), .ZN(n8231) );
  NAND2_X1 U6554 ( .A1(REGFILE_reg_out_21__0_), .A2(net77444), .ZN(n8241) );
  NAND2_X1 U6555 ( .A1(REGFILE_reg_out_13__0_), .A2(net77444), .ZN(n8251) );
  NAND2_X1 U6556 ( .A1(REGFILE_reg_out_29__1_), .A2(net77444), .ZN(n8187) );
  NAND2_X1 U6557 ( .A1(REGFILE_reg_out_21__1_), .A2(net77444), .ZN(n8197) );
  NAND2_X1 U6558 ( .A1(REGFILE_reg_out_13__1_), .A2(net77444), .ZN(n8207) );
  NAND2_X1 U6559 ( .A1(REGFILE_reg_out_5__1_), .A2(net77444), .ZN(n8217) );
  NAND2_X1 U6560 ( .A1(net77444), .A2(REGFILE_reg_out_29__27_), .ZN(n7042) );
  NAND2_X1 U6561 ( .A1(net77444), .A2(REGFILE_reg_out_13__27_), .ZN(n7062) );
  NAND2_X1 U6562 ( .A1(net77444), .A2(REGFILE_reg_out_5__27_), .ZN(n7072) );
  NAND2_X1 U6563 ( .A1(net77444), .A2(REGFILE_reg_out_13__28_), .ZN(n7018) );
  BUF_X32 U6564 ( .A(n5851), .Z(n5931) );
  INV_X16 U6565 ( .A(net77800), .ZN(net77798) );
  AOI22_X4 U6566 ( .A1(REGFILE_reg_out_9__15_), .A2(net77700), .B1(
        REGFILE_reg_out_8__15_), .B2(n4829), .ZN(n6596) );
  INV_X32 U6567 ( .A(net77856), .ZN(net77852) );
  AOI22_X4 U6568 ( .A1(REGFILE_reg_out_7__16_), .A2(net77714), .B1(n4860), 
        .B2(net75456), .ZN(n6575) );
  NAND2_X1 U6569 ( .A1(net77382), .A2(REGFILE_reg_out_12__16_), .ZN(n7555) );
  AOI22_X1 U6570 ( .A1(REGFILE_reg_out_7__4_), .A2(net75455), .B1(
        REGFILE_reg_out_6__4_), .B2(net75456), .ZN(n6821) );
  AOI22_X1 U6571 ( .A1(REGFILE_reg_out_7__5_), .A2(net75455), .B1(
        REGFILE_reg_out_6__5_), .B2(net75456), .ZN(n6799) );
  INV_X1 U6572 ( .A(n4864), .ZN(n5805) );
  INV_X4 U6573 ( .A(dmem_write_out[24]), .ZN(n6410) );
  INV_X4 U6574 ( .A(net77324), .ZN(net77312) );
  INV_X4 U6575 ( .A(net77324), .ZN(net77310) );
  INV_X4 U6576 ( .A(net77324), .ZN(net77308) );
  AOI22_X2 U6577 ( .A1(REGFILE_reg_out_17__24_), .A2(net77798), .B1(
        REGFILE_reg_out_18__24_), .B2(n5890), .ZN(net76034) );
  AOI22_X4 U6578 ( .A1(REGFILE_reg_out_29__18_), .A2(net77652), .B1(
        REGFILE_reg_out_28__18_), .B2(n5751), .ZN(n6547) );
  NAND2_X2 U6579 ( .A1(instruction[28]), .A2(net77276), .ZN(n5658) );
  NAND2_X4 U6580 ( .A1(n5657), .A2(n5658), .ZN(aluA[28]) );
  INV_X8 U6581 ( .A(net77464), .ZN(net77460) );
  BUF_X8 U6582 ( .A(net36470), .Z(net85047) );
  INV_X4 U6583 ( .A(n10909), .ZN(n5659) );
  OAI22_X4 U6584 ( .A1(n5823), .A2(net86238), .B1(n5999), .B2(net93763), .ZN(
        n5822) );
  AOI22_X4 U6585 ( .A1(REGFILE_reg_out_9__18_), .A2(net77700), .B1(
        REGFILE_reg_out_8__18_), .B2(n4829), .ZN(n6542) );
  AOI22_X4 U6586 ( .A1(REGFILE_reg_out_9__14_), .A2(net77700), .B1(
        REGFILE_reg_out_8__14_), .B2(net75454), .ZN(n6620) );
  NAND2_X2 U6587 ( .A1(n6807), .A2(n6806), .ZN(dmem_write_out[5]) );
  AOI22_X2 U6588 ( .A1(REGFILE_reg_out_11__5_), .A2(net77746), .B1(
        REGFILE_reg_out_12__5_), .B2(net75466), .ZN(n6791) );
  NAND2_X1 U6589 ( .A1(n5902), .A2(net75464), .ZN(n5946) );
  AOI22_X2 U6590 ( .A1(REGFILE_reg_out_0__14_), .A2(net82342), .B1(n5829), 
        .B2(net83203), .ZN(n6612) );
  INV_X8 U6591 ( .A(net77324), .ZN(net77306) );
  INV_X8 U6592 ( .A(net77324), .ZN(net77304) );
  INV_X8 U6593 ( .A(net77324), .ZN(net77302) );
  AOI22_X4 U6594 ( .A1(REGFILE_reg_out_9__17_), .A2(net77700), .B1(
        REGFILE_reg_out_8__17_), .B2(net75454), .ZN(n6560) );
  AOI21_X1 U6595 ( .B1(n10418), .B2(n10384), .A(n10383), .ZN(n10388) );
  INV_X16 U6596 ( .A(n6010), .ZN(n5663) );
  INV_X8 U6597 ( .A(n6010), .ZN(n6009) );
  AOI22_X2 U6598 ( .A1(REGFILE_reg_out_11__9_), .A2(net77746), .B1(
        REGFILE_reg_out_12__9_), .B2(net75466), .ZN(n6715) );
  NAND2_X4 U6599 ( .A1(REGFILE_reg_out_4__29_), .A2(net77386), .ZN(n6961) );
  INV_X2 U6600 ( .A(n5665), .ZN(n5666) );
  INV_X2 U6601 ( .A(n5667), .ZN(n5668) );
  NAND2_X1 U6602 ( .A1(net73708), .A2(n6007), .ZN(n8694) );
  NAND2_X1 U6603 ( .A1(n10542), .A2(n6007), .ZN(n8766) );
  AOI22_X1 U6604 ( .A1(n9297), .A2(net72962), .B1(n4912), .B2(n6007), .ZN(
        n9769) );
  NAND2_X1 U6605 ( .A1(net70720), .A2(n6007), .ZN(n9081) );
  NAND2_X1 U6606 ( .A1(n9065), .A2(n6007), .ZN(n8837) );
  NAND2_X1 U6607 ( .A1(net70719), .A2(n6007), .ZN(n9943) );
  NAND2_X1 U6608 ( .A1(n6040), .A2(n6007), .ZN(n8711) );
  NAND2_X1 U6609 ( .A1(n6007), .A2(n10315), .ZN(n10316) );
  AOI21_X1 U6610 ( .B1(n8593), .B2(n6007), .A(n8592), .ZN(n8884) );
  XNOR2_X1 U6611 ( .A(n8591), .B(n6007), .ZN(n8773) );
  INV_X1 U6612 ( .A(n6007), .ZN(n8638) );
  NAND3_X2 U6613 ( .A1(n8694), .A2(n8693), .A3(n8692), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  NOR2_X2 U6614 ( .A1(n9769), .A2(n9770), .ZN(n8983) );
  OAI22_X1 U6615 ( .A1(n9771), .A2(n9770), .B1(n9769), .B2(n9802), .ZN(n9772)
         );
  NAND3_X2 U6616 ( .A1(n9081), .A2(n9080), .A3(n9079), .ZN(n9621) );
  NAND3_X2 U6617 ( .A1(n9944), .A2(n9943), .A3(n9942), .ZN(n10541) );
  OAI21_X2 U6618 ( .B1(n8884), .B2(n8883), .A(n8595), .ZN(n9776) );
  NOR2_X2 U6619 ( .A1(n6428), .A2(n6429), .ZN(n6430) );
  INV_X8 U6620 ( .A(net76259), .ZN(net121496) );
  INV_X4 U6621 ( .A(net148091), .ZN(net76208) );
  AOI22_X4 U6622 ( .A1(REGFILE_reg_out_17__13_), .A2(net77796), .B1(
        REGFILE_reg_out_18__13_), .B2(n6896), .ZN(n6630) );
  INV_X4 U6623 ( .A(n10392), .ZN(n10911) );
  NAND2_X2 U6624 ( .A1(REGFILE_reg_out_15__6_), .A2(net77484), .ZN(n7988) );
  AND2_X2 U6625 ( .A1(REGFILE_reg_out_11__24_), .A2(net77750), .ZN(n5669) );
  AND2_X2 U6626 ( .A1(REGFILE_reg_out_12__24_), .A2(net75466), .ZN(n5670) );
  NOR2_X2 U6627 ( .A1(n5669), .A2(n5670), .ZN(n6393) );
  INV_X2 U6628 ( .A(n5671), .ZN(n5672) );
  INV_X2 U6629 ( .A(n5673), .ZN(n5674) );
  AOI22_X2 U6630 ( .A1(REGFILE_reg_out_24__13_), .A2(net75437), .B1(n5940), 
        .B2(net124970), .ZN(n6638) );
  INV_X8 U6631 ( .A(net76255), .ZN(net77834) );
  AOI22_X1 U6632 ( .A1(REGFILE_reg_out_9__28_), .A2(net77702), .B1(
        REGFILE_reg_out_8__28_), .B2(n4829), .ZN(n6309) );
  AOI22_X2 U6633 ( .A1(REGFILE_reg_out_16__15_), .A2(net75467), .B1(n5782), 
        .B2(net75468), .ZN(n6590) );
  AOI22_X2 U6634 ( .A1(REGFILE_reg_out_26__22_), .A2(net75439), .B1(
        REGFILE_reg_out_27__22_), .B2(net89184), .ZN(n6449) );
  BUF_X16 U6635 ( .A(n10385), .Z(n5758) );
  NAND2_X2 U6636 ( .A1(REGFILE_reg_out_6__7_), .A2(net75456), .ZN(n5698) );
  OAI21_X1 U6637 ( .B1(n4819), .B2(net73697), .A(n6504), .ZN(n5675) );
  NAND2_X1 U6638 ( .A1(REGFILE_reg_out_3__15_), .A2(net77418), .ZN(n7610) );
  AOI22_X2 U6639 ( .A1(REGFILE_reg_out_31__15_), .A2(net77668), .B1(
        REGFILE_reg_out_3__15_), .B2(net77676), .ZN(n6594) );
  INV_X2 U6640 ( .A(n5676), .ZN(n5677) );
  AOI22_X2 U6641 ( .A1(REGFILE_reg_out_7__24_), .A2(net77716), .B1(
        REGFILE_reg_out_6__24_), .B2(net75456), .ZN(n6400) );
  NOR2_X2 U6642 ( .A1(n6827), .A2(n6826), .ZN(n6828) );
  NAND3_X1 U6643 ( .A1(net71078), .A2(n6007), .A3(n10926), .ZN(n8776) );
  XNOR2_X1 U6644 ( .A(n6007), .B(n10926), .ZN(n10441) );
  INV_X2 U6645 ( .A(n10926), .ZN(n10315) );
  NOR2_X4 U6646 ( .A1(n6539), .A2(n6538), .ZN(n6551) );
  NOR2_X4 U6647 ( .A1(n6549), .A2(n6548), .ZN(n6550) );
  AOI22_X1 U6648 ( .A1(REGFILE_reg_out_4__26_), .A2(n5678), .B1(
        REGFILE_reg_out_5__26_), .B2(net75452), .ZN(n6355) );
  AOI22_X2 U6649 ( .A1(REGFILE_reg_out_4__14_), .A2(n5678), .B1(
        REGFILE_reg_out_5__14_), .B2(net84475), .ZN(n6619) );
  NAND2_X4 U6650 ( .A1(net76206), .A2(net76195), .ZN(net76205) );
  AOI22_X2 U6651 ( .A1(REGFILE_reg_out_29__19_), .A2(net77652), .B1(
        REGFILE_reg_out_28__19_), .B2(n5751), .ZN(n6523) );
  INV_X8 U6652 ( .A(net76219), .ZN(n5678) );
  INV_X8 U6653 ( .A(net76219), .ZN(n5679) );
  INV_X8 U6654 ( .A(net76219), .ZN(net75451) );
  INV_X16 U6655 ( .A(n6239), .ZN(n6911) );
  NAND2_X1 U6656 ( .A1(net77346), .A2(REGFILE_reg_out_2__15_), .ZN(n7608) );
  NAND2_X1 U6657 ( .A1(n4804), .A2(REGFILE_reg_out_15__16_), .ZN(n9218) );
  OAI21_X4 U6658 ( .B1(n7037), .B2(n7036), .A(net77290), .ZN(n7038) );
  AOI22_X2 U6659 ( .A1(REGFILE_reg_out_17__5_), .A2(net77794), .B1(
        REGFILE_reg_out_18__5_), .B2(n5890), .ZN(n6786) );
  AOI22_X4 U6660 ( .A1(REGFILE_reg_out_16__20_), .A2(net77762), .B1(
        REGFILE_reg_out_15__20_), .B2(n5579), .ZN(n6488) );
  NAND2_X1 U6661 ( .A1(REGFILE_reg_out_12__19_), .A2(net77384), .ZN(n7425) );
  AOI22_X2 U6662 ( .A1(REGFILE_reg_out_11__19_), .A2(net77748), .B1(
        REGFILE_reg_out_12__19_), .B2(net83168), .ZN(n6511) );
  AOI22_X1 U6663 ( .A1(REGFILE_reg_out_11__23_), .A2(net77750), .B1(
        REGFILE_reg_out_12__23_), .B2(net83168), .ZN(n6416) );
  AOI22_X2 U6664 ( .A1(REGFILE_reg_out_26__8_), .A2(net75439), .B1(
        REGFILE_reg_out_27__8_), .B2(net89184), .ZN(n6747) );
  AOI22_X1 U6665 ( .A1(REGFILE_reg_out_24__23_), .A2(net75437), .B1(
        REGFILE_reg_out_25__23_), .B2(net124970), .ZN(n6425) );
  NAND2_X1 U6666 ( .A1(net77526), .A2(REGFILE_reg_out_25__15_), .ZN(n7575) );
  INV_X16 U6667 ( .A(n6006), .ZN(n6007) );
  AOI22_X1 U6668 ( .A1(REGFILE_reg_out_30__4_), .A2(net77634), .B1(
        REGFILE_reg_out_2__4_), .B2(net75442), .ZN(n6824) );
  INV_X2 U6669 ( .A(n5857), .ZN(n5684) );
  NAND2_X4 U6670 ( .A1(n10215), .A2(n10214), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  INV_X16 U6671 ( .A(net77784), .ZN(net77778) );
  AOI22_X4 U6672 ( .A1(REGFILE_reg_out_11__15_), .A2(net77748), .B1(n4854), 
        .B2(net83167), .ZN(n6589) );
  AOI22_X2 U6673 ( .A1(REGFILE_reg_out_16__19_), .A2(net77762), .B1(
        REGFILE_reg_out_15__19_), .B2(net75468), .ZN(n6512) );
  AOI22_X4 U6674 ( .A1(REGFILE_reg_out_9__8_), .A2(net77698), .B1(
        REGFILE_reg_out_8__8_), .B2(n4829), .ZN(n6744) );
  INV_X2 U6675 ( .A(n5686), .ZN(n5687) );
  AOI22_X2 U6676 ( .A1(REGFILE_reg_out_0__25_), .A2(net82342), .B1(
        REGFILE_reg_out_10__25_), .B2(net81764), .ZN(n6372) );
  INV_X16 U6677 ( .A(net77800), .ZN(net77794) );
  NOR2_X2 U6678 ( .A1(net91561), .A2(n5754), .ZN(n5753) );
  NAND2_X2 U6680 ( .A1(net76488), .A2(REGFILE_reg_out_31__2_), .ZN(n5690) );
  INV_X16 U6681 ( .A(n5696), .ZN(net77116) );
  INV_X16 U6682 ( .A(n5696), .ZN(net77114) );
  NAND2_X4 U6683 ( .A1(n5691), .A2(reset), .ZN(n5689) );
  OAI211_X4 U6684 ( .C1(net71394), .C2(net76646), .A(net70740), .B(n5692), 
        .ZN(n5691) );
  INV_X4 U6685 ( .A(dmem_read_in[2]), .ZN(n5694) );
  AND2_X2 U6686 ( .A1(net80797), .A2(n5698), .ZN(net75623) );
  NAND2_X4 U6687 ( .A1(net76206), .A2(net83210), .ZN(n5697) );
  INV_X8 U6688 ( .A(net81164), .ZN(net83210) );
  NAND2_X4 U6689 ( .A1(net83210), .A2(net76202), .ZN(net76203) );
  NAND2_X4 U6690 ( .A1(net121496), .A2(net83210), .ZN(net76219) );
  NAND2_X4 U6691 ( .A1(net76238), .A2(net76206), .ZN(net76255) );
  NAND3_X4 U6692 ( .A1(net82738), .A2(instruction[14]), .A3(instruction[13]), 
        .ZN(net76256) );
  MUX2_X2 U6693 ( .A(net82738), .B(net73512), .S(net73509), .Z(net73510) );
  NAND2_X1 U6694 ( .A1(REGFILE_reg_out_7__7_), .A2(net75455), .ZN(net80797) );
  INV_X8 U6695 ( .A(net76224), .ZN(net75455) );
  NAND2_X2 U6696 ( .A1(REGFILE_reg_out_6__7_), .A2(net77556), .ZN(net74359) );
  NAND2_X2 U6697 ( .A1(n4889), .A2(REGFILE_reg_out_6__7_), .ZN(net71936) );
  NAND2_X2 U6698 ( .A1(REGFILE_reg_out_7__7_), .A2(net77484), .ZN(net74361) );
  NAND2_X2 U6699 ( .A1(n4886), .A2(REGFILE_reg_out_7__7_), .ZN(net71934) );
  NAND2_X4 U6700 ( .A1(net75615), .A2(net75616), .ZN(dmem_write_out[7]) );
  OAI21_X4 U6701 ( .B1(dmem_write_out[7]), .B2(net75427), .A(n10945), .ZN(
        net72015) );
  NOR2_X4 U6702 ( .A1(net75617), .A2(net75618), .ZN(net75616) );
  NAND4_X2 U6703 ( .A1(net75619), .A2(net75620), .A3(net75621), .A4(n5699), 
        .ZN(net75618) );
  AOI22_X2 U6704 ( .A1(REGFILE_reg_out_24__7_), .A2(net75437), .B1(
        REGFILE_reg_out_25__7_), .B2(net124970), .ZN(n5699) );
  NAND2_X4 U6705 ( .A1(net76196), .A2(n5576), .ZN(net76194) );
  AOI22_X2 U6706 ( .A1(REGFILE_reg_out_26__23_), .A2(net77618), .B1(
        REGFILE_reg_out_27__23_), .B2(net77630), .ZN(net75995) );
  INV_X8 U6707 ( .A(net72015), .ZN(net36479) );
  AOI22_X2 U6708 ( .A1(REGFILE_reg_out_31__7_), .A2(net77666), .B1(
        REGFILE_reg_out_3__7_), .B2(n5609), .ZN(net75626) );
  INV_X32 U6709 ( .A(n5704), .ZN(net77676) );
  INV_X8 U6710 ( .A(n5705), .ZN(n5704) );
  NOR2_X4 U6711 ( .A1(net85731), .A2(n5706), .ZN(n5705) );
  INV_X8 U6712 ( .A(n5700), .ZN(n5703) );
  NOR2_X4 U6713 ( .A1(n4844), .A2(net87489), .ZN(n5700) );
  AOI22_X2 U6714 ( .A1(REGFILE_reg_out_4__7_), .A2(n5678), .B1(
        REGFILE_reg_out_5__7_), .B2(net84475), .ZN(net75625) );
  INV_X16 U6715 ( .A(n5702), .ZN(net84475) );
  NAND2_X4 U6716 ( .A1(net76204), .A2(n5701), .ZN(n5702) );
  INV_X8 U6717 ( .A(n4821), .ZN(n5701) );
  NAND2_X2 U6718 ( .A1(net76204), .A2(n5701), .ZN(net91311) );
  NAND2_X2 U6719 ( .A1(n5701), .A2(net76195), .ZN(net76209) );
  NAND2_X2 U6720 ( .A1(net76238), .A2(n5701), .ZN(net76260) );
  INV_X4 U6721 ( .A(net70868), .ZN(net70720) );
  INV_X4 U6722 ( .A(net72163), .ZN(net70697) );
  INV_X4 U6723 ( .A(net71027), .ZN(net36488) );
  INV_X4 U6724 ( .A(net71300), .ZN(net70696) );
  NAND2_X2 U6725 ( .A1(n5707), .A2(net73543), .ZN(net78014) );
  INV_X4 U6726 ( .A(aluA[16]), .ZN(n5708) );
  INV_X4 U6727 ( .A(net70706), .ZN(net105349) );
  AOI21_X4 U6728 ( .B1(n5709), .B2(net105360), .A(net70714), .ZN(net105352) );
  INV_X4 U6729 ( .A(net70845), .ZN(n5707) );
  INV_X4 U6730 ( .A(net70703), .ZN(n5710) );
  INV_X4 U6731 ( .A(net78014), .ZN(net70701) );
  NAND2_X2 U6732 ( .A1(net70719), .A2(net36391), .ZN(n5711) );
  OAI211_X2 U6733 ( .C1(net70868), .C2(n5708), .A(n5711), .B(net70717), .ZN(
        n5709) );
  NAND2_X1 U6734 ( .A1(REGFILE_reg_out_12__15_), .A2(net77382), .ZN(n7599) );
  NAND2_X1 U6735 ( .A1(REGFILE_reg_out_26__13_), .A2(net77344), .ZN(n7666) );
  NAND2_X1 U6736 ( .A1(n4893), .A2(REGFILE_reg_out_26__13_), .ZN(n9463) );
  AOI22_X2 U6737 ( .A1(REGFILE_reg_out_26__13_), .A2(net75439), .B1(n5938), 
        .B2(net75440), .ZN(n6639) );
  INV_X1 U6738 ( .A(n4828), .ZN(n5713) );
  NAND2_X4 U6739 ( .A1(n9637), .A2(net76270), .ZN(n9646) );
  OAI211_X4 U6740 ( .C1(n9636), .C2(net76646), .A(net70740), .B(n9635), .ZN(
        n9637) );
  INV_X2 U6741 ( .A(n5715), .ZN(n5716) );
  AOI22_X1 U6742 ( .A1(REGFILE_reg_out_9__1_), .A2(net77698), .B1(
        REGFILE_reg_out_8__1_), .B2(n4829), .ZN(n6886) );
  AOI22_X1 U6743 ( .A1(REGFILE_reg_out_9__3_), .A2(net77698), .B1(
        REGFILE_reg_out_8__3_), .B2(n4829), .ZN(n6842) );
  AOI22_X1 U6744 ( .A1(REGFILE_reg_out_9__0_), .A2(net77698), .B1(
        REGFILE_reg_out_8__0_), .B2(n4829), .ZN(n6909) );
  AOI22_X1 U6745 ( .A1(REGFILE_reg_out_9__2_), .A2(net77698), .B1(
        REGFILE_reg_out_8__2_), .B2(n4829), .ZN(n6864) );
  AOI22_X1 U6746 ( .A1(REGFILE_reg_out_9__26_), .A2(net77702), .B1(
        REGFILE_reg_out_8__26_), .B2(n4829), .ZN(n6356) );
  AOI22_X1 U6747 ( .A1(REGFILE_reg_out_9__29_), .A2(net77702), .B1(
        REGFILE_reg_out_8__29_), .B2(n4829), .ZN(n6285) );
  AOI22_X1 U6748 ( .A1(REGFILE_reg_out_9__25_), .A2(net77702), .B1(
        REGFILE_reg_out_8__25_), .B2(n4829), .ZN(n6380) );
  AOI22_X2 U6749 ( .A1(REGFILE_reg_out_0__24_), .A2(net82342), .B1(
        REGFILE_reg_out_10__24_), .B2(net75464), .ZN(n6392) );
  INV_X2 U6750 ( .A(n8810), .ZN(n8599) );
  NAND2_X1 U6751 ( .A1(net36391), .A2(n10331), .ZN(n10332) );
  NOR3_X1 U6752 ( .A1(n10331), .A2(net72312), .A3(net78003), .ZN(n8644) );
  XNOR2_X1 U6753 ( .A(net36391), .B(n8599), .ZN(n8808) );
  NOR3_X2 U6754 ( .A1(n8646), .A2(n8645), .A3(n8644), .ZN(n8647) );
  INV_X1 U6755 ( .A(n10430), .ZN(n8601) );
  NAND2_X2 U6757 ( .A1(net77422), .A2(REGFILE_reg_out_27__20_), .ZN(n7362) );
  AOI22_X2 U6758 ( .A1(REGFILE_reg_out_31__13_), .A2(net77668), .B1(n5802), 
        .B2(net77676), .ZN(n6634) );
  OAI21_X4 U6759 ( .B1(n6553), .B2(net78056), .A(n6552), .ZN(n5759) );
  INV_X2 U6760 ( .A(n5717), .ZN(n5718) );
  INV_X8 U6761 ( .A(net90830), .ZN(net84754) );
  AOI22_X4 U6762 ( .A1(REGFILE_reg_out_17__17_), .A2(net77796), .B1(
        REGFILE_reg_out_18__17_), .B2(n6896), .ZN(n6554) );
  AOI22_X1 U6763 ( .A1(REGFILE_reg_out_29__31_), .A2(net77650), .B1(
        REGFILE_reg_out_28__31_), .B2(n6911), .ZN(n6243) );
  AOI22_X1 U6764 ( .A1(REGFILE_reg_out_29__0_), .A2(net77650), .B1(
        REGFILE_reg_out_28__0_), .B2(n6911), .ZN(n6915) );
  AOI22_X1 U6765 ( .A1(REGFILE_reg_out_29__30_), .A2(net77650), .B1(
        REGFILE_reg_out_28__30_), .B2(n6911), .ZN(n6268) );
  AOI22_X1 U6766 ( .A1(REGFILE_reg_out_29__28_), .A2(net77650), .B1(
        REGFILE_reg_out_28__28_), .B2(n6911), .ZN(n6314) );
  AOI22_X1 U6767 ( .A1(REGFILE_reg_out_29__26_), .A2(net77650), .B1(
        REGFILE_reg_out_28__26_), .B2(n6911), .ZN(n6361) );
  AOI22_X1 U6768 ( .A1(REGFILE_reg_out_29__27_), .A2(net77650), .B1(
        REGFILE_reg_out_28__27_), .B2(n6911), .ZN(n6338) );
  AOI22_X1 U6769 ( .A1(REGFILE_reg_out_29__3_), .A2(net77650), .B1(
        REGFILE_reg_out_28__3_), .B2(n6911), .ZN(n6847) );
  INV_X2 U6770 ( .A(n5719), .ZN(n5720) );
  NAND2_X1 U6771 ( .A1(REGFILE_reg_out_10__19_), .A2(net77348), .ZN(n7424) );
  AOI22_X2 U6772 ( .A1(REGFILE_reg_out_19__2_), .A2(net77810), .B1(
        REGFILE_reg_out_1__2_), .B2(net82631), .ZN(n6853) );
  AOI22_X2 U6773 ( .A1(REGFILE_reg_out_16__11_), .A2(net75467), .B1(n5909), 
        .B2(net75468), .ZN(n6672) );
  NAND2_X1 U6774 ( .A1(REGFILE_reg_out_18__15_), .A2(net77346), .ZN(n7588) );
  NAND2_X1 U6775 ( .A1(REGFILE_reg_out_22__15_), .A2(net77562), .ZN(n7586) );
  OAI21_X2 U6776 ( .B1(n10403), .B2(n10402), .A(n10401), .ZN(n10406) );
  NAND2_X4 U6777 ( .A1(REGFILE_reg_out_27__29_), .A2(net77426), .ZN(n6986) );
  AOI21_X2 U6778 ( .B1(n10391), .B2(n10390), .A(n10389), .ZN(n10395) );
  OAI21_X1 U6779 ( .B1(n9692), .B2(n9854), .A(n9691), .ZN(n9693) );
  NOR2_X2 U6780 ( .A1(n9694), .A2(n9693), .ZN(n9695) );
  AOI22_X2 U6781 ( .A1(REGFILE_reg_out_4__4_), .A2(net75451), .B1(
        REGFILE_reg_out_5__4_), .B2(net75452), .ZN(n6819) );
  AOI22_X2 U6782 ( .A1(REGFILE_reg_out_16__25_), .A2(net75467), .B1(
        REGFILE_reg_out_15__25_), .B2(net77774), .ZN(n6374) );
  AOI22_X1 U6783 ( .A1(REGFILE_reg_out_11__25_), .A2(net77750), .B1(
        REGFILE_reg_out_12__25_), .B2(net75466), .ZN(n6373) );
  AOI22_X2 U6784 ( .A1(REGFILE_reg_out_11__8_), .A2(net77746), .B1(n5951), 
        .B2(net75466), .ZN(n6737) );
  NAND2_X1 U6785 ( .A1(REGFILE_reg_out_6__13_), .A2(net77560), .ZN(n7694) );
  NAND2_X1 U6786 ( .A1(net77308), .A2(REGFILE_reg_out_8__13_), .ZN(n7685) );
  NAND2_X4 U6787 ( .A1(net77100), .A2(n10607), .ZN(n10209) );
  NAND2_X4 U6788 ( .A1(net77102), .A2(n10614), .ZN(n10213) );
  INV_X16 U6789 ( .A(n10052), .ZN(n6074) );
  NAND4_X1 U6790 ( .A1(n6996), .A2(n4858), .A3(n6997), .A4(n6995), .ZN(n5748)
         );
  OR2_X4 U6791 ( .A1(n10115), .A2(n5571), .ZN(n5749) );
  OAI22_X2 U6792 ( .A1(n10114), .A2(net70691), .B1(n10113), .B2(n10408), .ZN(
        n10115) );
  NAND2_X4 U6793 ( .A1(net77104), .A2(net70574), .ZN(n10215) );
  NAND2_X4 U6794 ( .A1(n10213), .A2(n10212), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X4 U6795 ( .A1(n10209), .A2(n10208), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  INV_X16 U6796 ( .A(n6069), .ZN(n6067) );
  INV_X16 U6797 ( .A(n6069), .ZN(n6068) );
  INV_X1 U6798 ( .A(n9967), .ZN(dmem_addr_out[4]) );
  INV_X32 U6799 ( .A(instruction[15]), .ZN(net92447) );
  INV_X16 U6800 ( .A(net77392), .ZN(net77388) );
  NAND2_X2 U6801 ( .A1(net77478), .A2(REGFILE_reg_out_7__28_), .ZN(n7029) );
  INV_X4 U6802 ( .A(net73585), .ZN(net92392) );
  INV_X8 U6803 ( .A(n6239), .ZN(n5751) );
  OAI21_X1 U6804 ( .B1(dmem_write_out[3]), .B2(net75427), .A(n10945), .ZN(
        n5752) );
  INV_X2 U6805 ( .A(n5755), .ZN(n5756) );
  NAND2_X1 U6806 ( .A1(REGFILE_reg_out_3__16_), .A2(n4871), .ZN(n9256) );
  AOI22_X2 U6807 ( .A1(REGFILE_reg_out_23__5_), .A2(net77826), .B1(
        REGFILE_reg_out_22__5_), .B2(net77834), .ZN(n6788) );
  AOI22_X4 U6808 ( .A1(n5812), .A2(net77452), .B1(n5894), .B2(net77388), .ZN(
        n6926) );
  INV_X8 U6809 ( .A(net91311), .ZN(net75452) );
  BUF_X4 U6810 ( .A(n10392), .Z(n5757) );
  AOI22_X4 U6811 ( .A1(REGFILE_reg_out_31__16_), .A2(net77668), .B1(n5677), 
        .B2(net77676), .ZN(n6572) );
  AOI22_X1 U6812 ( .A1(REGFILE_reg_out_23__4_), .A2(net77826), .B1(
        REGFILE_reg_out_22__4_), .B2(net77834), .ZN(n6810) );
  AOI22_X2 U6813 ( .A1(REGFILE_reg_out_23__0_), .A2(net77826), .B1(
        REGFILE_reg_out_22__0_), .B2(net77834), .ZN(n6899) );
  AOI22_X2 U6814 ( .A1(REGFILE_reg_out_23__6_), .A2(net77826), .B1(
        REGFILE_reg_out_22__6_), .B2(net77834), .ZN(n6766) );
  AOI22_X2 U6815 ( .A1(REGFILE_reg_out_7__6_), .A2(net77714), .B1(
        REGFILE_reg_out_6__6_), .B2(net75456), .ZN(n6777) );
  AOI22_X2 U6816 ( .A1(REGFILE_reg_out_7__21_), .A2(net77714), .B1(
        REGFILE_reg_out_6__21_), .B2(net75456), .ZN(n6471) );
  AOI22_X1 U6817 ( .A1(REGFILE_reg_out_7__1_), .A2(net75455), .B1(
        REGFILE_reg_out_6__1_), .B2(net75456), .ZN(n6887) );
  AOI22_X4 U6818 ( .A1(n5960), .A2(net77406), .B1(n5997), .B2(n6014), .ZN(
        n6947) );
  AOI22_X1 U6819 ( .A1(REGFILE_reg_out_11__2_), .A2(net77746), .B1(
        REGFILE_reg_out_12__2_), .B2(net83168), .ZN(n6857) );
  NAND4_X2 U6820 ( .A1(n6673), .A2(n6671), .A3(n6670), .A4(n6672), .ZN(n6674)
         );
  AOI22_X2 U6821 ( .A1(REGFILE_reg_out_4__20_), .A2(n5679), .B1(
        REGFILE_reg_out_5__20_), .B2(net84475), .ZN(n6493) );
  AOI22_X2 U6822 ( .A1(REGFILE_reg_out_4__8_), .A2(net75451), .B1(n5687), .B2(
        net84475), .ZN(n6743) );
  AOI22_X4 U6823 ( .A1(REGFILE_reg_out_29__9_), .A2(net77650), .B1(
        REGFILE_reg_out_28__9_), .B2(n5751), .ZN(n6727) );
  NAND2_X4 U6824 ( .A1(instruction[11]), .A2(instruction[12]), .ZN(net87489)
         );
  INV_X8 U6825 ( .A(aluA[27]), .ZN(n5760) );
  INV_X16 U6826 ( .A(n5760), .ZN(n5761) );
  OAI21_X4 U6827 ( .B1(n6974), .B2(n6975), .A(n6019), .ZN(n6996) );
  INV_X16 U6828 ( .A(net74051), .ZN(net77548) );
  INV_X16 U6829 ( .A(net77542), .ZN(net77516) );
  INV_X32 U6830 ( .A(instruction[8]), .ZN(net90864) );
  AOI22_X4 U6831 ( .A1(REGFILE_reg_out_4__17_), .A2(net75451), .B1(
        REGFILE_reg_out_5__17_), .B2(net75452), .ZN(n6559) );
  AOI22_X4 U6832 ( .A1(n5796), .A2(net77406), .B1(n5972), .B2(n6014), .ZN(
        n6935) );
  NOR2_X2 U6835 ( .A1(n6260), .A2(n6259), .ZN(n6272) );
  INV_X2 U6836 ( .A(n5765), .ZN(n5766) );
  AOI22_X2 U6837 ( .A1(REGFILE_reg_out_24__16_), .A2(net75437), .B1(n5613), 
        .B2(net124970), .ZN(n6576) );
  INV_X1 U6838 ( .A(n10420), .ZN(n9836) );
  NAND4_X2 U6839 ( .A1(n6591), .A2(n6589), .A3(n6588), .A4(n6590), .ZN(n6592)
         );
  AOI22_X2 U6840 ( .A1(REGFILE_reg_out_19__14_), .A2(net77812), .B1(
        REGFILE_reg_out_1__14_), .B2(net75478), .ZN(n6609) );
  AOI22_X2 U6841 ( .A1(REGFILE_reg_out_19__11_), .A2(net77812), .B1(
        REGFILE_reg_out_1__11_), .B2(net75478), .ZN(n6667) );
  INV_X2 U6842 ( .A(n5767), .ZN(n5768) );
  NAND2_X1 U6843 ( .A1(REGFILE_reg_out_1__13_), .A2(net77524), .ZN(n7693) );
  NAND2_X1 U6844 ( .A1(n4877), .A2(REGFILE_reg_out_1__13_), .ZN(n9449) );
  OAI21_X2 U6845 ( .B1(n9100), .B2(n9854), .A(n9099), .ZN(n9101) );
  INV_X2 U6846 ( .A(n5847), .ZN(n5769) );
  NOR2_X2 U6847 ( .A1(n10447), .A2(net78014), .ZN(n9181) );
  INV_X2 U6848 ( .A(n9054), .ZN(n9055) );
  XNOR2_X1 U6849 ( .A(n9054), .B(aluA[16]), .ZN(n9178) );
  OAI21_X2 U6850 ( .B1(n9196), .B2(n9854), .A(n9195), .ZN(n9197) );
  XNOR2_X1 U6851 ( .A(n10930), .B(n8989), .ZN(n10435) );
  XNOR2_X1 U6852 ( .A(n10930), .B(n4808), .ZN(n8988) );
  NOR3_X2 U6853 ( .A1(n10437), .A2(n10436), .A3(n10435), .ZN(n10438) );
  NAND2_X1 U6854 ( .A1(net70701), .A2(n10435), .ZN(n8991) );
  AOI21_X2 U6855 ( .B1(net71271), .B2(n8993), .A(n8992), .ZN(n8995) );
  NAND2_X1 U6856 ( .A1(n8816), .A2(aluA[20]), .ZN(n8817) );
  NOR3_X2 U6857 ( .A1(n10451), .A2(n10450), .A3(n10449), .ZN(n10452) );
  AOI21_X2 U6858 ( .B1(net71271), .B2(n10056), .A(n10055), .ZN(n10077) );
  NOR3_X2 U6859 ( .A1(n10074), .A2(n10073), .A3(n10072), .ZN(n10075) );
  AOI22_X2 U6860 ( .A1(REGFILE_reg_out_26__30_), .A2(net77620), .B1(
        REGFILE_reg_out_27__30_), .B2(net77630), .ZN(n6266) );
  INV_X8 U6861 ( .A(net76199), .ZN(net89184) );
  INV_X1 U6862 ( .A(n10922), .ZN(n9306) );
  AOI22_X4 U6863 ( .A1(REGFILE_reg_out_21__13_), .A2(net77844), .B1(n5720), 
        .B2(net77852), .ZN(n6633) );
  NAND2_X4 U6864 ( .A1(instruction[5]), .A2(net73170), .ZN(net73532) );
  NAND2_X1 U6865 ( .A1(n4966), .A2(net73170), .ZN(net73780) );
  INV_X32 U6866 ( .A(instruction[3]), .ZN(net73170) );
  INV_X4 U6867 ( .A(n8410), .ZN(n5815) );
  INV_X8 U6868 ( .A(n10036), .ZN(n10908) );
  AOI22_X2 U6869 ( .A1(REGFILE_reg_out_11__3_), .A2(net77746), .B1(
        REGFILE_reg_out_12__3_), .B2(net83167), .ZN(n6835) );
  AOI22_X1 U6870 ( .A1(REGFILE_reg_out_30__25_), .A2(net77638), .B1(
        REGFILE_reg_out_2__25_), .B2(net75442), .ZN(n6384) );
  NAND2_X1 U6871 ( .A1(REGFILE_reg_out_0__14_), .A2(net77310), .ZN(n7651) );
  NAND2_X1 U6872 ( .A1(REGFILE_reg_out_12__16_), .A2(n4873), .ZN(n9212) );
  INV_X2 U6873 ( .A(n5771), .ZN(n5772) );
  AOI22_X2 U6874 ( .A1(REGFILE_reg_out_26__15_), .A2(net75439), .B1(n4839), 
        .B2(net75440), .ZN(n6599) );
  NAND4_X2 U6875 ( .A1(n6945), .A2(n6942), .A3(n6944), .A4(n6943), .ZN(n8410)
         );
  AOI22_X1 U6876 ( .A1(REGFILE_reg_out_23__31_), .A2(net77828), .B1(
        REGFILE_reg_out_22__31_), .B2(net77836), .ZN(n6227) );
  AOI22_X2 U6877 ( .A1(n5825), .A2(net77406), .B1(n5828), .B2(n6014), .ZN(
        n6925) );
  INV_X32 U6878 ( .A(instruction[14]), .ZN(net86794) );
  NOR2_X4 U6879 ( .A1(n6763), .A2(n6762), .ZN(net75615) );
  NAND2_X4 U6880 ( .A1(REGFILE_reg_out_25__29_), .A2(net77514), .ZN(n6984) );
  INV_X2 U6881 ( .A(n5776), .ZN(n5777) );
  INV_X2 U6882 ( .A(n5778), .ZN(n5779) );
  INV_X2 U6883 ( .A(n5780), .ZN(n5781) );
  NAND4_X2 U6884 ( .A1(n6547), .A2(n6546), .A3(n6544), .A4(n6545), .ZN(n6548)
         );
  NOR2_X4 U6885 ( .A1(n6580), .A2(n6581), .ZN(n6582) );
  OAI22_X1 U6886 ( .A1(n9961), .A2(net70691), .B1(n9960), .B2(n5659), .ZN(
        n9962) );
  XNOR2_X1 U6887 ( .A(n5659), .B(net77040), .ZN(n10033) );
  NAND2_X1 U6888 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_4__MUX_N1), .A2(n5659), .ZN(
        n10401) );
  XNOR2_X1 U6889 ( .A(n5659), .B(n9954), .ZN(n10306) );
  INV_X8 U6890 ( .A(net76203), .ZN(net75442) );
  AOI22_X2 U6891 ( .A1(REGFILE_reg_out_26__2_), .A2(net77620), .B1(
        REGFILE_reg_out_27__2_), .B2(net77630), .ZN(n6867) );
  AOI22_X2 U6892 ( .A1(REGFILE_reg_out_17__19_), .A2(net77796), .B1(
        REGFILE_reg_out_18__19_), .B2(n6896), .ZN(n6506) );
  NAND2_X1 U6893 ( .A1(net77298), .A2(REGFILE_reg_out_16__27_), .ZN(n7056) );
  AOI22_X2 U6894 ( .A1(n5793), .A2(net77514), .B1(n5892), .B2(net77298), .ZN(
        n6928) );
  NOR2_X4 U6896 ( .A1(n6729), .A2(n6728), .ZN(n6730) );
  AOI22_X2 U6897 ( .A1(REGFILE_reg_out_16__21_), .A2(net87506), .B1(
        REGFILE_reg_out_15__21_), .B2(n5579), .ZN(n6464) );
  AOI22_X1 U6898 ( .A1(REGFILE_reg_out_16__28_), .A2(net87506), .B1(
        REGFILE_reg_out_15__28_), .B2(n5579), .ZN(n6303) );
  AOI22_X2 U6899 ( .A1(REGFILE_reg_out_0__16_), .A2(net82342), .B1(n5772), 
        .B2(net83203), .ZN(n6566) );
  NAND2_X2 U6900 ( .A1(n6431), .A2(n6430), .ZN(dmem_write_out[23]) );
  AOI22_X2 U6901 ( .A1(REGFILE_reg_out_26__3_), .A2(net77620), .B1(
        REGFILE_reg_out_27__3_), .B2(net77630), .ZN(n6845) );
  INV_X2 U6902 ( .A(n5866), .ZN(n5782) );
  OAI21_X1 U6903 ( .B1(n6481), .B2(net78056), .A(n6480), .ZN(n5783) );
  NAND2_X1 U6904 ( .A1(REGFILE_reg_out_18__13_), .A2(net77344), .ZN(n7676) );
  NAND2_X1 U6905 ( .A1(REGFILE_reg_out_10__22_), .A2(n6015), .ZN(n7286) );
  INV_X1 U6906 ( .A(n10923), .ZN(n10331) );
  INV_X4 U6907 ( .A(net77624), .ZN(net77618) );
  INV_X8 U6908 ( .A(n5931), .ZN(n5870) );
  OAI21_X2 U6909 ( .B1(n7538), .B2(n7537), .A(n6012), .ZN(n7572) );
  INV_X2 U6910 ( .A(n5786), .ZN(n5787) );
  OAI22_X2 U6911 ( .A1(n5948), .A2(net77506), .B1(n5949), .B2(net75424), .ZN(
        n5947) );
  NAND2_X4 U6912 ( .A1(n5916), .A2(n6929), .ZN(n8403) );
  INV_X4 U6913 ( .A(net77608), .ZN(net77602) );
  AOI22_X2 U6914 ( .A1(REGFILE_reg_out_26__21_), .A2(net75439), .B1(
        REGFILE_reg_out_27__21_), .B2(net89184), .ZN(n6473) );
  INV_X2 U6915 ( .A(n5788), .ZN(n5789) );
  INV_X2 U6916 ( .A(n5790), .ZN(n5791) );
  NOR2_X1 U6917 ( .A1(net73850), .A2(net73836), .ZN(n8406) );
  INV_X2 U6918 ( .A(n5792), .ZN(n5793) );
  INV_X1 U6919 ( .A(n5672), .ZN(n10936) );
  INV_X2 U6920 ( .A(n5794), .ZN(n5795) );
  OAI21_X2 U6921 ( .B1(n6223), .B2(net76480), .A(n8755), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  INV_X4 U6922 ( .A(n5898), .ZN(n5796) );
  AND2_X2 U6923 ( .A1(n5899), .A2(n5900), .ZN(n5797) );
  NAND2_X2 U6924 ( .A1(instruction[29]), .A2(net77276), .ZN(n5900) );
  AOI22_X2 U6925 ( .A1(REGFILE_reg_out_17__11_), .A2(net77796), .B1(
        REGFILE_reg_out_18__11_), .B2(n6896), .ZN(n6666) );
  AOI22_X1 U6926 ( .A1(REGFILE_reg_out_7__25_), .A2(net77714), .B1(
        REGFILE_reg_out_6__25_), .B2(net75456), .ZN(n6381) );
  NOR2_X2 U6927 ( .A1(n6467), .A2(n6466), .ZN(n6479) );
  AOI22_X2 U6928 ( .A1(REGFILE_reg_out_0__22_), .A2(net82342), .B1(
        REGFILE_reg_out_10__22_), .B2(net83203), .ZN(n6438) );
  AOI22_X2 U6929 ( .A1(REGFILE_reg_out_30__21_), .A2(net84761), .B1(
        REGFILE_reg_out_2__21_), .B2(net75442), .ZN(n6474) );
  INV_X2 U6930 ( .A(REGFILE_reg_out_15__31_), .ZN(n10522) );
  NAND4_X2 U6931 ( .A1(n6641), .A2(n6640), .A3(n6638), .A4(n6639), .ZN(n6642)
         );
  AOI22_X2 U6932 ( .A1(REGFILE_reg_out_23__11_), .A2(net77828), .B1(
        REGFILE_reg_out_22__11_), .B2(net77836), .ZN(n6668) );
  AOI22_X1 U6933 ( .A1(REGFILE_reg_out_0__27_), .A2(net82342), .B1(
        REGFILE_reg_out_10__27_), .B2(net75464), .ZN(n6325) );
  AOI22_X2 U6934 ( .A1(REGFILE_reg_out_19__12_), .A2(net77812), .B1(
        REGFILE_reg_out_1__12_), .B2(net75478), .ZN(n6645) );
  BUF_X32 U6935 ( .A(aluA[30]), .Z(n5798) );
  INV_X32 U6936 ( .A(instruction[9]), .ZN(net87098) );
  OAI22_X2 U6937 ( .A1(n6002), .A2(net77440), .B1(n6003), .B2(net85371), .ZN(
        n6001) );
  NAND4_X2 U6938 ( .A1(n6451), .A2(n6450), .A3(n6449), .A4(n6448), .ZN(n6452)
         );
  INV_X8 U6939 ( .A(net75425), .ZN(net86304) );
  INV_X4 U6940 ( .A(n5947), .ZN(n6931) );
  INV_X1 U6941 ( .A(REGFILE_reg_out_20__31_), .ZN(n10525) );
  AOI22_X1 U6942 ( .A1(REGFILE_reg_out_21__31_), .A2(net77846), .B1(
        REGFILE_reg_out_20__31_), .B2(net77854), .ZN(n6228) );
  INV_X2 U6943 ( .A(n5799), .ZN(n5800) );
  INV_X2 U6944 ( .A(n5801), .ZN(n5802) );
  INV_X2 U6945 ( .A(n5803), .ZN(n5804) );
  AOI22_X2 U6946 ( .A1(REGFILE_reg_out_0__13_), .A2(net82342), .B1(n5814), 
        .B2(net75464), .ZN(net75764) );
  NOR2_X2 U6948 ( .A1(n6477), .A2(n6476), .ZN(n6478) );
  NOR2_X1 U6949 ( .A1(n4856), .A2(n10334), .ZN(n10335) );
  AOI22_X1 U6950 ( .A1(REGFILE_reg_out_11__27_), .A2(net77750), .B1(
        REGFILE_reg_out_12__27_), .B2(net75466), .ZN(n6326) );
  INV_X4 U6951 ( .A(dmem_write_out[23]), .ZN(n6433) );
  INV_X2 U6952 ( .A(n10323), .ZN(n5806) );
  NAND2_X1 U6953 ( .A1(REGFILE_reg_out_25__21_), .A2(net77530), .ZN(n7316) );
  AOI22_X2 U6954 ( .A1(REGFILE_reg_out_24__21_), .A2(net75437), .B1(
        REGFILE_reg_out_25__21_), .B2(net75438), .ZN(n6472) );
  INV_X2 U6955 ( .A(REGFILE_reg_out_18__31_), .ZN(n10524) );
  INV_X2 U6956 ( .A(n5808), .ZN(n5809) );
  INV_X2 U6957 ( .A(n5811), .ZN(n5812) );
  INV_X2 U6958 ( .A(n5813), .ZN(n5814) );
  AOI22_X2 U6959 ( .A1(REGFILE_reg_out_30__11_), .A2(net84761), .B1(n5874), 
        .B2(net82613), .ZN(n6682) );
  INV_X2 U6960 ( .A(n5816), .ZN(n5817) );
  INV_X4 U6961 ( .A(n5924), .ZN(n5818) );
  NOR2_X2 U6963 ( .A1(n6443), .A2(n6442), .ZN(n6455) );
  INV_X8 U6964 ( .A(net77632), .ZN(net77626) );
  NAND2_X1 U6965 ( .A1(REGFILE_reg_out_27__19_), .A2(net77422), .ZN(n7406) );
  OAI21_X2 U6966 ( .B1(n10388), .B2(n10387), .A(n10386), .ZN(n10390) );
  AND2_X2 U6967 ( .A1(n5916), .A2(n6929), .ZN(n5820) );
  INV_X8 U6968 ( .A(n5822), .ZN(n6929) );
  AOI22_X2 U6969 ( .A1(REGFILE_reg_out_21__8_), .A2(net77842), .B1(
        REGFILE_reg_out_20__8_), .B2(net77850), .ZN(n6735) );
  NOR2_X4 U6970 ( .A1(n6719), .A2(n6718), .ZN(n6731) );
  NAND2_X1 U6971 ( .A1(net77346), .A2(REGFILE_reg_out_2__14_), .ZN(n7652) );
  INV_X1 U6972 ( .A(REGFILE_reg_out_13__31_), .ZN(n10518) );
  INV_X2 U6973 ( .A(n5824), .ZN(n5825) );
  INV_X1 U6974 ( .A(REGFILE_reg_out_9__31_), .ZN(n10537) );
  AOI22_X1 U6975 ( .A1(REGFILE_reg_out_9__31_), .A2(net77702), .B1(
        REGFILE_reg_out_8__31_), .B2(n4829), .ZN(n6237) );
  INV_X4 U6976 ( .A(n6946), .ZN(n6932) );
  AOI22_X2 U6977 ( .A1(REGFILE_reg_out_24__12_), .A2(net75437), .B1(n5865), 
        .B2(net124970), .ZN(n6658) );
  AOI22_X2 U6978 ( .A1(REGFILE_reg_out_24__11_), .A2(net75437), .B1(n5882), 
        .B2(net124970), .ZN(n6680) );
  INV_X1 U6979 ( .A(n10913), .ZN(n5826) );
  NAND2_X1 U6980 ( .A1(REGFILE_reg_out_3__8_), .A2(net77414), .ZN(n7918) );
  NAND2_X2 U6981 ( .A1(REGFILE_reg_out_25__20_), .A2(net77530), .ZN(n7357) );
  NAND4_X2 U6982 ( .A1(n6495), .A2(n6494), .A3(n6493), .A4(n6492), .ZN(n6501)
         );
  AOI22_X2 U6983 ( .A1(REGFILE_reg_out_7__19_), .A2(net77714), .B1(
        REGFILE_reg_out_6__19_), .B2(net75456), .ZN(n6519) );
  NOR3_X1 U6985 ( .A1(n10352), .A2(n8849), .A3(net78003), .ZN(n8865) );
  AOI22_X1 U6986 ( .A1(REGFILE_reg_out_7__30_), .A2(net77714), .B1(
        REGFILE_reg_out_6__30_), .B2(net75456), .ZN(n6264) );
  AOI22_X1 U6987 ( .A1(REGFILE_reg_out_7__28_), .A2(net77716), .B1(
        REGFILE_reg_out_6__28_), .B2(net75456), .ZN(n6310) );
  AOI22_X1 U6988 ( .A1(REGFILE_reg_out_7__27_), .A2(net77716), .B1(
        REGFILE_reg_out_6__27_), .B2(net75456), .ZN(n6334) );
  AOI22_X2 U6989 ( .A1(REGFILE_reg_out_26__20_), .A2(net75439), .B1(
        REGFILE_reg_out_27__20_), .B2(net89184), .ZN(n6497) );
  AOI22_X1 U6990 ( .A1(REGFILE_reg_out_24__30_), .A2(net77602), .B1(
        REGFILE_reg_out_25__30_), .B2(net77610), .ZN(n6265) );
  NAND2_X1 U6991 ( .A1(REGFILE_reg_out_27__21_), .A2(net77422), .ZN(n7313) );
  AOI22_X2 U6992 ( .A1(REGFILE_reg_out_17__12_), .A2(net77796), .B1(
        REGFILE_reg_out_18__12_), .B2(n6896), .ZN(n6644) );
  NOR2_X2 U6993 ( .A1(n6377), .A2(n6376), .ZN(n6389) );
  NAND2_X4 U6994 ( .A1(n5990), .A2(net77462), .ZN(n6988) );
  XNOR2_X1 U6995 ( .A(n5806), .B(aluA[26]), .ZN(n10444) );
  INV_X1 U6996 ( .A(n10925), .ZN(n10323) );
  XNOR2_X1 U6997 ( .A(n5806), .B(net77040), .ZN(n8596) );
  AOI22_X1 U6998 ( .A1(REGFILE_reg_out_0__5_), .A2(net82342), .B1(
        REGFILE_reg_out_10__5_), .B2(net75464), .ZN(n6790) );
  AOI22_X2 U6999 ( .A1(REGFILE_reg_out_26__25_), .A2(net77620), .B1(
        REGFILE_reg_out_27__25_), .B2(net77626), .ZN(n6383) );
  NAND4_X2 U7000 ( .A1(n6499), .A2(n6497), .A3(n6498), .A4(n6496), .ZN(n6500)
         );
  NAND2_X1 U7001 ( .A1(REGFILE_reg_out_8__14_), .A2(net77310), .ZN(n7641) );
  NAND2_X1 U7002 ( .A1(n5781), .A2(net77382), .ZN(n7633) );
  NAND2_X1 U7003 ( .A1(REGFILE_reg_out_28__14_), .A2(n6175), .ZN(n10271) );
  NAND2_X1 U7004 ( .A1(REGFILE_reg_out_28__14_), .A2(net77382), .ZN(n7623) );
  OAI21_X4 U7005 ( .B1(n6296), .B2(net73697), .A(n6295), .ZN(n10927) );
  INV_X16 U7006 ( .A(n10927), .ZN(n6004) );
  NAND2_X1 U7007 ( .A1(net76488), .A2(REGFILE_reg_out_31__30_), .ZN(n8755) );
  AOI22_X1 U7008 ( .A1(REGFILE_reg_out_31__30_), .A2(net77670), .B1(
        REGFILE_reg_out_3__30_), .B2(n5609), .ZN(n6261) );
  NAND2_X1 U7009 ( .A1(REGFILE_reg_out_1__15_), .A2(net77526), .ZN(n7605) );
  AOI22_X2 U7010 ( .A1(REGFILE_reg_out_0__7_), .A2(net82342), .B1(
        REGFILE_reg_out_10__7_), .B2(net75464), .ZN(n6758) );
  INV_X2 U7011 ( .A(n5827), .ZN(n5828) );
  INV_X8 U7012 ( .A(net77506), .ZN(net77480) );
  INV_X4 U7013 ( .A(n5844), .ZN(n5829) );
  NAND4_X2 U7014 ( .A1(n6637), .A2(n6636), .A3(n6635), .A4(n6634), .ZN(n6643)
         );
  NAND2_X1 U7015 ( .A1(n10926), .A2(n5652), .ZN(n9094) );
  NAND2_X1 U7016 ( .A1(n5652), .A2(n10315), .ZN(n9581) );
  XNOR2_X1 U7017 ( .A(n5761), .B(n5652), .ZN(n10436) );
  XNOR2_X1 U7018 ( .A(net77040), .B(n5652), .ZN(n8594) );
  INV_X4 U7019 ( .A(n5918), .ZN(n5830) );
  NAND2_X1 U7020 ( .A1(REGFILE_reg_out_3__14_), .A2(net77418), .ZN(n7654) );
  INV_X4 U7021 ( .A(n5831), .ZN(n5832) );
  INV_X2 U7022 ( .A(n5833), .ZN(n5834) );
  AOI22_X2 U7023 ( .A1(REGFILE_reg_out_26__4_), .A2(net77620), .B1(
        REGFILE_reg_out_27__4_), .B2(net77626), .ZN(n6823) );
  NAND2_X1 U7024 ( .A1(n4890), .A2(REGFILE_reg_out_8__13_), .ZN(n9487) );
  INV_X2 U7025 ( .A(n5835), .ZN(n5836) );
  AOI22_X2 U7026 ( .A1(REGFILE_reg_out_0__11_), .A2(net82342), .B1(
        REGFILE_reg_out_10__11_), .B2(net75464), .ZN(n6670) );
  AOI22_X2 U7027 ( .A1(REGFILE_reg_out_0__19_), .A2(net82342), .B1(
        REGFILE_reg_out_10__19_), .B2(net83203), .ZN(n6510) );
  INV_X16 U7028 ( .A(net77500), .ZN(net77496) );
  INV_X16 U7029 ( .A(net77500), .ZN(net77494) );
  AOI22_X4 U7030 ( .A1(REGFILE_reg_out_23__13_), .A2(net77828), .B1(n5800), 
        .B2(net77836), .ZN(n6632) );
  NAND3_X1 U7031 ( .A1(n10929), .A2(n5761), .A3(net71078), .ZN(n8886) );
  NAND2_X1 U7032 ( .A1(n10929), .A2(net70696), .ZN(n9093) );
  NAND2_X1 U7033 ( .A1(n10929), .A2(n10926), .ZN(net70866) );
  NAND2_X1 U7034 ( .A1(n10929), .A2(n10315), .ZN(net70868) );
  NOR2_X1 U7035 ( .A1(n10929), .A2(n10319), .ZN(n10320) );
  NAND2_X1 U7036 ( .A1(net73708), .A2(aluA[26]), .ZN(n8683) );
  NAND3_X1 U7037 ( .A1(net71078), .A2(aluA[26]), .A3(n5806), .ZN(n9780) );
  NOR2_X1 U7038 ( .A1(n8449), .A2(n8448), .ZN(n8453) );
  NAND2_X1 U7039 ( .A1(n8937), .A2(aluA[26]), .ZN(n8938) );
  NAND2_X1 U7040 ( .A1(n9065), .A2(aluA[26]), .ZN(n8843) );
  NAND2_X1 U7041 ( .A1(net70720), .A2(aluA[26]), .ZN(n9359) );
  NAND2_X1 U7042 ( .A1(net70719), .A2(aluA[26]), .ZN(n10097) );
  NAND2_X1 U7043 ( .A1(n6040), .A2(aluA[26]), .ZN(n8714) );
  INV_X2 U7044 ( .A(aluA[26]), .ZN(n8597) );
  XNOR2_X1 U7045 ( .A(n8596), .B(aluA[26]), .ZN(n9777) );
  NAND2_X1 U7046 ( .A1(REGFILE_reg_out_28__13_), .A2(n6177), .ZN(n9467) );
  NAND2_X1 U7047 ( .A1(REGFILE_reg_out_28__13_), .A2(net77380), .ZN(n7667) );
  NAND2_X1 U7048 ( .A1(REGFILE_reg_out_2__20_), .A2(n6015), .ZN(n7390) );
  AOI22_X4 U7049 ( .A1(REGFILE_reg_out_29__14_), .A2(net77652), .B1(n4832), 
        .B2(n6911), .ZN(n6625) );
  INV_X2 U7050 ( .A(n5839), .ZN(n5840) );
  AOI22_X4 U7051 ( .A1(REGFILE_reg_out_23__14_), .A2(net77828), .B1(
        REGFILE_reg_out_22__14_), .B2(net77836), .ZN(n6610) );
  AOI22_X2 U7052 ( .A1(REGFILE_reg_out_30__24_), .A2(net77638), .B1(
        REGFILE_reg_out_2__24_), .B2(net75442), .ZN(n6403) );
  AOI22_X2 U7053 ( .A1(REGFILE_reg_out_30__19_), .A2(net84761), .B1(
        REGFILE_reg_out_2__19_), .B2(net75442), .ZN(n6522) );
  XNOR2_X1 U7054 ( .A(n10923), .B(net77038), .ZN(n8810) );
  XNOR2_X1 U7055 ( .A(n10408), .B(net77040), .ZN(n10165) );
  NAND2_X1 U7056 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_2__MUX_N1), .A2(n10408), .ZN(
        n10409) );
  XNOR2_X1 U7057 ( .A(n10408), .B(n10109), .ZN(n10104) );
  AOI22_X4 U7058 ( .A1(REGFILE_reg_out_17__14_), .A2(net77796), .B1(n10953), 
        .B2(n5890), .ZN(n6608) );
  XNOR2_X1 U7059 ( .A(n5752), .B(net77040), .ZN(n10110) );
  XNOR2_X1 U7060 ( .A(n5752), .B(n10404), .ZN(n10407) );
  INV_X8 U7061 ( .A(net76205), .ZN(net75441) );
  NAND4_X2 U7062 ( .A1(n6661), .A2(n6659), .A3(n6660), .A4(n6658), .ZN(n6662)
         );
  INV_X8 U7063 ( .A(net76248), .ZN(net76202) );
  INV_X1 U7064 ( .A(n10917), .ZN(n5847) );
  NAND2_X1 U7065 ( .A1(net77550), .A2(REGFILE_reg_out_22__27_), .ZN(n7055) );
  NAND2_X1 U7066 ( .A1(net77348), .A2(REGFILE_reg_out_2__17_), .ZN(n7520) );
  NAND2_X1 U7067 ( .A1(REGFILE_reg_out_25__17_), .A2(net77528), .ZN(n7489) );
  AOI22_X1 U7068 ( .A1(REGFILE_reg_out_11__0_), .A2(net77746), .B1(
        REGFILE_reg_out_12__0_), .B2(net75466), .ZN(n6902) );
  AOI22_X2 U7069 ( .A1(REGFILE_reg_out_26__27_), .A2(net77620), .B1(
        REGFILE_reg_out_27__27_), .B2(net77630), .ZN(n6336) );
  AOI22_X2 U7070 ( .A1(REGFILE_reg_out_17__21_), .A2(net77796), .B1(
        REGFILE_reg_out_18__21_), .B2(n6896), .ZN(n6458) );
  AOI22_X2 U7071 ( .A1(REGFILE_reg_out_4__9_), .A2(n5678), .B1(
        REGFILE_reg_out_5__9_), .B2(net84475), .ZN(n6721) );
  NOR2_X2 U7072 ( .A1(n6387), .A2(n6386), .ZN(n6388) );
  NAND2_X1 U7073 ( .A1(net73878), .A2(net88253), .ZN(n8306) );
  AOI22_X2 U7074 ( .A1(REGFILE_reg_out_17__20_), .A2(net77796), .B1(
        REGFILE_reg_out_18__20_), .B2(n6896), .ZN(n6482) );
  AOI22_X2 U7075 ( .A1(REGFILE_reg_out_30__18_), .A2(net84761), .B1(
        REGFILE_reg_out_2__18_), .B2(net82613), .ZN(n6546) );
  AOI22_X1 U7076 ( .A1(REGFILE_reg_out_7__31_), .A2(net77716), .B1(
        REGFILE_reg_out_6__31_), .B2(net75456), .ZN(n6238) );
  AOI22_X1 U7077 ( .A1(REGFILE_reg_out_7__29_), .A2(net77714), .B1(
        REGFILE_reg_out_6__29_), .B2(net75456), .ZN(n6286) );
  AOI22_X1 U7078 ( .A1(REGFILE_reg_out_7__26_), .A2(net77714), .B1(
        REGFILE_reg_out_6__26_), .B2(net75456), .ZN(n6357) );
  AOI22_X1 U7079 ( .A1(REGFILE_reg_out_7__23_), .A2(net77714), .B1(
        REGFILE_reg_out_6__23_), .B2(net75456), .ZN(n6424) );
  INV_X8 U7080 ( .A(net76234), .ZN(net75466) );
  INV_X2 U7081 ( .A(n10352), .ZN(n5848) );
  NAND4_X2 U7082 ( .A1(n6441), .A2(n6440), .A3(n6439), .A4(n6438), .ZN(n6442)
         );
  AOI22_X4 U7083 ( .A1(REGFILE_reg_out_14__14_), .A2(net77780), .B1(n4853), 
        .B2(n5664), .ZN(n6615) );
  AOI22_X2 U7084 ( .A1(REGFILE_reg_out_26__5_), .A2(net77620), .B1(
        REGFILE_reg_out_27__5_), .B2(net77626), .ZN(n6801) );
  AOI22_X1 U7085 ( .A1(REGFILE_reg_out_4__5_), .A2(net75451), .B1(
        REGFILE_reg_out_5__5_), .B2(net75452), .ZN(n6797) );
  NAND2_X1 U7086 ( .A1(net77344), .A2(REGFILE_reg_out_2__13_), .ZN(n7696) );
  INV_X2 U7087 ( .A(n5849), .ZN(n5850) );
  INV_X16 U7088 ( .A(net75475), .ZN(net77800) );
  AOI22_X1 U7089 ( .A1(REGFILE_reg_out_11__1_), .A2(net77746), .B1(
        REGFILE_reg_out_12__1_), .B2(net75466), .ZN(n6879) );
  AOI22_X2 U7090 ( .A1(REGFILE_reg_out_11__7_), .A2(net77746), .B1(
        REGFILE_reg_out_12__7_), .B2(net75466), .ZN(n6759) );
  AOI22_X2 U7091 ( .A1(REGFILE_reg_out_11__20_), .A2(net77748), .B1(
        REGFILE_reg_out_12__20_), .B2(net83168), .ZN(n6487) );
  INV_X8 U7092 ( .A(net75441), .ZN(net77640) );
  INV_X2 U7093 ( .A(n5852), .ZN(n5853) );
  INV_X2 U7094 ( .A(n5854), .ZN(n5855) );
  AOI22_X4 U7095 ( .A1(REGFILE_reg_out_29__15_), .A2(net77652), .B1(n10951), 
        .B2(n6911), .ZN(n6601) );
  AOI22_X2 U7096 ( .A1(REGFILE_reg_out_30__10_), .A2(net77634), .B1(
        REGFILE_reg_out_2__10_), .B2(net82613), .ZN(n6704) );
  AOI22_X4 U7097 ( .A1(REGFILE_reg_out_29__13_), .A2(net77652), .B1(n5768), 
        .B2(n5751), .ZN(n6641) );
  NAND2_X1 U7098 ( .A1(REGFILE_reg_out_27__8_), .A2(net77414), .ZN(n7888) );
  INV_X1 U7099 ( .A(REGFILE_reg_out_27__14_), .ZN(n10270) );
  AOI22_X1 U7100 ( .A1(REGFILE_reg_out_26__31_), .A2(net77620), .B1(
        REGFILE_reg_out_27__31_), .B2(net89184), .ZN(n6241) );
  AOI22_X2 U7101 ( .A1(REGFILE_reg_out_0__21_), .A2(net120684), .B1(n5809), 
        .B2(net75464), .ZN(n6462) );
  AOI22_X2 U7102 ( .A1(REGFILE_reg_out_11__21_), .A2(net77748), .B1(
        REGFILE_reg_out_12__21_), .B2(net83168), .ZN(n6463) );
  INV_X1 U7103 ( .A(REGFILE_reg_out_16__31_), .ZN(n10523) );
  AOI22_X1 U7104 ( .A1(REGFILE_reg_out_16__31_), .A2(net75467), .B1(
        REGFILE_reg_out_15__31_), .B2(net77774), .ZN(n6231) );
  NAND2_X1 U7105 ( .A1(REGFILE_reg_out_2__18_), .A2(net77348), .ZN(n7478) );
  AOI22_X1 U7106 ( .A1(REGFILE_reg_out_30__23_), .A2(net77638), .B1(
        REGFILE_reg_out_2__23_), .B2(net75442), .ZN(n6426) );
  INV_X2 U7107 ( .A(n5858), .ZN(n5859) );
  INV_X2 U7108 ( .A(n5860), .ZN(n5861) );
  INV_X2 U7109 ( .A(n5862), .ZN(n5863) );
  INV_X2 U7110 ( .A(n5864), .ZN(n5865) );
  INV_X2 U7111 ( .A(REGFILE_reg_out_10__15_), .ZN(n10298) );
  INV_X2 U7112 ( .A(n9057), .ZN(n9058) );
  INV_X1 U7113 ( .A(n10424), .ZN(n10281) );
  AOI22_X1 U7114 ( .A1(REGFILE_reg_out_17__27_), .A2(net77798), .B1(
        REGFILE_reg_out_18__27_), .B2(n5890), .ZN(n6321) );
  AOI22_X1 U7115 ( .A1(REGFILE_reg_out_17__23_), .A2(net77798), .B1(
        REGFILE_reg_out_18__23_), .B2(n5890), .ZN(n6411) );
  AOI22_X2 U7116 ( .A1(REGFILE_reg_out_16__7_), .A2(net77762), .B1(
        REGFILE_reg_out_15__7_), .B2(net75468), .ZN(n6760) );
  INV_X32 U7117 ( .A(net77500), .ZN(net77498) );
  INV_X16 U7118 ( .A(net77856), .ZN(net77850) );
  INV_X1 U7119 ( .A(n10915), .ZN(n5867) );
  INV_X8 U7120 ( .A(net76258), .ZN(net75482) );
  AOI22_X2 U7121 ( .A1(REGFILE_reg_out_9__7_), .A2(net77698), .B1(
        REGFILE_reg_out_8__7_), .B2(n4829), .ZN(net75624) );
  NAND2_X1 U7122 ( .A1(REGFILE_reg_out_27__11_), .A2(n4872), .ZN(n9907) );
  NAND2_X1 U7123 ( .A1(REGFILE_reg_out_27__11_), .A2(net77416), .ZN(n7756) );
  INV_X1 U7124 ( .A(REGFILE_reg_out_15__10_), .ZN(n10144) );
  NAND2_X1 U7125 ( .A1(REGFILE_reg_out_15__10_), .A2(net77484), .ZN(n7814) );
  NAND2_X1 U7126 ( .A1(n6100), .A2(REGFILE_reg_out_13__11_), .ZN(n9877) );
  NAND2_X1 U7127 ( .A1(REGFILE_reg_out_13__11_), .A2(net77452), .ZN(n7769) );
  NAND2_X2 U7128 ( .A1(REGFILE_reg_out_25__8_), .A2(net77522), .ZN(n7883) );
  OAI22_X1 U7129 ( .A1(n8729), .A2(n8823), .B1(n6005), .B2(n8714), .ZN(n9297)
         );
  AOI22_X1 U7130 ( .A1(REGFILE_reg_out_26__28_), .A2(net77620), .B1(
        REGFILE_reg_out_27__28_), .B2(net89184), .ZN(n6312) );
  AOI22_X1 U7131 ( .A1(REGFILE_reg_out_26__0_), .A2(net77620), .B1(
        REGFILE_reg_out_27__0_), .B2(net89184), .ZN(n6913) );
  AOI22_X1 U7132 ( .A1(REGFILE_reg_out_26__1_), .A2(net77620), .B1(
        REGFILE_reg_out_27__1_), .B2(net77630), .ZN(n6889) );
  NAND4_X2 U7133 ( .A1(n6523), .A2(n6522), .A3(n6521), .A4(n6520), .ZN(n6524)
         );
  NAND2_X2 U7134 ( .A1(REGFILE_reg_out_10__14_), .A2(net77346), .ZN(n7642) );
  AOI22_X2 U7136 ( .A1(REGFILE_reg_out_16__9_), .A2(net87506), .B1(
        REGFILE_reg_out_15__9_), .B2(net75468), .ZN(n6716) );
  INV_X16 U7137 ( .A(net77640), .ZN(net77638) );
  INV_X8 U7138 ( .A(net76234), .ZN(net83168) );
  INV_X2 U7139 ( .A(n5871), .ZN(n5872) );
  INV_X2 U7140 ( .A(n5873), .ZN(n5874) );
  AOI22_X1 U7141 ( .A1(REGFILE_reg_out_0__23_), .A2(net82342), .B1(
        REGFILE_reg_out_10__23_), .B2(net75464), .ZN(n6415) );
  NAND2_X1 U7142 ( .A1(net77376), .A2(REGFILE_reg_out_12__10_), .ZN(n7819) );
  OAI21_X1 U7143 ( .B1(n9855), .B2(n9854), .A(n9853), .ZN(n9856) );
  OAI21_X2 U7144 ( .B1(n10381), .B2(n10380), .A(n10379), .ZN(n10384) );
  INV_X2 U7145 ( .A(n9029), .ZN(n9030) );
  XNOR2_X1 U7146 ( .A(n9029), .B(aluA[18]), .ZN(n9028) );
  NAND2_X1 U7147 ( .A1(aluA[18]), .A2(n10352), .ZN(n10353) );
  NOR2_X1 U7148 ( .A1(n5931), .A2(n10463), .ZN(n10362) );
  AOI21_X2 U7149 ( .B1(n10424), .B2(n10363), .A(n10362), .ZN(n10367) );
  INV_X2 U7150 ( .A(n5875), .ZN(n5876) );
  NAND2_X1 U7151 ( .A1(net73878), .A2(net73987), .ZN(n8301) );
  INV_X8 U7152 ( .A(n10371), .ZN(n5943) );
  NAND2_X4 U7153 ( .A1(net121496), .A2(net76195), .ZN(n6239) );
  NAND2_X1 U7154 ( .A1(REGFILE_reg_out_25__10_), .A2(net77522), .ZN(n7795) );
  NAND2_X1 U7155 ( .A1(REGFILE_reg_out_12__11_), .A2(net77380), .ZN(n7775) );
  NAND2_X1 U7156 ( .A1(REGFILE_reg_out_12__11_), .A2(n4873), .ZN(n9875) );
  INV_X2 U7157 ( .A(n5879), .ZN(n5880) );
  INV_X2 U7158 ( .A(n5881), .ZN(n5882) );
  NAND2_X1 U7159 ( .A1(n4878), .A2(REGFILE_reg_out_25__16_), .ZN(n9240) );
  NAND2_X1 U7160 ( .A1(net77528), .A2(REGFILE_reg_out_25__16_), .ZN(n7531) );
  INV_X2 U7161 ( .A(n5883), .ZN(n5884) );
  NOR2_X2 U7162 ( .A1(n9857), .A2(n9856), .ZN(n9858) );
  INV_X1 U7163 ( .A(n10422), .ZN(n9402) );
  AOI21_X2 U7164 ( .B1(n10422), .B2(n10370), .A(n10369), .ZN(n10374) );
  NAND3_X1 U7165 ( .A1(net71078), .A2(WIRE_ALU_A_MUX2TO1_32BIT_13__MUX_N1), 
        .A3(net85047), .ZN(n9413) );
  NOR2_X1 U7166 ( .A1(net85047), .A2(n10368), .ZN(n10369) );
  AOI22_X4 U7167 ( .A1(REGFILE_reg_out_31__18_), .A2(net77668), .B1(
        REGFILE_reg_out_3__18_), .B2(net77676), .ZN(n6540) );
  AOI22_X2 U7168 ( .A1(REGFILE_reg_out_7__10_), .A2(net75455), .B1(
        REGFILE_reg_out_6__10_), .B2(net75456), .ZN(n6701) );
  AOI22_X1 U7169 ( .A1(REGFILE_reg_out_24__0_), .A2(net77602), .B1(
        REGFILE_reg_out_25__0_), .B2(net77614), .ZN(n6912) );
  AOI22_X1 U7170 ( .A1(REGFILE_reg_out_24__1_), .A2(net77602), .B1(
        REGFILE_reg_out_25__1_), .B2(net77610), .ZN(n6888) );
  AOI22_X1 U7171 ( .A1(REGFILE_reg_out_24__28_), .A2(net75437), .B1(
        REGFILE_reg_out_25__28_), .B2(net77610), .ZN(n6311) );
  NAND4_X2 U7172 ( .A1(n6427), .A2(n6426), .A3(net75995), .A4(n6425), .ZN(
        n6428) );
  OAI21_X1 U7173 ( .B1(net148116), .B2(net73697), .A(net75843), .ZN(n5885) );
  NAND2_X1 U7174 ( .A1(REGFILE_reg_out_25__9_), .A2(net77522), .ZN(n7839) );
  NAND2_X1 U7175 ( .A1(REGFILE_reg_out_2__9_), .A2(net77342), .ZN(n7872) );
  NAND2_X1 U7176 ( .A1(REGFILE_reg_out_12__18_), .A2(net77384), .ZN(n7469) );
  AOI22_X1 U7177 ( .A1(REGFILE_reg_out_29__1_), .A2(net77650), .B1(
        REGFILE_reg_out_28__1_), .B2(n6911), .ZN(n6891) );
  NAND4_X2 U7178 ( .A1(n6891), .A2(n6890), .A3(n6889), .A4(n6888), .ZN(n6892)
         );
  INV_X16 U7179 ( .A(n5649), .ZN(n5890) );
  NOR2_X2 U7180 ( .A1(net76261), .A2(net88131), .ZN(n6000) );
  AOI22_X2 U7181 ( .A1(REGFILE_reg_out_26__12_), .A2(net75439), .B1(n5861), 
        .B2(net75440), .ZN(n6659) );
  AOI22_X2 U7182 ( .A1(REGFILE_reg_out_26__16_), .A2(net75439), .B1(
        REGFILE_reg_out_27__16_), .B2(net89184), .ZN(n6577) );
  INV_X8 U7183 ( .A(n8885), .ZN(n10929) );
  INV_X2 U7184 ( .A(n5891), .ZN(n5892) );
  AOI22_X2 U7185 ( .A1(REGFILE_reg_out_17__22_), .A2(net77798), .B1(
        REGFILE_reg_out_18__22_), .B2(n5890), .ZN(n6434) );
  INV_X2 U7186 ( .A(n5893), .ZN(n5894) );
  INV_X2 U7187 ( .A(n5895), .ZN(n5896) );
  INV_X2 U7188 ( .A(net82499), .ZN(net82500) );
  INV_X16 U7189 ( .A(net77106), .ZN(net77100) );
  NAND4_X2 U7190 ( .A1(n6465), .A2(n6464), .A3(n6462), .A4(n6463), .ZN(n6466)
         );
  NAND2_X4 U7191 ( .A1(n6342), .A2(n6341), .ZN(dmem_write_out[27]) );
  INV_X1 U7192 ( .A(n5762), .ZN(n8989) );
  NOR2_X1 U7193 ( .A1(n5762), .A2(n10327), .ZN(n10328) );
  NAND3_X1 U7194 ( .A1(n10930), .A2(n5762), .A3(net71078), .ZN(n8990) );
  OAI21_X1 U7195 ( .B1(n6457), .B2(net78055), .A(n6456), .ZN(n5897) );
  NOR2_X2 U7196 ( .A1(n6406), .A2(n6405), .ZN(n6407) );
  INV_X8 U7197 ( .A(net76222), .ZN(net75453) );
  INV_X8 U7198 ( .A(net76209), .ZN(net75443) );
  NAND2_X4 U7199 ( .A1(n6583), .A2(n6582), .ZN(dmem_write_out[16]) );
  AOI22_X1 U7200 ( .A1(REGFILE_reg_out_17__25_), .A2(net77798), .B1(
        REGFILE_reg_out_18__25_), .B2(n5890), .ZN(n6368) );
  AOI22_X2 U7201 ( .A1(REGFILE_reg_out_17__8_), .A2(net77794), .B1(
        REGFILE_reg_out_18__8_), .B2(n6896), .ZN(n6732) );
  INV_X8 U7202 ( .A(aluA[28]), .ZN(n6006) );
  AOI22_X4 U7203 ( .A1(REGFILE_reg_out_4__13_), .A2(n5679), .B1(n5817), .B2(
        net84475), .ZN(n6635) );
  XNOR2_X1 U7204 ( .A(n5870), .B(net77038), .ZN(n9057) );
  XNOR2_X1 U7205 ( .A(n5870), .B(n10463), .ZN(n10424) );
  INV_X16 U7206 ( .A(net76255), .ZN(net77836) );
  XNOR2_X1 U7207 ( .A(n9615), .B(n9656), .ZN(n9664) );
  OAI21_X2 U7208 ( .B1(n10395), .B2(n10394), .A(n10393), .ZN(n10398) );
  NAND2_X4 U7209 ( .A1(n5936), .A2(net123282), .ZN(n5899) );
  NAND2_X4 U7210 ( .A1(n5899), .A2(n5900), .ZN(aluA[29]) );
  NAND3_X2 U7211 ( .A1(n6980), .A2(n6981), .A3(n5753), .ZN(n6982) );
  NAND2_X1 U7212 ( .A1(REGFILE_reg_out_21__29_), .A2(net77462), .ZN(n6980) );
  NAND2_X1 U7214 ( .A1(REGFILE_reg_out_12__13_), .A2(n4873), .ZN(n9433) );
  NAND2_X1 U7215 ( .A1(REGFILE_reg_out_12__13_), .A2(net77380), .ZN(n7687) );
  AOI22_X1 U7216 ( .A1(REGFILE_reg_out_4__29_), .A2(n5678), .B1(
        REGFILE_reg_out_5__29_), .B2(net84475), .ZN(n6284) );
  NAND2_X1 U7217 ( .A1(n6093), .A2(REGFILE_reg_out_10__13_), .ZN(n9429) );
  NAND2_X1 U7218 ( .A1(REGFILE_reg_out_10__13_), .A2(net77344), .ZN(n7686) );
  INV_X4 U7219 ( .A(n5903), .ZN(n5904) );
  INV_X1 U7220 ( .A(n10910), .ZN(n5905) );
  NAND2_X1 U7221 ( .A1(n5904), .A2(n4872), .ZN(n9244) );
  NAND2_X1 U7222 ( .A1(REGFILE_reg_out_5__5_), .A2(net77456), .ZN(n8041) );
  NAND2_X1 U7223 ( .A1(REGFILE_reg_out_27__16_), .A2(net77420), .ZN(n7536) );
  NAND2_X1 U7224 ( .A1(aluA[16]), .A2(n5847), .ZN(n10359) );
  NAND2_X1 U7225 ( .A1(REGFILE_reg_out_10__5_), .A2(net77338), .ZN(n8036) );
  NAND2_X1 U7226 ( .A1(REGFILE_reg_out_2__5_), .A2(net77338), .ZN(n8046) );
  INV_X2 U7227 ( .A(n9050), .ZN(n9051) );
  XNOR2_X1 U7228 ( .A(n9050), .B(aluA[17]), .ZN(n9052) );
  AOI21_X2 U7229 ( .B1(n10448), .B2(n10358), .A(n10357), .ZN(n10361) );
  NOR2_X2 U7230 ( .A1(n10448), .A2(net78014), .ZN(n9023) );
  NAND2_X1 U7231 ( .A1(n6180), .A2(n5850), .ZN(n9473) );
  NAND2_X1 U7232 ( .A1(n5850), .A2(net77560), .ZN(n7664) );
  INV_X4 U7233 ( .A(n5906), .ZN(n5907) );
  INV_X2 U7234 ( .A(n5908), .ZN(n5909) );
  INV_X1 U7235 ( .A(n5897), .ZN(n10338) );
  AOI22_X1 U7236 ( .A1(REGFILE_reg_out_11__30_), .A2(net77750), .B1(
        REGFILE_reg_out_12__30_), .B2(net83168), .ZN(n6256) );
  AOI22_X1 U7237 ( .A1(REGFILE_reg_out_11__28_), .A2(net77750), .B1(
        REGFILE_reg_out_12__28_), .B2(net83168), .ZN(n6302) );
  AOI22_X1 U7238 ( .A1(REGFILE_reg_out_11__29_), .A2(net77750), .B1(
        REGFILE_reg_out_12__29_), .B2(net83168), .ZN(n6278) );
  AOI22_X1 U7239 ( .A1(REGFILE_reg_out_11__26_), .A2(net77750), .B1(
        REGFILE_reg_out_12__26_), .B2(net83168), .ZN(n6349) );
  XNOR2_X1 U7240 ( .A(n5905), .B(n10396), .ZN(n10399) );
  XNOR2_X1 U7241 ( .A(n5905), .B(net77038), .ZN(n9956) );
  NOR3_X1 U7242 ( .A1(net78003), .A2(n5905), .A3(n10396), .ZN(n9591) );
  NOR2_X1 U7243 ( .A1(n10910), .A2(n10396), .ZN(n10397) );
  AOI21_X2 U7244 ( .B1(n10399), .B2(n10398), .A(n10397), .ZN(n10403) );
  NOR2_X1 U7245 ( .A1(n10399), .A2(net78014), .ZN(n9607) );
  NAND2_X1 U7246 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_5__MUX_N1), .A2(n9956), .ZN(
        n9957) );
  AOI21_X2 U7247 ( .B1(n9592), .B2(net70697), .A(n9591), .ZN(n9632) );
  AOI22_X4 U7248 ( .A1(REGFILE_reg_out_31__8_), .A2(net77666), .B1(
        REGFILE_reg_out_3__8_), .B2(n5609), .ZN(n6742) );
  INV_X2 U7249 ( .A(n5911), .ZN(n5912) );
  XNOR2_X1 U7250 ( .A(n10933), .B(n9559), .ZN(n10431) );
  NOR2_X2 U7251 ( .A1(n10432), .A2(n10431), .ZN(n10439) );
  INV_X2 U7252 ( .A(REGFILE_reg_out_2__8_), .ZN(n9524) );
  NAND2_X1 U7253 ( .A1(REGFILE_reg_out_2__8_), .A2(net77342), .ZN(n7916) );
  INV_X4 U7254 ( .A(net36479), .ZN(net81810) );
  AOI21_X2 U7255 ( .B1(n10344), .B2(n10343), .A(n10342), .ZN(n10348) );
  NOR3_X1 U7256 ( .A1(n9559), .A2(n10341), .A3(net78003), .ZN(n9560) );
  XNOR2_X1 U7257 ( .A(n10933), .B(n4810), .ZN(n9543) );
  OAI21_X2 U7258 ( .B1(n10348), .B2(n10347), .A(n10346), .ZN(n10351) );
  NOR3_X2 U7259 ( .A1(n9562), .A2(n9561), .A3(n9560), .ZN(n9563) );
  INV_X1 U7260 ( .A(n5783), .ZN(n9559) );
  AOI22_X1 U7261 ( .A1(REGFILE_reg_out_30__0_), .A2(net77634), .B1(
        REGFILE_reg_out_2__0_), .B2(net75442), .ZN(n6914) );
  AOI22_X1 U7262 ( .A1(REGFILE_reg_out_30__29_), .A2(net77638), .B1(
        REGFILE_reg_out_2__29_), .B2(net75442), .ZN(n6289) );
  AOI22_X1 U7263 ( .A1(REGFILE_reg_out_30__28_), .A2(net77638), .B1(
        REGFILE_reg_out_2__28_), .B2(net75442), .ZN(n6313) );
  XNOR2_X1 U7264 ( .A(n5897), .B(net77038), .ZN(n8813) );
  AOI22_X1 U7265 ( .A1(REGFILE_reg_out_7__0_), .A2(net77716), .B1(
        REGFILE_reg_out_6__0_), .B2(net75456), .ZN(n6910) );
  AOI22_X2 U7266 ( .A1(REGFILE_reg_out_7__15_), .A2(net77714), .B1(
        REGFILE_reg_out_6__15_), .B2(net75456), .ZN(n6597) );
  AOI22_X2 U7267 ( .A1(REGFILE_reg_out_17__9_), .A2(net77794), .B1(
        REGFILE_reg_out_18__9_), .B2(n6896), .ZN(n6710) );
  AOI22_X2 U7268 ( .A1(REGFILE_reg_out_19__9_), .A2(net77810), .B1(
        REGFILE_reg_out_1__9_), .B2(net75478), .ZN(n6711) );
  AOI22_X1 U7269 ( .A1(REGFILE_reg_out_0__2_), .A2(net82342), .B1(
        REGFILE_reg_out_10__2_), .B2(net75464), .ZN(n6856) );
  AOI22_X1 U7270 ( .A1(REGFILE_reg_out_17__31_), .A2(net77798), .B1(
        REGFILE_reg_out_18__31_), .B2(n5890), .ZN(n6225) );
  AOI22_X1 U7271 ( .A1(REGFILE_reg_out_17__30_), .A2(net77798), .B1(
        REGFILE_reg_out_18__30_), .B2(n5890), .ZN(n6251) );
  AOI22_X1 U7272 ( .A1(REGFILE_reg_out_17__29_), .A2(net77798), .B1(
        REGFILE_reg_out_18__29_), .B2(n5890), .ZN(n6273) );
  AOI22_X1 U7273 ( .A1(REGFILE_reg_out_17__28_), .A2(net77798), .B1(
        REGFILE_reg_out_18__28_), .B2(n5890), .ZN(n6297) );
  AOI22_X1 U7274 ( .A1(REGFILE_reg_out_17__26_), .A2(net77798), .B1(
        REGFILE_reg_out_18__26_), .B2(n5890), .ZN(n6344) );
  INV_X1 U7275 ( .A(n4852), .ZN(n10352) );
  NAND2_X4 U7276 ( .A1(n10046), .A2(net76270), .ZN(n10052) );
  NAND2_X1 U7277 ( .A1(n6093), .A2(REGFILE_reg_out_10__7_), .ZN(n9707) );
  NAND2_X1 U7278 ( .A1(REGFILE_reg_out_10__7_), .A2(net77338), .ZN(n7950) );
  INV_X2 U7279 ( .A(n5846), .ZN(n10266) );
  NAND2_X1 U7280 ( .A1(n5846), .A2(net77382), .ZN(n7643) );
  NAND2_X1 U7281 ( .A1(REGFILE_reg_out_27__14_), .A2(net77418), .ZN(n7624) );
  NAND2_X1 U7282 ( .A1(n4879), .A2(REGFILE_reg_out_2__7_), .ZN(n9749) );
  NAND2_X1 U7283 ( .A1(REGFILE_reg_out_2__7_), .A2(net77338), .ZN(n7958) );
  NAND2_X1 U7284 ( .A1(REGFILE_reg_out_27__7_), .A2(n4872), .ZN(n9743) );
  OR2_X2 U7285 ( .A1(n5914), .A2(net77506), .ZN(n6970) );
  INV_X2 U7286 ( .A(REGFILE_reg_out_25__14_), .ZN(n10269) );
  NAND2_X1 U7287 ( .A1(REGFILE_reg_out_25__14_), .A2(net77526), .ZN(n7619) );
  INV_X2 U7288 ( .A(REGFILE_reg_out_14__31_), .ZN(n10520) );
  AOI22_X1 U7289 ( .A1(REGFILE_reg_out_14__31_), .A2(net77778), .B1(
        REGFILE_reg_out_13__31_), .B2(n6009), .ZN(n6232) );
  INV_X1 U7290 ( .A(n5619), .ZN(net73850) );
  INV_X2 U7291 ( .A(REGFILE_reg_out_12__31_), .ZN(n10515) );
  AOI22_X1 U7292 ( .A1(REGFILE_reg_out_11__31_), .A2(net77750), .B1(
        REGFILE_reg_out_12__31_), .B2(net83167), .ZN(n6230) );
  NAND2_X2 U7293 ( .A1(REGFILE_reg_out_8__29_), .A2(net77318), .ZN(n6973) );
  AOI21_X2 U7294 ( .B1(n10446), .B2(n10351), .A(n10350), .ZN(n10355) );
  NAND4_X1 U7295 ( .A1(n10448), .A2(n10447), .A3(n10446), .A4(n10445), .ZN(
        n10449) );
  NOR2_X2 U7296 ( .A1(n10446), .A2(net78014), .ZN(n9985) );
  INV_X2 U7297 ( .A(n8819), .ZN(n8820) );
  XNOR2_X1 U7298 ( .A(n8819), .B(aluA[19]), .ZN(n9992) );
  AOI22_X2 U7299 ( .A1(REGFILE_reg_out_17__7_), .A2(net77794), .B1(
        REGFILE_reg_out_18__7_), .B2(n5890), .ZN(n6754) );
  INV_X1 U7300 ( .A(n5650), .ZN(n9995) );
  NOR2_X1 U7301 ( .A1(n5783), .A2(n10341), .ZN(n10342) );
  INV_X2 U7302 ( .A(n8815), .ZN(n8816) );
  XNOR2_X1 U7303 ( .A(n8815), .B(aluA[20]), .ZN(n10053) );
  NAND4_X1 U7304 ( .A1(n10444), .A2(n10443), .A3(n10442), .A4(n10441), .ZN(
        n10450) );
  NOR2_X2 U7305 ( .A1(n10443), .A2(net78014), .ZN(n10055) );
  NAND2_X1 U7306 ( .A1(aluA[20]), .A2(n10345), .ZN(n10346) );
  NOR3_X2 U7307 ( .A1(n10345), .A2(n10071), .A3(net78003), .ZN(n10072) );
  AOI22_X1 U7308 ( .A1(REGFILE_reg_out_17__0_), .A2(net77794), .B1(
        REGFILE_reg_out_18__0_), .B2(n5890), .ZN(n6897) );
  AOI22_X1 U7309 ( .A1(REGFILE_reg_out_17__1_), .A2(net77794), .B1(
        REGFILE_reg_out_18__1_), .B2(n5890), .ZN(n6874) );
  AOI22_X1 U7310 ( .A1(REGFILE_reg_out_17__2_), .A2(net77794), .B1(
        REGFILE_reg_out_18__2_), .B2(n5890), .ZN(n6852) );
  AOI22_X1 U7311 ( .A1(REGFILE_reg_out_17__4_), .A2(net77794), .B1(
        REGFILE_reg_out_18__4_), .B2(n5890), .ZN(n6808) );
  AOI22_X1 U7312 ( .A1(REGFILE_reg_out_17__3_), .A2(net77794), .B1(
        REGFILE_reg_out_18__3_), .B2(n5890), .ZN(n6830) );
  XNOR2_X1 U7313 ( .A(n5675), .B(net77038), .ZN(n8815) );
  XNOR2_X1 U7314 ( .A(n5675), .B(aluA[20]), .ZN(n10443) );
  INV_X1 U7315 ( .A(n5675), .ZN(n10345) );
  XNOR2_X1 U7316 ( .A(n5848), .B(aluA[18]), .ZN(n10445) );
  XNOR2_X1 U7317 ( .A(n5848), .B(net77038), .ZN(n9029) );
  NOR2_X1 U7318 ( .A1(n5650), .A2(n10349), .ZN(n10350) );
  XNOR2_X1 U7319 ( .A(n5650), .B(aluA[19]), .ZN(n10446) );
  XNOR2_X1 U7320 ( .A(n5650), .B(net77038), .ZN(n8819) );
  NAND2_X1 U7321 ( .A1(REGFILE_reg_out_27__7_), .A2(net77410), .ZN(n7932) );
  NAND2_X1 U7322 ( .A1(net77418), .A2(REGFILE_reg_out_27__15_), .ZN(n7580) );
  NAND2_X2 U7323 ( .A1(REGFILE_reg_out_0__6_), .A2(net120684), .ZN(n5945) );
  NOR2_X2 U7324 ( .A1(n6839), .A2(n6838), .ZN(n6851) );
  AOI22_X1 U7325 ( .A1(REGFILE_reg_out_30__3_), .A2(net77634), .B1(
        REGFILE_reg_out_2__3_), .B2(net82613), .ZN(n6846) );
  NOR2_X1 U7326 ( .A1(net36479), .A2(n10464), .ZN(n10389) );
  NAND3_X1 U7327 ( .A1(net71078), .A2(WIRE_ALU_A_MUX2TO1_32BIT_7__MUX_N1), 
        .A3(net36479), .ZN(n9691) );
  AOI22_X2 U7328 ( .A1(REGFILE_reg_out_4__6_), .A2(n5678), .B1(
        REGFILE_reg_out_5__6_), .B2(net84475), .ZN(n6775) );
  NAND2_X1 U7329 ( .A1(n4878), .A2(REGFILE_reg_out_25__7_), .ZN(n9739) );
  NAND2_X1 U7330 ( .A1(REGFILE_reg_out_25__7_), .A2(net77520), .ZN(n7927) );
  AOI22_X1 U7331 ( .A1(net73838), .A2(n10949), .B1(n6019), .B2(n5998), .ZN(
        n8413) );
  INV_X4 U7332 ( .A(n5958), .ZN(n5919) );
  INV_X2 U7333 ( .A(n5920), .ZN(n5921) );
  INV_X2 U7334 ( .A(n5922), .ZN(n5923) );
  INV_X2 U7335 ( .A(n5925), .ZN(n5926) );
  INV_X2 U7336 ( .A(n5927), .ZN(n5928) );
  INV_X2 U7337 ( .A(n5929), .ZN(n5930) );
  NAND2_X1 U7338 ( .A1(n10423), .A2(n10422), .ZN(n10427) );
  AOI22_X4 U7339 ( .A1(REGFILE_reg_out_4__10_), .A2(net75451), .B1(n4798), 
        .B2(net84475), .ZN(n6699) );
  XNOR2_X1 U7340 ( .A(n5885), .B(net77038), .ZN(n9050) );
  XNOR2_X1 U7341 ( .A(n5885), .B(aluA[17]), .ZN(n10448) );
  NOR2_X1 U7342 ( .A1(n5885), .A2(n10356), .ZN(n10357) );
  INV_X1 U7343 ( .A(n5885), .ZN(n9035) );
  NAND3_X4 U7344 ( .A1(net75368), .A2(n6955), .A3(net75367), .ZN(aluA[30]) );
  AOI22_X1 U7345 ( .A1(REGFILE_reg_out_4__1_), .A2(n5678), .B1(
        REGFILE_reg_out_5__1_), .B2(net84475), .ZN(n6885) );
  AOI22_X1 U7346 ( .A1(REGFILE_reg_out_4__2_), .A2(n5679), .B1(
        REGFILE_reg_out_5__2_), .B2(net75452), .ZN(n6863) );
  AOI22_X1 U7347 ( .A1(REGFILE_reg_out_4__3_), .A2(net75451), .B1(
        REGFILE_reg_out_5__3_), .B2(net75452), .ZN(n6841) );
  NOR2_X4 U7348 ( .A1(n6571), .A2(n6570), .ZN(n6583) );
  OAI22_X1 U7349 ( .A1(n10290), .A2(net70691), .B1(n10289), .B2(n5870), .ZN(
        n10291) );
  INV_X4 U7350 ( .A(net77386), .ZN(net77396) );
  INV_X4 U7351 ( .A(net77386), .ZN(net77394) );
  AOI22_X1 U7352 ( .A1(REGFILE_reg_out_16__1_), .A2(net87506), .B1(
        REGFILE_reg_out_15__1_), .B2(n5579), .ZN(n6880) );
  XNOR2_X1 U7353 ( .A(net81810), .B(net77040), .ZN(n9612) );
  XNOR2_X1 U7354 ( .A(net81810), .B(n10464), .ZN(n10391) );
  AOI22_X1 U7355 ( .A1(REGFILE_reg_out_14__0_), .A2(net77778), .B1(
        REGFILE_reg_out_13__0_), .B2(n6009), .ZN(n6904) );
  AOI22_X1 U7356 ( .A1(REGFILE_reg_out_14__1_), .A2(net77778), .B1(
        REGFILE_reg_out_13__1_), .B2(n5663), .ZN(n6881) );
  AOI22_X1 U7357 ( .A1(REGFILE_reg_out_14__2_), .A2(net77778), .B1(
        REGFILE_reg_out_13__2_), .B2(n5663), .ZN(n6859) );
  AOI22_X1 U7358 ( .A1(REGFILE_reg_out_14__3_), .A2(net77778), .B1(
        REGFILE_reg_out_13__3_), .B2(n5664), .ZN(n6837) );
  AOI22_X1 U7359 ( .A1(REGFILE_reg_out_14__4_), .A2(net77778), .B1(
        REGFILE_reg_out_13__4_), .B2(n6009), .ZN(n6815) );
  AOI22_X4 U7360 ( .A1(REGFILE_reg_out_31__17_), .A2(net77668), .B1(
        REGFILE_reg_out_3__17_), .B2(net77676), .ZN(n6558) );
  XNOR2_X1 U7361 ( .A(n5805), .B(net77038), .ZN(n9059) );
  XNOR2_X1 U7362 ( .A(n5805), .B(n10247), .ZN(n10425) );
  AND3_X4 U7364 ( .A1(instruction[16]), .A2(net77272), .A3(net78056), .ZN(
        n5933) );
  AOI22_X1 U7365 ( .A1(REGFILE_reg_out_19__30_), .A2(net77814), .B1(
        REGFILE_reg_out_1__30_), .B2(net82631), .ZN(n6252) );
  INV_X2 U7366 ( .A(n5934), .ZN(n5935) );
  XNOR2_X1 U7367 ( .A(n5867), .B(n10375), .ZN(n10420) );
  XNOR2_X1 U7368 ( .A(n5867), .B(net77040), .ZN(n9354) );
  NAND4_X1 U7369 ( .A1(n10421), .A2(n10420), .A3(n10419), .A4(n10418), .ZN(
        n10428) );
  AOI21_X2 U7370 ( .B1(n10420), .B2(n10377), .A(n10376), .ZN(n10381) );
  NAND2_X1 U7371 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_11__MUX_N1), .A2(n9354), .ZN(
        n9355) );
  INV_X2 U7372 ( .A(REGFILE_reg_out_9__30_), .ZN(n8757) );
  INV_X2 U7373 ( .A(REGFILE_reg_out_1__31_), .ZN(net70780) );
  AOI22_X1 U7374 ( .A1(REGFILE_reg_out_19__31_), .A2(net77814), .B1(
        REGFILE_reg_out_1__31_), .B2(net82631), .ZN(n6226) );
  NAND2_X1 U7375 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_14__MUX_N1), .A2(n5805), .ZN(
        n10365) );
  AOI22_X4 U7376 ( .A1(REGFILE_reg_out_31__9_), .A2(net77666), .B1(
        REGFILE_reg_out_3__9_), .B2(net77676), .ZN(n6720) );
  INV_X8 U7377 ( .A(n9616), .ZN(n10910) );
  AOI22_X1 U7378 ( .A1(REGFILE_reg_out_7__2_), .A2(net75455), .B1(
        REGFILE_reg_out_6__2_), .B2(net75456), .ZN(n6865) );
  NOR2_X1 U7379 ( .A1(n10375), .A2(n10915), .ZN(n10376) );
  NAND3_X1 U7380 ( .A1(net71078), .A2(WIRE_ALU_A_MUX2TO1_32BIT_11__MUX_N1), 
        .A3(n5868), .ZN(n9853) );
  XNOR2_X1 U7381 ( .A(net84663), .B(net77040), .ZN(n9060) );
  XNOR2_X1 U7382 ( .A(net84663), .B(n10368), .ZN(n10422) );
  NAND2_X1 U7383 ( .A1(n4879), .A2(REGFILE_reg_out_2__13_), .ZN(n9471) );
  INV_X2 U7384 ( .A(n5937), .ZN(n5938) );
  INV_X2 U7385 ( .A(n5939), .ZN(n5940) );
  AND2_X2 U7386 ( .A1(n5942), .A2(n5941), .ZN(n6640) );
  NAND3_X1 U7387 ( .A1(net71078), .A2(aluA[16]), .A3(n5769), .ZN(n9195) );
  XNOR2_X1 U7388 ( .A(n5769), .B(net77038), .ZN(n9054) );
  XNOR2_X1 U7389 ( .A(n5769), .B(aluA[16]), .ZN(n10447) );
  NAND2_X4 U7390 ( .A1(n6604), .A2(n6605), .ZN(dmem_write_out[15]) );
  AOI22_X1 U7391 ( .A1(REGFILE_reg_out_31__1_), .A2(net77666), .B1(
        REGFILE_reg_out_3__1_), .B2(n5609), .ZN(n6884) );
  AOI22_X1 U7392 ( .A1(REGFILE_reg_out_31__3_), .A2(net77666), .B1(
        REGFILE_reg_out_3__3_), .B2(n5609), .ZN(n6840) );
  NAND2_X4 U7393 ( .A1(n6628), .A2(n6629), .ZN(dmem_write_out[14]) );
  NAND2_X1 U7394 ( .A1(n10615), .A2(REGFILE_reg_out_30__30_), .ZN(n8754) );
  AOI22_X1 U7395 ( .A1(REGFILE_reg_out_30__30_), .A2(net77638), .B1(
        REGFILE_reg_out_2__30_), .B2(net75442), .ZN(n6267) );
  AND2_X2 U7396 ( .A1(n5946), .A2(n5945), .ZN(n6768) );
  AOI22_X2 U7397 ( .A1(REGFILE_reg_out_30__6_), .A2(net77634), .B1(
        REGFILE_reg_out_2__6_), .B2(net75442), .ZN(n6780) );
  INV_X16 U7398 ( .A(n10946), .ZN(net77104) );
  NAND3_X1 U7399 ( .A1(net71078), .A2(WIRE_ALU_A_MUX2TO1_32BIT_12__MUX_N1), 
        .A3(n5577), .ZN(n9099) );
  AOI22_X1 U7400 ( .A1(REGFILE_reg_out_0__30_), .A2(net82342), .B1(
        REGFILE_reg_out_10__30_), .B2(net81764), .ZN(n6255) );
  AOI22_X1 U7401 ( .A1(REGFILE_reg_out_0__28_), .A2(net82342), .B1(
        REGFILE_reg_out_10__28_), .B2(net75464), .ZN(n6301) );
  AOI22_X1 U7402 ( .A1(REGFILE_reg_out_0__29_), .A2(net82342), .B1(
        REGFILE_reg_out_10__29_), .B2(net75464), .ZN(n6277) );
  AOI22_X1 U7403 ( .A1(REGFILE_reg_out_0__26_), .A2(net82342), .B1(
        REGFILE_reg_out_10__26_), .B2(net75464), .ZN(n6348) );
  AOI22_X1 U7404 ( .A1(REGFILE_reg_out_0__0_), .A2(net82342), .B1(
        REGFILE_reg_out_10__0_), .B2(net81764), .ZN(n6901) );
  OAI22_X1 U7405 ( .A1(n10256), .A2(net70691), .B1(n10255), .B2(n5805), .ZN(
        n10257) );
  INV_X8 U7406 ( .A(n10364), .ZN(n10916) );
  INV_X2 U7407 ( .A(REGFILE_reg_out_10__31_), .ZN(n10513) );
  AOI22_X1 U7408 ( .A1(REGFILE_reg_out_0__31_), .A2(net82342), .B1(
        REGFILE_reg_out_10__31_), .B2(net81764), .ZN(n6229) );
  AOI22_X2 U7409 ( .A1(REGFILE_reg_out_16__8_), .A2(net87506), .B1(
        REGFILE_reg_out_15__8_), .B2(net75468), .ZN(n6738) );
  INV_X2 U7410 ( .A(n5950), .ZN(n5951) );
  XNOR2_X1 U7411 ( .A(n5826), .B(net77040), .ZN(n9508) );
  XNOR2_X1 U7412 ( .A(n5826), .B(n10382), .ZN(n10418) );
  NOR3_X1 U7413 ( .A1(net78003), .A2(n5826), .A3(n10382), .ZN(n9337) );
  NOR2_X1 U7414 ( .A1(n10913), .A2(n10382), .ZN(n10383) );
  AOI22_X2 U7415 ( .A1(REGFILE_reg_out_0__8_), .A2(net120684), .B1(
        REGFILE_reg_out_10__8_), .B2(net75464), .ZN(n6736) );
  NOR2_X2 U7416 ( .A1(n6849), .A2(n6848), .ZN(n6850) );
  AOI22_X1 U7417 ( .A1(REGFILE_reg_out_30__1_), .A2(net77634), .B1(
        REGFILE_reg_out_2__1_), .B2(net75442), .ZN(n6890) );
  AOI22_X1 U7418 ( .A1(REGFILE_reg_out_0__1_), .A2(net82342), .B1(
        REGFILE_reg_out_10__1_), .B2(net81764), .ZN(n6878) );
  XNOR2_X1 U7419 ( .A(n5944), .B(net77038), .ZN(n9351) );
  NAND2_X1 U7420 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_12__MUX_N1), .A2(n5944), .ZN(
        n10372) );
  XNOR2_X1 U7421 ( .A(n5944), .B(n9075), .ZN(n10423) );
  OAI22_X1 U7422 ( .A1(n10134), .A2(net70691), .B1(n10133), .B2(n5713), .ZN(
        n10135) );
  XNOR2_X1 U7423 ( .A(n5713), .B(net77040), .ZN(n9357) );
  NAND2_X1 U7424 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_10__MUX_N1), .A2(n5713), .ZN(
        n10379) );
  XNOR2_X1 U7425 ( .A(n5713), .B(n10125), .ZN(n10421) );
  INV_X1 U7426 ( .A(n5815), .ZN(n5952) );
  INV_X4 U7427 ( .A(net78235), .ZN(net80443) );
  AOI22_X2 U7429 ( .A1(REGFILE_reg_out_19__5_), .A2(net77810), .B1(
        REGFILE_reg_out_1__5_), .B2(net82631), .ZN(n6787) );
  AOI22_X2 U7430 ( .A1(REGFILE_reg_out_31__5_), .A2(net77666), .B1(
        REGFILE_reg_out_3__5_), .B2(n5609), .ZN(n6796) );
  INV_X2 U7431 ( .A(n5956), .ZN(n5957) );
  INV_X1 U7432 ( .A(REGFILE_reg_out_16__30_), .ZN(n8745) );
  XNOR2_X1 U7433 ( .A(n8587), .B(n5955), .ZN(n9809) );
  NAND2_X1 U7434 ( .A1(net73708), .A2(n5955), .ZN(n8696) );
  NAND2_X1 U7435 ( .A1(n6040), .A2(n5955), .ZN(n8726) );
  NAND2_X1 U7436 ( .A1(n10542), .A2(n5955), .ZN(n8768) );
  NAND2_X1 U7437 ( .A1(n9065), .A2(n5955), .ZN(n8822) );
  AOI22_X1 U7438 ( .A1(n8974), .A2(net72962), .B1(n4912), .B2(n5955), .ZN(
        n9771) );
  NAND2_X1 U7439 ( .A1(net70720), .A2(n5955), .ZN(n9070) );
  NAND2_X1 U7440 ( .A1(net70719), .A2(n5955), .ZN(n9599) );
  INV_X1 U7441 ( .A(n5955), .ZN(n10312) );
  XNOR2_X1 U7442 ( .A(n5955), .B(n6005), .ZN(n10442) );
  NAND2_X1 U7443 ( .A1(n8588), .A2(n5955), .ZN(n8589) );
  AOI22_X2 U7444 ( .A1(REGFILE_reg_out_19__1_), .A2(net77810), .B1(
        REGFILE_reg_out_1__1_), .B2(net82631), .ZN(n6875) );
  INV_X16 U7445 ( .A(net75455), .ZN(net77720) );
  INV_X8 U7446 ( .A(n10408), .ZN(n10907) );
  AOI21_X2 U7447 ( .B1(n10407), .B2(n10406), .A(n10405), .ZN(n10410) );
  OAI21_X2 U7448 ( .B1(n10410), .B2(n10414), .A(n10409), .ZN(n10411) );
  AOI22_X2 U7449 ( .A1(REGFILE_reg_out_21__2_), .A2(net77842), .B1(
        REGFILE_reg_out_20__2_), .B2(net77850), .ZN(n6855) );
  NOR2_X1 U7450 ( .A1(n10908), .A2(n10404), .ZN(n10405) );
  NAND4_X2 U7451 ( .A1(n6868), .A2(n6869), .A3(n6867), .A4(n6866), .ZN(n6870)
         );
  NAND2_X4 U7452 ( .A1(n8539), .A2(net73496), .ZN(net73622) );
  INV_X8 U7453 ( .A(net76249), .ZN(net75475) );
  NOR2_X4 U7454 ( .A1(n6883), .A2(n6882), .ZN(n6895) );
  NAND2_X4 U7455 ( .A1(n6665), .A2(n6664), .ZN(dmem_write_out[12]) );
  NAND2_X4 U7456 ( .A1(n6687), .A2(n6686), .ZN(dmem_write_out[11]) );
  NAND2_X4 U7457 ( .A1(n6708), .A2(n6709), .ZN(dmem_write_out[10]) );
  INV_X2 U7458 ( .A(n5959), .ZN(n5960) );
  OAI22_X1 U7459 ( .A1(net73608), .A2(n8823), .B1(n10319), .B2(n8634), .ZN(
        n8974) );
  AOI21_X1 U7460 ( .B1(n10305), .B2(n10304), .A(net73608), .ZN(n10461) );
  INV_X2 U7461 ( .A(n5961), .ZN(n5962) );
  AOI21_X1 U7462 ( .B1(n6019), .B2(n8401), .A(n8400), .ZN(n8415) );
  NOR2_X4 U7463 ( .A1(n6952), .A2(n6951), .ZN(n6953) );
  INV_X2 U7464 ( .A(n5963), .ZN(n5964) );
  INV_X2 U7465 ( .A(n5965), .ZN(n5966) );
  INV_X2 U7466 ( .A(n5967), .ZN(n5968) );
  INV_X2 U7467 ( .A(n5969), .ZN(n5970) );
  XNOR2_X1 U7468 ( .A(n5758), .B(n9535), .ZN(n10419) );
  XNOR2_X1 U7469 ( .A(n5758), .B(net77040), .ZN(n9609) );
  OAI22_X1 U7470 ( .A1(n9513), .A2(net70691), .B1(n9512), .B2(n5758), .ZN(
        n9514) );
  NAND2_X1 U7471 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_8__MUX_N1), .A2(n5758), .ZN(
        n10386) );
  XNOR2_X1 U7472 ( .A(n9609), .B(n9535), .ZN(n9610) );
  INV_X2 U7473 ( .A(n5971), .ZN(n5972) );
  NOR2_X1 U7474 ( .A1(net73842), .A2(net73848), .ZN(n8405) );
  NOR3_X2 U7475 ( .A1(n8406), .A2(n8405), .A3(n8404), .ZN(n8414) );
  INV_X2 U7476 ( .A(n5973), .ZN(n5974) );
  AOI22_X4 U7477 ( .A1(n5923), .A2(net77444), .B1(n5966), .B2(net77400), .ZN(
        n6936) );
  INV_X1 U7478 ( .A(net80390), .ZN(net73848) );
  AOI22_X1 U7479 ( .A1(REGFILE_reg_out_4__0_), .A2(n5678), .B1(
        REGFILE_reg_out_5__0_), .B2(net84475), .ZN(n6908) );
  AOI22_X4 U7480 ( .A1(REGFILE_reg_out_29__8_), .A2(net77650), .B1(
        REGFILE_reg_out_28__8_), .B2(n6911), .ZN(n6749) );
  OAI22_X1 U7481 ( .A1(n9666), .A2(net70691), .B1(n9665), .B2(n5757), .ZN(
        n9667) );
  XNOR2_X1 U7482 ( .A(n5757), .B(net77040), .ZN(n9615) );
  NAND2_X1 U7483 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_6__MUX_N1), .A2(n5757), .ZN(
        n10393) );
  XNOR2_X1 U7484 ( .A(n5757), .B(n9656), .ZN(n9657) );
  NAND2_X2 U7485 ( .A1(REGFILE_reg_out_19__4_), .A2(net77810), .ZN(n5975) );
  NAND2_X1 U7486 ( .A1(REGFILE_reg_out_1__4_), .A2(net75478), .ZN(n5976) );
  AND2_X2 U7487 ( .A1(n5975), .A2(n5976), .ZN(n6809) );
  NOR2_X4 U7488 ( .A1(n5815), .A2(n6946), .ZN(n6954) );
  INV_X2 U7489 ( .A(REGFILE_reg_out_8__30_), .ZN(n8756) );
  AOI22_X1 U7490 ( .A1(REGFILE_reg_out_9__30_), .A2(net77702), .B1(
        REGFILE_reg_out_8__30_), .B2(n4829), .ZN(n6263) );
  NAND2_X1 U7491 ( .A1(REGFILE_reg_out_3__3_), .A2(net77410), .ZN(n8136) );
  NAND2_X1 U7493 ( .A1(REGFILE_reg_out_1__4_), .A2(net77518), .ZN(n8087) );
  INV_X2 U7496 ( .A(n5985), .ZN(n5986) );
  OR2_X2 U7497 ( .A1(n5987), .A2(net77542), .ZN(n6972) );
  INV_X16 U7498 ( .A(net74051), .ZN(net77542) );
  NAND2_X1 U7499 ( .A1(net76488), .A2(REGFILE_reg_out_31__29_), .ZN(n9831) );
  AOI22_X1 U7500 ( .A1(REGFILE_reg_out_31__29_), .A2(net77670), .B1(
        REGFILE_reg_out_3__29_), .B2(n5609), .ZN(n6283) );
  INV_X1 U7501 ( .A(REGFILE_reg_out_23__29_), .ZN(net71824) );
  AOI22_X1 U7502 ( .A1(REGFILE_reg_out_23__29_), .A2(net77826), .B1(
        REGFILE_reg_out_22__29_), .B2(net77834), .ZN(n6275) );
  INV_X2 U7503 ( .A(n5989), .ZN(n5990) );
  INV_X1 U7504 ( .A(REGFILE_reg_out_15__29_), .ZN(n9828) );
  AOI22_X1 U7505 ( .A1(REGFILE_reg_out_21__29_), .A2(net77846), .B1(
        REGFILE_reg_out_20__29_), .B2(net77854), .ZN(n6276) );
  INV_X1 U7506 ( .A(REGFILE_reg_out_28__29_), .ZN(n10934) );
  AOI22_X1 U7507 ( .A1(REGFILE_reg_out_29__29_), .A2(net77650), .B1(
        REGFILE_reg_out_28__29_), .B2(n6911), .ZN(n6290) );
  AOI22_X1 U7508 ( .A1(REGFILE_reg_out_19__0_), .A2(net77810), .B1(
        REGFILE_reg_out_1__0_), .B2(net82631), .ZN(n6898) );
  AOI22_X1 U7509 ( .A1(REGFILE_reg_out_31__0_), .A2(net77666), .B1(
        REGFILE_reg_out_3__0_), .B2(n5609), .ZN(n6907) );
  AOI22_X1 U7510 ( .A1(REGFILE_reg_out_31__2_), .A2(net77666), .B1(
        REGFILE_reg_out_3__2_), .B2(n5609), .ZN(n6862) );
  AOI22_X1 U7511 ( .A1(REGFILE_reg_out_31__4_), .A2(net77666), .B1(n5982), 
        .B2(n5609), .ZN(n6818) );
  INV_X8 U7512 ( .A(n9358), .ZN(n10913) );
  AOI22_X2 U7513 ( .A1(REGFILE_reg_out_31__6_), .A2(net77666), .B1(
        REGFILE_reg_out_3__6_), .B2(n5609), .ZN(n6774) );
  AOI22_X2 U7514 ( .A1(REGFILE_reg_out_17__6_), .A2(net77794), .B1(
        REGFILE_reg_out_18__6_), .B2(n5890), .ZN(n6764) );
  NOR2_X4 U7515 ( .A1(n6817), .A2(n6816), .ZN(n6829) );
  NAND2_X4 U7516 ( .A1(n6248), .A2(n4865), .ZN(net73629) );
  INV_X32 U7517 ( .A(instruction[4]), .ZN(net73498) );
  INV_X8 U7518 ( .A(net76211), .ZN(net76195) );
  NAND2_X4 U7519 ( .A1(REGFILE_reg_out_24__29_), .A2(net77318), .ZN(n6985) );
  NAND2_X4 U7520 ( .A1(n6785), .A2(n6784), .ZN(dmem_write_out[6]) );
  NAND2_X4 U7521 ( .A1(n6873), .A2(n6872), .ZN(dmem_write_out[2]) );
  NOR3_X1 U7522 ( .A1(n8451), .A2(n5748), .A3(n8450), .ZN(n8452) );
  AOI22_X1 U7523 ( .A1(REGFILE_reg_out_24__31_), .A2(net77602), .B1(
        REGFILE_reg_out_25__31_), .B2(net77610), .ZN(n6240) );
  XNOR2_X1 U7524 ( .A(n8584), .B(net80189), .ZN(n8583) );
  INV_X4 U7525 ( .A(net78107), .ZN(net75401) );
  INV_X2 U7526 ( .A(n5992), .ZN(n5993) );
  AOI22_X1 U7527 ( .A1(net77588), .A2(n4834), .B1(n8411), .B2(n5952), .ZN(
        n8412) );
  AOI22_X4 U7528 ( .A1(n5830), .A2(net77478), .B1(n5993), .B2(net77550), .ZN(
        n6949) );
  INV_X1 U7529 ( .A(n6952), .ZN(n5998) );
  NAND2_X1 U7530 ( .A1(net73708), .A2(net80189), .ZN(n10655) );
  NAND3_X2 U7531 ( .A1(n10470), .A2(net80189), .A3(n10542), .ZN(n10471) );
  NAND2_X1 U7532 ( .A1(n9065), .A2(net80189), .ZN(n8827) );
  NAND2_X1 U7533 ( .A1(n4912), .A2(net80189), .ZN(n8767) );
  INV_X4 U7534 ( .A(n6001), .ZN(n6930) );
  INV_X2 U7535 ( .A(REGFILE_reg_out_4__31_), .ZN(net70757) );
  AOI22_X1 U7536 ( .A1(REGFILE_reg_out_4__31_), .A2(net75451), .B1(
        REGFILE_reg_out_5__31_), .B2(net75452), .ZN(n6236) );
  INV_X1 U7537 ( .A(REGFILE_reg_out_2__31_), .ZN(net70761) );
  AOI22_X1 U7538 ( .A1(REGFILE_reg_out_30__31_), .A2(net84761), .B1(
        REGFILE_reg_out_2__31_), .B2(net75442), .ZN(n6242) );
  INV_X16 U7539 ( .A(net70537), .ZN(net76508) );
  INV_X16 U7540 ( .A(net75419), .ZN(net74051) );
  NAND2_X4 U7541 ( .A1(n5574), .A2(instruction[12]), .ZN(net76242) );
  NOR2_X4 U7542 ( .A1(n6893), .A2(n6892), .ZN(n6894) );
  NOR2_X2 U7543 ( .A1(n8409), .A2(n5820), .ZN(n8404) );
  NAND4_X2 U7544 ( .A1(n6881), .A2(n6880), .A3(n6879), .A4(n6878), .ZN(n6882)
         );
  NAND2_X4 U7545 ( .A1(instruction[11]), .A2(instruction[12]), .ZN(net76211)
         );
  XNOR2_X1 U7546 ( .A(net70921), .B(net77040), .ZN(net70734) );
  NAND2_X1 U7547 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_1__MUX_N1), .A2(net70921), 
        .ZN(n10412) );
  XNOR2_X1 U7548 ( .A(net70921), .B(net71273), .ZN(n10164) );
  NAND2_X1 U7549 ( .A1(n5798), .A2(net71026), .ZN(n10309) );
  NAND2_X1 U7550 ( .A1(net70719), .A2(n5798), .ZN(n9619) );
  NAND2_X1 U7551 ( .A1(net70720), .A2(n5798), .ZN(n9078) );
  NAND2_X1 U7552 ( .A1(n9065), .A2(n5798), .ZN(n8841) );
  NAND2_X1 U7553 ( .A1(n4912), .A2(n5798), .ZN(n8765) );
  INV_X1 U7554 ( .A(n5798), .ZN(n8729) );
  NAND2_X1 U7555 ( .A1(net73708), .A2(n5798), .ZN(n8703) );
  XNOR2_X1 U7556 ( .A(n8585), .B(n5798), .ZN(n8706) );
  AOI22_X4 U7557 ( .A1(n8401), .A2(n6933), .B1(n8403), .B2(n6932), .ZN(
        net75397) );
  NAND3_X4 U7558 ( .A1(net74011), .A2(net73503), .A3(net73170), .ZN(net78055)
         );
  NAND3_X4 U7559 ( .A1(net74011), .A2(net73503), .A3(net73170), .ZN(net78056)
         );
  INV_X32 U7560 ( .A(n6004), .ZN(n6005) );
  INV_X16 U7561 ( .A(n10327), .ZN(n10930) );
  NAND2_X4 U7562 ( .A1(net74009), .A2(instruction[16]), .ZN(net73878) );
  NAND4_X4 U7563 ( .A1(n8572), .A2(n8571), .A3(n8570), .A4(n8569), .ZN(n10494)
         );
  INV_X16 U7564 ( .A(n6005), .ZN(n10099) );
  INV_X16 U7565 ( .A(net78051), .ZN(net71026) );
  INV_X8 U7566 ( .A(n9803), .ZN(n10058) );
  INV_X16 U7567 ( .A(n9094), .ZN(n9065) );
  INV_X8 U7568 ( .A(net70866), .ZN(net70719) );
  NAND2_X4 U7569 ( .A1(n10494), .A2(n10470), .ZN(n10472) );
  INV_X8 U7570 ( .A(net70710), .ZN(n10064) );
  INV_X8 U7571 ( .A(n9606), .ZN(n10066) );
  INV_X8 U7572 ( .A(net70710), .ZN(net71094) );
  INV_X8 U7573 ( .A(n9854), .ZN(net71092) );
  INV_X8 U7574 ( .A(n9012), .ZN(n10280) );
  INV_X32 U7575 ( .A(net75482), .ZN(net77856) );
  INV_X32 U7576 ( .A(net77704), .ZN(net77700) );
  INV_X32 U7577 ( .A(net77656), .ZN(net77650) );
  INV_X32 U7578 ( .A(net77656), .ZN(net77652) );
  INV_X32 U7579 ( .A(n6013), .ZN(n6011) );
  INV_X32 U7580 ( .A(net77548), .ZN(net77544) );
  INV_X32 U7581 ( .A(net77542), .ZN(net77514) );
  INV_X32 U7582 ( .A(net77540), .ZN(net77518) );
  INV_X32 U7583 ( .A(net77540), .ZN(net77520) );
  INV_X32 U7584 ( .A(net77540), .ZN(net77522) );
  INV_X32 U7585 ( .A(net77538), .ZN(net77524) );
  INV_X32 U7586 ( .A(net77538), .ZN(net77526) );
  INV_X32 U7587 ( .A(net77538), .ZN(net77528) );
  INV_X32 U7588 ( .A(net77538), .ZN(net77530) );
  INV_X32 U7589 ( .A(net77548), .ZN(net77532) );
  INV_X32 U7590 ( .A(net77544), .ZN(net77538) );
  INV_X32 U7591 ( .A(net77544), .ZN(net77540) );
  INV_X32 U7592 ( .A(net77502), .ZN(net77488) );
  INV_X32 U7593 ( .A(net77502), .ZN(net77490) );
  INV_X32 U7594 ( .A(net77502), .ZN(net77492) );
  INV_X32 U7595 ( .A(net77508), .ZN(net77500) );
  INV_X32 U7596 ( .A(net77464), .ZN(net77462) );
  INV_X32 U7597 ( .A(net77474), .ZN(net77464) );
  INV_X32 U7598 ( .A(net77428), .ZN(net77426) );
  INV_X32 U7599 ( .A(net77396), .ZN(net77376) );
  INV_X32 U7600 ( .A(net77360), .ZN(net77342) );
  INV_X32 U7601 ( .A(net77358), .ZN(net77344) );
  INV_X32 U7602 ( .A(net77358), .ZN(net77346) );
  INV_X32 U7603 ( .A(net77358), .ZN(net77348) );
  INV_X32 U7604 ( .A(n6018), .ZN(n6015) );
  INV_X32 U7605 ( .A(n6018), .ZN(n6016) );
  INV_X32 U7606 ( .A(n6018), .ZN(n6017) );
  INV_X32 U7607 ( .A(n6014), .ZN(n6018) );
  INV_X32 U7608 ( .A(n6020), .ZN(n6019) );
  INV_X32 U7609 ( .A(n6022), .ZN(n6021) );
  INV_X32 U7610 ( .A(n6028), .ZN(n6027) );
  INV_X32 U7611 ( .A(n6031), .ZN(n6029) );
  INV_X32 U7612 ( .A(n6031), .ZN(n6030) );
  INV_X32 U7613 ( .A(n4964), .ZN(n6032) );
  INV_X32 U7614 ( .A(n6039), .ZN(n6038) );
  INV_X32 U7615 ( .A(n6052), .ZN(n6051) );
  INV_X32 U7616 ( .A(n6061), .ZN(n6059) );
  INV_X32 U7617 ( .A(n6061), .ZN(n6060) );
  INV_X32 U7618 ( .A(n6064), .ZN(n6062) );
  INV_X32 U7619 ( .A(n6064), .ZN(n6063) );
  INV_X32 U7620 ( .A(n6077), .ZN(n6075) );
  INV_X32 U7621 ( .A(n6077), .ZN(n6076) );
  INV_X32 U7622 ( .A(n4965), .ZN(n6087) );
  INV_X32 U7623 ( .A(net77042), .ZN(net77038) );
  INV_X32 U7624 ( .A(net77042), .ZN(net77040) );
  INV_X32 U7625 ( .A(net76514), .ZN(net76510) );
  INV_X32 U7627 ( .A(net76508), .ZN(net76506) );
  INV_X32 U7628 ( .A(n10511), .ZN(n6191) );
  INV_X32 U7629 ( .A(n5012), .ZN(n6221) );
  INV_X32 U7630 ( .A(n5013), .ZN(n6222) );
  INV_X32 U7631 ( .A(n5011), .ZN(n6223) );
  NAND3_X4 U7632 ( .A1(net92447), .A2(net86793), .A3(instruction[13]), .ZN(
        net76259) );
  NAND3_X4 U7633 ( .A1(instruction[15]), .A2(instruction[14]), .A3(
        instruction[13]), .ZN(net76217) );
  NAND3_X4 U7634 ( .A1(net87495), .A2(net82739), .A3(instruction[14]), .ZN(
        net76248) );
  NAND4_X2 U7635 ( .A1(n6228), .A2(n6227), .A3(n6226), .A4(n6225), .ZN(n6234)
         );
  NAND4_X2 U7636 ( .A1(n6232), .A2(n6231), .A3(n6230), .A4(n6229), .ZN(n6233)
         );
  NOR2_X4 U7637 ( .A1(n6234), .A2(n6233), .ZN(n6247) );
  AOI22_X2 U7638 ( .A1(REGFILE_reg_out_31__31_), .A2(net77670), .B1(
        REGFILE_reg_out_3__31_), .B2(n5609), .ZN(n6235) );
  NAND4_X2 U7639 ( .A1(n6238), .A2(n6237), .A3(n6236), .A4(n6235), .ZN(n6245)
         );
  NAND4_X2 U7640 ( .A1(n6243), .A2(n6242), .A3(n6241), .A4(n6240), .ZN(n6244)
         );
  NOR2_X4 U7641 ( .A1(n6245), .A2(n6244), .ZN(n6246) );
  NAND2_X2 U7642 ( .A1(n6247), .A2(n6246), .ZN(dmem_write_out[31]) );
  INV_X4 U7643 ( .A(dmem_write_out[31]), .ZN(n6250) );
  NOR2_X4 U7644 ( .A1(instruction[1]), .A2(instruction[0]), .ZN(n6248) );
  NAND3_X4 U7645 ( .A1(net74011), .A2(net73503), .A3(net73170), .ZN(net73697)
         );
  NAND2_X2 U7646 ( .A1(instruction[31]), .A2(net75844), .ZN(n6249) );
  OAI21_X4 U7647 ( .B1(n6250), .B2(net78055), .A(n6249), .ZN(n10928) );
  AOI22_X2 U7648 ( .A1(REGFILE_reg_out_21__30_), .A2(net77846), .B1(
        REGFILE_reg_out_20__30_), .B2(net77854), .ZN(n6254) );
  AOI22_X2 U7649 ( .A1(REGFILE_reg_out_23__30_), .A2(net77826), .B1(
        REGFILE_reg_out_22__30_), .B2(net77836), .ZN(n6253) );
  NAND4_X2 U7650 ( .A1(n6254), .A2(n6253), .A3(n6252), .A4(n6251), .ZN(n6260)
         );
  AOI22_X2 U7651 ( .A1(REGFILE_reg_out_14__30_), .A2(net77778), .B1(
        REGFILE_reg_out_13__30_), .B2(n6009), .ZN(n6258) );
  NAND4_X2 U7652 ( .A1(n6255), .A2(n6257), .A3(n6256), .A4(n6258), .ZN(n6259)
         );
  AOI22_X2 U7653 ( .A1(n5672), .A2(n5679), .B1(REGFILE_reg_out_5__30_), .B2(
        net84475), .ZN(n6262) );
  NAND4_X2 U7654 ( .A1(n6264), .A2(n6263), .A3(n6262), .A4(n6261), .ZN(n6270)
         );
  NAND4_X2 U7655 ( .A1(n6265), .A2(n6267), .A3(n6266), .A4(n6268), .ZN(n6269)
         );
  NOR2_X4 U7656 ( .A1(n6270), .A2(n6269), .ZN(n6271) );
  NAND2_X2 U7657 ( .A1(n6272), .A2(n6271), .ZN(dmem_write_out[30]) );
  INV_X4 U7658 ( .A(dmem_write_out[30]), .ZN(net76154) );
  NAND4_X2 U7659 ( .A1(n6276), .A2(n6275), .A3(n6274), .A4(n6273), .ZN(n6282)
         );
  AOI22_X2 U7660 ( .A1(REGFILE_reg_out_14__29_), .A2(net77778), .B1(
        REGFILE_reg_out_13__29_), .B2(n5663), .ZN(n6280) );
  NAND4_X2 U7661 ( .A1(n6280), .A2(n6279), .A3(n6278), .A4(n6277), .ZN(n6281)
         );
  NOR2_X4 U7662 ( .A1(n6282), .A2(n6281), .ZN(n6294) );
  NAND4_X2 U7663 ( .A1(n6286), .A2(n6285), .A3(n6284), .A4(n6283), .ZN(n6292)
         );
  NAND4_X2 U7664 ( .A1(n6288), .A2(n6289), .A3(n6290), .A4(n6287), .ZN(n6291)
         );
  NOR2_X4 U7665 ( .A1(n6292), .A2(n6291), .ZN(n6293) );
  NAND2_X2 U7666 ( .A1(n6294), .A2(n6293), .ZN(dmem_write_out[29]) );
  INV_X4 U7667 ( .A(dmem_write_out[29]), .ZN(n6296) );
  NAND2_X2 U7668 ( .A1(net75844), .A2(instruction[29]), .ZN(n6295) );
  AOI22_X2 U7669 ( .A1(REGFILE_reg_out_21__28_), .A2(net77846), .B1(
        REGFILE_reg_out_20__28_), .B2(net77854), .ZN(n6300) );
  AOI22_X2 U7670 ( .A1(REGFILE_reg_out_23__28_), .A2(net77828), .B1(
        REGFILE_reg_out_22__28_), .B2(net77834), .ZN(n6299) );
  NAND4_X2 U7671 ( .A1(n6300), .A2(n6299), .A3(n6298), .A4(n6297), .ZN(n6306)
         );
  NAND4_X2 U7672 ( .A1(n6304), .A2(n6303), .A3(n6302), .A4(n6301), .ZN(n6305)
         );
  NOR2_X4 U7673 ( .A1(n6306), .A2(n6305), .ZN(n6318) );
  AOI22_X2 U7674 ( .A1(REGFILE_reg_out_4__28_), .A2(net75451), .B1(
        REGFILE_reg_out_5__28_), .B2(net84475), .ZN(n6308) );
  AOI22_X2 U7675 ( .A1(REGFILE_reg_out_31__28_), .A2(net77670), .B1(
        REGFILE_reg_out_3__28_), .B2(n5609), .ZN(n6307) );
  NAND4_X2 U7676 ( .A1(n6310), .A2(n6309), .A3(n6308), .A4(n6307), .ZN(n6316)
         );
  NAND4_X2 U7677 ( .A1(n6312), .A2(n6311), .A3(n6314), .A4(n6313), .ZN(n6315)
         );
  NOR2_X4 U7678 ( .A1(n6316), .A2(n6315), .ZN(n6317) );
  NAND2_X2 U7679 ( .A1(n6318), .A2(n6317), .ZN(dmem_write_out[28]) );
  INV_X4 U7680 ( .A(dmem_write_out[28]), .ZN(n6320) );
  NAND2_X2 U7681 ( .A1(net75844), .A2(instruction[28]), .ZN(n6319) );
  OAI21_X4 U7682 ( .B1(n6320), .B2(net78055), .A(n6319), .ZN(n10926) );
  AOI22_X2 U7683 ( .A1(REGFILE_reg_out_21__27_), .A2(net77846), .B1(
        REGFILE_reg_out_20__27_), .B2(net77854), .ZN(n6324) );
  AOI22_X2 U7684 ( .A1(REGFILE_reg_out_23__27_), .A2(net77826), .B1(
        REGFILE_reg_out_22__27_), .B2(net77836), .ZN(n6323) );
  NAND4_X2 U7685 ( .A1(n6324), .A2(n6323), .A3(n6322), .A4(n6321), .ZN(n6330)
         );
  AOI22_X2 U7686 ( .A1(REGFILE_reg_out_14__27_), .A2(net77778), .B1(
        REGFILE_reg_out_13__27_), .B2(n5663), .ZN(n6328) );
  NAND4_X2 U7687 ( .A1(n6328), .A2(n6327), .A3(n6326), .A4(n6325), .ZN(n6329)
         );
  NOR2_X4 U7688 ( .A1(n6330), .A2(n6329), .ZN(n6342) );
  AOI22_X2 U7689 ( .A1(REGFILE_reg_out_9__27_), .A2(net77702), .B1(
        REGFILE_reg_out_8__27_), .B2(n4829), .ZN(n6333) );
  AOI22_X2 U7690 ( .A1(REGFILE_reg_out_4__27_), .A2(n5679), .B1(
        REGFILE_reg_out_5__27_), .B2(net84475), .ZN(n6332) );
  AOI22_X2 U7691 ( .A1(REGFILE_reg_out_31__27_), .A2(net77670), .B1(
        REGFILE_reg_out_3__27_), .B2(n5609), .ZN(n6331) );
  NAND4_X2 U7692 ( .A1(n6334), .A2(n6333), .A3(n6332), .A4(n6331), .ZN(n6340)
         );
  AOI22_X2 U7693 ( .A1(REGFILE_reg_out_24__27_), .A2(net77602), .B1(
        REGFILE_reg_out_25__27_), .B2(net77614), .ZN(n6335) );
  NAND4_X2 U7694 ( .A1(n6335), .A2(n6337), .A3(n6336), .A4(n6338), .ZN(n6339)
         );
  INV_X4 U7695 ( .A(instruction[27]), .ZN(net73696) );
  NAND2_X2 U7696 ( .A1(net75844), .A2(net73696), .ZN(n6343) );
  OAI21_X4 U7697 ( .B1(dmem_write_out[27]), .B2(net78056), .A(n6343), .ZN(
        n8885) );
  AOI22_X2 U7698 ( .A1(REGFILE_reg_out_21__26_), .A2(net77846), .B1(
        REGFILE_reg_out_20__26_), .B2(net77854), .ZN(n6347) );
  AOI22_X2 U7699 ( .A1(REGFILE_reg_out_23__26_), .A2(net77826), .B1(
        REGFILE_reg_out_22__26_), .B2(net77834), .ZN(n6346) );
  NAND4_X2 U7700 ( .A1(n6347), .A2(n6346), .A3(n6345), .A4(n6344), .ZN(n6353)
         );
  AOI22_X2 U7701 ( .A1(REGFILE_reg_out_14__26_), .A2(net77778), .B1(
        REGFILE_reg_out_13__26_), .B2(n5663), .ZN(n6351) );
  NAND4_X2 U7702 ( .A1(n6351), .A2(n6350), .A3(n6349), .A4(n6348), .ZN(n6352)
         );
  NOR2_X4 U7703 ( .A1(n6353), .A2(n6352), .ZN(n6365) );
  AOI22_X2 U7704 ( .A1(REGFILE_reg_out_31__26_), .A2(net77670), .B1(
        REGFILE_reg_out_3__26_), .B2(n5609), .ZN(n6354) );
  NAND4_X2 U7705 ( .A1(n6357), .A2(n6356), .A3(n6355), .A4(n6354), .ZN(n6363)
         );
  NAND4_X2 U7706 ( .A1(n6361), .A2(n6360), .A3(n6359), .A4(n6358), .ZN(n6362)
         );
  NAND2_X2 U7707 ( .A1(n6365), .A2(n6364), .ZN(dmem_write_out[26]) );
  INV_X4 U7708 ( .A(dmem_write_out[26]), .ZN(n6367) );
  NAND2_X2 U7709 ( .A1(net75844), .A2(instruction[26]), .ZN(n6366) );
  OAI21_X4 U7710 ( .B1(n6367), .B2(net73697), .A(n6366), .ZN(n10925) );
  AOI22_X2 U7711 ( .A1(REGFILE_reg_out_21__25_), .A2(net77846), .B1(
        REGFILE_reg_out_20__25_), .B2(net77854), .ZN(n6371) );
  AOI22_X2 U7712 ( .A1(REGFILE_reg_out_23__25_), .A2(net77826), .B1(
        REGFILE_reg_out_22__25_), .B2(net77836), .ZN(n6370) );
  NAND4_X2 U7713 ( .A1(n6371), .A2(n6370), .A3(n6369), .A4(n6368), .ZN(n6377)
         );
  AOI22_X2 U7714 ( .A1(REGFILE_reg_out_14__25_), .A2(net77778), .B1(
        REGFILE_reg_out_13__25_), .B2(n5663), .ZN(n6375) );
  NAND4_X2 U7715 ( .A1(n6372), .A2(n6373), .A3(n6375), .A4(n6374), .ZN(n6376)
         );
  AOI22_X2 U7716 ( .A1(REGFILE_reg_out_4__25_), .A2(n5679), .B1(
        REGFILE_reg_out_5__25_), .B2(net84475), .ZN(n6379) );
  AOI22_X2 U7717 ( .A1(REGFILE_reg_out_31__25_), .A2(net77670), .B1(
        REGFILE_reg_out_3__25_), .B2(n5609), .ZN(n6378) );
  NAND4_X2 U7718 ( .A1(n6380), .A2(n6381), .A3(n6379), .A4(n6378), .ZN(n6387)
         );
  NAND4_X2 U7719 ( .A1(n6384), .A2(n6385), .A3(n6383), .A4(n6382), .ZN(n6386)
         );
  NAND2_X2 U7720 ( .A1(n6389), .A2(n6388), .ZN(dmem_write_out[25]) );
  INV_X4 U7721 ( .A(dmem_write_out[25]), .ZN(n6391) );
  NAND2_X2 U7722 ( .A1(instruction[25]), .A2(net75844), .ZN(n6390) );
  OAI21_X4 U7723 ( .B1(n6391), .B2(net78055), .A(n6390), .ZN(n10924) );
  AOI22_X2 U7724 ( .A1(REGFILE_reg_out_21__24_), .A2(net77846), .B1(
        REGFILE_reg_out_20__24_), .B2(net77854), .ZN(net76031) );
  AOI22_X2 U7725 ( .A1(REGFILE_reg_out_23__24_), .A2(net77826), .B1(
        REGFILE_reg_out_22__24_), .B2(net77836), .ZN(net76032) );
  AOI22_X2 U7726 ( .A1(REGFILE_reg_out_14__24_), .A2(net77778), .B1(
        REGFILE_reg_out_13__24_), .B2(n5663), .ZN(n6395) );
  AOI22_X2 U7727 ( .A1(REGFILE_reg_out_16__24_), .A2(net77764), .B1(
        REGFILE_reg_out_15__24_), .B2(n5579), .ZN(n6394) );
  NOR2_X4 U7728 ( .A1(net76025), .A2(n6396), .ZN(n6408) );
  AOI22_X2 U7729 ( .A1(REGFILE_reg_out_9__24_), .A2(net77702), .B1(
        REGFILE_reg_out_8__24_), .B2(n4829), .ZN(n6399) );
  AOI22_X2 U7730 ( .A1(REGFILE_reg_out_4__24_), .A2(n5678), .B1(
        REGFILE_reg_out_5__24_), .B2(net84475), .ZN(n6398) );
  AOI22_X2 U7731 ( .A1(REGFILE_reg_out_31__24_), .A2(net77670), .B1(
        REGFILE_reg_out_3__24_), .B2(n5609), .ZN(n6397) );
  NAND4_X2 U7732 ( .A1(n6400), .A2(n6399), .A3(n6398), .A4(n6397), .ZN(n6406)
         );
  AOI22_X2 U7733 ( .A1(REGFILE_reg_out_29__24_), .A2(net77650), .B1(
        REGFILE_reg_out_28__24_), .B2(n6911), .ZN(n6404) );
  AOI22_X2 U7734 ( .A1(REGFILE_reg_out_24__24_), .A2(net75437), .B1(
        REGFILE_reg_out_25__24_), .B2(net75438), .ZN(n6401) );
  NAND4_X2 U7735 ( .A1(n6404), .A2(n6403), .A3(n6402), .A4(n6401), .ZN(n6405)
         );
  NAND2_X2 U7736 ( .A1(instruction[24]), .A2(net75844), .ZN(n6409) );
  OAI21_X4 U7737 ( .B1(n6410), .B2(net78056), .A(n6409), .ZN(n10923) );
  AOI22_X2 U7738 ( .A1(REGFILE_reg_out_21__23_), .A2(net77846), .B1(
        REGFILE_reg_out_20__23_), .B2(net77854), .ZN(n6414) );
  AOI22_X2 U7739 ( .A1(REGFILE_reg_out_23__23_), .A2(net77826), .B1(
        REGFILE_reg_out_22__23_), .B2(net77836), .ZN(n6413) );
  AOI22_X2 U7740 ( .A1(REGFILE_reg_out_19__23_), .A2(net77814), .B1(
        REGFILE_reg_out_1__23_), .B2(net82631), .ZN(n6412) );
  NAND4_X2 U7741 ( .A1(n6414), .A2(n6413), .A3(n6412), .A4(n6411), .ZN(n6420)
         );
  AOI22_X2 U7742 ( .A1(REGFILE_reg_out_16__23_), .A2(net87506), .B1(
        REGFILE_reg_out_15__23_), .B2(n5579), .ZN(n6417) );
  NAND4_X2 U7743 ( .A1(n6415), .A2(n6417), .A3(n6416), .A4(n6418), .ZN(n6419)
         );
  AOI22_X2 U7744 ( .A1(REGFILE_reg_out_9__23_), .A2(net77702), .B1(
        REGFILE_reg_out_8__23_), .B2(n4829), .ZN(n6423) );
  AOI22_X2 U7745 ( .A1(REGFILE_reg_out_4__23_), .A2(n5679), .B1(
        REGFILE_reg_out_5__23_), .B2(net84475), .ZN(n6422) );
  AOI22_X2 U7746 ( .A1(REGFILE_reg_out_31__23_), .A2(net77670), .B1(
        REGFILE_reg_out_3__23_), .B2(n5609), .ZN(n6421) );
  NAND4_X2 U7747 ( .A1(n6424), .A2(n6423), .A3(n6422), .A4(n6421), .ZN(n6429)
         );
  AOI22_X2 U7748 ( .A1(REGFILE_reg_out_29__23_), .A2(net77650), .B1(
        REGFILE_reg_out_28__23_), .B2(n6911), .ZN(n6427) );
  NAND2_X2 U7749 ( .A1(instruction[23]), .A2(net75844), .ZN(n6432) );
  OAI21_X4 U7750 ( .B1(n6433), .B2(net73697), .A(n6432), .ZN(n10922) );
  AOI22_X2 U7751 ( .A1(REGFILE_reg_out_21__22_), .A2(net77846), .B1(
        REGFILE_reg_out_20__22_), .B2(net77854), .ZN(n6437) );
  AOI22_X2 U7752 ( .A1(REGFILE_reg_out_23__22_), .A2(net77826), .B1(
        REGFILE_reg_out_22__22_), .B2(net77836), .ZN(n6436) );
  AOI22_X2 U7753 ( .A1(REGFILE_reg_out_19__22_), .A2(net77814), .B1(
        REGFILE_reg_out_1__22_), .B2(net75478), .ZN(n6435) );
  NAND4_X2 U7754 ( .A1(n6437), .A2(n6436), .A3(n6435), .A4(n6434), .ZN(n6443)
         );
  AOI22_X2 U7755 ( .A1(REGFILE_reg_out_14__22_), .A2(net77778), .B1(
        REGFILE_reg_out_13__22_), .B2(n5663), .ZN(n6441) );
  AOI22_X2 U7756 ( .A1(REGFILE_reg_out_7__22_), .A2(net77716), .B1(
        REGFILE_reg_out_6__22_), .B2(net75456), .ZN(n6447) );
  AOI22_X2 U7757 ( .A1(REGFILE_reg_out_9__22_), .A2(net77702), .B1(
        REGFILE_reg_out_8__22_), .B2(n4829), .ZN(n6446) );
  AOI22_X2 U7758 ( .A1(REGFILE_reg_out_4__22_), .A2(n5679), .B1(
        REGFILE_reg_out_5__22_), .B2(net84475), .ZN(n6445) );
  AOI22_X2 U7759 ( .A1(REGFILE_reg_out_31__22_), .A2(net77670), .B1(
        REGFILE_reg_out_3__22_), .B2(n5609), .ZN(n6444) );
  NAND4_X2 U7760 ( .A1(n6447), .A2(n6446), .A3(n6444), .A4(n6445), .ZN(n6453)
         );
  AOI22_X2 U7761 ( .A1(REGFILE_reg_out_29__22_), .A2(net77650), .B1(
        REGFILE_reg_out_28__22_), .B2(n6911), .ZN(n6451) );
  AOI22_X2 U7762 ( .A1(REGFILE_reg_out_30__22_), .A2(net77638), .B1(
        REGFILE_reg_out_2__22_), .B2(net82613), .ZN(n6450) );
  NAND2_X2 U7763 ( .A1(instruction[22]), .A2(net75844), .ZN(n6456) );
  OAI21_X4 U7764 ( .B1(n6457), .B2(net78055), .A(n6456), .ZN(n10921) );
  AOI22_X2 U7765 ( .A1(REGFILE_reg_out_21__21_), .A2(net77844), .B1(
        REGFILE_reg_out_20__21_), .B2(net77852), .ZN(n6461) );
  AOI22_X2 U7766 ( .A1(REGFILE_reg_out_23__21_), .A2(net77828), .B1(
        REGFILE_reg_out_22__21_), .B2(net77836), .ZN(n6460) );
  NAND4_X2 U7767 ( .A1(n6461), .A2(n6460), .A3(n6459), .A4(n6458), .ZN(n6467)
         );
  AOI22_X2 U7768 ( .A1(REGFILE_reg_out_14__21_), .A2(net77780), .B1(
        REGFILE_reg_out_13__21_), .B2(n5663), .ZN(n6465) );
  AOI22_X2 U7769 ( .A1(REGFILE_reg_out_9__21_), .A2(net77700), .B1(
        REGFILE_reg_out_8__21_), .B2(n4829), .ZN(n6470) );
  AOI22_X2 U7770 ( .A1(REGFILE_reg_out_4__21_), .A2(n5679), .B1(
        REGFILE_reg_out_5__21_), .B2(net84475), .ZN(n6469) );
  AOI22_X2 U7771 ( .A1(REGFILE_reg_out_31__21_), .A2(net77668), .B1(
        REGFILE_reg_out_3__21_), .B2(n5609), .ZN(n6468) );
  NAND4_X2 U7772 ( .A1(n6471), .A2(n6470), .A3(n6469), .A4(n6468), .ZN(n6477)
         );
  NAND4_X2 U7773 ( .A1(n6474), .A2(n6473), .A3(n6475), .A4(n6472), .ZN(n6476)
         );
  NAND2_X2 U7774 ( .A1(instruction[21]), .A2(net75844), .ZN(n6480) );
  OAI21_X4 U7775 ( .B1(n6481), .B2(net78056), .A(n6480), .ZN(n10920) );
  AOI22_X2 U7776 ( .A1(REGFILE_reg_out_21__20_), .A2(net77844), .B1(
        REGFILE_reg_out_20__20_), .B2(net77852), .ZN(n6485) );
  AOI22_X2 U7777 ( .A1(REGFILE_reg_out_23__20_), .A2(net77828), .B1(
        REGFILE_reg_out_22__20_), .B2(net77836), .ZN(n6484) );
  AOI22_X2 U7778 ( .A1(REGFILE_reg_out_19__20_), .A2(net77812), .B1(
        REGFILE_reg_out_1__20_), .B2(net75478), .ZN(n6483) );
  NAND4_X2 U7779 ( .A1(n6485), .A2(n6484), .A3(n6483), .A4(n6482), .ZN(n6491)
         );
  AOI22_X2 U7780 ( .A1(REGFILE_reg_out_14__20_), .A2(net77780), .B1(
        REGFILE_reg_out_13__20_), .B2(n5664), .ZN(n6489) );
  AOI22_X2 U7781 ( .A1(REGFILE_reg_out_7__20_), .A2(net77716), .B1(
        REGFILE_reg_out_6__20_), .B2(net75456), .ZN(n6495) );
  AOI22_X2 U7782 ( .A1(REGFILE_reg_out_31__20_), .A2(net77668), .B1(
        REGFILE_reg_out_3__20_), .B2(net77676), .ZN(n6492) );
  AOI22_X2 U7783 ( .A1(REGFILE_reg_out_29__20_), .A2(net77652), .B1(
        REGFILE_reg_out_28__20_), .B2(n5751), .ZN(n6499) );
  NAND2_X2 U7784 ( .A1(net75844), .A2(instruction[20]), .ZN(n6504) );
  OAI21_X4 U7785 ( .B1(n6505), .B2(net73697), .A(n6504), .ZN(n10919) );
  AOI22_X2 U7786 ( .A1(REGFILE_reg_out_21__19_), .A2(net77844), .B1(
        REGFILE_reg_out_20__19_), .B2(net77852), .ZN(n6509) );
  AOI22_X2 U7787 ( .A1(REGFILE_reg_out_23__19_), .A2(net77828), .B1(
        REGFILE_reg_out_22__19_), .B2(net77836), .ZN(n6508) );
  NAND4_X2 U7788 ( .A1(n6509), .A2(n6508), .A3(n6506), .A4(n6507), .ZN(n6515)
         );
  AOI22_X2 U7789 ( .A1(REGFILE_reg_out_14__19_), .A2(net77780), .B1(
        REGFILE_reg_out_13__19_), .B2(n5663), .ZN(n6513) );
  NAND4_X2 U7790 ( .A1(n6513), .A2(n6512), .A3(n6511), .A4(n6510), .ZN(n6514)
         );
  AOI22_X2 U7791 ( .A1(REGFILE_reg_out_9__19_), .A2(net77700), .B1(
        REGFILE_reg_out_8__19_), .B2(net75454), .ZN(n6518) );
  AOI22_X2 U7792 ( .A1(REGFILE_reg_out_4__19_), .A2(n5679), .B1(
        REGFILE_reg_out_5__19_), .B2(net84475), .ZN(n6517) );
  AOI22_X2 U7793 ( .A1(REGFILE_reg_out_31__19_), .A2(net77668), .B1(
        REGFILE_reg_out_3__19_), .B2(net77676), .ZN(n6516) );
  NAND4_X2 U7794 ( .A1(n6519), .A2(n6518), .A3(n6517), .A4(n6516), .ZN(n6525)
         );
  NAND2_X2 U7795 ( .A1(net75844), .A2(instruction[19]), .ZN(n6528) );
  OAI21_X4 U7796 ( .B1(n6529), .B2(net78055), .A(n6528), .ZN(n10918) );
  AOI22_X2 U7797 ( .A1(REGFILE_reg_out_21__18_), .A2(net77844), .B1(
        REGFILE_reg_out_20__18_), .B2(net77852), .ZN(n6533) );
  AOI22_X2 U7798 ( .A1(REGFILE_reg_out_19__18_), .A2(net77812), .B1(
        REGFILE_reg_out_1__18_), .B2(net75478), .ZN(n6531) );
  NAND4_X2 U7799 ( .A1(n6533), .A2(n6532), .A3(n6531), .A4(n6530), .ZN(n6539)
         );
  NAND4_X2 U7800 ( .A1(n6537), .A2(n6535), .A3(n6536), .A4(n6534), .ZN(n6538)
         );
  AOI22_X2 U7801 ( .A1(REGFILE_reg_out_7__18_), .A2(net77714), .B1(
        REGFILE_reg_out_6__18_), .B2(net75456), .ZN(n6543) );
  NAND2_X2 U7802 ( .A1(net75844), .A2(instruction[18]), .ZN(n6552) );
  AOI22_X2 U7803 ( .A1(REGFILE_reg_out_21__17_), .A2(net77844), .B1(
        REGFILE_reg_out_20__17_), .B2(net77852), .ZN(n6557) );
  NAND2_X2 U7804 ( .A1(net75844), .A2(instruction[17]), .ZN(net75843) );
  AOI22_X2 U7805 ( .A1(REGFILE_reg_out_21__16_), .A2(net77844), .B1(
        REGFILE_reg_out_20__16_), .B2(net77852), .ZN(n6565) );
  AOI22_X2 U7806 ( .A1(REGFILE_reg_out_23__16_), .A2(net77828), .B1(
        REGFILE_reg_out_22__16_), .B2(net77836), .ZN(n6564) );
  NAND4_X2 U7807 ( .A1(n6565), .A2(n6564), .A3(n6563), .A4(n6562), .ZN(n6571)
         );
  NAND4_X2 U7808 ( .A1(n6568), .A2(n6567), .A3(n6569), .A4(n6566), .ZN(n6570)
         );
  AOI22_X2 U7809 ( .A1(REGFILE_reg_out_30__16_), .A2(net77638), .B1(
        REGFILE_reg_out_2__16_), .B2(net82613), .ZN(n6578) );
  NAND4_X2 U7810 ( .A1(n6578), .A2(n6579), .A3(n6577), .A4(n6576), .ZN(n6580)
         );
  AOI22_X2 U7811 ( .A1(REGFILE_reg_out_21__15_), .A2(net77844), .B1(
        REGFILE_reg_out_20__15_), .B2(net77852), .ZN(n6587) );
  NAND4_X2 U7812 ( .A1(n6587), .A2(n6585), .A3(n6586), .A4(n6584), .ZN(n6593)
         );
  NOR2_X4 U7813 ( .A1(n6593), .A2(n6592), .ZN(n6605) );
  NAND4_X2 U7814 ( .A1(n6597), .A2(n6596), .A3(n6595), .A4(n6594), .ZN(n6603)
         );
  NAND4_X2 U7815 ( .A1(n6601), .A2(n6600), .A3(n6598), .A4(n6599), .ZN(n6602)
         );
  NOR2_X4 U7816 ( .A1(n6603), .A2(n6602), .ZN(n6604) );
  INV_X4 U7817 ( .A(instruction[0]), .ZN(net73499) );
  NAND2_X2 U7818 ( .A1(instruction[2]), .A2(net73499), .ZN(n6606) );
  INV_X4 U7819 ( .A(n6606), .ZN(n8539) );
  NOR2_X4 U7820 ( .A1(instruction[3]), .A2(instruction[0]), .ZN(n6607) );
  OAI21_X4 U7821 ( .B1(dmem_write_out[15]), .B2(net75427), .A(net78042), .ZN(
        n10288) );
  NAND4_X2 U7822 ( .A1(n6609), .A2(n6610), .A3(n6611), .A4(n6608), .ZN(n6617)
         );
  NAND4_X2 U7823 ( .A1(n6612), .A2(n6615), .A3(n6613), .A4(n6614), .ZN(n6616)
         );
  NOR2_X4 U7824 ( .A1(n6617), .A2(n6616), .ZN(n6629) );
  NAND4_X2 U7825 ( .A1(n6621), .A2(n6620), .A3(n6618), .A4(n6619), .ZN(n6627)
         );
  NOR2_X4 U7826 ( .A1(n6627), .A2(n6626), .ZN(n6628) );
  OAI21_X4 U7827 ( .B1(dmem_write_out[14]), .B2(net75427), .A(net78042), .ZN(
        n10364) );
  NOR2_X4 U7828 ( .A1(n6643), .A2(n6642), .ZN(net75748) );
  AOI22_X2 U7829 ( .A1(REGFILE_reg_out_21__12_), .A2(net77844), .B1(
        REGFILE_reg_out_20__12_), .B2(net77852), .ZN(n6647) );
  AOI22_X2 U7830 ( .A1(REGFILE_reg_out_23__12_), .A2(net77828), .B1(
        REGFILE_reg_out_22__12_), .B2(net77836), .ZN(n6646) );
  NAND4_X2 U7831 ( .A1(n6647), .A2(n6646), .A3(n6645), .A4(n6644), .ZN(n6653)
         );
  AOI22_X2 U7832 ( .A1(REGFILE_reg_out_14__12_), .A2(net77780), .B1(
        REGFILE_reg_out_13__12_), .B2(n5664), .ZN(n6651) );
  AOI22_X2 U7833 ( .A1(REGFILE_reg_out_0__12_), .A2(net82342), .B1(n5674), 
        .B2(net83203), .ZN(n6648) );
  NAND4_X2 U7834 ( .A1(n6651), .A2(n6650), .A3(n6649), .A4(n6648), .ZN(n6652)
         );
  NOR2_X4 U7835 ( .A1(n6653), .A2(n6652), .ZN(n6665) );
  AOI22_X2 U7836 ( .A1(REGFILE_reg_out_7__12_), .A2(net77714), .B1(
        REGFILE_reg_out_6__12_), .B2(net75456), .ZN(n6657) );
  AOI22_X2 U7837 ( .A1(REGFILE_reg_out_9__12_), .A2(net77700), .B1(
        REGFILE_reg_out_8__12_), .B2(net75454), .ZN(n6656) );
  NAND4_X2 U7838 ( .A1(n6657), .A2(n6656), .A3(n6655), .A4(n6654), .ZN(n6663)
         );
  AOI22_X2 U7839 ( .A1(REGFILE_reg_out_29__12_), .A2(net77652), .B1(
        REGFILE_reg_out_28__12_), .B2(n6911), .ZN(n6661) );
  NOR2_X4 U7840 ( .A1(n6663), .A2(n6662), .ZN(n6664) );
  OAI21_X4 U7841 ( .B1(dmem_write_out[12]), .B2(net75427), .A(net78042), .ZN(
        n10371) );
  AOI22_X2 U7842 ( .A1(REGFILE_reg_out_21__11_), .A2(net77844), .B1(
        REGFILE_reg_out_20__11_), .B2(net77852), .ZN(n6669) );
  NAND4_X2 U7843 ( .A1(n6669), .A2(n6666), .A3(n6667), .A4(n6668), .ZN(n6675)
         );
  NOR2_X4 U7844 ( .A1(n6675), .A2(n6674), .ZN(n6687) );
  AOI22_X2 U7845 ( .A1(REGFILE_reg_out_7__11_), .A2(net77716), .B1(
        REGFILE_reg_out_6__11_), .B2(net75456), .ZN(n6679) );
  AOI22_X2 U7846 ( .A1(REGFILE_reg_out_9__11_), .A2(net77700), .B1(
        REGFILE_reg_out_8__11_), .B2(net75454), .ZN(n6678) );
  NAND4_X2 U7847 ( .A1(n6679), .A2(n6678), .A3(n6677), .A4(n6676), .ZN(n6685)
         );
  NAND4_X2 U7848 ( .A1(n6683), .A2(n6682), .A3(n6681), .A4(n6680), .ZN(n6684)
         );
  NOR2_X4 U7849 ( .A1(n6685), .A2(n6684), .ZN(n6686) );
  OAI21_X4 U7850 ( .B1(dmem_write_out[11]), .B2(net75427), .A(net78042), .ZN(
        n9835) );
  AOI22_X2 U7851 ( .A1(REGFILE_reg_out_21__10_), .A2(net77842), .B1(
        REGFILE_reg_out_20__10_), .B2(net77850), .ZN(n6691) );
  NAND4_X2 U7852 ( .A1(n6691), .A2(n6690), .A3(n6689), .A4(n6688), .ZN(n6697)
         );
  NAND4_X2 U7853 ( .A1(n6695), .A2(n6694), .A3(n6693), .A4(n6692), .ZN(n6696)
         );
  NOR2_X4 U7854 ( .A1(n6697), .A2(n6696), .ZN(n6709) );
  NAND4_X2 U7855 ( .A1(n6701), .A2(n6700), .A3(n6699), .A4(n6698), .ZN(n6707)
         );
  NAND4_X2 U7856 ( .A1(n6705), .A2(n6702), .A3(n6704), .A4(n6703), .ZN(n6706)
         );
  NOR2_X4 U7857 ( .A1(n6706), .A2(n6707), .ZN(n6708) );
  OAI21_X4 U7858 ( .B1(dmem_write_out[10]), .B2(net75427), .A(net78042), .ZN(
        n10378) );
  AOI22_X2 U7859 ( .A1(REGFILE_reg_out_21__9_), .A2(net77842), .B1(
        REGFILE_reg_out_20__9_), .B2(net77850), .ZN(n6713) );
  AOI22_X2 U7860 ( .A1(REGFILE_reg_out_23__9_), .A2(net77826), .B1(
        REGFILE_reg_out_22__9_), .B2(net77834), .ZN(n6712) );
  NAND4_X2 U7861 ( .A1(n6713), .A2(n6712), .A3(n6711), .A4(n6710), .ZN(n6719)
         );
  AOI22_X2 U7862 ( .A1(REGFILE_reg_out_14__9_), .A2(net77778), .B1(
        REGFILE_reg_out_13__9_), .B2(n5664), .ZN(n6717) );
  NAND4_X2 U7863 ( .A1(n6717), .A2(n6716), .A3(n6715), .A4(n6714), .ZN(n6718)
         );
  AOI22_X2 U7864 ( .A1(REGFILE_reg_out_7__9_), .A2(net75455), .B1(
        REGFILE_reg_out_6__9_), .B2(net75456), .ZN(n6723) );
  AOI22_X2 U7865 ( .A1(REGFILE_reg_out_9__9_), .A2(net77698), .B1(
        REGFILE_reg_out_8__9_), .B2(n4829), .ZN(n6722) );
  NAND4_X2 U7866 ( .A1(n6723), .A2(n6722), .A3(n6721), .A4(n6720), .ZN(n6729)
         );
  AOI22_X2 U7867 ( .A1(REGFILE_reg_out_26__9_), .A2(net75439), .B1(
        REGFILE_reg_out_27__9_), .B2(net89184), .ZN(n6725) );
  NAND4_X2 U7868 ( .A1(n6727), .A2(n6725), .A3(n6726), .A4(n6724), .ZN(n6728)
         );
  OAI21_X4 U7869 ( .B1(dmem_write_out[9]), .B2(net75427), .A(n10945), .ZN(
        n9358) );
  AOI22_X2 U7870 ( .A1(REGFILE_reg_out_23__8_), .A2(net77826), .B1(
        REGFILE_reg_out_22__8_), .B2(net77834), .ZN(n6734) );
  NAND4_X2 U7871 ( .A1(n6733), .A2(n6734), .A3(n6735), .A4(n6732), .ZN(n6741)
         );
  NAND4_X2 U7872 ( .A1(n6739), .A2(n6738), .A3(n6737), .A4(n6736), .ZN(n6740)
         );
  NOR2_X4 U7873 ( .A1(n6741), .A2(n6740), .ZN(n6753) );
  NAND4_X2 U7874 ( .A1(n6745), .A2(n6744), .A3(n6743), .A4(n6742), .ZN(n6751)
         );
  NAND4_X2 U7875 ( .A1(n6749), .A2(n6748), .A3(n6746), .A4(n6747), .ZN(n6750)
         );
  OAI21_X4 U7876 ( .B1(dmem_write_out[8]), .B2(net75427), .A(net78042), .ZN(
        n10385) );
  AOI22_X2 U7877 ( .A1(REGFILE_reg_out_21__7_), .A2(net77842), .B1(
        REGFILE_reg_out_20__7_), .B2(net77850), .ZN(n6757) );
  AOI22_X2 U7878 ( .A1(REGFILE_reg_out_23__7_), .A2(net77826), .B1(
        REGFILE_reg_out_22__7_), .B2(net77834), .ZN(n6756) );
  AOI22_X2 U7879 ( .A1(REGFILE_reg_out_19__7_), .A2(net77810), .B1(
        REGFILE_reg_out_1__7_), .B2(net75478), .ZN(n6755) );
  NAND4_X2 U7880 ( .A1(n6757), .A2(n6756), .A3(n6755), .A4(n6754), .ZN(n6763)
         );
  AOI22_X2 U7881 ( .A1(REGFILE_reg_out_14__7_), .A2(net77778), .B1(
        REGFILE_reg_out_13__7_), .B2(n5664), .ZN(n6761) );
  NAND4_X2 U7882 ( .A1(n6759), .A2(n6760), .A3(n6761), .A4(n6758), .ZN(n6762)
         );
  AOI22_X2 U7883 ( .A1(REGFILE_reg_out_29__7_), .A2(net77650), .B1(
        REGFILE_reg_out_28__7_), .B2(n5751), .ZN(net75619) );
  AOI22_X2 U7884 ( .A1(REGFILE_reg_out_21__6_), .A2(net77842), .B1(
        REGFILE_reg_out_20__6_), .B2(net77850), .ZN(n6767) );
  AOI22_X2 U7885 ( .A1(REGFILE_reg_out_19__6_), .A2(net77810), .B1(
        REGFILE_reg_out_1__6_), .B2(net75478), .ZN(n6765) );
  NAND4_X2 U7886 ( .A1(n6767), .A2(n6766), .A3(n6765), .A4(n6764), .ZN(n6773)
         );
  AOI22_X2 U7887 ( .A1(REGFILE_reg_out_14__6_), .A2(net77778), .B1(
        REGFILE_reg_out_13__6_), .B2(n6009), .ZN(n6771) );
  NAND4_X2 U7888 ( .A1(n6770), .A2(n6771), .A3(n6769), .A4(n6768), .ZN(n6772)
         );
  NOR2_X4 U7889 ( .A1(n6772), .A2(n6773), .ZN(n6785) );
  AOI22_X2 U7890 ( .A1(REGFILE_reg_out_9__6_), .A2(net77698), .B1(
        REGFILE_reg_out_8__6_), .B2(n4829), .ZN(n6776) );
  NAND4_X2 U7891 ( .A1(n6777), .A2(n6776), .A3(n6775), .A4(n6774), .ZN(n6783)
         );
  AOI22_X2 U7892 ( .A1(REGFILE_reg_out_29__6_), .A2(net77650), .B1(
        REGFILE_reg_out_28__6_), .B2(n6911), .ZN(n6781) );
  NAND4_X2 U7893 ( .A1(n6780), .A2(n6781), .A3(n6779), .A4(n6778), .ZN(n6782)
         );
  NOR2_X4 U7894 ( .A1(n6783), .A2(n6782), .ZN(n6784) );
  OAI21_X4 U7895 ( .B1(dmem_write_out[6]), .B2(net75427), .A(n10945), .ZN(
        n10392) );
  AOI22_X2 U7896 ( .A1(REGFILE_reg_out_21__5_), .A2(net77842), .B1(
        REGFILE_reg_out_20__5_), .B2(net77850), .ZN(n6789) );
  NAND4_X2 U7897 ( .A1(n6789), .A2(n6788), .A3(n6787), .A4(n6786), .ZN(n6795)
         );
  AOI22_X2 U7898 ( .A1(REGFILE_reg_out_14__5_), .A2(net77778), .B1(
        REGFILE_reg_out_13__5_), .B2(n6009), .ZN(n6793) );
  NAND4_X2 U7899 ( .A1(n6790), .A2(n6792), .A3(n6791), .A4(n6793), .ZN(n6794)
         );
  AOI22_X2 U7900 ( .A1(REGFILE_reg_out_9__5_), .A2(net77698), .B1(
        REGFILE_reg_out_8__5_), .B2(n4829), .ZN(n6798) );
  NAND4_X2 U7901 ( .A1(n6799), .A2(n6798), .A3(n6797), .A4(n6796), .ZN(n6805)
         );
  AOI22_X2 U7902 ( .A1(REGFILE_reg_out_29__5_), .A2(net77650), .B1(
        REGFILE_reg_out_28__5_), .B2(n6911), .ZN(n6803) );
  NAND4_X2 U7903 ( .A1(n6803), .A2(n6802), .A3(n6801), .A4(n6800), .ZN(n6804)
         );
  OAI21_X4 U7904 ( .B1(dmem_write_out[5]), .B2(net75427), .A(n10945), .ZN(
        n9616) );
  AOI22_X2 U7905 ( .A1(REGFILE_reg_out_21__4_), .A2(net77842), .B1(
        REGFILE_reg_out_20__4_), .B2(net77850), .ZN(n6811) );
  NAND4_X2 U7906 ( .A1(n6811), .A2(n6810), .A3(n6809), .A4(n6808), .ZN(n6817)
         );
  NAND4_X2 U7907 ( .A1(n6815), .A2(n6812), .A3(n6813), .A4(n6814), .ZN(n6816)
         );
  AOI22_X2 U7908 ( .A1(REGFILE_reg_out_9__4_), .A2(net77698), .B1(
        REGFILE_reg_out_8__4_), .B2(n4829), .ZN(n6820) );
  NAND4_X2 U7909 ( .A1(n6821), .A2(n6820), .A3(n6819), .A4(n6818), .ZN(n6827)
         );
  AOI22_X2 U7910 ( .A1(REGFILE_reg_out_29__4_), .A2(net77650), .B1(
        REGFILE_reg_out_28__4_), .B2(n6911), .ZN(n6825) );
  NAND4_X2 U7911 ( .A1(n6824), .A2(n6825), .A3(n6823), .A4(n6822), .ZN(n6826)
         );
  AOI22_X2 U7912 ( .A1(REGFILE_reg_out_21__3_), .A2(net77842), .B1(
        REGFILE_reg_out_20__3_), .B2(net77850), .ZN(n6833) );
  NAND4_X2 U7913 ( .A1(n6833), .A2(n6832), .A3(n6830), .A4(n6831), .ZN(n6839)
         );
  NAND4_X2 U7914 ( .A1(n6836), .A2(n6834), .A3(n6835), .A4(n6837), .ZN(n6838)
         );
  NAND4_X2 U7915 ( .A1(n6840), .A2(n6842), .A3(n6841), .A4(n6843), .ZN(n6849)
         );
  NAND4_X2 U7916 ( .A1(n6847), .A2(n6846), .A3(n6845), .A4(n6844), .ZN(n6848)
         );
  OAI21_X4 U7917 ( .B1(dmem_write_out[3]), .B2(net75427), .A(n10945), .ZN(
        n10036) );
  AOI22_X2 U7918 ( .A1(REGFILE_reg_out_23__2_), .A2(net77826), .B1(
        REGFILE_reg_out_22__2_), .B2(net77834), .ZN(n6854) );
  NAND4_X2 U7919 ( .A1(n6853), .A2(n6854), .A3(n6855), .A4(n6852), .ZN(n6861)
         );
  NAND4_X2 U7920 ( .A1(n6859), .A2(n6858), .A3(n6857), .A4(n6856), .ZN(n6860)
         );
  NOR2_X4 U7921 ( .A1(n6861), .A2(n6860), .ZN(n6873) );
  NAND4_X2 U7922 ( .A1(n6862), .A2(n6864), .A3(n6863), .A4(n6865), .ZN(n6871)
         );
  AOI22_X2 U7923 ( .A1(REGFILE_reg_out_29__2_), .A2(net77650), .B1(
        REGFILE_reg_out_28__2_), .B2(n6911), .ZN(n6869) );
  NOR2_X4 U7924 ( .A1(n6871), .A2(n6870), .ZN(n6872) );
  OAI21_X4 U7925 ( .B1(dmem_write_out[2]), .B2(net75427), .A(n10945), .ZN(
        n10408) );
  AOI22_X2 U7926 ( .A1(REGFILE_reg_out_21__1_), .A2(net77842), .B1(
        REGFILE_reg_out_20__1_), .B2(net77850), .ZN(n6877) );
  AOI22_X2 U7927 ( .A1(REGFILE_reg_out_23__1_), .A2(net77826), .B1(
        REGFILE_reg_out_22__1_), .B2(net77834), .ZN(n6876) );
  NAND4_X2 U7928 ( .A1(n6877), .A2(n6876), .A3(n6875), .A4(n6874), .ZN(n6883)
         );
  NAND4_X2 U7929 ( .A1(n6884), .A2(n6886), .A3(n6885), .A4(n6887), .ZN(n6893)
         );
  AOI22_X2 U7930 ( .A1(REGFILE_reg_out_21__0_), .A2(net77842), .B1(
        REGFILE_reg_out_20__0_), .B2(net77850), .ZN(n6900) );
  NAND4_X2 U7931 ( .A1(n6900), .A2(n6899), .A3(n6898), .A4(n6897), .ZN(n6906)
         );
  NAND4_X2 U7932 ( .A1(n6901), .A2(n6903), .A3(n6902), .A4(n6904), .ZN(n6905)
         );
  NOR2_X4 U7933 ( .A1(n6906), .A2(n6905), .ZN(n6919) );
  NAND4_X2 U7934 ( .A1(n6910), .A2(n6909), .A3(n6908), .A4(n6907), .ZN(n6917)
         );
  NAND4_X2 U7935 ( .A1(n6915), .A2(n6914), .A3(n6913), .A4(n6912), .ZN(n6916)
         );
  NOR2_X4 U7936 ( .A1(n6917), .A2(n6916), .ZN(n6918) );
  NAND2_X2 U7937 ( .A1(n6919), .A2(n6918), .ZN(dmem_write_out[0]) );
  INV_X4 U7938 ( .A(instruction[7]), .ZN(n8295) );
  INV_X4 U7939 ( .A(instruction[6]), .ZN(n8287) );
  NAND2_X2 U7940 ( .A1(n8295), .A2(n8287), .ZN(net73842) );
  NAND3_X4 U7941 ( .A1(instruction[10]), .A2(instruction[8]), .A3(
        instruction[9]), .ZN(net75425) );
  NAND3_X4 U7942 ( .A1(instruction[8]), .A2(net73987), .A3(instruction[9]), 
        .ZN(net75424) );
  NAND3_X4 U7943 ( .A1(net90864), .A2(net73987), .A3(instruction[9]), .ZN(
        n6920) );
  NAND3_X4 U7944 ( .A1(net123932), .A2(net87098), .A3(instruction[10]), .ZN(
        net75419) );
  NAND3_X4 U7945 ( .A1(net73987), .A2(net87098), .A3(net73879), .ZN(net75418)
         );
  NAND2_X2 U7946 ( .A1(instruction[6]), .A2(n8295), .ZN(net73836) );
  NAND2_X2 U7947 ( .A1(instruction[7]), .A2(n8287), .ZN(n8407) );
  INV_X4 U7948 ( .A(n8407), .ZN(n8402) );
  NAND2_X2 U7949 ( .A1(n8402), .A2(net77272), .ZN(n6951) );
  INV_X4 U7950 ( .A(n6951), .ZN(n6933) );
  NAND2_X2 U7951 ( .A1(instruction[7]), .A2(instruction[6]), .ZN(n8409) );
  NOR2_X4 U7952 ( .A1(n6954), .A2(n6953), .ZN(n6955) );
  NAND2_X2 U7953 ( .A1(REGFILE_reg_out_2__29_), .A2(net77336), .ZN(n6959) );
  NAND2_X2 U7954 ( .A1(REGFILE_reg_out_3__29_), .A2(net77406), .ZN(n6958) );
  NAND2_X2 U7955 ( .A1(REGFILE_reg_out_0__29_), .A2(net77300), .ZN(n6957) );
  NAND2_X2 U7956 ( .A1(REGFILE_reg_out_7__29_), .A2(net77480), .ZN(n6962) );
  NAND2_X2 U7957 ( .A1(REGFILE_reg_out_12__29_), .A2(net77388), .ZN(n6969) );
  NAND2_X2 U7958 ( .A1(REGFILE_reg_out_13__29_), .A2(net77462), .ZN(n6968) );
  NAND2_X2 U7959 ( .A1(REGFILE_reg_out_10__29_), .A2(n6017), .ZN(n6967) );
  NAND2_X2 U7960 ( .A1(REGFILE_reg_out_11__29_), .A2(net77426), .ZN(n6966) );
  NAND2_X2 U7961 ( .A1(REGFILE_reg_out_18__29_), .A2(n6017), .ZN(n6979) );
  NAND2_X2 U7962 ( .A1(REGFILE_reg_out_19__29_), .A2(net77426), .ZN(n6978) );
  NAND2_X2 U7963 ( .A1(REGFILE_reg_out_16__29_), .A2(net77318), .ZN(n6977) );
  NAND4_X2 U7964 ( .A1(n6979), .A2(n6978), .A3(n6977), .A4(n6976), .ZN(n6983)
         );
  NAND2_X2 U7965 ( .A1(REGFILE_reg_out_26__29_), .A2(n6017), .ZN(n6987) );
  NAND2_X2 U7966 ( .A1(REGFILE_reg_out_30__29_), .A2(net77550), .ZN(n6991) );
  NAND2_X2 U7967 ( .A1(n5986), .A2(net77400), .ZN(n6989) );
  NAND2_X2 U7968 ( .A1(net77478), .A2(REGFILE_reg_out_31__28_), .ZN(n6999) );
  NAND2_X2 U7969 ( .A1(net77456), .A2(REGFILE_reg_out_29__28_), .ZN(n6998) );
  NAND4_X2 U7970 ( .A1(n7001), .A2(n7000), .A3(n6999), .A4(n6998), .ZN(n7007)
         );
  NAND2_X2 U7971 ( .A1(net77388), .A2(REGFILE_reg_out_28__28_), .ZN(n7004) );
  NAND2_X2 U7972 ( .A1(n6014), .A2(REGFILE_reg_out_26__28_), .ZN(n7003) );
  NAND4_X2 U7973 ( .A1(n7005), .A2(n7004), .A3(n7003), .A4(n7002), .ZN(n7006)
         );
  NAND2_X2 U7974 ( .A1(net77478), .A2(REGFILE_reg_out_23__28_), .ZN(n7009) );
  NAND2_X2 U7975 ( .A1(net77388), .A2(REGFILE_reg_out_20__28_), .ZN(n7014) );
  NAND2_X2 U7976 ( .A1(n6014), .A2(REGFILE_reg_out_18__28_), .ZN(n7013) );
  NAND4_X2 U7977 ( .A1(n7015), .A2(n7014), .A3(n7013), .A4(n7012), .ZN(n7016)
         );
  OAI21_X4 U7978 ( .B1(n7017), .B2(n7016), .A(net77588), .ZN(n7040) );
  NAND2_X2 U7979 ( .A1(net77516), .A2(REGFILE_reg_out_9__28_), .ZN(n7020) );
  NAND2_X2 U7980 ( .A1(net77480), .A2(REGFILE_reg_out_15__28_), .ZN(n7019) );
  NAND4_X2 U7981 ( .A1(n7021), .A2(n7020), .A3(n7019), .A4(n7018), .ZN(n7027)
         );
  NAND2_X2 U7982 ( .A1(net77422), .A2(REGFILE_reg_out_11__28_), .ZN(n7025) );
  NAND2_X2 U7983 ( .A1(net77336), .A2(REGFILE_reg_out_10__28_), .ZN(n7023) );
  NAND2_X2 U7984 ( .A1(net77300), .A2(REGFILE_reg_out_8__28_), .ZN(n7022) );
  NAND4_X2 U7985 ( .A1(n7025), .A2(n7024), .A3(n7023), .A4(n7022), .ZN(n7026)
         );
  NAND2_X2 U7986 ( .A1(net77514), .A2(REGFILE_reg_out_1__28_), .ZN(n7030) );
  NAND4_X2 U7987 ( .A1(n7031), .A2(n7030), .A3(n7029), .A4(n7028), .ZN(n7037)
         );
  NAND2_X2 U7988 ( .A1(net77388), .A2(REGFILE_reg_out_4__28_), .ZN(n7034) );
  NAND2_X2 U7989 ( .A1(n6014), .A2(REGFILE_reg_out_2__28_), .ZN(n7033) );
  NAND4_X2 U7990 ( .A1(n7035), .A2(n7034), .A3(n7033), .A4(n7032), .ZN(n7036)
         );
  NAND2_X2 U7991 ( .A1(net77516), .A2(REGFILE_reg_out_25__27_), .ZN(n7044) );
  NAND2_X2 U7992 ( .A1(net77480), .A2(REGFILE_reg_out_31__27_), .ZN(n7043) );
  NAND4_X2 U7993 ( .A1(n7045), .A2(n7044), .A3(n7043), .A4(n7042), .ZN(n7051)
         );
  NAND2_X2 U7994 ( .A1(net77414), .A2(REGFILE_reg_out_27__27_), .ZN(n7049) );
  NAND2_X2 U7995 ( .A1(net77336), .A2(REGFILE_reg_out_26__27_), .ZN(n7047) );
  NAND2_X2 U7996 ( .A1(net77300), .A2(REGFILE_reg_out_24__27_), .ZN(n7046) );
  NAND4_X2 U7997 ( .A1(n7049), .A2(n7048), .A3(n7047), .A4(n7046), .ZN(n7050)
         );
  OAI21_X4 U7998 ( .B1(n7051), .B2(n7050), .A(n6012), .ZN(n7085) );
  NAND2_X2 U7999 ( .A1(net77478), .A2(REGFILE_reg_out_23__27_), .ZN(n7053) );
  NAND2_X2 U8000 ( .A1(net77456), .A2(REGFILE_reg_out_21__27_), .ZN(n7052) );
  NAND4_X2 U8001 ( .A1(n7055), .A2(n7054), .A3(n7053), .A4(n7052), .ZN(n7061)
         );
  NAND2_X2 U8003 ( .A1(n6014), .A2(REGFILE_reg_out_18__27_), .ZN(n7057) );
  NAND4_X2 U8004 ( .A1(n7059), .A2(n7058), .A3(n7057), .A4(n7056), .ZN(n7060)
         );
  OAI21_X4 U8005 ( .B1(n7061), .B2(n7060), .A(net77588), .ZN(n7084) );
  NAND2_X2 U8006 ( .A1(net77516), .A2(REGFILE_reg_out_9__27_), .ZN(n7064) );
  NAND2_X2 U8007 ( .A1(net77480), .A2(REGFILE_reg_out_15__27_), .ZN(n7063) );
  NAND4_X2 U8008 ( .A1(n7065), .A2(n7064), .A3(n7063), .A4(n7062), .ZN(n7071)
         );
  NAND2_X2 U8009 ( .A1(net77420), .A2(REGFILE_reg_out_11__27_), .ZN(n7069) );
  NAND2_X2 U8010 ( .A1(net77336), .A2(REGFILE_reg_out_10__27_), .ZN(n7067) );
  NAND2_X2 U8011 ( .A1(net77300), .A2(REGFILE_reg_out_8__27_), .ZN(n7066) );
  NAND4_X2 U8012 ( .A1(n7069), .A2(n7068), .A3(n7067), .A4(n7066), .ZN(n7070)
         );
  OAI21_X4 U8013 ( .B1(n7071), .B2(n7070), .A(n6019), .ZN(n7083) );
  NAND2_X2 U8014 ( .A1(net77516), .A2(REGFILE_reg_out_1__27_), .ZN(n7074) );
  NAND2_X2 U8015 ( .A1(net77480), .A2(REGFILE_reg_out_7__27_), .ZN(n7073) );
  NAND4_X2 U8016 ( .A1(n7075), .A2(n7074), .A3(n7073), .A4(n7072), .ZN(n7081)
         );
  NAND2_X2 U8017 ( .A1(net77418), .A2(REGFILE_reg_out_3__27_), .ZN(n7079) );
  NAND2_X2 U8018 ( .A1(net77336), .A2(REGFILE_reg_out_2__27_), .ZN(n7077) );
  NAND4_X2 U8020 ( .A1(n7079), .A2(n7078), .A3(n7077), .A4(n7076), .ZN(n7080)
         );
  OAI21_X4 U8021 ( .B1(n7081), .B2(n7080), .A(net77292), .ZN(n7082) );
  MUX2_X2 U8022 ( .A(n8450), .B(instruction[27]), .S(net77276), .Z(aluA[27])
         );
  NAND2_X2 U8023 ( .A1(REGFILE_reg_out_30__26_), .A2(net77564), .ZN(n7089) );
  NAND2_X2 U8024 ( .A1(REGFILE_reg_out_31__26_), .A2(net77498), .ZN(n7087) );
  NAND2_X2 U8025 ( .A1(REGFILE_reg_out_29__26_), .A2(net77462), .ZN(n7086) );
  NAND4_X2 U8026 ( .A1(n7089), .A2(n7088), .A3(n7087), .A4(n7086), .ZN(n7095)
         );
  NAND2_X2 U8027 ( .A1(REGFILE_reg_out_27__26_), .A2(net77426), .ZN(n7093) );
  NAND2_X2 U8028 ( .A1(REGFILE_reg_out_28__26_), .A2(net77376), .ZN(n7092) );
  NAND2_X2 U8029 ( .A1(REGFILE_reg_out_26__26_), .A2(n6017), .ZN(n7091) );
  NAND2_X2 U8030 ( .A1(REGFILE_reg_out_24__26_), .A2(net77318), .ZN(n7090) );
  NAND4_X2 U8031 ( .A1(n7093), .A2(n7092), .A3(n7091), .A4(n7090), .ZN(n7094)
         );
  NAND2_X2 U8032 ( .A1(REGFILE_reg_out_22__26_), .A2(net77566), .ZN(n7099) );
  NAND2_X2 U8033 ( .A1(REGFILE_reg_out_23__26_), .A2(net77498), .ZN(n7097) );
  NAND2_X2 U8034 ( .A1(REGFILE_reg_out_21__26_), .A2(net77462), .ZN(n7096) );
  NAND4_X2 U8035 ( .A1(n7099), .A2(n7098), .A3(n7097), .A4(n7096), .ZN(n7105)
         );
  NAND2_X2 U8036 ( .A1(REGFILE_reg_out_19__26_), .A2(net77426), .ZN(n7103) );
  NAND2_X2 U8037 ( .A1(REGFILE_reg_out_20__26_), .A2(net77384), .ZN(n7102) );
  NAND2_X2 U8038 ( .A1(REGFILE_reg_out_18__26_), .A2(n6017), .ZN(n7101) );
  NAND2_X2 U8039 ( .A1(REGFILE_reg_out_16__26_), .A2(net77318), .ZN(n7100) );
  NAND4_X2 U8040 ( .A1(n7103), .A2(n7102), .A3(n7101), .A4(n7100), .ZN(n7104)
         );
  NAND2_X2 U8041 ( .A1(REGFILE_reg_out_14__26_), .A2(net77568), .ZN(n7109) );
  NAND2_X2 U8042 ( .A1(REGFILE_reg_out_15__26_), .A2(net77498), .ZN(n7107) );
  NAND2_X2 U8043 ( .A1(REGFILE_reg_out_13__26_), .A2(net77462), .ZN(n7106) );
  NAND4_X2 U8044 ( .A1(n7109), .A2(n7108), .A3(n7107), .A4(n7106), .ZN(n7115)
         );
  NAND2_X2 U8045 ( .A1(REGFILE_reg_out_11__26_), .A2(net77426), .ZN(n7113) );
  NAND2_X2 U8046 ( .A1(REGFILE_reg_out_12__26_), .A2(net77380), .ZN(n7112) );
  NAND2_X2 U8047 ( .A1(REGFILE_reg_out_10__26_), .A2(n6017), .ZN(n7111) );
  NAND2_X2 U8048 ( .A1(REGFILE_reg_out_8__26_), .A2(net77318), .ZN(n7110) );
  NAND4_X2 U8049 ( .A1(n7113), .A2(n7112), .A3(n7111), .A4(n7110), .ZN(n7114)
         );
  NAND2_X2 U8050 ( .A1(REGFILE_reg_out_6__26_), .A2(net77560), .ZN(n7119) );
  NAND2_X2 U8051 ( .A1(REGFILE_reg_out_7__26_), .A2(net77498), .ZN(n7117) );
  NAND2_X2 U8052 ( .A1(REGFILE_reg_out_5__26_), .A2(net77462), .ZN(n7116) );
  NAND4_X2 U8053 ( .A1(n7119), .A2(n7118), .A3(n7117), .A4(n7116), .ZN(n7125)
         );
  NAND2_X2 U8054 ( .A1(REGFILE_reg_out_3__26_), .A2(net77426), .ZN(n7123) );
  NAND2_X2 U8055 ( .A1(REGFILE_reg_out_4__26_), .A2(net77382), .ZN(n7122) );
  NAND2_X2 U8056 ( .A1(REGFILE_reg_out_2__26_), .A2(n6017), .ZN(n7121) );
  NAND2_X2 U8057 ( .A1(REGFILE_reg_out_0__26_), .A2(net77318), .ZN(n7120) );
  NAND4_X2 U8058 ( .A1(n7123), .A2(n7122), .A3(n7121), .A4(n7120), .ZN(n7124)
         );
  NAND4_X2 U8059 ( .A1(n7129), .A2(n7128), .A3(n7127), .A4(n7126), .ZN(n8448)
         );
  MUX2_X2 U8060 ( .A(n8448), .B(instruction[26]), .S(net77276), .Z(aluA[26])
         );
  NAND2_X2 U8061 ( .A1(REGFILE_reg_out_27__25_), .A2(net77426), .ZN(n7133) );
  NAND2_X2 U8062 ( .A1(REGFILE_reg_out_28__25_), .A2(net77376), .ZN(n7132) );
  NAND2_X2 U8063 ( .A1(REGFILE_reg_out_26__25_), .A2(n6017), .ZN(n7131) );
  NAND2_X2 U8064 ( .A1(REGFILE_reg_out_24__25_), .A2(net77318), .ZN(n7130) );
  NAND4_X2 U8065 ( .A1(n7133), .A2(n7132), .A3(n7131), .A4(n7130), .ZN(n7139)
         );
  NAND2_X2 U8066 ( .A1(REGFILE_reg_out_30__25_), .A2(net77558), .ZN(n7137) );
  NAND2_X2 U8067 ( .A1(REGFILE_reg_out_25__25_), .A2(net77544), .ZN(n7136) );
  NAND2_X2 U8068 ( .A1(REGFILE_reg_out_31__25_), .A2(net77498), .ZN(n7135) );
  NAND2_X2 U8069 ( .A1(REGFILE_reg_out_29__25_), .A2(net77462), .ZN(n7134) );
  NAND4_X2 U8070 ( .A1(n7137), .A2(n7136), .A3(n7135), .A4(n7134), .ZN(n7138)
         );
  NAND2_X2 U8071 ( .A1(REGFILE_reg_out_3__25_), .A2(net77424), .ZN(n7143) );
  NAND2_X2 U8073 ( .A1(REGFILE_reg_out_2__25_), .A2(n6016), .ZN(n7141) );
  NAND2_X2 U8074 ( .A1(REGFILE_reg_out_0__25_), .A2(net77316), .ZN(n7140) );
  NAND4_X2 U8075 ( .A1(n7143), .A2(n7142), .A3(n7141), .A4(n7140), .ZN(n7149)
         );
  NAND2_X2 U8076 ( .A1(REGFILE_reg_out_6__25_), .A2(net77568), .ZN(n7147) );
  NAND2_X2 U8077 ( .A1(REGFILE_reg_out_1__25_), .A2(net77532), .ZN(n7146) );
  NAND2_X2 U8078 ( .A1(REGFILE_reg_out_7__25_), .A2(net77496), .ZN(n7145) );
  NAND2_X2 U8079 ( .A1(REGFILE_reg_out_5__25_), .A2(net77460), .ZN(n7144) );
  NAND4_X2 U8080 ( .A1(n7147), .A2(n7146), .A3(n7145), .A4(n7144), .ZN(n7148)
         );
  NAND2_X2 U8081 ( .A1(REGFILE_reg_out_11__25_), .A2(net77424), .ZN(n7153) );
  NAND2_X2 U8083 ( .A1(REGFILE_reg_out_10__25_), .A2(n6016), .ZN(n7151) );
  NAND2_X2 U8084 ( .A1(REGFILE_reg_out_8__25_), .A2(net77316), .ZN(n7150) );
  NAND4_X2 U8085 ( .A1(n7153), .A2(n7152), .A3(n7151), .A4(n7150), .ZN(n7159)
         );
  NAND2_X2 U8086 ( .A1(REGFILE_reg_out_14__25_), .A2(net77568), .ZN(n7157) );
  NAND2_X2 U8087 ( .A1(REGFILE_reg_out_9__25_), .A2(net77532), .ZN(n7156) );
  NAND2_X2 U8088 ( .A1(REGFILE_reg_out_15__25_), .A2(net77496), .ZN(n7155) );
  NAND2_X2 U8089 ( .A1(REGFILE_reg_out_13__25_), .A2(net77460), .ZN(n7154) );
  NAND4_X2 U8090 ( .A1(n7157), .A2(n7156), .A3(n7155), .A4(n7154), .ZN(n7158)
         );
  NAND2_X2 U8091 ( .A1(REGFILE_reg_out_19__25_), .A2(net77424), .ZN(n7163) );
  NAND2_X2 U8093 ( .A1(REGFILE_reg_out_18__25_), .A2(n6016), .ZN(n7161) );
  NAND2_X2 U8094 ( .A1(REGFILE_reg_out_16__25_), .A2(net77316), .ZN(n7160) );
  NAND4_X2 U8095 ( .A1(n7163), .A2(n7162), .A3(n7161), .A4(n7160), .ZN(n7169)
         );
  NAND2_X2 U8096 ( .A1(REGFILE_reg_out_22__25_), .A2(net77568), .ZN(n7167) );
  NAND2_X2 U8097 ( .A1(REGFILE_reg_out_17__25_), .A2(net77532), .ZN(n7166) );
  NAND2_X2 U8098 ( .A1(REGFILE_reg_out_23__25_), .A2(net77496), .ZN(n7165) );
  NAND2_X2 U8099 ( .A1(REGFILE_reg_out_21__25_), .A2(net77460), .ZN(n7164) );
  NAND4_X2 U8100 ( .A1(n7167), .A2(n7166), .A3(n7165), .A4(n7164), .ZN(n7168)
         );
  NAND4_X2 U8101 ( .A1(n7173), .A2(n7172), .A3(n7171), .A4(n7170), .ZN(n8419)
         );
  INV_X4 U8102 ( .A(n8419), .ZN(n7174) );
  INV_X4 U8103 ( .A(instruction[25]), .ZN(n8329) );
  MUX2_X2 U8104 ( .A(n7174), .B(n8329), .S(net77276), .Z(n10327) );
  NAND2_X2 U8105 ( .A1(REGFILE_reg_out_27__24_), .A2(net77424), .ZN(n7178) );
  NAND2_X2 U8107 ( .A1(REGFILE_reg_out_26__24_), .A2(n6016), .ZN(n7176) );
  NAND2_X2 U8108 ( .A1(REGFILE_reg_out_24__24_), .A2(net77316), .ZN(n7175) );
  NAND4_X2 U8109 ( .A1(n7178), .A2(n7177), .A3(n7176), .A4(n7175), .ZN(n7184)
         );
  NAND2_X2 U8110 ( .A1(REGFILE_reg_out_30__24_), .A2(net77568), .ZN(n7182) );
  NAND2_X2 U8111 ( .A1(REGFILE_reg_out_25__24_), .A2(net77532), .ZN(n7181) );
  NAND2_X2 U8112 ( .A1(REGFILE_reg_out_31__24_), .A2(net77496), .ZN(n7180) );
  NAND2_X2 U8113 ( .A1(REGFILE_reg_out_29__24_), .A2(net77460), .ZN(n7179) );
  NAND4_X2 U8114 ( .A1(n7182), .A2(n7181), .A3(n7180), .A4(n7179), .ZN(n7183)
         );
  NAND2_X2 U8115 ( .A1(REGFILE_reg_out_3__24_), .A2(net77424), .ZN(n7188) );
  NAND2_X2 U8117 ( .A1(REGFILE_reg_out_2__24_), .A2(n6016), .ZN(n7186) );
  NAND2_X2 U8118 ( .A1(REGFILE_reg_out_0__24_), .A2(net77316), .ZN(n7185) );
  NAND4_X2 U8119 ( .A1(n7188), .A2(n7187), .A3(n7186), .A4(n7185), .ZN(n7194)
         );
  NAND2_X2 U8120 ( .A1(REGFILE_reg_out_6__24_), .A2(net77568), .ZN(n7192) );
  NAND2_X2 U8121 ( .A1(REGFILE_reg_out_1__24_), .A2(net77532), .ZN(n7191) );
  NAND2_X2 U8122 ( .A1(REGFILE_reg_out_7__24_), .A2(net77496), .ZN(n7190) );
  NAND2_X2 U8123 ( .A1(REGFILE_reg_out_5__24_), .A2(net77460), .ZN(n7189) );
  NAND4_X2 U8124 ( .A1(n7192), .A2(n7191), .A3(n7190), .A4(n7189), .ZN(n7193)
         );
  NAND2_X2 U8125 ( .A1(REGFILE_reg_out_11__24_), .A2(net77424), .ZN(n7198) );
  NAND2_X2 U8127 ( .A1(REGFILE_reg_out_10__24_), .A2(n6016), .ZN(n7196) );
  NAND2_X2 U8128 ( .A1(REGFILE_reg_out_8__24_), .A2(net77316), .ZN(n7195) );
  NAND4_X2 U8129 ( .A1(n7198), .A2(n7197), .A3(n7196), .A4(n7195), .ZN(n7204)
         );
  NAND2_X2 U8130 ( .A1(REGFILE_reg_out_14__24_), .A2(net77568), .ZN(n7202) );
  NAND2_X2 U8131 ( .A1(REGFILE_reg_out_9__24_), .A2(net77532), .ZN(n7201) );
  NAND2_X2 U8132 ( .A1(REGFILE_reg_out_15__24_), .A2(net77496), .ZN(n7200) );
  NAND2_X2 U8133 ( .A1(REGFILE_reg_out_13__24_), .A2(net77460), .ZN(n7199) );
  NAND4_X2 U8134 ( .A1(n7202), .A2(n7201), .A3(n7200), .A4(n7199), .ZN(n7203)
         );
  NAND2_X2 U8135 ( .A1(REGFILE_reg_out_19__24_), .A2(net77424), .ZN(n7208) );
  NAND2_X2 U8137 ( .A1(REGFILE_reg_out_18__24_), .A2(n6016), .ZN(n7206) );
  NAND2_X2 U8138 ( .A1(REGFILE_reg_out_16__24_), .A2(net77316), .ZN(n7205) );
  NAND4_X2 U8139 ( .A1(n7208), .A2(n7207), .A3(n7206), .A4(n7205), .ZN(n7214)
         );
  NAND2_X2 U8140 ( .A1(REGFILE_reg_out_22__24_), .A2(net77568), .ZN(n7212) );
  NAND2_X2 U8141 ( .A1(REGFILE_reg_out_17__24_), .A2(net77532), .ZN(n7211) );
  NAND2_X2 U8142 ( .A1(REGFILE_reg_out_23__24_), .A2(net77496), .ZN(n7210) );
  NAND2_X2 U8143 ( .A1(REGFILE_reg_out_21__24_), .A2(net77460), .ZN(n7209) );
  NAND4_X2 U8144 ( .A1(n7212), .A2(n7211), .A3(n7210), .A4(n7209), .ZN(n7213)
         );
  NAND4_X2 U8145 ( .A1(n7218), .A2(n7217), .A3(n7216), .A4(n7215), .ZN(n8420)
         );
  INV_X4 U8146 ( .A(n8420), .ZN(n7219) );
  INV_X4 U8147 ( .A(instruction[24]), .ZN(n8351) );
  MUX2_X2 U8148 ( .A(n7219), .B(n8351), .S(net77276), .Z(net72312) );
  INV_X4 U8149 ( .A(net72312), .ZN(net36391) );
  NAND2_X2 U8150 ( .A1(REGFILE_reg_out_27__23_), .A2(net77424), .ZN(n7223) );
  NAND2_X2 U8152 ( .A1(REGFILE_reg_out_26__23_), .A2(n6016), .ZN(n7221) );
  NAND2_X2 U8153 ( .A1(REGFILE_reg_out_24__23_), .A2(net77316), .ZN(n7220) );
  NAND4_X2 U8154 ( .A1(n7223), .A2(n7222), .A3(n7221), .A4(n7220), .ZN(n7229)
         );
  NAND2_X2 U8155 ( .A1(REGFILE_reg_out_30__23_), .A2(net77568), .ZN(n7227) );
  NAND2_X2 U8156 ( .A1(REGFILE_reg_out_25__23_), .A2(net77532), .ZN(n7226) );
  NAND2_X2 U8157 ( .A1(REGFILE_reg_out_31__23_), .A2(net77496), .ZN(n7225) );
  NAND2_X2 U8158 ( .A1(REGFILE_reg_out_29__23_), .A2(net77460), .ZN(n7224) );
  NAND4_X2 U8159 ( .A1(n7227), .A2(n7226), .A3(n7225), .A4(n7224), .ZN(n7228)
         );
  NAND2_X2 U8160 ( .A1(REGFILE_reg_out_3__23_), .A2(net77424), .ZN(n7233) );
  NAND2_X2 U8162 ( .A1(REGFILE_reg_out_2__23_), .A2(n6016), .ZN(n7231) );
  NAND2_X2 U8163 ( .A1(REGFILE_reg_out_0__23_), .A2(net77316), .ZN(n7230) );
  NAND4_X2 U8164 ( .A1(n7233), .A2(n7232), .A3(n7231), .A4(n7230), .ZN(n7239)
         );
  NAND2_X2 U8165 ( .A1(REGFILE_reg_out_6__23_), .A2(net77568), .ZN(n7237) );
  NAND2_X2 U8166 ( .A1(REGFILE_reg_out_1__23_), .A2(net77532), .ZN(n7236) );
  NAND2_X2 U8167 ( .A1(REGFILE_reg_out_7__23_), .A2(net77496), .ZN(n7235) );
  NAND2_X2 U8168 ( .A1(REGFILE_reg_out_5__23_), .A2(net77460), .ZN(n7234) );
  NAND4_X2 U8169 ( .A1(n7237), .A2(n7236), .A3(n7235), .A4(n7234), .ZN(n7238)
         );
  NAND2_X2 U8170 ( .A1(REGFILE_reg_out_11__23_), .A2(net77424), .ZN(n7243) );
  NAND2_X2 U8172 ( .A1(REGFILE_reg_out_10__23_), .A2(n6016), .ZN(n7241) );
  NAND2_X2 U8173 ( .A1(REGFILE_reg_out_8__23_), .A2(net77316), .ZN(n7240) );
  NAND4_X2 U8174 ( .A1(n7243), .A2(n7242), .A3(n7241), .A4(n7240), .ZN(n7249)
         );
  NAND2_X2 U8175 ( .A1(REGFILE_reg_out_14__23_), .A2(net77568), .ZN(n7247) );
  NAND2_X2 U8176 ( .A1(REGFILE_reg_out_9__23_), .A2(net77532), .ZN(n7246) );
  NAND2_X2 U8177 ( .A1(REGFILE_reg_out_15__23_), .A2(net77496), .ZN(n7245) );
  NAND2_X2 U8178 ( .A1(REGFILE_reg_out_13__23_), .A2(net77460), .ZN(n7244) );
  NAND4_X2 U8179 ( .A1(n7247), .A2(n7246), .A3(n7245), .A4(n7244), .ZN(n7248)
         );
  NAND2_X2 U8180 ( .A1(REGFILE_reg_out_19__23_), .A2(net77424), .ZN(n7253) );
  NAND2_X2 U8182 ( .A1(REGFILE_reg_out_18__23_), .A2(n6016), .ZN(n7251) );
  NAND2_X2 U8183 ( .A1(REGFILE_reg_out_16__23_), .A2(net77316), .ZN(n7250) );
  NAND4_X2 U8184 ( .A1(n7253), .A2(n7252), .A3(n7251), .A4(n7250), .ZN(n7259)
         );
  NAND2_X2 U8185 ( .A1(REGFILE_reg_out_22__23_), .A2(net77568), .ZN(n7257) );
  NAND2_X2 U8186 ( .A1(REGFILE_reg_out_17__23_), .A2(net77532), .ZN(n7256) );
  NAND2_X2 U8187 ( .A1(REGFILE_reg_out_23__23_), .A2(net77496), .ZN(n7255) );
  NAND2_X2 U8188 ( .A1(REGFILE_reg_out_21__23_), .A2(net77460), .ZN(n7254) );
  NAND4_X2 U8189 ( .A1(n7257), .A2(n7256), .A3(n7255), .A4(n7254), .ZN(n7258)
         );
  NAND4_X2 U8190 ( .A1(n7263), .A2(n7262), .A3(n7261), .A4(n7260), .ZN(n8418)
         );
  INV_X4 U8191 ( .A(n8418), .ZN(n7264) );
  INV_X4 U8192 ( .A(instruction[23]), .ZN(n8324) );
  MUX2_X2 U8193 ( .A(n7264), .B(n8324), .S(net77276), .Z(n10334) );
  INV_X4 U8194 ( .A(n10334), .ZN(n10931) );
  NAND2_X2 U8195 ( .A1(REGFILE_reg_out_27__22_), .A2(net77424), .ZN(n7268) );
  NAND2_X2 U8197 ( .A1(REGFILE_reg_out_26__22_), .A2(n6016), .ZN(n7266) );
  NAND2_X2 U8198 ( .A1(REGFILE_reg_out_24__22_), .A2(net77316), .ZN(n7265) );
  NAND4_X2 U8199 ( .A1(n7268), .A2(n7267), .A3(n7266), .A4(n7265), .ZN(n7274)
         );
  NAND2_X2 U8200 ( .A1(REGFILE_reg_out_30__22_), .A2(net77568), .ZN(n7272) );
  NAND2_X2 U8201 ( .A1(REGFILE_reg_out_25__22_), .A2(net77532), .ZN(n7271) );
  NAND2_X2 U8202 ( .A1(REGFILE_reg_out_31__22_), .A2(net77496), .ZN(n7270) );
  NAND2_X2 U8203 ( .A1(REGFILE_reg_out_29__22_), .A2(net77460), .ZN(n7269) );
  NAND4_X2 U8204 ( .A1(n7272), .A2(n7271), .A3(n7270), .A4(n7269), .ZN(n7273)
         );
  NAND2_X2 U8205 ( .A1(REGFILE_reg_out_3__22_), .A2(net77422), .ZN(n7278) );
  NAND2_X2 U8206 ( .A1(REGFILE_reg_out_2__22_), .A2(n6015), .ZN(n7276) );
  NAND2_X2 U8207 ( .A1(REGFILE_reg_out_0__22_), .A2(net77314), .ZN(n7275) );
  NAND4_X2 U8208 ( .A1(n7278), .A2(n7277), .A3(n7276), .A4(n7275), .ZN(n7284)
         );
  NAND2_X2 U8209 ( .A1(REGFILE_reg_out_6__22_), .A2(net77566), .ZN(n7282) );
  NAND2_X2 U8210 ( .A1(REGFILE_reg_out_1__22_), .A2(net77530), .ZN(n7281) );
  NAND2_X2 U8211 ( .A1(REGFILE_reg_out_7__22_), .A2(net77494), .ZN(n7280) );
  NAND2_X2 U8212 ( .A1(REGFILE_reg_out_5__22_), .A2(net77458), .ZN(n7279) );
  NAND4_X2 U8213 ( .A1(n7282), .A2(n7281), .A3(n7280), .A4(n7279), .ZN(n7283)
         );
  NAND2_X2 U8214 ( .A1(REGFILE_reg_out_11__22_), .A2(net77422), .ZN(n7288) );
  NAND2_X2 U8215 ( .A1(REGFILE_reg_out_8__22_), .A2(net77314), .ZN(n7285) );
  NAND4_X2 U8216 ( .A1(n7288), .A2(n7287), .A3(n7286), .A4(n7285), .ZN(n7294)
         );
  NAND2_X2 U8217 ( .A1(REGFILE_reg_out_14__22_), .A2(net77566), .ZN(n7292) );
  NAND2_X2 U8218 ( .A1(REGFILE_reg_out_9__22_), .A2(net77530), .ZN(n7291) );
  NAND2_X2 U8219 ( .A1(REGFILE_reg_out_15__22_), .A2(net77494), .ZN(n7290) );
  NAND2_X2 U8220 ( .A1(REGFILE_reg_out_13__22_), .A2(net77458), .ZN(n7289) );
  NAND4_X2 U8221 ( .A1(n7292), .A2(n7291), .A3(n7290), .A4(n7289), .ZN(n7293)
         );
  NAND2_X2 U8222 ( .A1(REGFILE_reg_out_19__22_), .A2(net77422), .ZN(n7298) );
  NAND2_X2 U8223 ( .A1(REGFILE_reg_out_18__22_), .A2(n6015), .ZN(n7296) );
  NAND2_X2 U8224 ( .A1(REGFILE_reg_out_16__22_), .A2(net77314), .ZN(n7295) );
  NAND4_X2 U8225 ( .A1(n7298), .A2(n7297), .A3(n7296), .A4(n7295), .ZN(n7304)
         );
  NAND2_X2 U8226 ( .A1(REGFILE_reg_out_22__22_), .A2(net77566), .ZN(n7302) );
  NAND2_X2 U8227 ( .A1(REGFILE_reg_out_17__22_), .A2(net77530), .ZN(n7301) );
  NAND2_X2 U8228 ( .A1(REGFILE_reg_out_23__22_), .A2(net77494), .ZN(n7300) );
  NAND2_X2 U8229 ( .A1(REGFILE_reg_out_21__22_), .A2(net77458), .ZN(n7299) );
  NAND4_X2 U8230 ( .A1(n7302), .A2(n7301), .A3(n7300), .A4(n7299), .ZN(n7303)
         );
  NAND4_X2 U8231 ( .A1(n7308), .A2(n7307), .A3(n7306), .A4(n7305), .ZN(n8400)
         );
  INV_X4 U8232 ( .A(n8400), .ZN(n7309) );
  INV_X4 U8233 ( .A(instruction[22]), .ZN(n8355) );
  MUX2_X2 U8234 ( .A(n7309), .B(n8355), .S(net77276), .Z(n8967) );
  INV_X4 U8235 ( .A(n8967), .ZN(n10932) );
  NAND2_X2 U8236 ( .A1(REGFILE_reg_out_26__21_), .A2(n6015), .ZN(n7311) );
  NAND2_X2 U8237 ( .A1(REGFILE_reg_out_24__21_), .A2(net77314), .ZN(n7310) );
  NAND4_X2 U8238 ( .A1(n7313), .A2(n7312), .A3(n7311), .A4(n7310), .ZN(n7319)
         );
  NAND2_X2 U8239 ( .A1(REGFILE_reg_out_30__21_), .A2(net77566), .ZN(n7317) );
  NAND2_X2 U8240 ( .A1(REGFILE_reg_out_31__21_), .A2(net77494), .ZN(n7315) );
  NAND2_X2 U8241 ( .A1(REGFILE_reg_out_29__21_), .A2(net77458), .ZN(n7314) );
  NAND4_X2 U8242 ( .A1(n7317), .A2(n7316), .A3(n7315), .A4(n7314), .ZN(n7318)
         );
  NAND2_X2 U8243 ( .A1(REGFILE_reg_out_3__21_), .A2(net77422), .ZN(n7323) );
  NAND2_X2 U8244 ( .A1(REGFILE_reg_out_2__21_), .A2(n6015), .ZN(n7321) );
  NAND2_X2 U8245 ( .A1(REGFILE_reg_out_0__21_), .A2(net77314), .ZN(n7320) );
  NAND4_X2 U8246 ( .A1(n7323), .A2(n7322), .A3(n7321), .A4(n7320), .ZN(n7329)
         );
  NAND2_X2 U8247 ( .A1(REGFILE_reg_out_6__21_), .A2(net77566), .ZN(n7327) );
  NAND2_X2 U8248 ( .A1(REGFILE_reg_out_1__21_), .A2(net77530), .ZN(n7326) );
  NAND2_X2 U8249 ( .A1(REGFILE_reg_out_7__21_), .A2(net77494), .ZN(n7325) );
  NAND2_X2 U8250 ( .A1(REGFILE_reg_out_5__21_), .A2(net77458), .ZN(n7324) );
  NAND4_X2 U8251 ( .A1(n7327), .A2(n7326), .A3(n7325), .A4(n7324), .ZN(n7328)
         );
  NAND2_X2 U8252 ( .A1(REGFILE_reg_out_11__21_), .A2(net77422), .ZN(n7333) );
  NAND2_X2 U8253 ( .A1(REGFILE_reg_out_10__21_), .A2(n6015), .ZN(n7331) );
  NAND2_X2 U8254 ( .A1(REGFILE_reg_out_8__21_), .A2(net77314), .ZN(n7330) );
  NAND4_X2 U8255 ( .A1(n7333), .A2(n7332), .A3(n7331), .A4(n7330), .ZN(n7339)
         );
  NAND2_X2 U8256 ( .A1(REGFILE_reg_out_14__21_), .A2(net77566), .ZN(n7337) );
  NAND2_X2 U8257 ( .A1(REGFILE_reg_out_9__21_), .A2(net77530), .ZN(n7336) );
  NAND2_X2 U8258 ( .A1(REGFILE_reg_out_15__21_), .A2(net77494), .ZN(n7335) );
  NAND2_X2 U8259 ( .A1(REGFILE_reg_out_13__21_), .A2(net77458), .ZN(n7334) );
  NAND4_X2 U8260 ( .A1(n7337), .A2(n7336), .A3(n7335), .A4(n7334), .ZN(n7338)
         );
  NAND2_X2 U8261 ( .A1(REGFILE_reg_out_19__21_), .A2(net77422), .ZN(n7343) );
  NAND2_X2 U8262 ( .A1(REGFILE_reg_out_18__21_), .A2(n6015), .ZN(n7341) );
  NAND2_X2 U8263 ( .A1(REGFILE_reg_out_16__21_), .A2(net77314), .ZN(n7340) );
  NAND4_X2 U8264 ( .A1(n7343), .A2(n7342), .A3(n7341), .A4(n7340), .ZN(n7349)
         );
  NAND2_X2 U8265 ( .A1(REGFILE_reg_out_22__21_), .A2(net77566), .ZN(n7347) );
  NAND2_X2 U8266 ( .A1(REGFILE_reg_out_17__21_), .A2(net77530), .ZN(n7346) );
  NAND2_X2 U8267 ( .A1(REGFILE_reg_out_23__21_), .A2(net77494), .ZN(n7345) );
  NAND2_X2 U8268 ( .A1(REGFILE_reg_out_21__21_), .A2(net77458), .ZN(n7344) );
  NAND4_X2 U8269 ( .A1(n7347), .A2(n7346), .A3(n7345), .A4(n7344), .ZN(n7348)
         );
  NAND4_X2 U8270 ( .A1(n7353), .A2(n7352), .A3(n7351), .A4(n7350), .ZN(n8417)
         );
  INV_X4 U8271 ( .A(n8417), .ZN(n7354) );
  INV_X4 U8272 ( .A(instruction[21]), .ZN(n8319) );
  MUX2_X2 U8273 ( .A(n7354), .B(n8319), .S(net77276), .Z(n10341) );
  INV_X4 U8274 ( .A(n10341), .ZN(n10933) );
  NAND2_X2 U8275 ( .A1(REGFILE_reg_out_30__20_), .A2(net77566), .ZN(n7358) );
  NAND2_X2 U8276 ( .A1(REGFILE_reg_out_31__20_), .A2(net77494), .ZN(n7356) );
  NAND2_X2 U8277 ( .A1(REGFILE_reg_out_29__20_), .A2(net77458), .ZN(n7355) );
  NAND4_X2 U8278 ( .A1(n7358), .A2(n7357), .A3(n7356), .A4(n7355), .ZN(n7364)
         );
  NAND2_X2 U8279 ( .A1(REGFILE_reg_out_26__20_), .A2(n6015), .ZN(n7360) );
  NAND2_X2 U8280 ( .A1(REGFILE_reg_out_24__20_), .A2(net77314), .ZN(n7359) );
  NAND4_X2 U8281 ( .A1(n7362), .A2(n7361), .A3(n7360), .A4(n7359), .ZN(n7363)
         );
  NAND2_X2 U8282 ( .A1(REGFILE_reg_out_22__20_), .A2(net77566), .ZN(n7368) );
  NAND2_X2 U8283 ( .A1(REGFILE_reg_out_17__20_), .A2(net77530), .ZN(n7367) );
  NAND2_X2 U8284 ( .A1(REGFILE_reg_out_23__20_), .A2(net77494), .ZN(n7366) );
  NAND2_X2 U8285 ( .A1(REGFILE_reg_out_21__20_), .A2(net77458), .ZN(n7365) );
  NAND4_X2 U8286 ( .A1(n7368), .A2(n7367), .A3(n7366), .A4(n7365), .ZN(n7374)
         );
  NAND2_X2 U8287 ( .A1(REGFILE_reg_out_19__20_), .A2(net77422), .ZN(n7372) );
  NAND2_X2 U8288 ( .A1(REGFILE_reg_out_18__20_), .A2(n6015), .ZN(n7370) );
  NAND2_X2 U8289 ( .A1(REGFILE_reg_out_16__20_), .A2(net77314), .ZN(n7369) );
  NAND4_X2 U8290 ( .A1(n7372), .A2(n7371), .A3(n7370), .A4(n7369), .ZN(n7373)
         );
  NAND2_X2 U8291 ( .A1(REGFILE_reg_out_14__20_), .A2(net77566), .ZN(n7378) );
  NAND2_X2 U8292 ( .A1(REGFILE_reg_out_9__20_), .A2(net77530), .ZN(n7377) );
  NAND2_X2 U8293 ( .A1(REGFILE_reg_out_15__20_), .A2(net77494), .ZN(n7376) );
  NAND2_X2 U8294 ( .A1(REGFILE_reg_out_13__20_), .A2(net77458), .ZN(n7375) );
  NAND4_X2 U8295 ( .A1(n7378), .A2(n7377), .A3(n7376), .A4(n7375), .ZN(n7384)
         );
  NAND2_X2 U8296 ( .A1(REGFILE_reg_out_11__20_), .A2(net77422), .ZN(n7382) );
  NAND2_X2 U8297 ( .A1(REGFILE_reg_out_10__20_), .A2(n6015), .ZN(n7380) );
  NAND2_X2 U8298 ( .A1(REGFILE_reg_out_8__20_), .A2(net77314), .ZN(n7379) );
  NAND4_X2 U8299 ( .A1(n7382), .A2(n7381), .A3(n7380), .A4(n7379), .ZN(n7383)
         );
  NAND2_X2 U8300 ( .A1(REGFILE_reg_out_6__20_), .A2(net77566), .ZN(n7388) );
  NAND2_X2 U8301 ( .A1(REGFILE_reg_out_1__20_), .A2(net77530), .ZN(n7387) );
  NAND2_X2 U8302 ( .A1(REGFILE_reg_out_7__20_), .A2(net77494), .ZN(n7386) );
  NAND2_X2 U8303 ( .A1(REGFILE_reg_out_5__20_), .A2(net77458), .ZN(n7385) );
  NAND4_X2 U8304 ( .A1(n7388), .A2(n7387), .A3(n7386), .A4(n7385), .ZN(n7394)
         );
  NAND2_X2 U8305 ( .A1(REGFILE_reg_out_0__20_), .A2(net77314), .ZN(n7389) );
  NAND4_X2 U8306 ( .A1(n7392), .A2(n7391), .A3(n7390), .A4(n7389), .ZN(n7393)
         );
  NAND4_X2 U8307 ( .A1(n7398), .A2(n7397), .A3(n7396), .A4(n7395), .ZN(n8449)
         );
  MUX2_X2 U8308 ( .A(n8449), .B(instruction[20]), .S(net77276), .Z(aluA[20])
         );
  NAND2_X2 U8309 ( .A1(REGFILE_reg_out_30__19_), .A2(net77566), .ZN(n7402) );
  NAND2_X2 U8310 ( .A1(REGFILE_reg_out_25__19_), .A2(net77530), .ZN(n7401) );
  NAND2_X2 U8311 ( .A1(REGFILE_reg_out_31__19_), .A2(net77494), .ZN(n7400) );
  NAND2_X2 U8312 ( .A1(REGFILE_reg_out_29__19_), .A2(net77458), .ZN(n7399) );
  NAND4_X2 U8313 ( .A1(n7402), .A2(n7401), .A3(n7400), .A4(n7399), .ZN(n7408)
         );
  NAND2_X2 U8314 ( .A1(REGFILE_reg_out_26__19_), .A2(n6015), .ZN(n7404) );
  NAND2_X2 U8315 ( .A1(REGFILE_reg_out_24__19_), .A2(net77314), .ZN(n7403) );
  NAND4_X2 U8316 ( .A1(n7406), .A2(n7405), .A3(n7404), .A4(n7403), .ZN(n7407)
         );
  NAND2_X2 U8317 ( .A1(REGFILE_reg_out_22__19_), .A2(net77564), .ZN(n7412) );
  NAND2_X2 U8318 ( .A1(REGFILE_reg_out_17__19_), .A2(net77528), .ZN(n7411) );
  NAND2_X2 U8319 ( .A1(REGFILE_reg_out_23__19_), .A2(net77492), .ZN(n7410) );
  NAND2_X2 U8320 ( .A1(REGFILE_reg_out_21__19_), .A2(net77456), .ZN(n7409) );
  NAND4_X2 U8321 ( .A1(n7412), .A2(n7411), .A3(n7410), .A4(n7409), .ZN(n7418)
         );
  NAND2_X2 U8322 ( .A1(REGFILE_reg_out_19__19_), .A2(net77420), .ZN(n7416) );
  NAND2_X2 U8323 ( .A1(REGFILE_reg_out_20__19_), .A2(net77384), .ZN(n7415) );
  NAND2_X2 U8324 ( .A1(REGFILE_reg_out_18__19_), .A2(net77348), .ZN(n7414) );
  NAND2_X2 U8325 ( .A1(REGFILE_reg_out_16__19_), .A2(net77312), .ZN(n7413) );
  NAND4_X2 U8326 ( .A1(n7416), .A2(n7415), .A3(n7414), .A4(n7413), .ZN(n7417)
         );
  NAND2_X2 U8327 ( .A1(REGFILE_reg_out_14__19_), .A2(net77564), .ZN(n7422) );
  NAND2_X2 U8328 ( .A1(REGFILE_reg_out_9__19_), .A2(net77528), .ZN(n7421) );
  NAND2_X2 U8329 ( .A1(REGFILE_reg_out_15__19_), .A2(net77492), .ZN(n7420) );
  NAND2_X2 U8330 ( .A1(REGFILE_reg_out_13__19_), .A2(net77456), .ZN(n7419) );
  NAND4_X2 U8331 ( .A1(n7422), .A2(n7421), .A3(n7420), .A4(n7419), .ZN(n7428)
         );
  NAND2_X2 U8332 ( .A1(REGFILE_reg_out_11__19_), .A2(net77420), .ZN(n7426) );
  NAND2_X2 U8333 ( .A1(REGFILE_reg_out_8__19_), .A2(net77312), .ZN(n7423) );
  NAND4_X2 U8334 ( .A1(n7426), .A2(n7425), .A3(n7424), .A4(n7423), .ZN(n7427)
         );
  NAND2_X2 U8335 ( .A1(REGFILE_reg_out_6__19_), .A2(net77564), .ZN(n7432) );
  NAND2_X2 U8336 ( .A1(REGFILE_reg_out_1__19_), .A2(net77528), .ZN(n7431) );
  NAND2_X2 U8337 ( .A1(REGFILE_reg_out_7__19_), .A2(net77492), .ZN(n7430) );
  NAND2_X2 U8338 ( .A1(REGFILE_reg_out_5__19_), .A2(net77456), .ZN(n7429) );
  NAND4_X2 U8339 ( .A1(n7432), .A2(n7431), .A3(n7430), .A4(n7429), .ZN(n7438)
         );
  NAND2_X2 U8340 ( .A1(REGFILE_reg_out_3__19_), .A2(net77420), .ZN(n7436) );
  NAND2_X2 U8341 ( .A1(REGFILE_reg_out_4__19_), .A2(net77384), .ZN(n7435) );
  NAND2_X2 U8342 ( .A1(REGFILE_reg_out_2__19_), .A2(net77348), .ZN(n7434) );
  NAND2_X2 U8343 ( .A1(REGFILE_reg_out_0__19_), .A2(net77312), .ZN(n7433) );
  NAND4_X2 U8344 ( .A1(n7436), .A2(n7435), .A3(n7434), .A4(n7433), .ZN(n7437)
         );
  NAND4_X2 U8345 ( .A1(n7442), .A2(n7441), .A3(n7440), .A4(n7439), .ZN(n8444)
         );
  MUX2_X2 U8346 ( .A(n8444), .B(instruction[19]), .S(net77276), .Z(aluA[19])
         );
  NAND2_X2 U8347 ( .A1(REGFILE_reg_out_30__18_), .A2(net77564), .ZN(n7446) );
  NAND2_X2 U8348 ( .A1(net77528), .A2(REGFILE_reg_out_25__18_), .ZN(n7445) );
  NAND2_X2 U8349 ( .A1(REGFILE_reg_out_31__18_), .A2(net77492), .ZN(n7444) );
  NAND2_X2 U8350 ( .A1(REGFILE_reg_out_29__18_), .A2(net77456), .ZN(n7443) );
  NAND4_X2 U8351 ( .A1(n7446), .A2(n7445), .A3(n7444), .A4(n7443), .ZN(n7452)
         );
  NAND2_X2 U8352 ( .A1(REGFILE_reg_out_26__18_), .A2(net77348), .ZN(n7448) );
  NAND2_X2 U8353 ( .A1(REGFILE_reg_out_24__18_), .A2(net77312), .ZN(n7447) );
  NAND4_X2 U8354 ( .A1(n7450), .A2(n7449), .A3(n7448), .A4(n7447), .ZN(n7451)
         );
  NAND2_X2 U8355 ( .A1(REGFILE_reg_out_22__18_), .A2(net77564), .ZN(n7456) );
  NAND2_X2 U8356 ( .A1(REGFILE_reg_out_17__18_), .A2(net77528), .ZN(n7455) );
  NAND2_X2 U8357 ( .A1(REGFILE_reg_out_23__18_), .A2(net77492), .ZN(n7454) );
  NAND2_X2 U8358 ( .A1(REGFILE_reg_out_21__18_), .A2(net77456), .ZN(n7453) );
  NAND4_X2 U8359 ( .A1(n7456), .A2(n7455), .A3(n7454), .A4(n7453), .ZN(n7462)
         );
  NAND2_X2 U8360 ( .A1(REGFILE_reg_out_19__18_), .A2(net77420), .ZN(n7460) );
  NAND2_X2 U8361 ( .A1(REGFILE_reg_out_20__18_), .A2(net77384), .ZN(n7459) );
  NAND2_X2 U8362 ( .A1(REGFILE_reg_out_18__18_), .A2(net77348), .ZN(n7458) );
  NAND2_X2 U8363 ( .A1(REGFILE_reg_out_16__18_), .A2(net77312), .ZN(n7457) );
  NAND4_X2 U8364 ( .A1(n7460), .A2(n7459), .A3(n7458), .A4(n7457), .ZN(n7461)
         );
  NAND2_X2 U8365 ( .A1(REGFILE_reg_out_14__18_), .A2(net77564), .ZN(n7466) );
  NAND2_X2 U8366 ( .A1(REGFILE_reg_out_9__18_), .A2(net77528), .ZN(n7465) );
  NAND2_X2 U8367 ( .A1(REGFILE_reg_out_15__18_), .A2(net77492), .ZN(n7464) );
  NAND2_X2 U8368 ( .A1(REGFILE_reg_out_13__18_), .A2(net77456), .ZN(n7463) );
  NAND4_X2 U8369 ( .A1(n7466), .A2(n7465), .A3(n7464), .A4(n7463), .ZN(n7472)
         );
  NAND2_X2 U8370 ( .A1(REGFILE_reg_out_11__18_), .A2(net77420), .ZN(n7470) );
  NAND2_X2 U8371 ( .A1(REGFILE_reg_out_10__18_), .A2(net77348), .ZN(n7468) );
  NAND2_X2 U8372 ( .A1(REGFILE_reg_out_8__18_), .A2(net77312), .ZN(n7467) );
  NAND4_X2 U8373 ( .A1(n7470), .A2(n7469), .A3(n7468), .A4(n7467), .ZN(n7471)
         );
  NAND2_X2 U8374 ( .A1(REGFILE_reg_out_6__18_), .A2(net77564), .ZN(n7476) );
  NAND2_X2 U8375 ( .A1(REGFILE_reg_out_1__18_), .A2(net77528), .ZN(n7475) );
  NAND2_X2 U8376 ( .A1(REGFILE_reg_out_7__18_), .A2(net77492), .ZN(n7474) );
  NAND4_X2 U8377 ( .A1(n7476), .A2(n7475), .A3(n7474), .A4(n7473), .ZN(n7482)
         );
  NAND2_X2 U8378 ( .A1(REGFILE_reg_out_3__18_), .A2(net77420), .ZN(n7480) );
  NAND2_X2 U8379 ( .A1(REGFILE_reg_out_4__18_), .A2(net77384), .ZN(n7479) );
  NAND2_X2 U8380 ( .A1(REGFILE_reg_out_0__18_), .A2(net77312), .ZN(n7477) );
  NAND4_X2 U8381 ( .A1(n7480), .A2(n7479), .A3(n7478), .A4(n7477), .ZN(n7481)
         );
  NAND4_X2 U8382 ( .A1(n7486), .A2(n7485), .A3(n7484), .A4(n7483), .ZN(n8443)
         );
  MUX2_X2 U8383 ( .A(n8443), .B(instruction[18]), .S(net77276), .Z(aluA[18])
         );
  NAND2_X2 U8384 ( .A1(REGFILE_reg_out_30__17_), .A2(net77564), .ZN(n7490) );
  NAND2_X2 U8385 ( .A1(REGFILE_reg_out_31__17_), .A2(net77492), .ZN(n7488) );
  NAND2_X2 U8386 ( .A1(REGFILE_reg_out_29__17_), .A2(net77456), .ZN(n7487) );
  NAND4_X2 U8387 ( .A1(n7490), .A2(n7489), .A3(n7488), .A4(n7487), .ZN(n7496)
         );
  NAND2_X2 U8388 ( .A1(REGFILE_reg_out_28__17_), .A2(net77384), .ZN(n7493) );
  NAND2_X2 U8389 ( .A1(REGFILE_reg_out_26__17_), .A2(net77348), .ZN(n7492) );
  NAND2_X2 U8390 ( .A1(REGFILE_reg_out_24__17_), .A2(net77312), .ZN(n7491) );
  NAND4_X2 U8391 ( .A1(n7494), .A2(n7493), .A3(n7492), .A4(n7491), .ZN(n7495)
         );
  NAND2_X2 U8392 ( .A1(REGFILE_reg_out_22__17_), .A2(net77564), .ZN(n7500) );
  NAND2_X2 U8393 ( .A1(REGFILE_reg_out_17__17_), .A2(net77528), .ZN(n7499) );
  NAND2_X2 U8394 ( .A1(REGFILE_reg_out_23__17_), .A2(net77492), .ZN(n7498) );
  NAND2_X2 U8395 ( .A1(REGFILE_reg_out_21__17_), .A2(net77456), .ZN(n7497) );
  NAND4_X2 U8396 ( .A1(n7500), .A2(n7499), .A3(n7498), .A4(n7497), .ZN(n7506)
         );
  NAND2_X2 U8397 ( .A1(REGFILE_reg_out_19__17_), .A2(net77420), .ZN(n7504) );
  NAND2_X2 U8398 ( .A1(REGFILE_reg_out_20__17_), .A2(net77384), .ZN(n7503) );
  NAND2_X2 U8399 ( .A1(REGFILE_reg_out_18__17_), .A2(net77348), .ZN(n7502) );
  NAND2_X2 U8400 ( .A1(REGFILE_reg_out_16__17_), .A2(net77312), .ZN(n7501) );
  NAND4_X2 U8401 ( .A1(n7504), .A2(n7503), .A3(n7502), .A4(n7501), .ZN(n7505)
         );
  NAND2_X2 U8402 ( .A1(REGFILE_reg_out_14__17_), .A2(net77564), .ZN(n7510) );
  NAND2_X2 U8403 ( .A1(REGFILE_reg_out_9__17_), .A2(net77528), .ZN(n7509) );
  NAND2_X2 U8404 ( .A1(REGFILE_reg_out_15__17_), .A2(net77492), .ZN(n7508) );
  NAND2_X2 U8405 ( .A1(REGFILE_reg_out_13__17_), .A2(net77456), .ZN(n7507) );
  NAND4_X2 U8406 ( .A1(n7510), .A2(n7509), .A3(n7508), .A4(n7507), .ZN(n7515)
         );
  NAND2_X2 U8407 ( .A1(REGFILE_reg_out_11__17_), .A2(net77420), .ZN(n7513) );
  NAND2_X2 U8408 ( .A1(REGFILE_reg_out_12__17_), .A2(net77384), .ZN(n7512) );
  NAND2_X2 U8409 ( .A1(REGFILE_reg_out_8__17_), .A2(net77312), .ZN(n7511) );
  NAND4_X2 U8410 ( .A1(n7513), .A2(n7512), .A3(net74808), .A4(n7511), .ZN(
        n7514) );
  NAND2_X2 U8411 ( .A1(REGFILE_reg_out_6__17_), .A2(net77564), .ZN(n7519) );
  NAND2_X2 U8412 ( .A1(REGFILE_reg_out_1__17_), .A2(net77528), .ZN(n7518) );
  NAND2_X2 U8413 ( .A1(REGFILE_reg_out_7__17_), .A2(net77492), .ZN(n7517) );
  NAND2_X2 U8414 ( .A1(REGFILE_reg_out_5__17_), .A2(net77456), .ZN(n7516) );
  NAND4_X2 U8415 ( .A1(n7519), .A2(n7518), .A3(n7517), .A4(n7516), .ZN(n7524)
         );
  NAND2_X2 U8416 ( .A1(REGFILE_reg_out_3__17_), .A2(net77420), .ZN(n7522) );
  NAND2_X2 U8417 ( .A1(REGFILE_reg_out_4__17_), .A2(net77384), .ZN(n7521) );
  NAND4_X2 U8418 ( .A1(n7522), .A2(n7521), .A3(n7520), .A4(net74799), .ZN(
        n7523) );
  NAND4_X2 U8419 ( .A1(n7528), .A2(n7527), .A3(n7526), .A4(n7525), .ZN(n8447)
         );
  MUX2_X2 U8420 ( .A(n8447), .B(instruction[17]), .S(net77276), .Z(aluA[17])
         );
  NAND2_X2 U8421 ( .A1(REGFILE_reg_out_30__16_), .A2(net77564), .ZN(n7532) );
  NAND2_X2 U8422 ( .A1(REGFILE_reg_out_31__16_), .A2(net77492), .ZN(n7530) );
  NAND2_X2 U8423 ( .A1(REGFILE_reg_out_29__16_), .A2(net77456), .ZN(n7529) );
  NAND4_X2 U8424 ( .A1(n7532), .A2(n7531), .A3(n7530), .A4(n7529), .ZN(n7538)
         );
  NAND2_X2 U8425 ( .A1(REGFILE_reg_out_28__16_), .A2(net77384), .ZN(n7535) );
  NAND2_X2 U8426 ( .A1(REGFILE_reg_out_26__16_), .A2(net77348), .ZN(n7534) );
  NAND2_X2 U8427 ( .A1(REGFILE_reg_out_24__16_), .A2(net77312), .ZN(n7533) );
  NAND4_X2 U8428 ( .A1(n7536), .A2(n7535), .A3(n7534), .A4(n7533), .ZN(n7537)
         );
  NAND2_X2 U8429 ( .A1(REGFILE_reg_out_22__16_), .A2(net77562), .ZN(n7542) );
  NAND2_X2 U8430 ( .A1(REGFILE_reg_out_17__16_), .A2(net77526), .ZN(n7541) );
  NAND2_X2 U8431 ( .A1(REGFILE_reg_out_23__16_), .A2(net77490), .ZN(n7540) );
  NAND2_X2 U8432 ( .A1(REGFILE_reg_out_21__16_), .A2(net77454), .ZN(n7539) );
  NAND4_X2 U8433 ( .A1(n7542), .A2(n7541), .A3(n7540), .A4(n7539), .ZN(n7548)
         );
  NAND2_X2 U8434 ( .A1(REGFILE_reg_out_19__16_), .A2(net77418), .ZN(n7546) );
  NAND2_X2 U8435 ( .A1(REGFILE_reg_out_20__16_), .A2(net77382), .ZN(n7545) );
  NAND2_X2 U8436 ( .A1(REGFILE_reg_out_16__16_), .A2(net77310), .ZN(n7543) );
  NAND4_X2 U8437 ( .A1(n7546), .A2(n7545), .A3(n7544), .A4(n7543), .ZN(n7547)
         );
  NAND2_X2 U8438 ( .A1(REGFILE_reg_out_14__16_), .A2(net77562), .ZN(n7552) );
  NAND2_X2 U8439 ( .A1(REGFILE_reg_out_9__16_), .A2(net77526), .ZN(n7551) );
  NAND2_X2 U8440 ( .A1(REGFILE_reg_out_15__16_), .A2(net77490), .ZN(n7550) );
  NAND2_X2 U8441 ( .A1(REGFILE_reg_out_13__16_), .A2(net77454), .ZN(n7549) );
  NAND4_X2 U8442 ( .A1(n7552), .A2(n7551), .A3(n7550), .A4(n7549), .ZN(n7558)
         );
  NAND2_X2 U8443 ( .A1(REGFILE_reg_out_11__16_), .A2(net77418), .ZN(n7556) );
  NAND2_X2 U8444 ( .A1(REGFILE_reg_out_10__16_), .A2(net77346), .ZN(n7554) );
  NAND2_X2 U8445 ( .A1(REGFILE_reg_out_8__16_), .A2(net77310), .ZN(n7553) );
  NAND4_X2 U8446 ( .A1(n7556), .A2(n7555), .A3(n7554), .A4(n7553), .ZN(n7557)
         );
  NAND2_X2 U8447 ( .A1(REGFILE_reg_out_7__16_), .A2(net77490), .ZN(n7560) );
  NAND2_X2 U8448 ( .A1(REGFILE_reg_out_5__16_), .A2(net77454), .ZN(n7559) );
  NAND4_X2 U8449 ( .A1(n7562), .A2(n7561), .A3(n7560), .A4(n7559), .ZN(n7568)
         );
  NAND2_X2 U8450 ( .A1(REGFILE_reg_out_3__16_), .A2(net77418), .ZN(n7566) );
  NAND2_X2 U8451 ( .A1(REGFILE_reg_out_4__16_), .A2(net77382), .ZN(n7565) );
  NAND2_X2 U8452 ( .A1(REGFILE_reg_out_2__16_), .A2(net77346), .ZN(n7564) );
  NAND2_X2 U8453 ( .A1(REGFILE_reg_out_0__16_), .A2(net77310), .ZN(n7563) );
  NAND4_X2 U8454 ( .A1(n7566), .A2(n7565), .A3(n7564), .A4(n7563), .ZN(n7567)
         );
  NAND4_X2 U8455 ( .A1(n7572), .A2(n7571), .A3(n7570), .A4(n7569), .ZN(n8445)
         );
  MUX2_X2 U8456 ( .A(n8445), .B(instruction[16]), .S(net77276), .Z(aluA[16])
         );
  NAND2_X2 U8457 ( .A1(REGFILE_reg_out_30__15_), .A2(net77562), .ZN(n7576) );
  NAND2_X2 U8458 ( .A1(REGFILE_reg_out_31__15_), .A2(net77490), .ZN(n7574) );
  NAND2_X2 U8459 ( .A1(REGFILE_reg_out_29__15_), .A2(net77454), .ZN(n7573) );
  NAND4_X2 U8460 ( .A1(n7576), .A2(n7575), .A3(n7574), .A4(n7573), .ZN(n7582)
         );
  NAND2_X2 U8461 ( .A1(REGFILE_reg_out_26__15_), .A2(net77346), .ZN(n7578) );
  NAND2_X2 U8462 ( .A1(REGFILE_reg_out_24__15_), .A2(net77310), .ZN(n7577) );
  NAND4_X2 U8463 ( .A1(n7580), .A2(n7579), .A3(n7578), .A4(n7577), .ZN(n7581)
         );
  NAND2_X2 U8464 ( .A1(REGFILE_reg_out_17__15_), .A2(net77526), .ZN(n7585) );
  NAND2_X2 U8465 ( .A1(REGFILE_reg_out_23__15_), .A2(net77490), .ZN(n7584) );
  NAND2_X2 U8466 ( .A1(REGFILE_reg_out_21__15_), .A2(net77454), .ZN(n7583) );
  NAND4_X2 U8467 ( .A1(n7586), .A2(n7585), .A3(n7584), .A4(n7583), .ZN(n7592)
         );
  NAND2_X2 U8468 ( .A1(REGFILE_reg_out_19__15_), .A2(net77418), .ZN(n7590) );
  NAND2_X2 U8469 ( .A1(REGFILE_reg_out_20__15_), .A2(net77382), .ZN(n7589) );
  NAND4_X2 U8470 ( .A1(n7590), .A2(n7589), .A3(n7588), .A4(n7587), .ZN(n7591)
         );
  NAND2_X2 U8471 ( .A1(REGFILE_reg_out_14__15_), .A2(net77562), .ZN(n7596) );
  NAND2_X2 U8472 ( .A1(REGFILE_reg_out_9__15_), .A2(net77526), .ZN(n7595) );
  NAND2_X2 U8473 ( .A1(REGFILE_reg_out_15__15_), .A2(net77490), .ZN(n7594) );
  NAND4_X2 U8474 ( .A1(n7596), .A2(n7595), .A3(n7594), .A4(n7593), .ZN(n7602)
         );
  NAND2_X2 U8475 ( .A1(REGFILE_reg_out_11__15_), .A2(net77418), .ZN(n7600) );
  NAND2_X2 U8476 ( .A1(REGFILE_reg_out_10__15_), .A2(net77346), .ZN(n7598) );
  NAND2_X2 U8477 ( .A1(REGFILE_reg_out_8__15_), .A2(net77310), .ZN(n7597) );
  NAND4_X2 U8478 ( .A1(n7600), .A2(n7599), .A3(n7598), .A4(n7597), .ZN(n7601)
         );
  NAND2_X2 U8479 ( .A1(REGFILE_reg_out_6__15_), .A2(net77562), .ZN(n7606) );
  NAND2_X2 U8480 ( .A1(REGFILE_reg_out_7__15_), .A2(net77490), .ZN(n7604) );
  NAND4_X2 U8481 ( .A1(n7606), .A2(n7605), .A3(n7604), .A4(n7603), .ZN(n7612)
         );
  NAND2_X2 U8482 ( .A1(REGFILE_reg_out_4__15_), .A2(net77382), .ZN(n7609) );
  NAND2_X2 U8483 ( .A1(REGFILE_reg_out_0__15_), .A2(net77310), .ZN(n7607) );
  NAND4_X2 U8484 ( .A1(n7610), .A2(n7609), .A3(n7608), .A4(n7607), .ZN(n7611)
         );
  NAND4_X2 U8485 ( .A1(n7616), .A2(n7615), .A3(n7614), .A4(n7613), .ZN(n8446)
         );
  NAND2_X2 U8486 ( .A1(n8446), .A2(net77272), .ZN(n10463) );
  INV_X4 U8487 ( .A(n10463), .ZN(WIRE_ALU_A_MUX2TO1_32BIT_15__MUX_N1) );
  NAND2_X2 U8488 ( .A1(REGFILE_reg_out_30__14_), .A2(net77562), .ZN(n7620) );
  NAND2_X2 U8489 ( .A1(REGFILE_reg_out_31__14_), .A2(net77490), .ZN(n7618) );
  NAND2_X2 U8490 ( .A1(REGFILE_reg_out_29__14_), .A2(net77454), .ZN(n7617) );
  NAND4_X2 U8491 ( .A1(n7620), .A2(n7619), .A3(n7618), .A4(n7617), .ZN(n7626)
         );
  NAND2_X2 U8492 ( .A1(net77346), .A2(REGFILE_reg_out_26__14_), .ZN(n7622) );
  NAND2_X2 U8493 ( .A1(REGFILE_reg_out_24__14_), .A2(net77310), .ZN(n7621) );
  NAND4_X2 U8494 ( .A1(n7624), .A2(n7623), .A3(n7622), .A4(n7621), .ZN(n7625)
         );
  NAND2_X2 U8495 ( .A1(REGFILE_reg_out_22__14_), .A2(net77562), .ZN(n7630) );
  NAND2_X2 U8496 ( .A1(REGFILE_reg_out_17__14_), .A2(net77526), .ZN(n7629) );
  NAND2_X2 U8497 ( .A1(REGFILE_reg_out_23__14_), .A2(net77490), .ZN(n7628) );
  NAND2_X2 U8498 ( .A1(REGFILE_reg_out_21__14_), .A2(net77454), .ZN(n7627) );
  NAND4_X2 U8499 ( .A1(n7630), .A2(n7629), .A3(n7628), .A4(n7627), .ZN(n7636)
         );
  NAND2_X2 U8500 ( .A1(REGFILE_reg_out_19__14_), .A2(net77418), .ZN(n7634) );
  NAND2_X2 U8501 ( .A1(REGFILE_reg_out_16__14_), .A2(net77310), .ZN(n7631) );
  NAND4_X2 U8502 ( .A1(n7634), .A2(n7633), .A3(n7632), .A4(n7631), .ZN(n7635)
         );
  NAND2_X2 U8503 ( .A1(REGFILE_reg_out_14__14_), .A2(net77562), .ZN(n7640) );
  NAND2_X2 U8504 ( .A1(REGFILE_reg_out_9__14_), .A2(net77526), .ZN(n7639) );
  NAND2_X2 U8505 ( .A1(REGFILE_reg_out_15__14_), .A2(net77490), .ZN(n7638) );
  NAND2_X2 U8506 ( .A1(REGFILE_reg_out_13__14_), .A2(net77454), .ZN(n7637) );
  NAND4_X2 U8507 ( .A1(n7640), .A2(n7639), .A3(n7638), .A4(n7637), .ZN(n7646)
         );
  NAND2_X2 U8508 ( .A1(net77418), .A2(n5777), .ZN(n7644) );
  NAND4_X2 U8509 ( .A1(n7644), .A2(n7643), .A3(n7642), .A4(n7641), .ZN(n7645)
         );
  NAND2_X2 U8510 ( .A1(REGFILE_reg_out_6__14_), .A2(net77562), .ZN(n7650) );
  NAND2_X2 U8511 ( .A1(REGFILE_reg_out_1__14_), .A2(net77526), .ZN(n7649) );
  NAND2_X2 U8512 ( .A1(REGFILE_reg_out_7__14_), .A2(net77490), .ZN(n7648) );
  NAND2_X2 U8513 ( .A1(n5832), .A2(net77454), .ZN(n7647) );
  NAND4_X2 U8514 ( .A1(n7650), .A2(n7649), .A3(n7648), .A4(n7647), .ZN(n7656)
         );
  NAND2_X2 U8515 ( .A1(REGFILE_reg_out_4__14_), .A2(net77382), .ZN(n7653) );
  NAND4_X2 U8516 ( .A1(n7654), .A2(n7653), .A3(n7652), .A4(n7651), .ZN(n7655)
         );
  NAND4_X2 U8517 ( .A1(n7660), .A2(n7659), .A3(n7658), .A4(n7657), .ZN(n8438)
         );
  NAND2_X2 U8518 ( .A1(n8438), .A2(net77272), .ZN(n10247) );
  INV_X4 U8519 ( .A(n10247), .ZN(WIRE_ALU_A_MUX2TO1_32BIT_14__MUX_N1) );
  NAND2_X2 U8520 ( .A1(REGFILE_reg_out_25__13_), .A2(net77524), .ZN(n7663) );
  NAND2_X2 U8521 ( .A1(REGFILE_reg_out_31__13_), .A2(net77488), .ZN(n7662) );
  NAND2_X2 U8522 ( .A1(REGFILE_reg_out_29__13_), .A2(net77452), .ZN(n7661) );
  NAND4_X2 U8523 ( .A1(n7664), .A2(n7663), .A3(n7662), .A4(n7661), .ZN(n7670)
         );
  NAND2_X2 U8524 ( .A1(REGFILE_reg_out_27__13_), .A2(net77416), .ZN(n7668) );
  NAND4_X2 U8525 ( .A1(n7668), .A2(n7667), .A3(n7666), .A4(n7665), .ZN(n7669)
         );
  NAND2_X2 U8526 ( .A1(REGFILE_reg_out_22__13_), .A2(net77560), .ZN(n7674) );
  NAND2_X2 U8527 ( .A1(REGFILE_reg_out_17__13_), .A2(net77524), .ZN(n7673) );
  NAND2_X2 U8528 ( .A1(REGFILE_reg_out_23__13_), .A2(net77488), .ZN(n7672) );
  NAND2_X2 U8529 ( .A1(REGFILE_reg_out_21__13_), .A2(net77452), .ZN(n7671) );
  NAND4_X2 U8530 ( .A1(n7674), .A2(n7673), .A3(n7672), .A4(n7671), .ZN(n7680)
         );
  NAND2_X2 U8531 ( .A1(REGFILE_reg_out_19__13_), .A2(net77416), .ZN(n7678) );
  NAND2_X2 U8532 ( .A1(REGFILE_reg_out_20__13_), .A2(net77380), .ZN(n7677) );
  NAND4_X2 U8533 ( .A1(n7678), .A2(n7677), .A3(n7676), .A4(n7675), .ZN(n7679)
         );
  NAND2_X2 U8534 ( .A1(REGFILE_reg_out_9__13_), .A2(net77524), .ZN(n7683) );
  NAND2_X2 U8535 ( .A1(REGFILE_reg_out_15__13_), .A2(net77488), .ZN(n7682) );
  NAND2_X2 U8536 ( .A1(REGFILE_reg_out_13__13_), .A2(net77452), .ZN(n7681) );
  NAND4_X2 U8537 ( .A1(n7684), .A2(n7683), .A3(n7682), .A4(n7681), .ZN(n7690)
         );
  NAND2_X2 U8538 ( .A1(net148736), .A2(net77416), .ZN(n7688) );
  NAND4_X2 U8539 ( .A1(n7688), .A2(n7687), .A3(n7686), .A4(n7685), .ZN(n7689)
         );
  NAND2_X2 U8540 ( .A1(REGFILE_reg_out_7__13_), .A2(net77488), .ZN(n7692) );
  NAND2_X2 U8541 ( .A1(REGFILE_reg_out_5__13_), .A2(net77452), .ZN(n7691) );
  NAND4_X2 U8542 ( .A1(n7694), .A2(n7693), .A3(n7692), .A4(n7691), .ZN(n7700)
         );
  NAND2_X2 U8543 ( .A1(REGFILE_reg_out_3__13_), .A2(net77416), .ZN(n7698) );
  NAND2_X2 U8544 ( .A1(REGFILE_reg_out_4__13_), .A2(net77380), .ZN(n7697) );
  NAND2_X2 U8545 ( .A1(REGFILE_reg_out_0__13_), .A2(net77308), .ZN(n7695) );
  NAND4_X2 U8546 ( .A1(n7698), .A2(n7697), .A3(n7696), .A4(n7695), .ZN(n7699)
         );
  NAND4_X2 U8547 ( .A1(n7704), .A2(n7703), .A3(n7702), .A4(n7701), .ZN(n8437)
         );
  NAND2_X2 U8548 ( .A1(n8437), .A2(net77272), .ZN(n10368) );
  INV_X4 U8549 ( .A(n10368), .ZN(WIRE_ALU_A_MUX2TO1_32BIT_13__MUX_N1) );
  NAND2_X2 U8550 ( .A1(REGFILE_reg_out_30__12_), .A2(net77560), .ZN(n7708) );
  NAND2_X2 U8551 ( .A1(REGFILE_reg_out_25__12_), .A2(net77524), .ZN(n7707) );
  NAND2_X2 U8552 ( .A1(REGFILE_reg_out_31__12_), .A2(net77488), .ZN(n7706) );
  NAND2_X2 U8553 ( .A1(REGFILE_reg_out_29__12_), .A2(net77452), .ZN(n7705) );
  NAND4_X2 U8554 ( .A1(n7708), .A2(n7707), .A3(n7706), .A4(n7705), .ZN(n7714)
         );
  NAND2_X2 U8555 ( .A1(REGFILE_reg_out_27__12_), .A2(net77416), .ZN(n7712) );
  NAND2_X2 U8556 ( .A1(REGFILE_reg_out_26__12_), .A2(net77344), .ZN(n7710) );
  NAND2_X2 U8557 ( .A1(REGFILE_reg_out_24__12_), .A2(net77308), .ZN(n7709) );
  NAND4_X2 U8558 ( .A1(n7712), .A2(n7711), .A3(n7710), .A4(n7709), .ZN(n7713)
         );
  NAND2_X2 U8559 ( .A1(REGFILE_reg_out_22__12_), .A2(net77560), .ZN(n7718) );
  NAND2_X2 U8560 ( .A1(REGFILE_reg_out_17__12_), .A2(net77524), .ZN(n7717) );
  NAND2_X2 U8561 ( .A1(REGFILE_reg_out_23__12_), .A2(net77488), .ZN(n7716) );
  NAND2_X2 U8562 ( .A1(REGFILE_reg_out_21__12_), .A2(net77452), .ZN(n7715) );
  NAND4_X2 U8563 ( .A1(n7718), .A2(n7717), .A3(n7716), .A4(n7715), .ZN(n7724)
         );
  NAND2_X2 U8564 ( .A1(REGFILE_reg_out_19__12_), .A2(net77416), .ZN(n7722) );
  NAND2_X2 U8565 ( .A1(REGFILE_reg_out_20__12_), .A2(net77380), .ZN(n7721) );
  NAND2_X2 U8566 ( .A1(REGFILE_reg_out_18__12_), .A2(net77344), .ZN(n7720) );
  NAND2_X2 U8567 ( .A1(REGFILE_reg_out_16__12_), .A2(net77308), .ZN(n7719) );
  NAND4_X2 U8568 ( .A1(n7722), .A2(n7721), .A3(n7720), .A4(n7719), .ZN(n7723)
         );
  NAND2_X2 U8569 ( .A1(REGFILE_reg_out_14__12_), .A2(net77560), .ZN(n7728) );
  NAND2_X2 U8570 ( .A1(REGFILE_reg_out_9__12_), .A2(net77524), .ZN(n7727) );
  NAND4_X2 U8571 ( .A1(n7728), .A2(n7727), .A3(n7726), .A4(n7725), .ZN(n7734)
         );
  NAND2_X2 U8572 ( .A1(REGFILE_reg_out_11__12_), .A2(net77416), .ZN(n7732) );
  NAND2_X2 U8573 ( .A1(REGFILE_reg_out_10__12_), .A2(net77344), .ZN(n7730) );
  NAND4_X2 U8575 ( .A1(n7732), .A2(n7731), .A3(n7730), .A4(n7729), .ZN(n7733)
         );
  NAND2_X2 U8576 ( .A1(REGFILE_reg_out_6__12_), .A2(net77560), .ZN(n7738) );
  NAND2_X2 U8577 ( .A1(REGFILE_reg_out_1__12_), .A2(net77524), .ZN(n7737) );
  NAND2_X2 U8578 ( .A1(REGFILE_reg_out_7__12_), .A2(net77488), .ZN(n7736) );
  NAND2_X2 U8579 ( .A1(REGFILE_reg_out_5__12_), .A2(net77452), .ZN(n7735) );
  NAND4_X2 U8580 ( .A1(n7738), .A2(n7737), .A3(n7736), .A4(n7735), .ZN(n7744)
         );
  NAND2_X2 U8582 ( .A1(REGFILE_reg_out_4__12_), .A2(net77380), .ZN(n7741) );
  NAND2_X2 U8583 ( .A1(REGFILE_reg_out_2__12_), .A2(net77344), .ZN(n7740) );
  NAND2_X2 U8584 ( .A1(REGFILE_reg_out_0__12_), .A2(net77308), .ZN(n7739) );
  NAND4_X2 U8585 ( .A1(n7742), .A2(n7741), .A3(n7740), .A4(n7739), .ZN(n7743)
         );
  NAND4_X2 U8586 ( .A1(n7748), .A2(n7747), .A3(n7746), .A4(n7745), .ZN(n8436)
         );
  NAND2_X2 U8587 ( .A1(n8436), .A2(net77272), .ZN(n9075) );
  INV_X4 U8588 ( .A(n9075), .ZN(WIRE_ALU_A_MUX2TO1_32BIT_12__MUX_N1) );
  NAND2_X2 U8589 ( .A1(REGFILE_reg_out_30__11_), .A2(net77560), .ZN(n7752) );
  NAND2_X2 U8590 ( .A1(REGFILE_reg_out_25__11_), .A2(net77524), .ZN(n7751) );
  NAND2_X2 U8591 ( .A1(REGFILE_reg_out_31__11_), .A2(net77488), .ZN(n7750) );
  NAND2_X2 U8592 ( .A1(REGFILE_reg_out_29__11_), .A2(net77452), .ZN(n7749) );
  NAND4_X2 U8593 ( .A1(n7752), .A2(n7751), .A3(n7750), .A4(n7749), .ZN(n7758)
         );
  NAND2_X2 U8594 ( .A1(REGFILE_reg_out_26__11_), .A2(net77344), .ZN(n7754) );
  NAND2_X2 U8595 ( .A1(REGFILE_reg_out_24__11_), .A2(net77308), .ZN(n7753) );
  NAND4_X2 U8596 ( .A1(n7756), .A2(n7755), .A3(n7754), .A4(n7753), .ZN(n7757)
         );
  NAND2_X2 U8597 ( .A1(REGFILE_reg_out_22__11_), .A2(net77560), .ZN(n7762) );
  NAND2_X2 U8598 ( .A1(REGFILE_reg_out_17__11_), .A2(net77524), .ZN(n7761) );
  NAND2_X2 U8599 ( .A1(REGFILE_reg_out_23__11_), .A2(net77488), .ZN(n7760) );
  NAND2_X2 U8600 ( .A1(REGFILE_reg_out_21__11_), .A2(net77452), .ZN(n7759) );
  NAND4_X2 U8601 ( .A1(n7762), .A2(n7761), .A3(n7760), .A4(n7759), .ZN(n7768)
         );
  NAND2_X2 U8602 ( .A1(REGFILE_reg_out_19__11_), .A2(net77416), .ZN(n7766) );
  NAND2_X2 U8603 ( .A1(REGFILE_reg_out_20__11_), .A2(net77380), .ZN(n7765) );
  NAND2_X2 U8604 ( .A1(REGFILE_reg_out_18__11_), .A2(net77344), .ZN(n7764) );
  NAND2_X2 U8605 ( .A1(REGFILE_reg_out_16__11_), .A2(net77308), .ZN(n7763) );
  NAND4_X2 U8606 ( .A1(n7766), .A2(n7765), .A3(n7764), .A4(n7763), .ZN(n7767)
         );
  NAND2_X2 U8607 ( .A1(REGFILE_reg_out_14__11_), .A2(net77560), .ZN(n7772) );
  NAND2_X2 U8608 ( .A1(REGFILE_reg_out_9__11_), .A2(net77524), .ZN(n7771) );
  NAND2_X2 U8609 ( .A1(REGFILE_reg_out_15__11_), .A2(net77488), .ZN(n7770) );
  NAND4_X2 U8610 ( .A1(n7772), .A2(n7771), .A3(n7770), .A4(n7769), .ZN(n7778)
         );
  NAND2_X2 U8611 ( .A1(REGFILE_reg_out_11__11_), .A2(net77416), .ZN(n7776) );
  NAND2_X2 U8612 ( .A1(n5907), .A2(net77344), .ZN(n7774) );
  NAND2_X2 U8613 ( .A1(REGFILE_reg_out_8__11_), .A2(net77308), .ZN(n7773) );
  NAND4_X2 U8614 ( .A1(n7776), .A2(n7775), .A3(n7774), .A4(n7773), .ZN(n7777)
         );
  NAND2_X2 U8615 ( .A1(REGFILE_reg_out_6__11_), .A2(net77560), .ZN(n7782) );
  NAND2_X2 U8616 ( .A1(REGFILE_reg_out_1__11_), .A2(net77524), .ZN(n7781) );
  NAND2_X2 U8617 ( .A1(REGFILE_reg_out_7__11_), .A2(net77488), .ZN(n7780) );
  NAND2_X2 U8618 ( .A1(REGFILE_reg_out_5__11_), .A2(net77452), .ZN(n7779) );
  NAND4_X2 U8619 ( .A1(n7782), .A2(n7781), .A3(n7780), .A4(n7779), .ZN(n7788)
         );
  NAND2_X2 U8620 ( .A1(REGFILE_reg_out_3__11_), .A2(net77416), .ZN(n7786) );
  NAND2_X2 U8621 ( .A1(REGFILE_reg_out_4__11_), .A2(net77380), .ZN(n7785) );
  NAND2_X2 U8622 ( .A1(net77344), .A2(REGFILE_reg_out_2__11_), .ZN(n7784) );
  NAND2_X2 U8623 ( .A1(REGFILE_reg_out_0__11_), .A2(net77308), .ZN(n7783) );
  NAND4_X2 U8624 ( .A1(n7786), .A2(n7785), .A3(n7784), .A4(n7783), .ZN(n7787)
         );
  NAND4_X2 U8625 ( .A1(n7792), .A2(n7791), .A3(n7790), .A4(n7789), .ZN(n8435)
         );
  NAND2_X2 U8626 ( .A1(n8435), .A2(net77272), .ZN(n10375) );
  INV_X4 U8627 ( .A(n10375), .ZN(WIRE_ALU_A_MUX2TO1_32BIT_11__MUX_N1) );
  NAND2_X2 U8628 ( .A1(REGFILE_reg_out_30__10_), .A2(net77558), .ZN(n7796) );
  NAND2_X2 U8629 ( .A1(REGFILE_reg_out_31__10_), .A2(net77482), .ZN(n7794) );
  NAND2_X2 U8630 ( .A1(REGFILE_reg_out_29__10_), .A2(net77456), .ZN(n7793) );
  NAND4_X2 U8631 ( .A1(n7796), .A2(n7795), .A3(n7794), .A4(n7793), .ZN(n7802)
         );
  NAND2_X2 U8632 ( .A1(REGFILE_reg_out_27__10_), .A2(net77414), .ZN(n7800) );
  NAND2_X2 U8633 ( .A1(REGFILE_reg_out_28__10_), .A2(net77376), .ZN(n7799) );
  NAND2_X2 U8634 ( .A1(REGFILE_reg_out_26__10_), .A2(net77342), .ZN(n7798) );
  NAND2_X2 U8635 ( .A1(REGFILE_reg_out_24__10_), .A2(net77306), .ZN(n7797) );
  NAND4_X2 U8636 ( .A1(n7800), .A2(n7799), .A3(n7798), .A4(n7797), .ZN(n7801)
         );
  NAND2_X2 U8637 ( .A1(REGFILE_reg_out_22__10_), .A2(net77558), .ZN(n7806) );
  NAND2_X2 U8638 ( .A1(REGFILE_reg_out_17__10_), .A2(net77522), .ZN(n7805) );
  NAND2_X2 U8639 ( .A1(REGFILE_reg_out_23__10_), .A2(net77482), .ZN(n7804) );
  NAND2_X2 U8640 ( .A1(REGFILE_reg_out_21__10_), .A2(net77456), .ZN(n7803) );
  NAND4_X2 U8641 ( .A1(n7806), .A2(n7805), .A3(n7804), .A4(n7803), .ZN(n7812)
         );
  NAND2_X2 U8642 ( .A1(REGFILE_reg_out_19__10_), .A2(net77414), .ZN(n7810) );
  NAND2_X2 U8643 ( .A1(REGFILE_reg_out_20__10_), .A2(net77376), .ZN(n7809) );
  NAND2_X2 U8644 ( .A1(REGFILE_reg_out_18__10_), .A2(net77342), .ZN(n7808) );
  NAND2_X2 U8645 ( .A1(REGFILE_reg_out_16__10_), .A2(net77306), .ZN(n7807) );
  NAND4_X2 U8646 ( .A1(n7810), .A2(n7809), .A3(n7808), .A4(n7807), .ZN(n7811)
         );
  NAND2_X2 U8647 ( .A1(REGFILE_reg_out_14__10_), .A2(net77558), .ZN(n7816) );
  NAND2_X2 U8648 ( .A1(REGFILE_reg_out_9__10_), .A2(net77522), .ZN(n7815) );
  NAND4_X2 U8649 ( .A1(n7816), .A2(n7815), .A3(n7814), .A4(n7813), .ZN(n7822)
         );
  NAND2_X2 U8650 ( .A1(REGFILE_reg_out_11__10_), .A2(net77414), .ZN(n7820) );
  NAND2_X2 U8651 ( .A1(REGFILE_reg_out_10__10_), .A2(net77342), .ZN(n7818) );
  NAND2_X2 U8652 ( .A1(REGFILE_reg_out_8__10_), .A2(net77306), .ZN(n7817) );
  NAND4_X2 U8653 ( .A1(n7820), .A2(n7819), .A3(n7818), .A4(n7817), .ZN(n7821)
         );
  NAND2_X2 U8654 ( .A1(REGFILE_reg_out_6__10_), .A2(net77558), .ZN(n7826) );
  NAND2_X2 U8655 ( .A1(REGFILE_reg_out_1__10_), .A2(net77522), .ZN(n7825) );
  NAND2_X2 U8656 ( .A1(REGFILE_reg_out_7__10_), .A2(net77482), .ZN(n7824) );
  NAND2_X2 U8657 ( .A1(REGFILE_reg_out_5__10_), .A2(net77456), .ZN(n7823) );
  NAND4_X2 U8658 ( .A1(n7826), .A2(n7825), .A3(n7824), .A4(n7823), .ZN(n7832)
         );
  NAND2_X2 U8659 ( .A1(REGFILE_reg_out_4__10_), .A2(net77376), .ZN(n7829) );
  NAND2_X2 U8660 ( .A1(REGFILE_reg_out_0__10_), .A2(net77306), .ZN(n7827) );
  NAND4_X2 U8661 ( .A1(n7830), .A2(n7829), .A3(n7828), .A4(n7827), .ZN(n7831)
         );
  NAND4_X2 U8662 ( .A1(n7836), .A2(n7835), .A3(n7834), .A4(n7833), .ZN(n8434)
         );
  NAND2_X2 U8663 ( .A1(n8434), .A2(net77272), .ZN(n10125) );
  INV_X4 U8664 ( .A(n10125), .ZN(WIRE_ALU_A_MUX2TO1_32BIT_10__MUX_N1) );
  NAND2_X2 U8665 ( .A1(REGFILE_reg_out_30__9_), .A2(net77558), .ZN(n7840) );
  NAND2_X2 U8666 ( .A1(REGFILE_reg_out_31__9_), .A2(net77482), .ZN(n7838) );
  NAND2_X2 U8667 ( .A1(REGFILE_reg_out_29__9_), .A2(net77456), .ZN(n7837) );
  NAND4_X2 U8668 ( .A1(n7840), .A2(n7839), .A3(n7838), .A4(n7837), .ZN(n7846)
         );
  NAND2_X2 U8669 ( .A1(REGFILE_reg_out_27__9_), .A2(net77414), .ZN(n7844) );
  NAND2_X2 U8670 ( .A1(REGFILE_reg_out_28__9_), .A2(net77376), .ZN(n7843) );
  NAND2_X2 U8671 ( .A1(REGFILE_reg_out_26__9_), .A2(net77342), .ZN(n7842) );
  NAND2_X2 U8672 ( .A1(REGFILE_reg_out_24__9_), .A2(net77306), .ZN(n7841) );
  NAND4_X2 U8673 ( .A1(n7844), .A2(n7843), .A3(n7842), .A4(n7841), .ZN(n7845)
         );
  NAND2_X2 U8674 ( .A1(REGFILE_reg_out_22__9_), .A2(net77558), .ZN(n7850) );
  NAND2_X2 U8675 ( .A1(REGFILE_reg_out_17__9_), .A2(net77522), .ZN(n7849) );
  NAND2_X2 U8676 ( .A1(REGFILE_reg_out_23__9_), .A2(net77482), .ZN(n7848) );
  NAND2_X2 U8677 ( .A1(REGFILE_reg_out_21__9_), .A2(net77456), .ZN(n7847) );
  NAND4_X2 U8678 ( .A1(n7850), .A2(n7849), .A3(n7848), .A4(n7847), .ZN(n7856)
         );
  NAND2_X2 U8679 ( .A1(REGFILE_reg_out_19__9_), .A2(net77414), .ZN(n7854) );
  NAND2_X2 U8680 ( .A1(REGFILE_reg_out_20__9_), .A2(net77376), .ZN(n7853) );
  NAND2_X2 U8681 ( .A1(REGFILE_reg_out_18__9_), .A2(net77342), .ZN(n7852) );
  NAND2_X2 U8682 ( .A1(REGFILE_reg_out_16__9_), .A2(net77306), .ZN(n7851) );
  NAND4_X2 U8683 ( .A1(n7854), .A2(n7853), .A3(n7852), .A4(n7851), .ZN(n7855)
         );
  NAND2_X2 U8684 ( .A1(REGFILE_reg_out_14__9_), .A2(net77558), .ZN(n7860) );
  NAND2_X2 U8685 ( .A1(REGFILE_reg_out_9__9_), .A2(net77522), .ZN(n7859) );
  NAND2_X2 U8686 ( .A1(REGFILE_reg_out_15__9_), .A2(net77482), .ZN(n7858) );
  NAND2_X2 U8687 ( .A1(REGFILE_reg_out_13__9_), .A2(net77456), .ZN(n7857) );
  NAND4_X2 U8688 ( .A1(n7860), .A2(n7859), .A3(n7858), .A4(n7857), .ZN(n7866)
         );
  NAND2_X2 U8689 ( .A1(REGFILE_reg_out_11__9_), .A2(net77414), .ZN(n7864) );
  NAND2_X2 U8690 ( .A1(net77376), .A2(REGFILE_reg_out_12__9_), .ZN(n7863) );
  NAND2_X2 U8691 ( .A1(REGFILE_reg_out_10__9_), .A2(net77342), .ZN(n7862) );
  NAND2_X2 U8692 ( .A1(REGFILE_reg_out_8__9_), .A2(net77306), .ZN(n7861) );
  NAND4_X2 U8693 ( .A1(n7864), .A2(n7863), .A3(n7862), .A4(n7861), .ZN(n7865)
         );
  NAND2_X2 U8694 ( .A1(REGFILE_reg_out_6__9_), .A2(net77558), .ZN(n7870) );
  NAND2_X2 U8695 ( .A1(REGFILE_reg_out_1__9_), .A2(net77522), .ZN(n7869) );
  NAND2_X2 U8696 ( .A1(REGFILE_reg_out_7__9_), .A2(net77482), .ZN(n7868) );
  NAND2_X2 U8697 ( .A1(REGFILE_reg_out_5__9_), .A2(net77456), .ZN(n7867) );
  NAND4_X2 U8698 ( .A1(n7870), .A2(n7869), .A3(n7868), .A4(n7867), .ZN(n7876)
         );
  NAND2_X2 U8699 ( .A1(REGFILE_reg_out_3__9_), .A2(net77414), .ZN(n7874) );
  NAND2_X2 U8700 ( .A1(REGFILE_reg_out_4__9_), .A2(net77376), .ZN(n7873) );
  NAND2_X2 U8701 ( .A1(REGFILE_reg_out_0__9_), .A2(net77306), .ZN(n7871) );
  NAND4_X2 U8702 ( .A1(n7874), .A2(n7873), .A3(n7872), .A4(n7871), .ZN(n7875)
         );
  NAND4_X2 U8703 ( .A1(n7880), .A2(n7879), .A3(n7878), .A4(n7877), .ZN(n8430)
         );
  NAND2_X2 U8704 ( .A1(n8430), .A2(net77272), .ZN(n10382) );
  INV_X4 U8705 ( .A(n10382), .ZN(WIRE_ALU_A_MUX2TO1_32BIT_9__MUX_N1) );
  NAND2_X2 U8706 ( .A1(REGFILE_reg_out_30__8_), .A2(net77558), .ZN(n7884) );
  NAND2_X2 U8707 ( .A1(REGFILE_reg_out_31__8_), .A2(net77482), .ZN(n7882) );
  NAND2_X2 U8708 ( .A1(REGFILE_reg_out_29__8_), .A2(net77456), .ZN(n7881) );
  NAND4_X2 U8709 ( .A1(n7884), .A2(n7883), .A3(n7882), .A4(n7881), .ZN(n7890)
         );
  NAND2_X2 U8710 ( .A1(REGFILE_reg_out_28__8_), .A2(net77376), .ZN(n7887) );
  NAND2_X2 U8711 ( .A1(REGFILE_reg_out_26__8_), .A2(net77342), .ZN(n7886) );
  NAND2_X2 U8712 ( .A1(REGFILE_reg_out_24__8_), .A2(net77306), .ZN(n7885) );
  NAND4_X2 U8713 ( .A1(n7888), .A2(n7887), .A3(n7886), .A4(n7885), .ZN(n7889)
         );
  NAND2_X2 U8714 ( .A1(REGFILE_reg_out_22__8_), .A2(net77558), .ZN(n7894) );
  NAND2_X2 U8715 ( .A1(REGFILE_reg_out_17__8_), .A2(net77522), .ZN(n7893) );
  NAND2_X2 U8716 ( .A1(REGFILE_reg_out_23__8_), .A2(net77482), .ZN(n7892) );
  NAND2_X2 U8717 ( .A1(REGFILE_reg_out_21__8_), .A2(net77456), .ZN(n7891) );
  NAND4_X2 U8718 ( .A1(n7894), .A2(n7893), .A3(n7892), .A4(n7891), .ZN(n7900)
         );
  NAND2_X2 U8719 ( .A1(REGFILE_reg_out_19__8_), .A2(net77414), .ZN(n7898) );
  NAND2_X2 U8720 ( .A1(REGFILE_reg_out_20__8_), .A2(net77376), .ZN(n7897) );
  NAND2_X2 U8721 ( .A1(REGFILE_reg_out_18__8_), .A2(net77342), .ZN(n7896) );
  NAND2_X2 U8722 ( .A1(REGFILE_reg_out_16__8_), .A2(net77306), .ZN(n7895) );
  NAND4_X2 U8723 ( .A1(n7898), .A2(n7897), .A3(n7896), .A4(n7895), .ZN(n7899)
         );
  NAND2_X2 U8724 ( .A1(REGFILE_reg_out_14__8_), .A2(net77558), .ZN(n7904) );
  NAND2_X2 U8725 ( .A1(REGFILE_reg_out_9__8_), .A2(net77522), .ZN(n7903) );
  NAND2_X2 U8726 ( .A1(REGFILE_reg_out_15__8_), .A2(net77482), .ZN(n7902) );
  NAND2_X2 U8727 ( .A1(REGFILE_reg_out_13__8_), .A2(net77456), .ZN(n7901) );
  NAND4_X2 U8728 ( .A1(n7904), .A2(n7903), .A3(n7902), .A4(n7901), .ZN(n7910)
         );
  NAND2_X2 U8729 ( .A1(REGFILE_reg_out_11__8_), .A2(net77414), .ZN(n7908) );
  NAND2_X2 U8730 ( .A1(REGFILE_reg_out_12__8_), .A2(net77376), .ZN(n7907) );
  NAND2_X2 U8731 ( .A1(REGFILE_reg_out_10__8_), .A2(net77342), .ZN(n7906) );
  NAND2_X2 U8732 ( .A1(REGFILE_reg_out_8__8_), .A2(net77306), .ZN(n7905) );
  NAND4_X2 U8733 ( .A1(n7908), .A2(n7907), .A3(n7906), .A4(n7905), .ZN(n7909)
         );
  NAND2_X2 U8734 ( .A1(REGFILE_reg_out_6__8_), .A2(net77558), .ZN(n7914) );
  NAND2_X2 U8735 ( .A1(REGFILE_reg_out_1__8_), .A2(net77522), .ZN(n7913) );
  NAND2_X2 U8736 ( .A1(REGFILE_reg_out_7__8_), .A2(net77482), .ZN(n7912) );
  NAND2_X2 U8737 ( .A1(REGFILE_reg_out_5__8_), .A2(net77456), .ZN(n7911) );
  NAND4_X2 U8738 ( .A1(n7914), .A2(n7913), .A3(n7912), .A4(n7911), .ZN(n7920)
         );
  NAND2_X2 U8739 ( .A1(REGFILE_reg_out_4__8_), .A2(net77376), .ZN(n7917) );
  NAND2_X2 U8740 ( .A1(REGFILE_reg_out_0__8_), .A2(net77306), .ZN(n7915) );
  NAND4_X2 U8741 ( .A1(n7918), .A2(n7917), .A3(n7916), .A4(n7915), .ZN(n7919)
         );
  NAND4_X2 U8742 ( .A1(n7924), .A2(n7923), .A3(n7922), .A4(n7921), .ZN(n8431)
         );
  NAND2_X2 U8743 ( .A1(n8431), .A2(net77272), .ZN(n9535) );
  INV_X4 U8744 ( .A(n9535), .ZN(WIRE_ALU_A_MUX2TO1_32BIT_8__MUX_N1) );
  NAND2_X2 U8745 ( .A1(REGFILE_reg_out_30__7_), .A2(net77556), .ZN(n7928) );
  NAND2_X2 U8746 ( .A1(REGFILE_reg_out_31__7_), .A2(net77484), .ZN(n7926) );
  NAND2_X2 U8747 ( .A1(REGFILE_reg_out_29__7_), .A2(net77456), .ZN(n7925) );
  NAND4_X2 U8748 ( .A1(n7928), .A2(n7927), .A3(n7926), .A4(n7925), .ZN(n7934)
         );
  NAND2_X2 U8749 ( .A1(REGFILE_reg_out_28__7_), .A2(net77376), .ZN(n7931) );
  NAND2_X2 U8750 ( .A1(REGFILE_reg_out_26__7_), .A2(net77338), .ZN(n7930) );
  NAND2_X2 U8751 ( .A1(REGFILE_reg_out_24__7_), .A2(net77304), .ZN(n7929) );
  NAND4_X2 U8752 ( .A1(n7932), .A2(n7931), .A3(n7930), .A4(n7929), .ZN(n7933)
         );
  NAND2_X2 U8753 ( .A1(REGFILE_reg_out_22__7_), .A2(net77556), .ZN(n7938) );
  NAND2_X2 U8754 ( .A1(REGFILE_reg_out_17__7_), .A2(net77520), .ZN(n7937) );
  NAND2_X2 U8755 ( .A1(REGFILE_reg_out_23__7_), .A2(net77484), .ZN(n7936) );
  NAND2_X2 U8756 ( .A1(REGFILE_reg_out_21__7_), .A2(net77456), .ZN(n7935) );
  NAND4_X2 U8757 ( .A1(n7938), .A2(n7937), .A3(n7936), .A4(n7935), .ZN(n7944)
         );
  NAND2_X2 U8758 ( .A1(REGFILE_reg_out_19__7_), .A2(net77410), .ZN(n7942) );
  NAND2_X2 U8759 ( .A1(REGFILE_reg_out_20__7_), .A2(net77376), .ZN(n7941) );
  NAND2_X2 U8760 ( .A1(REGFILE_reg_out_18__7_), .A2(net77338), .ZN(n7940) );
  NAND2_X2 U8761 ( .A1(REGFILE_reg_out_16__7_), .A2(net77304), .ZN(n7939) );
  NAND4_X2 U8762 ( .A1(n7942), .A2(n7941), .A3(n7940), .A4(n7939), .ZN(n7943)
         );
  NAND2_X2 U8763 ( .A1(REGFILE_reg_out_14__7_), .A2(net77556), .ZN(n7948) );
  NAND2_X2 U8764 ( .A1(REGFILE_reg_out_9__7_), .A2(net77520), .ZN(n7947) );
  NAND2_X2 U8765 ( .A1(REGFILE_reg_out_15__7_), .A2(net77484), .ZN(n7946) );
  NAND2_X2 U8766 ( .A1(REGFILE_reg_out_13__7_), .A2(net77456), .ZN(n7945) );
  NAND4_X2 U8767 ( .A1(n7948), .A2(n7947), .A3(n7946), .A4(n7945), .ZN(n7954)
         );
  NAND2_X2 U8768 ( .A1(REGFILE_reg_out_11__7_), .A2(net77410), .ZN(n7952) );
  NAND2_X2 U8769 ( .A1(REGFILE_reg_out_12__7_), .A2(net77376), .ZN(n7951) );
  NAND2_X2 U8770 ( .A1(REGFILE_reg_out_8__7_), .A2(net77304), .ZN(n7949) );
  NAND4_X2 U8771 ( .A1(n7952), .A2(n7951), .A3(n7950), .A4(n7949), .ZN(n7953)
         );
  NAND2_X2 U8772 ( .A1(REGFILE_reg_out_1__7_), .A2(net77520), .ZN(n7956) );
  NAND2_X2 U8773 ( .A1(REGFILE_reg_out_5__7_), .A2(net77456), .ZN(n7955) );
  NAND4_X2 U8774 ( .A1(net74359), .A2(n7956), .A3(net74361), .A4(n7955), .ZN(
        n7962) );
  NAND2_X2 U8775 ( .A1(REGFILE_reg_out_3__7_), .A2(net77410), .ZN(n7960) );
  NAND2_X2 U8776 ( .A1(REGFILE_reg_out_4__7_), .A2(net77376), .ZN(n7959) );
  NAND2_X2 U8777 ( .A1(REGFILE_reg_out_0__7_), .A2(net77304), .ZN(n7957) );
  NAND4_X2 U8778 ( .A1(n7960), .A2(n7959), .A3(n7958), .A4(n7957), .ZN(n7961)
         );
  NAND4_X2 U8779 ( .A1(n7966), .A2(n7965), .A3(n7964), .A4(n7963), .ZN(n8432)
         );
  NAND2_X2 U8780 ( .A1(n8432), .A2(net77272), .ZN(n10464) );
  INV_X4 U8781 ( .A(n10464), .ZN(WIRE_ALU_A_MUX2TO1_32BIT_7__MUX_N1) );
  NAND2_X2 U8782 ( .A1(REGFILE_reg_out_30__6_), .A2(net77556), .ZN(n7970) );
  NAND2_X2 U8783 ( .A1(n5764), .A2(net77520), .ZN(n7969) );
  NAND2_X2 U8784 ( .A1(REGFILE_reg_out_31__6_), .A2(net77484), .ZN(n7968) );
  NAND2_X2 U8785 ( .A1(REGFILE_reg_out_29__6_), .A2(net77456), .ZN(n7967) );
  NAND4_X2 U8786 ( .A1(n7970), .A2(n7969), .A3(n7968), .A4(n7967), .ZN(n7976)
         );
  NAND2_X2 U8787 ( .A1(REGFILE_reg_out_27__6_), .A2(net77410), .ZN(n7974) );
  NAND2_X2 U8788 ( .A1(REGFILE_reg_out_28__6_), .A2(net77376), .ZN(n7973) );
  NAND2_X2 U8789 ( .A1(REGFILE_reg_out_26__6_), .A2(net77338), .ZN(n7972) );
  NAND2_X2 U8790 ( .A1(REGFILE_reg_out_24__6_), .A2(net77304), .ZN(n7971) );
  NAND4_X2 U8791 ( .A1(n7974), .A2(n7973), .A3(n7972), .A4(n7971), .ZN(n7975)
         );
  NAND2_X2 U8792 ( .A1(REGFILE_reg_out_22__6_), .A2(net77556), .ZN(n7980) );
  NAND2_X2 U8793 ( .A1(REGFILE_reg_out_17__6_), .A2(net77520), .ZN(n7979) );
  NAND2_X2 U8794 ( .A1(REGFILE_reg_out_23__6_), .A2(net77484), .ZN(n7978) );
  NAND2_X2 U8795 ( .A1(REGFILE_reg_out_21__6_), .A2(net77456), .ZN(n7977) );
  NAND4_X2 U8796 ( .A1(n7980), .A2(n7979), .A3(n7978), .A4(n7977), .ZN(n7986)
         );
  NAND2_X2 U8797 ( .A1(REGFILE_reg_out_19__6_), .A2(net77410), .ZN(n7984) );
  NAND2_X2 U8798 ( .A1(REGFILE_reg_out_20__6_), .A2(net77376), .ZN(n7983) );
  NAND2_X2 U8799 ( .A1(REGFILE_reg_out_18__6_), .A2(net77338), .ZN(n7982) );
  NAND2_X2 U8800 ( .A1(REGFILE_reg_out_16__6_), .A2(net77304), .ZN(n7981) );
  NAND4_X2 U8801 ( .A1(n7984), .A2(n7983), .A3(n7982), .A4(n7981), .ZN(n7985)
         );
  NAND2_X2 U8802 ( .A1(REGFILE_reg_out_14__6_), .A2(net77556), .ZN(n7990) );
  NAND2_X2 U8803 ( .A1(REGFILE_reg_out_9__6_), .A2(net77520), .ZN(n7989) );
  NAND2_X2 U8804 ( .A1(REGFILE_reg_out_13__6_), .A2(net77456), .ZN(n7987) );
  NAND4_X2 U8805 ( .A1(n7990), .A2(n7989), .A3(n7988), .A4(n7987), .ZN(n7996)
         );
  NAND2_X2 U8806 ( .A1(REGFILE_reg_out_11__6_), .A2(net77410), .ZN(n7994) );
  NAND2_X2 U8807 ( .A1(REGFILE_reg_out_12__6_), .A2(net77376), .ZN(n7993) );
  NAND2_X2 U8808 ( .A1(n5902), .A2(net77338), .ZN(n7992) );
  NAND2_X2 U8809 ( .A1(REGFILE_reg_out_8__6_), .A2(net77304), .ZN(n7991) );
  NAND4_X2 U8810 ( .A1(n7994), .A2(n7993), .A3(n7992), .A4(n7991), .ZN(n7995)
         );
  NAND2_X2 U8811 ( .A1(REGFILE_reg_out_6__6_), .A2(net77556), .ZN(n8000) );
  NAND2_X2 U8812 ( .A1(REGFILE_reg_out_1__6_), .A2(net77520), .ZN(n7999) );
  NAND2_X2 U8813 ( .A1(REGFILE_reg_out_7__6_), .A2(net77484), .ZN(n7998) );
  NAND2_X2 U8814 ( .A1(REGFILE_reg_out_5__6_), .A2(net77456), .ZN(n7997) );
  NAND4_X2 U8815 ( .A1(n8000), .A2(n7999), .A3(n7998), .A4(n7997), .ZN(n8006)
         );
  NAND2_X2 U8816 ( .A1(REGFILE_reg_out_3__6_), .A2(net77410), .ZN(n8004) );
  NAND2_X2 U8817 ( .A1(REGFILE_reg_out_4__6_), .A2(net77376), .ZN(n8003) );
  NAND2_X2 U8818 ( .A1(REGFILE_reg_out_2__6_), .A2(net77338), .ZN(n8002) );
  NAND2_X2 U8819 ( .A1(REGFILE_reg_out_0__6_), .A2(net77304), .ZN(n8001) );
  NAND4_X2 U8820 ( .A1(n8004), .A2(n8003), .A3(n8002), .A4(n8001), .ZN(n8005)
         );
  NAND4_X2 U8821 ( .A1(n8010), .A2(n8009), .A3(n8008), .A4(n8007), .ZN(n8433)
         );
  NAND2_X2 U8822 ( .A1(n8433), .A2(net77272), .ZN(n9656) );
  INV_X4 U8823 ( .A(n9656), .ZN(WIRE_ALU_A_MUX2TO1_32BIT_6__MUX_N1) );
  NAND2_X2 U8824 ( .A1(REGFILE_reg_out_30__5_), .A2(net77556), .ZN(n8014) );
  NAND2_X2 U8825 ( .A1(REGFILE_reg_out_25__5_), .A2(net77520), .ZN(n8013) );
  NAND2_X2 U8826 ( .A1(REGFILE_reg_out_31__5_), .A2(net77484), .ZN(n8012) );
  NAND2_X2 U8827 ( .A1(REGFILE_reg_out_29__5_), .A2(net77456), .ZN(n8011) );
  NAND4_X2 U8828 ( .A1(n8014), .A2(n8013), .A3(n8012), .A4(n8011), .ZN(n8020)
         );
  NAND2_X2 U8829 ( .A1(REGFILE_reg_out_27__5_), .A2(net77410), .ZN(n8018) );
  NAND2_X2 U8830 ( .A1(REGFILE_reg_out_28__5_), .A2(net77376), .ZN(n8017) );
  NAND2_X2 U8831 ( .A1(REGFILE_reg_out_26__5_), .A2(net77338), .ZN(n8016) );
  NAND2_X2 U8832 ( .A1(REGFILE_reg_out_24__5_), .A2(net77304), .ZN(n8015) );
  NAND4_X2 U8833 ( .A1(n8018), .A2(n8017), .A3(n8016), .A4(n8015), .ZN(n8019)
         );
  NAND2_X2 U8834 ( .A1(REGFILE_reg_out_22__5_), .A2(net77556), .ZN(n8024) );
  NAND2_X2 U8835 ( .A1(REGFILE_reg_out_17__5_), .A2(net77520), .ZN(n8023) );
  NAND2_X2 U8836 ( .A1(REGFILE_reg_out_23__5_), .A2(net77484), .ZN(n8022) );
  NAND2_X2 U8837 ( .A1(REGFILE_reg_out_21__5_), .A2(net77456), .ZN(n8021) );
  NAND4_X2 U8838 ( .A1(n8024), .A2(n8023), .A3(n8022), .A4(n8021), .ZN(n8030)
         );
  NAND2_X2 U8839 ( .A1(REGFILE_reg_out_19__5_), .A2(net77410), .ZN(n8028) );
  NAND2_X2 U8840 ( .A1(REGFILE_reg_out_20__5_), .A2(net77376), .ZN(n8027) );
  NAND2_X2 U8841 ( .A1(REGFILE_reg_out_18__5_), .A2(net77338), .ZN(n8026) );
  NAND2_X2 U8842 ( .A1(REGFILE_reg_out_16__5_), .A2(net77304), .ZN(n8025) );
  NAND4_X2 U8843 ( .A1(n8028), .A2(n8027), .A3(n8026), .A4(n8025), .ZN(n8029)
         );
  NAND2_X2 U8844 ( .A1(REGFILE_reg_out_14__5_), .A2(net77556), .ZN(n8034) );
  NAND2_X2 U8845 ( .A1(REGFILE_reg_out_9__5_), .A2(net77520), .ZN(n8033) );
  NAND2_X2 U8846 ( .A1(REGFILE_reg_out_15__5_), .A2(net77484), .ZN(n8032) );
  NAND2_X2 U8847 ( .A1(REGFILE_reg_out_13__5_), .A2(net77456), .ZN(n8031) );
  NAND4_X2 U8848 ( .A1(n8034), .A2(n8033), .A3(n8032), .A4(n8031), .ZN(n8040)
         );
  NAND2_X2 U8849 ( .A1(REGFILE_reg_out_11__5_), .A2(net77410), .ZN(n8038) );
  NAND2_X2 U8850 ( .A1(REGFILE_reg_out_12__5_), .A2(net77376), .ZN(n8037) );
  NAND2_X2 U8851 ( .A1(REGFILE_reg_out_8__5_), .A2(net77304), .ZN(n8035) );
  NAND4_X2 U8852 ( .A1(n8038), .A2(n8037), .A3(n8036), .A4(n8035), .ZN(n8039)
         );
  NAND2_X2 U8853 ( .A1(REGFILE_reg_out_6__5_), .A2(net77556), .ZN(n8044) );
  NAND2_X2 U8854 ( .A1(REGFILE_reg_out_1__5_), .A2(net77520), .ZN(n8043) );
  NAND2_X2 U8855 ( .A1(REGFILE_reg_out_7__5_), .A2(net77484), .ZN(n8042) );
  NAND4_X2 U8856 ( .A1(n8044), .A2(n8043), .A3(n8042), .A4(n8041), .ZN(n8050)
         );
  NAND2_X2 U8857 ( .A1(REGFILE_reg_out_3__5_), .A2(net77410), .ZN(n8048) );
  NAND2_X2 U8858 ( .A1(REGFILE_reg_out_4__5_), .A2(net77376), .ZN(n8047) );
  NAND2_X2 U8859 ( .A1(REGFILE_reg_out_0__5_), .A2(net77304), .ZN(n8045) );
  NAND4_X2 U8860 ( .A1(n8048), .A2(n8047), .A3(n8046), .A4(n8045), .ZN(n8049)
         );
  NAND4_X2 U8861 ( .A1(n8054), .A2(n8053), .A3(n8052), .A4(n8051), .ZN(n8424)
         );
  NAND2_X2 U8862 ( .A1(n8424), .A2(n4866), .ZN(n10396) );
  INV_X4 U8863 ( .A(n10396), .ZN(WIRE_ALU_A_MUX2TO1_32BIT_5__MUX_N1) );
  NAND2_X2 U8864 ( .A1(REGFILE_reg_out_30__4_), .A2(net77554), .ZN(n8058) );
  NAND2_X2 U8865 ( .A1(REGFILE_reg_out_25__4_), .A2(net77518), .ZN(n8057) );
  NAND2_X2 U8866 ( .A1(REGFILE_reg_out_31__4_), .A2(net77482), .ZN(n8056) );
  NAND2_X2 U8867 ( .A1(REGFILE_reg_out_29__4_), .A2(net77456), .ZN(n8055) );
  NAND4_X2 U8868 ( .A1(n8058), .A2(n8057), .A3(n8056), .A4(n8055), .ZN(n8064)
         );
  NAND2_X2 U8869 ( .A1(REGFILE_reg_out_27__4_), .A2(net77410), .ZN(n8062) );
  NAND2_X2 U8870 ( .A1(REGFILE_reg_out_28__4_), .A2(net77376), .ZN(n8061) );
  NAND2_X2 U8871 ( .A1(REGFILE_reg_out_26__4_), .A2(net77338), .ZN(n8060) );
  NAND2_X2 U8872 ( .A1(REGFILE_reg_out_24__4_), .A2(net77302), .ZN(n8059) );
  NAND4_X2 U8873 ( .A1(n8062), .A2(n8061), .A3(n8060), .A4(n8059), .ZN(n8063)
         );
  NAND2_X2 U8874 ( .A1(REGFILE_reg_out_22__4_), .A2(net77554), .ZN(n8068) );
  NAND2_X2 U8875 ( .A1(REGFILE_reg_out_17__4_), .A2(net77518), .ZN(n8067) );
  NAND2_X2 U8876 ( .A1(REGFILE_reg_out_23__4_), .A2(net77482), .ZN(n8066) );
  NAND2_X2 U8877 ( .A1(REGFILE_reg_out_21__4_), .A2(net77456), .ZN(n8065) );
  NAND4_X2 U8878 ( .A1(n8068), .A2(n8067), .A3(n8066), .A4(n8065), .ZN(n8074)
         );
  NAND2_X2 U8879 ( .A1(REGFILE_reg_out_19__4_), .A2(net77410), .ZN(n8072) );
  NAND2_X2 U8880 ( .A1(REGFILE_reg_out_20__4_), .A2(net77376), .ZN(n8071) );
  NAND2_X2 U8881 ( .A1(REGFILE_reg_out_18__4_), .A2(net77338), .ZN(n8070) );
  NAND2_X2 U8882 ( .A1(REGFILE_reg_out_16__4_), .A2(net77302), .ZN(n8069) );
  NAND4_X2 U8883 ( .A1(n8072), .A2(n8071), .A3(n8070), .A4(n8069), .ZN(n8073)
         );
  NAND2_X2 U8884 ( .A1(REGFILE_reg_out_14__4_), .A2(net77554), .ZN(n8078) );
  NAND2_X2 U8885 ( .A1(REGFILE_reg_out_9__4_), .A2(net77518), .ZN(n8077) );
  NAND2_X2 U8886 ( .A1(REGFILE_reg_out_15__4_), .A2(net77482), .ZN(n8076) );
  NAND2_X2 U8887 ( .A1(REGFILE_reg_out_13__4_), .A2(net77456), .ZN(n8075) );
  NAND4_X2 U8888 ( .A1(n8078), .A2(n8077), .A3(n8076), .A4(n8075), .ZN(n8084)
         );
  NAND2_X2 U8889 ( .A1(REGFILE_reg_out_11__4_), .A2(net77410), .ZN(n8082) );
  NAND2_X2 U8890 ( .A1(REGFILE_reg_out_12__4_), .A2(net77376), .ZN(n8081) );
  NAND2_X2 U8891 ( .A1(REGFILE_reg_out_10__4_), .A2(net77338), .ZN(n8080) );
  NAND2_X2 U8892 ( .A1(REGFILE_reg_out_8__4_), .A2(net77302), .ZN(n8079) );
  NAND4_X2 U8893 ( .A1(n8082), .A2(n8081), .A3(n8080), .A4(n8079), .ZN(n8083)
         );
  NAND2_X2 U8894 ( .A1(REGFILE_reg_out_6__4_), .A2(net77554), .ZN(n8088) );
  NAND2_X2 U8895 ( .A1(REGFILE_reg_out_7__4_), .A2(net77482), .ZN(n8086) );
  NAND2_X2 U8896 ( .A1(REGFILE_reg_out_5__4_), .A2(net77456), .ZN(n8085) );
  NAND4_X2 U8897 ( .A1(n8088), .A2(n8087), .A3(n8086), .A4(n8085), .ZN(n8094)
         );
  NAND2_X2 U8898 ( .A1(n5982), .A2(net77410), .ZN(n8092) );
  NAND2_X2 U8899 ( .A1(REGFILE_reg_out_4__4_), .A2(net77376), .ZN(n8091) );
  NAND2_X2 U8900 ( .A1(REGFILE_reg_out_2__4_), .A2(net77338), .ZN(n8090) );
  NAND2_X2 U8901 ( .A1(REGFILE_reg_out_0__4_), .A2(net77302), .ZN(n8089) );
  NAND4_X2 U8902 ( .A1(n8092), .A2(n8091), .A3(n8090), .A4(n8089), .ZN(n8093)
         );
  NAND4_X2 U8903 ( .A1(n8098), .A2(n8097), .A3(n8096), .A4(n8095), .ZN(n8425)
         );
  NAND2_X2 U8904 ( .A1(n8425), .A2(n4866), .ZN(n9954) );
  INV_X4 U8905 ( .A(n9954), .ZN(WIRE_ALU_A_MUX2TO1_32BIT_4__MUX_N1) );
  NAND2_X2 U8906 ( .A1(REGFILE_reg_out_30__3_), .A2(net77554), .ZN(n8102) );
  NAND2_X2 U8907 ( .A1(n5957), .A2(net77518), .ZN(n8101) );
  NAND2_X2 U8908 ( .A1(REGFILE_reg_out_31__3_), .A2(net77482), .ZN(n8100) );
  NAND2_X2 U8909 ( .A1(REGFILE_reg_out_29__3_), .A2(net77460), .ZN(n8099) );
  NAND4_X2 U8910 ( .A1(n8102), .A2(n8101), .A3(n8100), .A4(n8099), .ZN(n8108)
         );
  NAND2_X2 U8911 ( .A1(REGFILE_reg_out_27__3_), .A2(net77410), .ZN(n8106) );
  NAND2_X2 U8912 ( .A1(REGFILE_reg_out_28__3_), .A2(net77376), .ZN(n8105) );
  NAND2_X2 U8913 ( .A1(REGFILE_reg_out_26__3_), .A2(net77338), .ZN(n8104) );
  NAND2_X2 U8914 ( .A1(REGFILE_reg_out_24__3_), .A2(net77302), .ZN(n8103) );
  NAND4_X2 U8915 ( .A1(n8106), .A2(n8105), .A3(n8104), .A4(n8103), .ZN(n8107)
         );
  NAND2_X2 U8916 ( .A1(REGFILE_reg_out_22__3_), .A2(net77554), .ZN(n8112) );
  NAND2_X2 U8917 ( .A1(REGFILE_reg_out_17__3_), .A2(net77518), .ZN(n8111) );
  NAND2_X2 U8918 ( .A1(REGFILE_reg_out_23__3_), .A2(net77482), .ZN(n8110) );
  NAND2_X2 U8919 ( .A1(REGFILE_reg_out_21__3_), .A2(net77456), .ZN(n8109) );
  NAND4_X2 U8920 ( .A1(n8112), .A2(n8111), .A3(n8110), .A4(n8109), .ZN(n8118)
         );
  NAND2_X2 U8921 ( .A1(REGFILE_reg_out_19__3_), .A2(net77410), .ZN(n8116) );
  NAND2_X2 U8922 ( .A1(REGFILE_reg_out_20__3_), .A2(net77376), .ZN(n8115) );
  NAND2_X2 U8923 ( .A1(REGFILE_reg_out_18__3_), .A2(net77338), .ZN(n8114) );
  NAND2_X2 U8924 ( .A1(REGFILE_reg_out_16__3_), .A2(net77302), .ZN(n8113) );
  NAND4_X2 U8925 ( .A1(n8116), .A2(n8115), .A3(n8114), .A4(n8113), .ZN(n8117)
         );
  NAND2_X2 U8926 ( .A1(REGFILE_reg_out_14__3_), .A2(net77554), .ZN(n8122) );
  NAND2_X2 U8927 ( .A1(REGFILE_reg_out_9__3_), .A2(net77518), .ZN(n8121) );
  NAND2_X2 U8928 ( .A1(REGFILE_reg_out_15__3_), .A2(net77482), .ZN(n8120) );
  NAND2_X2 U8929 ( .A1(REGFILE_reg_out_13__3_), .A2(net77456), .ZN(n8119) );
  NAND4_X2 U8930 ( .A1(n8122), .A2(n8121), .A3(n8120), .A4(n8119), .ZN(n8128)
         );
  NAND2_X2 U8931 ( .A1(REGFILE_reg_out_11__3_), .A2(net77410), .ZN(n8126) );
  NAND2_X2 U8932 ( .A1(REGFILE_reg_out_12__3_), .A2(net77376), .ZN(n8125) );
  NAND2_X2 U8933 ( .A1(REGFILE_reg_out_10__3_), .A2(net77338), .ZN(n8124) );
  NAND2_X2 U8934 ( .A1(REGFILE_reg_out_8__3_), .A2(net77302), .ZN(n8123) );
  NAND4_X2 U8935 ( .A1(n8126), .A2(n8125), .A3(n8124), .A4(n8123), .ZN(n8127)
         );
  NAND2_X2 U8936 ( .A1(REGFILE_reg_out_6__3_), .A2(net77554), .ZN(n8132) );
  NAND2_X2 U8937 ( .A1(REGFILE_reg_out_1__3_), .A2(net77518), .ZN(n8131) );
  NAND2_X2 U8938 ( .A1(REGFILE_reg_out_7__3_), .A2(net77482), .ZN(n8130) );
  NAND2_X2 U8939 ( .A1(REGFILE_reg_out_5__3_), .A2(net77456), .ZN(n8129) );
  NAND4_X2 U8940 ( .A1(n8132), .A2(n8131), .A3(n8130), .A4(n8129), .ZN(n8138)
         );
  NAND2_X2 U8941 ( .A1(REGFILE_reg_out_4__3_), .A2(net77376), .ZN(n8135) );
  NAND2_X2 U8942 ( .A1(REGFILE_reg_out_0__3_), .A2(net77302), .ZN(n8133) );
  NAND4_X2 U8943 ( .A1(n8136), .A2(n8135), .A3(n8134), .A4(n8133), .ZN(n8137)
         );
  NAND4_X2 U8944 ( .A1(n8142), .A2(n8141), .A3(n8140), .A4(n8139), .ZN(n8423)
         );
  NAND2_X2 U8945 ( .A1(n8423), .A2(n4866), .ZN(n10404) );
  INV_X4 U8946 ( .A(n10404), .ZN(WIRE_ALU_A_MUX2TO1_32BIT_3__MUX_N1) );
  NAND2_X2 U8947 ( .A1(REGFILE_reg_out_30__2_), .A2(net77554), .ZN(n8146) );
  NAND2_X2 U8948 ( .A1(REGFILE_reg_out_25__2_), .A2(net77518), .ZN(n8145) );
  NAND2_X2 U8949 ( .A1(REGFILE_reg_out_31__2_), .A2(net77482), .ZN(n8144) );
  NAND2_X2 U8950 ( .A1(REGFILE_reg_out_29__2_), .A2(net77456), .ZN(n8143) );
  NAND4_X2 U8951 ( .A1(n8146), .A2(n8145), .A3(n8144), .A4(n8143), .ZN(n8152)
         );
  NAND2_X2 U8952 ( .A1(REGFILE_reg_out_27__2_), .A2(net77410), .ZN(n8150) );
  NAND2_X2 U8953 ( .A1(REGFILE_reg_out_28__2_), .A2(net77376), .ZN(n8149) );
  NAND2_X2 U8954 ( .A1(REGFILE_reg_out_26__2_), .A2(net77338), .ZN(n8148) );
  NAND2_X2 U8955 ( .A1(REGFILE_reg_out_24__2_), .A2(net77302), .ZN(n8147) );
  NAND4_X2 U8956 ( .A1(n8150), .A2(n8149), .A3(n8148), .A4(n8147), .ZN(n8151)
         );
  NAND2_X2 U8957 ( .A1(REGFILE_reg_out_22__2_), .A2(net77554), .ZN(n8156) );
  NAND2_X2 U8958 ( .A1(REGFILE_reg_out_17__2_), .A2(net77518), .ZN(n8155) );
  NAND2_X2 U8959 ( .A1(REGFILE_reg_out_23__2_), .A2(net77482), .ZN(n8154) );
  NAND2_X2 U8960 ( .A1(REGFILE_reg_out_21__2_), .A2(net77456), .ZN(n8153) );
  NAND4_X2 U8961 ( .A1(n8156), .A2(n8155), .A3(n8154), .A4(n8153), .ZN(n8162)
         );
  NAND2_X2 U8962 ( .A1(REGFILE_reg_out_19__2_), .A2(net77410), .ZN(n8160) );
  NAND2_X2 U8963 ( .A1(REGFILE_reg_out_20__2_), .A2(net77376), .ZN(n8159) );
  NAND2_X2 U8964 ( .A1(REGFILE_reg_out_18__2_), .A2(net77338), .ZN(n8158) );
  NAND2_X2 U8965 ( .A1(REGFILE_reg_out_16__2_), .A2(net77302), .ZN(n8157) );
  NAND4_X2 U8966 ( .A1(n8160), .A2(n8159), .A3(n8158), .A4(n8157), .ZN(n8161)
         );
  NAND2_X2 U8967 ( .A1(REGFILE_reg_out_14__2_), .A2(net77554), .ZN(n8166) );
  NAND2_X2 U8968 ( .A1(REGFILE_reg_out_9__2_), .A2(net77518), .ZN(n8165) );
  NAND2_X2 U8969 ( .A1(REGFILE_reg_out_15__2_), .A2(net77482), .ZN(n8164) );
  NAND2_X2 U8970 ( .A1(REGFILE_reg_out_13__2_), .A2(net77456), .ZN(n8163) );
  NAND4_X2 U8971 ( .A1(n8166), .A2(n8165), .A3(n8164), .A4(n8163), .ZN(n8172)
         );
  NAND2_X2 U8972 ( .A1(REGFILE_reg_out_11__2_), .A2(net77410), .ZN(n8170) );
  NAND2_X2 U8973 ( .A1(REGFILE_reg_out_12__2_), .A2(net77376), .ZN(n8169) );
  NAND2_X2 U8974 ( .A1(REGFILE_reg_out_10__2_), .A2(net77338), .ZN(n8168) );
  NAND2_X2 U8975 ( .A1(REGFILE_reg_out_8__2_), .A2(net77302), .ZN(n8167) );
  NAND4_X2 U8976 ( .A1(n8170), .A2(n8169), .A3(n8168), .A4(n8167), .ZN(n8171)
         );
  NAND2_X2 U8977 ( .A1(REGFILE_reg_out_6__2_), .A2(net77554), .ZN(n8176) );
  NAND2_X2 U8978 ( .A1(REGFILE_reg_out_1__2_), .A2(net77518), .ZN(n8175) );
  NAND2_X2 U8979 ( .A1(REGFILE_reg_out_7__2_), .A2(net77482), .ZN(n8174) );
  NAND2_X2 U8980 ( .A1(REGFILE_reg_out_5__2_), .A2(net77456), .ZN(n8173) );
  NAND4_X2 U8981 ( .A1(n8176), .A2(n8175), .A3(n8174), .A4(n8173), .ZN(n8182)
         );
  NAND2_X2 U8982 ( .A1(REGFILE_reg_out_3__2_), .A2(net77410), .ZN(n8180) );
  NAND2_X2 U8983 ( .A1(REGFILE_reg_out_4__2_), .A2(net77376), .ZN(n8179) );
  NAND2_X2 U8984 ( .A1(REGFILE_reg_out_2__2_), .A2(net77338), .ZN(n8178) );
  NAND2_X2 U8985 ( .A1(REGFILE_reg_out_0__2_), .A2(net77302), .ZN(n8177) );
  NAND4_X2 U8986 ( .A1(n8180), .A2(n8179), .A3(n8178), .A4(n8177), .ZN(n8181)
         );
  NAND4_X2 U8987 ( .A1(n8186), .A2(n8185), .A3(n8184), .A4(n8183), .ZN(n8421)
         );
  NAND2_X2 U8988 ( .A1(n8421), .A2(n4866), .ZN(n10109) );
  INV_X4 U8989 ( .A(n10109), .ZN(WIRE_ALU_A_MUX2TO1_32BIT_2__MUX_N1) );
  NAND2_X2 U8990 ( .A1(REGFILE_reg_out_25__1_), .A2(net77516), .ZN(n8189) );
  NAND2_X2 U8991 ( .A1(REGFILE_reg_out_31__1_), .A2(net77480), .ZN(n8188) );
  NAND4_X2 U8992 ( .A1(n8190), .A2(n8189), .A3(n8188), .A4(n8187), .ZN(n8196)
         );
  NAND2_X2 U8993 ( .A1(REGFILE_reg_out_27__1_), .A2(net77410), .ZN(n8194) );
  NAND2_X2 U8994 ( .A1(REGFILE_reg_out_28__1_), .A2(net77376), .ZN(n8193) );
  NAND2_X2 U8995 ( .A1(REGFILE_reg_out_26__1_), .A2(net77336), .ZN(n8192) );
  NAND4_X2 U8997 ( .A1(n8194), .A2(n8193), .A3(n8192), .A4(n8191), .ZN(n8195)
         );
  NAND2_X2 U8998 ( .A1(REGFILE_reg_out_17__1_), .A2(net77516), .ZN(n8199) );
  NAND2_X2 U8999 ( .A1(REGFILE_reg_out_23__1_), .A2(net77480), .ZN(n8198) );
  NAND4_X2 U9000 ( .A1(n8200), .A2(n8199), .A3(n8198), .A4(n8197), .ZN(n8206)
         );
  NAND2_X2 U9001 ( .A1(REGFILE_reg_out_19__1_), .A2(net77410), .ZN(n8204) );
  NAND2_X2 U9002 ( .A1(REGFILE_reg_out_18__1_), .A2(net77336), .ZN(n8202) );
  NAND4_X2 U9004 ( .A1(n8204), .A2(n8203), .A3(n8202), .A4(n8201), .ZN(n8205)
         );
  NAND2_X2 U9005 ( .A1(REGFILE_reg_out_9__1_), .A2(net77516), .ZN(n8209) );
  NAND2_X2 U9006 ( .A1(REGFILE_reg_out_15__1_), .A2(net77480), .ZN(n8208) );
  NAND4_X2 U9007 ( .A1(n8210), .A2(n8209), .A3(n8208), .A4(n8207), .ZN(n8216)
         );
  NAND2_X2 U9008 ( .A1(REGFILE_reg_out_11__1_), .A2(net77410), .ZN(n8214) );
  NAND2_X2 U9009 ( .A1(REGFILE_reg_out_12__1_), .A2(net77376), .ZN(n8213) );
  NAND2_X2 U9010 ( .A1(REGFILE_reg_out_10__1_), .A2(net77336), .ZN(n8212) );
  NAND4_X2 U9012 ( .A1(n8214), .A2(n8213), .A3(n8212), .A4(n8211), .ZN(n8215)
         );
  NAND2_X2 U9013 ( .A1(REGFILE_reg_out_1__1_), .A2(net77516), .ZN(n8219) );
  NAND2_X2 U9014 ( .A1(REGFILE_reg_out_7__1_), .A2(net77480), .ZN(n8218) );
  NAND4_X2 U9015 ( .A1(n8220), .A2(n8219), .A3(n8218), .A4(n8217), .ZN(n8226)
         );
  NAND2_X2 U9016 ( .A1(REGFILE_reg_out_3__1_), .A2(net77410), .ZN(n8224) );
  NAND2_X2 U9017 ( .A1(REGFILE_reg_out_4__1_), .A2(net77376), .ZN(n8223) );
  NAND2_X2 U9018 ( .A1(REGFILE_reg_out_2__1_), .A2(net77336), .ZN(n8222) );
  NAND4_X2 U9020 ( .A1(n8224), .A2(n8223), .A3(n8222), .A4(n8221), .ZN(n8225)
         );
  NAND4_X2 U9021 ( .A1(n8230), .A2(n8229), .A3(n8228), .A4(n8227), .ZN(n8422)
         );
  NAND2_X2 U9022 ( .A1(n8422), .A2(n4866), .ZN(net71273) );
  NAND2_X2 U9023 ( .A1(REGFILE_reg_out_25__0_), .A2(net77516), .ZN(n8233) );
  NAND2_X2 U9024 ( .A1(REGFILE_reg_out_31__0_), .A2(net77480), .ZN(n8232) );
  NAND4_X2 U9025 ( .A1(n8234), .A2(n8233), .A3(n8232), .A4(n8231), .ZN(n8240)
         );
  NAND2_X2 U9026 ( .A1(REGFILE_reg_out_27__0_), .A2(net77410), .ZN(n8238) );
  NAND2_X2 U9028 ( .A1(REGFILE_reg_out_26__0_), .A2(net77336), .ZN(n8236) );
  NAND2_X2 U9029 ( .A1(REGFILE_reg_out_24__0_), .A2(net77300), .ZN(n8235) );
  NAND4_X2 U9030 ( .A1(n8238), .A2(n8237), .A3(n8236), .A4(n8235), .ZN(n8239)
         );
  NAND2_X2 U9031 ( .A1(REGFILE_reg_out_17__0_), .A2(net77516), .ZN(n8243) );
  NAND2_X2 U9032 ( .A1(REGFILE_reg_out_23__0_), .A2(net77480), .ZN(n8242) );
  NAND4_X2 U9033 ( .A1(n8244), .A2(n8243), .A3(n8242), .A4(n8241), .ZN(n8250)
         );
  NAND2_X2 U9034 ( .A1(REGFILE_reg_out_19__0_), .A2(net77410), .ZN(n8248) );
  NAND2_X2 U9035 ( .A1(REGFILE_reg_out_18__0_), .A2(net77336), .ZN(n8246) );
  NAND2_X2 U9036 ( .A1(REGFILE_reg_out_16__0_), .A2(net77300), .ZN(n8245) );
  NAND4_X2 U9037 ( .A1(n8248), .A2(n8247), .A3(n8246), .A4(n8245), .ZN(n8249)
         );
  NAND2_X2 U9038 ( .A1(REGFILE_reg_out_9__0_), .A2(net77516), .ZN(n8253) );
  NAND2_X2 U9039 ( .A1(REGFILE_reg_out_15__0_), .A2(net77480), .ZN(n8252) );
  NAND4_X2 U9040 ( .A1(n8254), .A2(n8253), .A3(n8252), .A4(n8251), .ZN(n8260)
         );
  NAND2_X2 U9041 ( .A1(REGFILE_reg_out_11__0_), .A2(net77410), .ZN(n8258) );
  NAND2_X2 U9042 ( .A1(REGFILE_reg_out_12__0_), .A2(net77376), .ZN(n8257) );
  NAND2_X2 U9043 ( .A1(REGFILE_reg_out_10__0_), .A2(net77336), .ZN(n8256) );
  NAND4_X2 U9045 ( .A1(n8258), .A2(n8257), .A3(n8256), .A4(n8255), .ZN(n8259)
         );
  NAND2_X2 U9046 ( .A1(REGFILE_reg_out_6__0_), .A2(net77562), .ZN(n8264) );
  NAND2_X2 U9047 ( .A1(REGFILE_reg_out_1__0_), .A2(net77526), .ZN(n8263) );
  NAND2_X2 U9048 ( .A1(REGFILE_reg_out_7__0_), .A2(net77490), .ZN(n8262) );
  NAND2_X2 U9049 ( .A1(REGFILE_reg_out_5__0_), .A2(net77454), .ZN(n8261) );
  NAND4_X2 U9050 ( .A1(n8264), .A2(n8263), .A3(n8262), .A4(n8261), .ZN(n8270)
         );
  NAND2_X2 U9051 ( .A1(REGFILE_reg_out_3__0_), .A2(net77418), .ZN(n8268) );
  NAND2_X2 U9052 ( .A1(REGFILE_reg_out_4__0_), .A2(net77382), .ZN(n8267) );
  NAND2_X2 U9053 ( .A1(REGFILE_reg_out_2__0_), .A2(net77346), .ZN(n8266) );
  NAND2_X2 U9054 ( .A1(REGFILE_reg_out_0__0_), .A2(net77310), .ZN(n8265) );
  NAND4_X2 U9055 ( .A1(n8268), .A2(n8267), .A3(n8266), .A4(n8265), .ZN(n8269)
         );
  NAND4_X2 U9056 ( .A1(n8274), .A2(n8273), .A3(n8272), .A4(n8271), .ZN(n8416)
         );
  NAND2_X2 U9057 ( .A1(n8416), .A2(n4866), .ZN(net70535) );
  NAND2_X2 U9058 ( .A1(instructionAddr_out[28]), .A2(instructionAddr_out[29]), 
        .ZN(n8337) );
  NOR2_X4 U9059 ( .A1(n8337), .A2(n4969), .ZN(n8344) );
  NAND2_X2 U9060 ( .A1(instructionAddr_out[26]), .A2(n8344), .ZN(n8343) );
  INV_X4 U9061 ( .A(n8343), .ZN(n8275) );
  NAND2_X2 U9062 ( .A1(instructionAddr_out[25]), .A2(n8275), .ZN(n8326) );
  NAND2_X2 U9063 ( .A1(instructionAddr_out[24]), .A2(n8328), .ZN(n8327) );
  INV_X4 U9064 ( .A(n8327), .ZN(n8276) );
  NAND2_X2 U9065 ( .A1(instructionAddr_out[23]), .A2(n8276), .ZN(n8321) );
  NAND2_X2 U9066 ( .A1(instructionAddr_out[22]), .A2(n8323), .ZN(n8322) );
  INV_X4 U9067 ( .A(n8322), .ZN(n8277) );
  NAND2_X2 U9068 ( .A1(instructionAddr_out[21]), .A2(n8277), .ZN(n8316) );
  NAND2_X2 U9069 ( .A1(instructionAddr_out[20]), .A2(n8318), .ZN(n8317) );
  INV_X4 U9070 ( .A(n8317), .ZN(n8278) );
  NAND2_X2 U9071 ( .A1(instructionAddr_out[19]), .A2(n8278), .ZN(n8315) );
  INV_X4 U9072 ( .A(n8315), .ZN(n8279) );
  NAND2_X2 U9073 ( .A1(instructionAddr_out[18]), .A2(n8279), .ZN(n8314) );
  INV_X4 U9074 ( .A(n8314), .ZN(n8280) );
  NAND2_X2 U9075 ( .A1(instructionAddr_out[17]), .A2(n8280), .ZN(n8312) );
  INV_X4 U9076 ( .A(n8312), .ZN(n8281) );
  NAND2_X2 U9077 ( .A1(instructionAddr_out[16]), .A2(n8281), .ZN(n8364) );
  INV_X4 U9078 ( .A(n8364), .ZN(n8282) );
  NAND2_X2 U9079 ( .A1(instructionAddr_out[15]), .A2(n8282), .ZN(n8362) );
  INV_X4 U9080 ( .A(n8362), .ZN(n8310) );
  NAND3_X4 U9081 ( .A1(instructionAddr_out[13]), .A2(instructionAddr_out[14]), 
        .A3(n8310), .ZN(n8308) );
  INV_X4 U9082 ( .A(n8308), .ZN(n8283) );
  NAND3_X4 U9083 ( .A1(instructionAddr_out[11]), .A2(instructionAddr_out[12]), 
        .A3(n8283), .ZN(n8303) );
  INV_X4 U9084 ( .A(n8303), .ZN(n8302) );
  NAND3_X4 U9085 ( .A1(instructionAddr_out[10]), .A2(instructionAddr_out[9]), 
        .A3(n8302), .ZN(n8379) );
  INV_X4 U9086 ( .A(n8379), .ZN(n8284) );
  NAND3_X4 U9087 ( .A1(instructionAddr_out[7]), .A2(instructionAddr_out[8]), 
        .A3(n8284), .ZN(n8296) );
  INV_X4 U9088 ( .A(n8296), .ZN(n8389) );
  NAND3_X4 U9089 ( .A1(instructionAddr_out[6]), .A2(instructionAddr_out[5]), 
        .A3(n8389), .ZN(n8391) );
  INV_X4 U9090 ( .A(n8391), .ZN(n8285) );
  NAND2_X2 U9091 ( .A1(instructionAddr_out[4]), .A2(n8285), .ZN(n8293) );
  INV_X4 U9092 ( .A(n8293), .ZN(n8291) );
  NAND2_X2 U9093 ( .A1(instructionAddr_out[3]), .A2(n8291), .ZN(n8290) );
  INV_X4 U9094 ( .A(n8290), .ZN(n8286) );
  NAND2_X2 U9095 ( .A1(instructionAddr_out[2]), .A2(n8286), .ZN(n8289) );
  INV_X4 U9096 ( .A(n8289), .ZN(n10538) );
  XNOR2_X2 U9097 ( .A(instructionAddr_out[1]), .B(n10538), .ZN(net73771) );
  NAND2_X2 U9098 ( .A1(instruction[3]), .A2(net74011), .ZN(net73519) );
  INV_X4 U9099 ( .A(net73519), .ZN(net74009) );
  NAND2_X2 U9100 ( .A1(net73878), .A2(n8287), .ZN(n8288) );
  NAND2_X2 U9101 ( .A1(net74009), .A2(net73878), .ZN(net73877) );
  NAND2_X2 U9102 ( .A1(n8288), .A2(net73877), .ZN(net70531) );
  INV_X4 U9103 ( .A(net73778), .ZN(net73855) );
  AOI21_X4 U9104 ( .B1(n8290), .B2(n4923), .A(n10538), .ZN(net71396) );
  XNOR2_X2 U9105 ( .A(net73858), .B(net71396), .ZN(n8470) );
  XNOR2_X2 U9106 ( .A(instructionAddr_out[3]), .B(n8291), .ZN(n8292) );
  INV_X4 U9107 ( .A(n8292), .ZN(n10043) );
  NAND2_X2 U9108 ( .A1(n10043), .A2(net73858), .ZN(n8397) );
  AOI21_X4 U9109 ( .B1(n8391), .B2(n4924), .A(n8291), .ZN(n9965) );
  XNOR2_X2 U9110 ( .A(net73858), .B(n9965), .ZN(n8479) );
  XNOR2_X2 U9111 ( .A(instructionAddr_out[6]), .B(n8389), .ZN(n8294) );
  INV_X4 U9112 ( .A(n8294), .ZN(n9671) );
  NAND2_X2 U9113 ( .A1(net73858), .A2(n9671), .ZN(n8388) );
  NAND2_X2 U9114 ( .A1(n8297), .A2(n8296), .ZN(n8298) );
  INV_X4 U9115 ( .A(n8298), .ZN(n9700) );
  XNOR2_X2 U9116 ( .A(n8385), .B(n9700), .ZN(n8493) );
  AOI21_X4 U9117 ( .B1(n8302), .B2(instructionAddr_out[10]), .A(
        instructionAddr_out[9]), .ZN(n8299) );
  INV_X4 U9118 ( .A(n8299), .ZN(n8300) );
  NAND2_X2 U9119 ( .A1(n8300), .A2(n8379), .ZN(n8499) );
  NAND2_X2 U9120 ( .A1(net73988), .A2(net73877), .ZN(n8378) );
  XNOR2_X2 U9121 ( .A(n8499), .B(n8378), .ZN(n8497) );
  XNOR2_X2 U9122 ( .A(instructionAddr_out[10]), .B(n8302), .ZN(n8376) );
  NAND2_X2 U9123 ( .A1(n8304), .A2(n8303), .ZN(n8305) );
  INV_X4 U9124 ( .A(n8305), .ZN(n9864) );
  XNOR2_X2 U9125 ( .A(n8374), .B(n9864), .ZN(n8516) );
  XNOR2_X2 U9126 ( .A(n8308), .B(n4908), .ZN(n9107) );
  NAND2_X2 U9127 ( .A1(n8306), .A2(net73877), .ZN(n8372) );
  AOI21_X4 U9128 ( .B1(n8310), .B2(instructionAddr_out[14]), .A(
        instructionAddr_out[13]), .ZN(n8307) );
  INV_X4 U9129 ( .A(n8307), .ZN(n8309) );
  NAND2_X2 U9130 ( .A1(n8309), .A2(n8308), .ZN(n8368) );
  NAND2_X2 U9131 ( .A1(net73974), .A2(net73877), .ZN(n8367) );
  XNOR2_X2 U9132 ( .A(n8368), .B(n8367), .ZN(n9389) );
  XNOR2_X2 U9133 ( .A(instructionAddr_out[14]), .B(n8310), .ZN(n8311) );
  INV_X4 U9134 ( .A(n8311), .ZN(n10261) );
  XNOR2_X2 U9135 ( .A(net73900), .B(n10261), .ZN(n8502) );
  INV_X4 U9136 ( .A(instruction[16]), .ZN(net73908) );
  OAI21_X4 U9137 ( .B1(instructionAddr_out[16]), .B2(n8281), .A(n8364), .ZN(
        n8512) );
  XNOR2_X2 U9138 ( .A(n8314), .B(n5084), .ZN(n8313) );
  INV_X4 U9139 ( .A(n8313), .ZN(n9041) );
  INV_X4 U9140 ( .A(instruction[17]), .ZN(n8650) );
  XNOR2_X2 U9141 ( .A(n8313), .B(n8650), .ZN(n8796) );
  INV_X4 U9142 ( .A(n8796), .ZN(n8360) );
  OAI21_X4 U9143 ( .B1(instructionAddr_out[18]), .B2(n8279), .A(n8314), .ZN(
        n8804) );
  AOI21_X4 U9144 ( .B1(n8317), .B2(n5063), .A(n8279), .ZN(n10003) );
  INV_X4 U9145 ( .A(n8316), .ZN(n8318) );
  OAI21_X4 U9146 ( .B1(instructionAddr_out[20]), .B2(n8318), .A(n8317), .ZN(
        n9279) );
  XNOR2_X2 U9147 ( .A(n8322), .B(n5085), .ZN(n8320) );
  INV_X4 U9148 ( .A(n8320), .ZN(n9569) );
  XNOR2_X2 U9149 ( .A(n8320), .B(n8319), .ZN(n9536) );
  INV_X4 U9150 ( .A(n9536), .ZN(n8357) );
  INV_X4 U9151 ( .A(instruction[22]), .ZN(n8356) );
  INV_X4 U9152 ( .A(n8321), .ZN(n8323) );
  OAI21_X4 U9153 ( .B1(instructionAddr_out[22]), .B2(n8323), .A(n8322), .ZN(
        n8950) );
  XNOR2_X2 U9154 ( .A(n8327), .B(n5086), .ZN(n8325) );
  INV_X4 U9155 ( .A(n8325), .ZN(n9316) );
  XNOR2_X2 U9156 ( .A(n8325), .B(n8324), .ZN(n9283) );
  INV_X4 U9157 ( .A(n9283), .ZN(n8353) );
  INV_X4 U9158 ( .A(instruction[24]), .ZN(n8352) );
  INV_X4 U9159 ( .A(n8326), .ZN(n8328) );
  OAI21_X4 U9160 ( .B1(instructionAddr_out[24]), .B2(n8328), .A(n8327), .ZN(
        n8530) );
  XNOR2_X2 U9161 ( .A(n8343), .B(n5087), .ZN(n8330) );
  INV_X4 U9162 ( .A(n8330), .ZN(n9000) );
  XNOR2_X2 U9163 ( .A(n8330), .B(n8329), .ZN(n8968) );
  INV_X4 U9164 ( .A(n8968), .ZN(n8349) );
  INV_X4 U9165 ( .A(n8331), .ZN(n8788) );
  NAND2_X2 U9166 ( .A1(n8788), .A2(instruction[28]), .ZN(n8336) );
  INV_X4 U9167 ( .A(instruction[28]), .ZN(net73670) );
  XNOR2_X2 U9168 ( .A(n8331), .B(net73670), .ZN(n8690) );
  INV_X4 U9169 ( .A(n8690), .ZN(n8335) );
  NAND2_X2 U9170 ( .A1(instructionAddr_out[31]), .A2(instruction[31]), .ZN(
        n8699) );
  INV_X4 U9171 ( .A(n8699), .ZN(n8333) );
  XNOR2_X2 U9172 ( .A(instructionAddr_out[30]), .B(instruction[30]), .ZN(n8700) );
  INV_X4 U9173 ( .A(n8700), .ZN(n8332) );
  NAND2_X2 U9174 ( .A1(n8333), .A2(n8332), .ZN(n8702) );
  INV_X4 U9175 ( .A(n8702), .ZN(n8334) );
  AOI21_X4 U9176 ( .B1(instructionAddr_out[30]), .B2(instruction[30]), .A(
        n8334), .ZN(net73394) );
  XNOR2_X2 U9177 ( .A(instructionAddr_out[29]), .B(instruction[29]), .ZN(
        net73395) );
  INV_X4 U9178 ( .A(net73395), .ZN(net73938) );
  NAND2_X2 U9179 ( .A1(n8335), .A2(net73400), .ZN(n8691) );
  NAND2_X2 U9180 ( .A1(n8336), .A2(n8691), .ZN(n8686) );
  INV_X4 U9181 ( .A(n8686), .ZN(n8342) );
  INV_X4 U9182 ( .A(n8337), .ZN(n8339) );
  INV_X4 U9183 ( .A(n8344), .ZN(n8338) );
  OAI21_X4 U9184 ( .B1(instructionAddr_out[27]), .B2(n8339), .A(n8338), .ZN(
        n8340) );
  INV_X4 U9185 ( .A(n8340), .ZN(n8908) );
  XNOR2_X2 U9186 ( .A(instruction[27]), .B(n8908), .ZN(n8685) );
  NAND2_X2 U9187 ( .A1(n8908), .A2(instruction[27]), .ZN(n8341) );
  OAI21_X4 U9188 ( .B1(n8342), .B2(n8685), .A(n8341), .ZN(n8681) );
  INV_X4 U9189 ( .A(n8681), .ZN(n8348) );
  OAI21_X4 U9190 ( .B1(instructionAddr_out[26]), .B2(n8344), .A(n8343), .ZN(
        n8346) );
  INV_X4 U9191 ( .A(instruction[26]), .ZN(n8345) );
  XNOR2_X2 U9192 ( .A(n8346), .B(n8345), .ZN(n8680) );
  INV_X4 U9193 ( .A(n8346), .ZN(n9791) );
  NAND2_X2 U9194 ( .A1(n9791), .A2(instruction[26]), .ZN(n8347) );
  OAI21_X4 U9195 ( .B1(n8348), .B2(n8680), .A(n8347), .ZN(n8970) );
  NAND2_X2 U9196 ( .A1(n8349), .A2(n8970), .ZN(n8969) );
  INV_X4 U9197 ( .A(n8969), .ZN(n8350) );
  AOI21_X4 U9198 ( .B1(n9000), .B2(instruction[25]), .A(n8350), .ZN(n8528) );
  XNOR2_X2 U9199 ( .A(n8530), .B(n8351), .ZN(n8529) );
  OAI22_X2 U9200 ( .A1(n8352), .A2(n8530), .B1(n8528), .B2(n8529), .ZN(n9285)
         );
  NAND2_X2 U9201 ( .A1(n8353), .A2(n9285), .ZN(n9284) );
  INV_X4 U9202 ( .A(n9284), .ZN(n8354) );
  AOI21_X4 U9203 ( .B1(n9316), .B2(instruction[23]), .A(n8354), .ZN(n8963) );
  XNOR2_X2 U9204 ( .A(n8950), .B(n8355), .ZN(n8962) );
  OAI22_X2 U9205 ( .A1(n8356), .A2(n8950), .B1(n8963), .B2(n8962), .ZN(n9538)
         );
  NAND2_X2 U9206 ( .A1(n8357), .A2(n9538), .ZN(n9537) );
  INV_X4 U9207 ( .A(n9537), .ZN(n8358) );
  AOI21_X4 U9208 ( .B1(n9569), .B2(instruction[21]), .A(n8358), .ZN(n9278) );
  INV_X4 U9209 ( .A(instruction[20]), .ZN(net73512) );
  XNOR2_X2 U9210 ( .A(n9279), .B(net73512), .ZN(n9277) );
  OAI22_X2 U9211 ( .A1(net73512), .A2(n9279), .B1(n9278), .B2(n9277), .ZN(
        n9271) );
  NAND2_X2 U9212 ( .A1(n4968), .A2(n9271), .ZN(n9272) );
  INV_X4 U9213 ( .A(n9272), .ZN(n8359) );
  AOI21_X4 U9214 ( .B1(n10003), .B2(instruction[19]), .A(n8359), .ZN(n8803) );
  INV_X4 U9215 ( .A(instruction[18]), .ZN(net73529) );
  XNOR2_X2 U9216 ( .A(n8804), .B(net73529), .ZN(n8802) );
  OAI22_X2 U9217 ( .A1(net73529), .A2(n8804), .B1(n8803), .B2(n8802), .ZN(
        n8798) );
  NAND2_X2 U9218 ( .A1(n8360), .A2(n8798), .ZN(n8797) );
  INV_X4 U9219 ( .A(n8797), .ZN(n8361) );
  AOI21_X4 U9220 ( .B1(n9041), .B2(instruction[17]), .A(n8361), .ZN(n8511) );
  XNOR2_X2 U9221 ( .A(n8512), .B(net73908), .ZN(n8510) );
  OAI22_X2 U9222 ( .A1(net73908), .A2(n8512), .B1(n8511), .B2(n8510), .ZN(
        n8506) );
  INV_X4 U9223 ( .A(n8362), .ZN(n8363) );
  AOI21_X4 U9224 ( .B1(n8364), .B2(n5064), .A(n8363), .ZN(n10294) );
  XNOR2_X2 U9225 ( .A(net73902), .B(n10294), .ZN(n8507) );
  INV_X4 U9226 ( .A(n8507), .ZN(n8365) );
  AOI22_X2 U9227 ( .A1(n8506), .A2(n8365), .B1(net73902), .B2(n10294), .ZN(
        n8503) );
  NAND2_X2 U9228 ( .A1(net73900), .A2(n10261), .ZN(n8366) );
  INV_X4 U9229 ( .A(n9388), .ZN(n8371) );
  INV_X4 U9230 ( .A(n8367), .ZN(n8369) );
  INV_X4 U9231 ( .A(n8368), .ZN(n9422) );
  NAND2_X2 U9232 ( .A1(n8369), .A2(n9422), .ZN(n8370) );
  OAI21_X4 U9233 ( .B1(n9389), .B2(n8371), .A(n8370), .ZN(n8521) );
  XNOR2_X2 U9234 ( .A(n9107), .B(n8372), .ZN(n8520) );
  NAND2_X2 U9235 ( .A1(n8521), .A2(n8522), .ZN(n8523) );
  INV_X4 U9236 ( .A(n8373), .ZN(n8517) );
  NAND2_X2 U9237 ( .A1(n8374), .A2(n9864), .ZN(n8375) );
  OAI21_X4 U9238 ( .B1(n8516), .B2(n8517), .A(n8375), .ZN(n9384) );
  INV_X4 U9239 ( .A(n8376), .ZN(n10139) );
  XNOR2_X2 U9240 ( .A(n4921), .B(n10139), .ZN(n8377) );
  INV_X4 U9241 ( .A(n8377), .ZN(n9385) );
  AOI22_X2 U9242 ( .A1(n4921), .A2(n10139), .B1(n9384), .B2(n9385), .ZN(n8498)
         );
  OAI22_X2 U9243 ( .A1(n8499), .A2(n8378), .B1(n8497), .B2(n8498), .ZN(n9529)
         );
  XNOR2_X2 U9244 ( .A(n8379), .B(n4909), .ZN(n8382) );
  NAND2_X2 U9245 ( .A1(n8380), .A2(net73877), .ZN(n8381) );
  XNOR2_X2 U9246 ( .A(n8382), .B(n8381), .ZN(n9530) );
  INV_X4 U9247 ( .A(n9530), .ZN(n8384) );
  INV_X4 U9248 ( .A(n8381), .ZN(n8383) );
  INV_X4 U9249 ( .A(n8382), .ZN(n9531) );
  AOI22_X2 U9250 ( .A1(n9529), .A2(n8384), .B1(n8383), .B2(n9531), .ZN(n8494)
         );
  NAND2_X2 U9251 ( .A1(n8385), .A2(n9700), .ZN(n8386) );
  XNOR2_X2 U9252 ( .A(net73858), .B(n9671), .ZN(n8387) );
  INV_X4 U9253 ( .A(n8387), .ZN(n8488) );
  NAND2_X2 U9254 ( .A1(n8487), .A2(n8488), .ZN(n8489) );
  NAND2_X2 U9255 ( .A1(n8388), .A2(n8489), .ZN(n8483) );
  AOI21_X4 U9256 ( .B1(n8389), .B2(instructionAddr_out[6]), .A(
        instructionAddr_out[5]), .ZN(n8390) );
  INV_X4 U9257 ( .A(n8390), .ZN(n8392) );
  NAND2_X2 U9258 ( .A1(n8392), .A2(n8391), .ZN(n8393) );
  XNOR2_X2 U9259 ( .A(n8393), .B(net70531), .ZN(n8484) );
  INV_X4 U9260 ( .A(n8484), .ZN(n8394) );
  INV_X4 U9261 ( .A(n8393), .ZN(n9634) );
  AOI22_X2 U9262 ( .A1(n8483), .A2(n8394), .B1(n9634), .B2(net73858), .ZN(
        n8480) );
  NAND2_X2 U9263 ( .A1(n9965), .A2(net73858), .ZN(n8395) );
  XNOR2_X2 U9264 ( .A(net73858), .B(n10043), .ZN(n8396) );
  INV_X4 U9265 ( .A(n8396), .ZN(n8474) );
  NAND2_X2 U9266 ( .A1(n8473), .A2(n8474), .ZN(n8475) );
  NAND2_X2 U9267 ( .A1(n8397), .A2(n8475), .ZN(n8469) );
  INV_X4 U9268 ( .A(n8469), .ZN(n8399) );
  NAND2_X2 U9269 ( .A1(net71396), .A2(net73858), .ZN(n8398) );
  OAI21_X4 U9270 ( .B1(n8470), .B2(n8399), .A(n8398), .ZN(n8462) );
  INV_X4 U9271 ( .A(n10650), .ZN(n8464) );
  INV_X4 U9272 ( .A(net73842), .ZN(net73838) );
  INV_X4 U9273 ( .A(n8409), .ZN(n8411) );
  NAND4_X2 U9274 ( .A1(n8415), .A2(n8414), .A3(n8413), .A4(n8412), .ZN(n8459)
         );
  NAND4_X2 U9275 ( .A1(n8429), .A2(n8428), .A3(n8427), .A4(n8426), .ZN(n8458)
         );
  NAND4_X2 U9276 ( .A1(n8442), .A2(n8441), .A3(n8440), .A4(n8439), .ZN(n8457)
         );
  NOR4_X2 U9277 ( .A1(n8446), .A2(n8445), .A3(n8444), .A4(n8443), .ZN(n8455)
         );
  INV_X4 U9278 ( .A(n8447), .ZN(n8454) );
  NAND4_X2 U9279 ( .A1(n8455), .A2(n8454), .A3(n8453), .A4(n8452), .ZN(n8456)
         );
  NOR4_X2 U9280 ( .A1(n8459), .A2(n8458), .A3(n8457), .A4(n8456), .ZN(n8460)
         );
  XNOR2_X2 U9281 ( .A(n8460), .B(instruction[5]), .ZN(n8461) );
  NAND2_X2 U9282 ( .A1(n8462), .A2(net73855), .ZN(n10640) );
  NAND2_X2 U9283 ( .A1(n10649), .A2(n10640), .ZN(n8467) );
  INV_X4 U9284 ( .A(n8463), .ZN(n8465) );
  NAND2_X2 U9285 ( .A1(n8465), .A2(n8464), .ZN(n8527) );
  NAND2_X2 U9286 ( .A1(n6190), .A2(n5592), .ZN(n8466) );
  OAI221_X2 U9287 ( .B1(net71273), .B2(n4962), .C1(n8468), .C2(n8467), .A(
        n8466), .ZN(PCLOGIC_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  XOR2_X2 U9288 ( .A(n8470), .B(n8469), .Z(n8472) );
  NAND2_X2 U9289 ( .A1(n6190), .A2(net71396), .ZN(n8471) );
  OAI221_X2 U9290 ( .B1(n10109), .B2(n4962), .C1(n8472), .C2(n6008), .A(n8471), 
        .ZN(PCLOGIC_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9291 ( .A1(n10649), .A2(n8475), .ZN(n8477) );
  NAND2_X2 U9292 ( .A1(n6190), .A2(n10043), .ZN(n8476) );
  OAI221_X2 U9293 ( .B1(n10404), .B2(n4962), .C1(n8478), .C2(n8477), .A(n8476), 
        .ZN(PCLOGIC_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U9294 ( .A(n8480), .B(n8479), .ZN(n8482) );
  NAND2_X2 U9295 ( .A1(n6190), .A2(n9965), .ZN(n8481) );
  OAI221_X2 U9296 ( .B1(n9954), .B2(n4962), .C1(n6008), .C2(n8482), .A(n8481), 
        .ZN(PCLOGIC_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  XOR2_X2 U9297 ( .A(n8484), .B(n8483), .Z(n8486) );
  NAND2_X2 U9298 ( .A1(n6190), .A2(n9634), .ZN(n8485) );
  OAI221_X2 U9299 ( .B1(n10396), .B2(n4962), .C1(n8486), .C2(n9533), .A(n8485), 
        .ZN(PCLOGIC_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9300 ( .A1(n10649), .A2(n8489), .ZN(n8491) );
  NAND2_X2 U9301 ( .A1(n6190), .A2(n9671), .ZN(n8490) );
  OAI221_X2 U9302 ( .B1(n9656), .B2(n4962), .C1(n8492), .C2(n8491), .A(n8490), 
        .ZN(PCLOGIC_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U9303 ( .A(n8494), .B(n8493), .ZN(n8496) );
  NAND2_X2 U9304 ( .A1(n6190), .A2(n9700), .ZN(n8495) );
  OAI221_X2 U9305 ( .B1(n10464), .B2(n4962), .C1(n9533), .C2(n8496), .A(n8495), 
        .ZN(PCLOGIC_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U9306 ( .A(n8498), .B(n8497), .ZN(n8501) );
  INV_X4 U9307 ( .A(n8499), .ZN(n9375) );
  NAND2_X2 U9308 ( .A1(n6190), .A2(n9375), .ZN(n8500) );
  OAI221_X2 U9309 ( .B1(n10382), .B2(n4962), .C1(n6008), .C2(n8501), .A(n8500), 
        .ZN(PCLOGIC_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U9310 ( .A(n8503), .B(n8502), .ZN(n8505) );
  NAND2_X2 U9311 ( .A1(n6190), .A2(n10261), .ZN(n8504) );
  OAI221_X2 U9312 ( .B1(n10247), .B2(n4962), .C1(n9533), .C2(n8505), .A(n8504), 
        .ZN(PCLOGIC_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  XOR2_X2 U9313 ( .A(n8507), .B(n8506), .Z(n8509) );
  NAND2_X2 U9314 ( .A1(n6190), .A2(n10294), .ZN(n8508) );
  OAI221_X2 U9315 ( .B1(n10463), .B2(n4962), .C1(n8509), .C2(n6008), .A(n8508), 
        .ZN(PCLOGIC_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U9316 ( .A(n8511), .B(n8510), .ZN(n8515) );
  INV_X4 U9317 ( .A(n8512), .ZN(n9203) );
  NAND2_X2 U9318 ( .A1(n6190), .A2(n9203), .ZN(n8514) );
  NAND2_X2 U9319 ( .A1(net73708), .A2(aluA[16]), .ZN(n8513) );
  OAI211_X2 U9320 ( .C1(n8515), .C2(n9533), .A(n8514), .B(n8513), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U9321 ( .A(n8517), .B(n8516), .ZN(n8519) );
  NAND2_X2 U9322 ( .A1(n6190), .A2(n9864), .ZN(n8518) );
  OAI221_X2 U9323 ( .B1(n10375), .B2(n4962), .C1(n6008), .C2(n8519), .A(n8518), 
        .ZN(PCLOGIC_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9324 ( .A(n8520), .ZN(n8522) );
  NAND2_X2 U9325 ( .A1(n8523), .A2(n10649), .ZN(n8525) );
  INV_X4 U9326 ( .A(n4962), .ZN(net73708) );
  NAND2_X2 U9327 ( .A1(net73708), .A2(WIRE_ALU_A_MUX2TO1_32BIT_12__MUX_N1), 
        .ZN(n8524) );
  OAI221_X2 U9328 ( .B1(n9107), .B2(n8527), .C1(n8526), .C2(n8525), .A(n8524), 
        .ZN(PCLOGIC_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U9329 ( .A(n8529), .B(n8528), .ZN(n8533) );
  NAND2_X2 U9330 ( .A1(net73708), .A2(net36391), .ZN(n8532) );
  INV_X4 U9331 ( .A(n8530), .ZN(n8664) );
  NAND2_X2 U9332 ( .A1(n6190), .A2(n8664), .ZN(n8531) );
  OAI211_X2 U9333 ( .C1(n8533), .C2(n6008), .A(n8532), .B(n8531), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9335 ( .A(net73620), .ZN(net73684) );
  INV_X4 U9336 ( .A(net73695), .ZN(net73638) );
  NAND2_X2 U9337 ( .A1(net73638), .A2(net73619), .ZN(n8558) );
  INV_X4 U9338 ( .A(instruction[4]), .ZN(net73694) );
  NAND2_X2 U9339 ( .A1(n8576), .A2(net73694), .ZN(n8557) );
  INV_X4 U9340 ( .A(n8565), .ZN(n8576) );
  INV_X4 U9341 ( .A(instruction[31]), .ZN(net73652) );
  NAND3_X2 U9342 ( .A1(net73638), .A2(net73652), .A3(net73619), .ZN(n8534) );
  NAND2_X2 U9343 ( .A1(n8535), .A2(n8534), .ZN(n8582) );
  INV_X4 U9344 ( .A(n8582), .ZN(n8548) );
  NAND2_X2 U9345 ( .A1(instruction[4]), .A2(net73503), .ZN(n8655) );
  INV_X4 U9346 ( .A(n8655), .ZN(n8536) );
  NAND2_X2 U9347 ( .A1(n8536), .A2(instruction[3]), .ZN(n8538) );
  NAND2_X2 U9348 ( .A1(instruction[30]), .A2(net73652), .ZN(net73630) );
  NAND4_X2 U9349 ( .A1(net73646), .A2(instruction[29]), .A3(net73670), .A4(
        net73684), .ZN(n8537) );
  OAI21_X4 U9350 ( .B1(net73622), .B2(n8538), .A(n8537), .ZN(n8574) );
  INV_X4 U9351 ( .A(n8574), .ZN(n8547) );
  NAND3_X4 U9352 ( .A1(n8539), .A2(instruction[3]), .A3(net73498), .ZN(n8540)
         );
  INV_X4 U9353 ( .A(n8540), .ZN(n8564) );
  NAND3_X2 U9354 ( .A1(n4967), .A2(instruction[31]), .A3(net73670), .ZN(n8541)
         );
  NAND2_X2 U9355 ( .A1(n8542), .A2(n8541), .ZN(n8543) );
  INV_X4 U9356 ( .A(n8543), .ZN(n8579) );
  NOR2_X4 U9357 ( .A1(instruction[26]), .A2(instruction[27]), .ZN(n8544) );
  NAND4_X2 U9358 ( .A1(net73509), .A2(instruction[29]), .A3(net73670), .A4(
        n8544), .ZN(n8563) );
  INV_X4 U9359 ( .A(n8563), .ZN(n8545) );
  NAND2_X2 U9360 ( .A1(instruction[1]), .A2(instruction[3]), .ZN(n8559) );
  NAND4_X2 U9361 ( .A1(n8548), .A2(n8547), .A3(n8579), .A4(n8546), .ZN(n8549)
         );
  INV_X4 U9362 ( .A(n8549), .ZN(n8572) );
  NAND3_X2 U9363 ( .A1(n4967), .A2(net73670), .A3(net73652), .ZN(n8550) );
  NAND2_X2 U9364 ( .A1(n8551), .A2(n8550), .ZN(n8575) );
  NAND2_X2 U9365 ( .A1(n8552), .A2(net73619), .ZN(n8555) );
  NAND3_X2 U9366 ( .A1(n8555), .A2(n8554), .A3(net77272), .ZN(n8581) );
  NAND4_X2 U9367 ( .A1(n8558), .A2(n8557), .A3(n8572), .A4(n8556), .ZN(
        net73543) );
  INV_X4 U9368 ( .A(net73543), .ZN(net70821) );
  NAND2_X2 U9369 ( .A1(instruction[31]), .A2(instruction[30]), .ZN(n8562) );
  INV_X4 U9370 ( .A(n8559), .ZN(n8560) );
  NAND3_X2 U9371 ( .A1(n4966), .A2(instruction[5]), .A3(n8560), .ZN(n8561) );
  OAI21_X4 U9372 ( .B1(n8563), .B2(n8562), .A(n8561), .ZN(n8573) );
  INV_X4 U9373 ( .A(n8573), .ZN(n8571) );
  NAND2_X2 U9374 ( .A1(n4967), .A2(instruction[28]), .ZN(net73653) );
  INV_X4 U9375 ( .A(net73653), .ZN(net73616) );
  NAND2_X2 U9376 ( .A1(net73616), .A2(net73652), .ZN(n8570) );
  NAND2_X2 U9377 ( .A1(n8564), .A2(instruction[1]), .ZN(net73612) );
  INV_X4 U9378 ( .A(net73612), .ZN(net73637) );
  AOI21_X4 U9379 ( .B1(net73637), .B2(net73503), .A(n8566), .ZN(n8567) );
  INV_X4 U9380 ( .A(n8567), .ZN(n8568) );
  NOR3_X4 U9381 ( .A1(n8575), .A2(n8574), .A3(n8573), .ZN(net73611) );
  NAND4_X2 U9382 ( .A1(net73611), .A2(n8579), .A3(n8578), .A4(n8577), .ZN(
        net73541) );
  NOR2_X4 U9383 ( .A1(n8582), .A2(n8581), .ZN(net73613) );
  NOR2_X4 U9384 ( .A1(net73498), .A2(net73622), .ZN(net73615) );
  XNOR2_X2 U9385 ( .A(n10315), .B(net77042), .ZN(n8591) );
  INV_X4 U9386 ( .A(n8591), .ZN(n8593) );
  XNOR2_X2 U9387 ( .A(n10099), .B(net77042), .ZN(n8587) );
  INV_X4 U9388 ( .A(n9809), .ZN(n8590) );
  XNOR2_X2 U9389 ( .A(net71026), .B(net77042), .ZN(n8585) );
  XNOR2_X2 U9390 ( .A(n10928), .B(net77038), .ZN(n8584) );
  INV_X4 U9391 ( .A(n8583), .ZN(n10490) );
  OAI22_X2 U9392 ( .A1(net73608), .A2(n8584), .B1(net77042), .B2(n10490), .ZN(
        n8707) );
  INV_X4 U9393 ( .A(n8585), .ZN(n8586) );
  AOI22_X2 U9394 ( .A1(n8706), .A2(n8707), .B1(n8586), .B2(n5798), .ZN(n9810)
         );
  INV_X4 U9395 ( .A(n8587), .ZN(n8588) );
  OAI21_X4 U9396 ( .B1(n8590), .B2(n9810), .A(n8589), .ZN(n8772) );
  NAND2_X2 U9397 ( .A1(n8772), .A2(n8773), .ZN(n8771) );
  INV_X4 U9398 ( .A(n8771), .ZN(n8592) );
  XNOR2_X2 U9399 ( .A(n8594), .B(n5761), .ZN(n8883) );
  NAND2_X2 U9400 ( .A1(n8594), .A2(n5761), .ZN(n8595) );
  NAND2_X2 U9401 ( .A1(n9776), .A2(n9777), .ZN(n9774) );
  OAI21_X4 U9402 ( .B1(n8597), .B2(n8596), .A(n9774), .ZN(n8987) );
  INV_X4 U9403 ( .A(n8988), .ZN(n8598) );
  AOI22_X2 U9404 ( .A1(n8987), .A2(n8598), .B1(n10930), .B2(n4808), .ZN(n8809)
         );
  INV_X4 U9405 ( .A(n8808), .ZN(n8600) );
  XNOR2_X2 U9406 ( .A(n8809), .B(n8600), .ZN(n8603) );
  XNOR2_X2 U9407 ( .A(net36391), .B(n10331), .ZN(n10430) );
  NAND2_X2 U9408 ( .A1(n10494), .A2(net73541), .ZN(net70845) );
  NAND2_X2 U9409 ( .A1(multOut[24]), .A2(net81873), .ZN(n8648) );
  NAND2_X2 U9410 ( .A1(n10928), .A2(n10494), .ZN(n10474) );
  INV_X4 U9411 ( .A(n10474), .ZN(n8854) );
  INV_X4 U9412 ( .A(net73541), .ZN(net70826) );
  NAND2_X2 U9413 ( .A1(net77042), .A2(n10494), .ZN(n10304) );
  INV_X4 U9414 ( .A(n10494), .ZN(n10457) );
  NAND2_X2 U9415 ( .A1(n10457), .A2(net77040), .ZN(n8642) );
  NAND2_X2 U9416 ( .A1(n10304), .A2(n8642), .ZN(n10475) );
  NAND2_X2 U9417 ( .A1(net70826), .A2(n10475), .ZN(n8604) );
  MUX2_X2 U9418 ( .A(n8604), .B(net70845), .S(net70821), .Z(net72163) );
  NAND2_X2 U9419 ( .A1(n8854), .A2(net70697), .ZN(n9803) );
  NAND2_X2 U9420 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_5__MUX_N1), .A2(net70720), 
        .ZN(n8607) );
  INV_X4 U9421 ( .A(n9581), .ZN(n9330) );
  NAND2_X2 U9422 ( .A1(n10933), .A2(n6041), .ZN(n8821) );
  NAND2_X2 U9423 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_13__MUX_N1), .A2(n9065), .ZN(
        n9597) );
  INV_X4 U9424 ( .A(n9597), .ZN(n8605) );
  NAND2_X2 U9425 ( .A1(net70534), .A2(net73541), .ZN(net71300) );
  NAND2_X2 U9426 ( .A1(net70719), .A2(net70696), .ZN(n8855) );
  INV_X4 U9427 ( .A(n8855), .ZN(n8624) );
  NOR2_X4 U9428 ( .A1(n8605), .A2(n8624), .ZN(n8606) );
  NAND3_X4 U9429 ( .A1(n8607), .A2(n8821), .A3(n8606), .ZN(n8977) );
  NAND2_X2 U9430 ( .A1(n10102), .A2(n8977), .ZN(n8619) );
  NAND2_X2 U9431 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_7__MUX_N1), .A2(net70720), 
        .ZN(n8610) );
  NAND2_X2 U9432 ( .A1(n10931), .A2(n6041), .ZN(n8826) );
  NAND2_X2 U9433 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_15__MUX_N1), .A2(n9065), .ZN(
        n9593) );
  INV_X4 U9434 ( .A(n9593), .ZN(n8608) );
  NOR2_X4 U9435 ( .A1(n8608), .A2(n8624), .ZN(n8609) );
  NAND3_X4 U9436 ( .A1(n8610), .A2(n8826), .A3(n8609), .ZN(n8976) );
  NAND2_X2 U9437 ( .A1(net77086), .A2(n8976), .ZN(n8618) );
  NAND2_X2 U9438 ( .A1(n6040), .A2(aluA[19]), .ZN(n8828) );
  NAND2_X2 U9439 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_11__MUX_N1), .A2(n9065), .ZN(
        n10018) );
  INV_X4 U9440 ( .A(n10018), .ZN(n8612) );
  NOR2_X4 U9441 ( .A1(n8612), .A2(n8611), .ZN(n8613) );
  NAND3_X4 U9442 ( .A1(n8855), .A2(n8828), .A3(n8613), .ZN(n9976) );
  NAND2_X2 U9443 ( .A1(n6040), .A2(aluA[17]), .ZN(n9017) );
  NAND2_X2 U9444 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_9__MUX_N1), .A2(n9065), .ZN(
        n10155) );
  INV_X4 U9445 ( .A(n10155), .ZN(n8615) );
  NOR2_X4 U9446 ( .A1(n8615), .A2(n8614), .ZN(n8616) );
  NAND3_X4 U9447 ( .A1(n8855), .A2(n9017), .A3(n8616), .ZN(n9975) );
  AOI22_X2 U9448 ( .A1(n6082), .A2(n9976), .B1(n6083), .B2(n9975), .ZN(n8617)
         );
  NAND2_X2 U9449 ( .A1(n10058), .A2(n9294), .ZN(n8633) );
  INV_X4 U9450 ( .A(n10928), .ZN(n10470) );
  INV_X4 U9451 ( .A(n10472), .ZN(n8861) );
  INV_X4 U9452 ( .A(n9854), .ZN(n10060) );
  NAND2_X2 U9453 ( .A1(n6040), .A2(aluA[18]), .ZN(n8842) );
  NAND2_X2 U9454 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_10__MUX_N1), .A2(n9065), .ZN(
        n10095) );
  INV_X4 U9455 ( .A(n10095), .ZN(n8621) );
  NOR2_X4 U9456 ( .A1(n8621), .A2(n8620), .ZN(n8622) );
  NAND3_X4 U9457 ( .A1(n8855), .A2(n8842), .A3(n8622), .ZN(n9546) );
  NAND2_X2 U9458 ( .A1(n6083), .A2(n9546), .ZN(n8631) );
  NAND2_X2 U9459 ( .A1(n6040), .A2(aluA[20]), .ZN(n8836) );
  NAND2_X2 U9460 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_12__MUX_N1), .A2(n9065), .ZN(
        n9938) );
  NAND3_X4 U9461 ( .A1(n8836), .A2(n9938), .A3(n8625), .ZN(n9547) );
  NAND2_X2 U9462 ( .A1(n6082), .A2(n9547), .ZN(n8630) );
  NAND2_X2 U9463 ( .A1(n10932), .A2(n6041), .ZN(n8840) );
  NAND2_X2 U9464 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_14__MUX_N1), .A2(n9065), .ZN(
        n9617) );
  NAND2_X2 U9465 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_6__MUX_N1), .A2(net70720), 
        .ZN(n8626) );
  NAND4_X2 U9466 ( .A1(n8840), .A2(n9617), .A3(n8626), .A4(n8855), .ZN(n8928)
         );
  NAND2_X2 U9467 ( .A1(n8728), .A2(n8928), .ZN(n8629) );
  NAND2_X2 U9468 ( .A1(net36391), .A2(n6041), .ZN(n8637) );
  NAND2_X2 U9469 ( .A1(n9065), .A2(aluA[16]), .ZN(n9499) );
  AOI22_X2 U9470 ( .A1(net70719), .A2(net70534), .B1(net70720), .B2(
        WIRE_ALU_A_MUX2TO1_32BIT_8__MUX_N1), .ZN(n8627) );
  NAND2_X2 U9471 ( .A1(net77084), .A2(n8892), .ZN(n8628) );
  NAND4_X2 U9472 ( .A1(n8631), .A2(n8630), .A3(n8629), .A4(n8628), .ZN(n8975)
         );
  NAND2_X2 U9473 ( .A1(n10060), .A2(n8975), .ZN(n8632) );
  NAND2_X2 U9474 ( .A1(n8633), .A2(n8632), .ZN(n8646) );
  NAND2_X2 U9475 ( .A1(n10457), .A2(n10928), .ZN(n9770) );
  INV_X4 U9476 ( .A(n9770), .ZN(n10303) );
  NAND2_X2 U9477 ( .A1(n6040), .A2(n6005), .ZN(n8823) );
  INV_X4 U9478 ( .A(n5761), .ZN(n10319) );
  NAND2_X2 U9479 ( .A1(n6040), .A2(n10099), .ZN(n8634) );
  NAND2_X2 U9480 ( .A1(n10064), .A2(n8974), .ZN(n8636) );
  NAND2_X2 U9481 ( .A1(n10457), .A2(n10470), .ZN(n9802) );
  NAND2_X2 U9482 ( .A1(n10066), .A2(n9297), .ZN(n8635) );
  NAND2_X2 U9483 ( .A1(n8636), .A2(n8635), .ZN(n8641) );
  NAND2_X2 U9484 ( .A1(n10930), .A2(n6041), .ZN(n8724) );
  OAI22_X2 U9485 ( .A1(n10312), .A2(n8823), .B1(n6005), .B2(n8724), .ZN(n9298)
         );
  NAND2_X2 U9486 ( .A1(n10064), .A2(n9298), .ZN(n8640) );
  OAI22_X2 U9487 ( .A1(n8638), .A2(n8823), .B1(n6005), .B2(n8637), .ZN(n9301)
         );
  NAND2_X2 U9488 ( .A1(n10066), .A2(n9301), .ZN(n8639) );
  NAND2_X2 U9489 ( .A1(n8640), .A2(n8639), .ZN(n8942) );
  MUX2_X2 U9490 ( .A(n8641), .B(n8942), .S(net71026), .Z(n8645) );
  INV_X4 U9491 ( .A(n8642), .ZN(n10491) );
  NAND2_X2 U9492 ( .A1(n10491), .A2(net73543), .ZN(n8643) );
  NAND2_X2 U9493 ( .A1(n8643), .A2(n10304), .ZN(net70706) );
  NAND3_X2 U9494 ( .A1(n8649), .A2(n8648), .A3(n8647), .ZN(dmem_addr_out[24])
         );
  MUX2_X2 U9495 ( .A(net88253), .B(n8650), .S(net73509), .Z(n8651) );
  NAND2_X2 U9496 ( .A1(n8651), .A2(net70738), .ZN(net73443) );
  NAND2_X2 U9497 ( .A1(net73527), .A2(net70738), .ZN(net73429) );
  MUX2_X2 U9498 ( .A(n4820), .B(net73908), .S(net73509), .Z(n8652) );
  NAND2_X2 U9499 ( .A1(n8652), .A2(net70738), .ZN(net73468) );
  NAND2_X2 U9500 ( .A1(instruction[0]), .A2(instruction[2]), .ZN(n8653) );
  NAND2_X2 U9501 ( .A1(net73510), .A2(net70738), .ZN(n8671) );
  INV_X4 U9502 ( .A(n8671), .ZN(n8669) );
  INV_X4 U9503 ( .A(instruction[19]), .ZN(n8656) );
  MUX2_X2 U9504 ( .A(net86793), .B(n8656), .S(net73509), .Z(n8657) );
  NAND2_X2 U9505 ( .A1(n8657), .A2(net70738), .ZN(n8670) );
  INV_X4 U9506 ( .A(n8670), .ZN(n8672) );
  INV_X4 U9507 ( .A(dmem_addr_out[24]), .ZN(n8667) );
  INV_X4 U9508 ( .A(n8870), .ZN(dmem_dsize[1]) );
  INV_X4 U9509 ( .A(dmem_read_in[8]), .ZN(n9516) );
  NAND2_X2 U9510 ( .A1(n4899), .A2(n8870), .ZN(net70811) );
  INV_X4 U9511 ( .A(dmem_read_in[0]), .ZN(n10540) );
  INV_X4 U9512 ( .A(dmem_read_in[24]), .ZN(n8662) );
  OAI211_X2 U9513 ( .C1(n8667), .C2(net76646), .A(n8666), .B(n8665), .ZN(n8668) );
  OAI22_X2 U9514 ( .A1(n5128), .A2(n6088), .B1(net76660), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9515 ( .A1(n8669), .A2(n8670), .ZN(net73436) );
  INV_X4 U9516 ( .A(net73436), .ZN(net73423) );
  NAND2_X2 U9517 ( .A1(net76270), .A2(n6156), .ZN(n10512) );
  OAI22_X2 U9518 ( .A1(n5253), .A2(n6091), .B1(n6156), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9519 ( .A1(n8670), .A2(n8671), .ZN(net73434) );
  INV_X4 U9520 ( .A(net73434), .ZN(net73421) );
  OAI22_X2 U9521 ( .A1(n6192), .A2(n5563), .B1(n6195), .B2(n8679), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9522 ( .A1(n6196), .A2(n5564), .B1(n6199), .B2(n8679), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9523 ( .A1(n8672), .A2(n8671), .ZN(net73439) );
  NAND2_X2 U9524 ( .A1(n4894), .A2(net73416), .ZN(n10516) );
  NAND2_X2 U9525 ( .A1(net76270), .A2(n10516), .ZN(n10517) );
  OAI22_X2 U9526 ( .A1(n4946), .A2(n6097), .B1(n6095), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9527 ( .A1(n4894), .A2(net73423), .ZN(n10519) );
  OAI22_X2 U9528 ( .A1(n5129), .A2(n6103), .B1(n6102), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9529 ( .A1(n4894), .A2(net73421), .ZN(n10521) );
  OAI22_X2 U9530 ( .A1(n4947), .A2(n6108), .B1(n6106), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9531 ( .A1(n5130), .A2(n6112), .B1(n6158), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9532 ( .A1(n5131), .A2(n6115), .B1(n6160), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9533 ( .A1(n5254), .A2(n6118), .B1(n6162), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9534 ( .A1(n6200), .A2(n5363), .B1(n6204), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9535 ( .A1(n5255), .A2(net76862), .B1(net76616), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9536 ( .A1(n6205), .A2(n5398), .B1(n6208), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9537 ( .A1(n5132), .A2(n6121), .B1(n6164), .B2(n8679), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9538 ( .A1(n5256), .A2(n6124), .B1(n6166), .B2(n8679), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9539 ( .A1(n5133), .A2(n6127), .B1(n6168), .B2(n8679), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9540 ( .A1(n5134), .A2(n6129), .B1(n6170), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9541 ( .A1(n5257), .A2(n6132), .B1(n6172), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9542 ( .A1(n5135), .A2(n6136), .B1(n6174), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9543 ( .A1(n6209), .A2(n5399), .B1(n6212), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9544 ( .A(n8677), .ZN(n8673) );
  NAND2_X2 U9545 ( .A1(REGFILE_reg_out_28__24_), .A2(n6177), .ZN(n8674) );
  OAI21_X4 U9546 ( .B1(n6213), .B2(n6021), .A(n8674), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9547 ( .A(n10607), .ZN(n10532) );
  NAND2_X2 U9548 ( .A1(n6178), .A2(REGFILE_reg_out_29__24_), .ZN(n8675) );
  OAI21_X4 U9549 ( .B1(n6138), .B2(n6021), .A(n8675), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9550 ( .A1(n5258), .A2(n6139), .B1(net76550), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9551 ( .A(n10614), .ZN(n10534) );
  NAND2_X2 U9552 ( .A1(n6180), .A2(REGFILE_reg_out_30__24_), .ZN(n8676) );
  OAI21_X4 U9553 ( .B1(n6142), .B2(n6021), .A(n8676), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9554 ( .A(net70574), .ZN(net70509) );
  NAND2_X2 U9555 ( .A1(net76488), .A2(REGFILE_reg_out_31__24_), .ZN(n8678) );
  OAI21_X4 U9556 ( .B1(net76480), .B2(n6021), .A(n8678), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9557 ( .A1(n6215), .A2(n5400), .B1(net76320), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9558 ( .A1(n6217), .A2(n5364), .B1(n6220), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9559 ( .A1(n5259), .A2(n6144), .B1(n6183), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9560 ( .A1(net73423), .A2(n4895), .ZN(n10535) );
  OAI22_X2 U9561 ( .A1(n5260), .A2(net76706), .B1(n6147), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9562 ( .A1(n5136), .A2(net76692), .B1(n6185), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9563 ( .A1(n5261), .A2(n6150), .B1(n6187), .B2(n6021), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9564 ( .A1(n5137), .A2(n6153), .B1(n6189), .B2(n8679), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  XOR2_X2 U9565 ( .A(n8681), .B(n8680), .Z(n8684) );
  NAND2_X2 U9566 ( .A1(n6190), .A2(n9791), .ZN(n8682) );
  OAI211_X2 U9567 ( .C1(n8684), .C2(n9533), .A(n8683), .B(n8682), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  XOR2_X2 U9568 ( .A(n8686), .B(n8685), .Z(n8689) );
  NAND2_X2 U9569 ( .A1(net73708), .A2(n5761), .ZN(n8688) );
  NAND2_X2 U9570 ( .A1(n6190), .A2(n8908), .ZN(n8687) );
  OAI211_X2 U9571 ( .C1(n8689), .C2(n6008), .A(n8688), .B(n8687), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI211_X2 U9572 ( .C1(n8335), .C2(net73400), .A(n8691), .B(n10649), .ZN(
        n8693) );
  NAND2_X2 U9573 ( .A1(n6190), .A2(n8788), .ZN(n8692) );
  XOR2_X2 U9574 ( .A(net73394), .B(net73395), .Z(n8697) );
  NAND2_X2 U9575 ( .A1(n6190), .A2(n5016), .ZN(n8695) );
  OAI211_X2 U9576 ( .C1(n8697), .C2(n9533), .A(n8696), .B(n8695), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9578 ( .A1(n6190), .A2(instructionAddr_out[30]), .ZN(n8705) );
  NAND2_X2 U9579 ( .A1(n8700), .A2(n8699), .ZN(n8701) );
  XOR2_X2 U9580 ( .A(n8707), .B(n8706), .Z(n8719) );
  NAND2_X2 U9581 ( .A1(net77084), .A2(n6041), .ZN(n10159) );
  INV_X4 U9582 ( .A(n10159), .ZN(n10542) );
  NAND2_X2 U9583 ( .A1(n10542), .A2(n5798), .ZN(n9805) );
  NAND2_X2 U9584 ( .A1(n10932), .A2(n9065), .ZN(n9076) );
  OAI21_X4 U9585 ( .B1(n8709), .B2(n8708), .A(net77084), .ZN(n8717) );
  NAND2_X2 U9586 ( .A1(n9065), .A2(aluA[20]), .ZN(n9079) );
  AOI22_X2 U9587 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_4__MUX_N1), .A2(net70719), 
        .B1(WIRE_ALU_A_MUX2TO1_32BIT_12__MUX_N1), .B2(net70720), .ZN(n8710) );
  NAND3_X2 U9588 ( .A1(n9079), .A2(n8711), .A3(n8710), .ZN(n8712) );
  MUX2_X2 U9589 ( .A(n8892), .B(n8712), .S(n10099), .Z(n8758) );
  NAND2_X2 U9590 ( .A1(n8758), .A2(net78051), .ZN(n8716) );
  NAND2_X2 U9591 ( .A1(n9065), .A2(aluA[18]), .ZN(n9360) );
  AOI22_X2 U9592 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_2__MUX_N1), .A2(net70719), 
        .B1(WIRE_ALU_A_MUX2TO1_32BIT_10__MUX_N1), .B2(net70720), .ZN(n8713) );
  NAND3_X4 U9593 ( .A1(n9360), .A2(n8714), .A3(n8713), .ZN(n8891) );
  NAND2_X2 U9594 ( .A1(n6081), .A2(n8891), .ZN(n8715) );
  AOI21_X4 U9595 ( .B1(n4910), .B2(n8719), .A(n8718), .ZN(n8734) );
  XNOR2_X2 U9596 ( .A(n5798), .B(net78051), .ZN(n10433) );
  INV_X4 U9597 ( .A(n10433), .ZN(n10310) );
  NAND2_X2 U9598 ( .A1(net70701), .A2(n10310), .ZN(n8733) );
  INV_X4 U9599 ( .A(n10094), .ZN(n8728) );
  NAND2_X2 U9600 ( .A1(n6040), .A2(n5761), .ZN(n8722) );
  NAND2_X2 U9601 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_11__MUX_N1), .A2(net70720), 
        .ZN(n8721) );
  NAND2_X2 U9602 ( .A1(n9065), .A2(aluA[19]), .ZN(n9340) );
  NAND2_X2 U9603 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_3__MUX_N1), .A2(net70719), 
        .ZN(n8720) );
  NAND4_X2 U9604 ( .A1(n8722), .A2(n8721), .A3(n9340), .A4(n8720), .ZN(n10466)
         );
  NAND2_X2 U9605 ( .A1(n9065), .A2(aluA[17]), .ZN(n9343) );
  AOI22_X2 U9606 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_1__MUX_N1), .A2(net70719), 
        .B1(WIRE_ALU_A_MUX2TO1_32BIT_9__MUX_N1), .B2(net70720), .ZN(n8723) );
  NAND2_X2 U9607 ( .A1(n10933), .A2(n9065), .ZN(n9068) );
  AOI22_X2 U9608 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_5__MUX_N1), .A2(net70719), 
        .B1(WIRE_ALU_A_MUX2TO1_32BIT_13__MUX_N1), .B2(net70720), .ZN(n8725) );
  NAND3_X2 U9609 ( .A1(n9068), .A2(n8726), .A3(n8725), .ZN(n8727) );
  MUX2_X2 U9610 ( .A(n8978), .B(n8727), .S(n10099), .Z(n10465) );
  NAND2_X2 U9611 ( .A1(n8854), .A2(net70697), .ZN(n9012) );
  OAI22_X2 U9612 ( .A1(n9801), .A2(n9012), .B1(n9606), .B2(n9805), .ZN(n8731)
         );
  NOR3_X4 U9613 ( .A1(n8731), .A2(n8730), .A3(n5062), .ZN(n8732) );
  MUX2_X2 U9614 ( .A(n8735), .B(multOut[30]), .S(net76452), .Z(
        dmem_addr_out[30]) );
  INV_X4 U9615 ( .A(dmem_read_in[6]), .ZN(n9669) );
  INV_X4 U9616 ( .A(dmem_read_in[14]), .ZN(n10259) );
  OAI22_X2 U9617 ( .A1(net70811), .A2(n9669), .B1(net77999), .B2(n10259), .ZN(
        n8736) );
  AOI21_X4 U9618 ( .B1(net76650), .B2(dmem_addr_out[30]), .A(n8736), .ZN(n8741) );
  INV_X4 U9619 ( .A(dmem_read_in[30]), .ZN(n8737) );
  NAND2_X2 U9620 ( .A1(n8741), .A2(n8740), .ZN(n8742) );
  OAI22_X2 U9621 ( .A1(n4975), .A2(n6088), .B1(n6223), .B2(net76658), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9622 ( .A(REGFILE_reg_out_10__30_), .ZN(n8743) );
  OAI22_X2 U9623 ( .A1(n8743), .A2(n6091), .B1(n6223), .B2(n6155), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9624 ( .A1(n5958), .A2(n6097), .B1(n6223), .B2(n6094), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9625 ( .A(REGFILE_reg_out_14__30_), .ZN(n8744) );
  OAI22_X2 U9626 ( .A1(n8744), .A2(n6103), .B1(n6223), .B2(n6102), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9627 ( .A1(n5918), .A2(n6108), .B1(n6223), .B2(n6105), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9628 ( .A1(n8745), .A2(n6112), .B1(n6223), .B2(n6157), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9629 ( .A(REGFILE_reg_out_17__30_), .ZN(n8746) );
  OAI22_X2 U9630 ( .A1(n8746), .A2(n6115), .B1(n6223), .B2(n6159), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9631 ( .A(REGFILE_reg_out_18__30_), .ZN(n8747) );
  OAI22_X2 U9632 ( .A1(n8747), .A2(n6118), .B1(n6223), .B2(n6161), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9633 ( .A1(n5124), .A2(net76862), .B1(n6223), .B2(net76614), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9634 ( .A(REGFILE_reg_out_21__30_), .ZN(n8748) );
  OAI22_X2 U9635 ( .A1(n8748), .A2(n6121), .B1(n6223), .B2(n6163), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9636 ( .A(REGFILE_reg_out_22__30_), .ZN(n8749) );
  OAI22_X2 U9637 ( .A1(n8749), .A2(n6124), .B1(n6223), .B2(n6165), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9638 ( .A(REGFILE_reg_out_23__30_), .ZN(n8750) );
  OAI22_X2 U9639 ( .A1(n8750), .A2(n6127), .B1(n6223), .B2(n6167), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9640 ( .A(REGFILE_reg_out_24__30_), .ZN(n8751) );
  OAI22_X2 U9641 ( .A1(n8751), .A2(n6129), .B1(n6223), .B2(n6169), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9642 ( .A1(n5924), .A2(n6132), .B1(n6223), .B2(n6171), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9643 ( .A(REGFILE_reg_out_26__30_), .ZN(n8752) );
  OAI22_X2 U9644 ( .A1(n8752), .A2(n6136), .B1(n6223), .B2(n6173), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9645 ( .A1(n6178), .A2(REGFILE_reg_out_29__30_), .ZN(n8753) );
  OAI22_X2 U9646 ( .A1(n5680), .A2(n6139), .B1(n6223), .B2(net76548), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9647 ( .A1(n5070), .A2(n6144), .B1(n6223), .B2(n6182), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9648 ( .A1(n5440), .A2(net76706), .B1(n6223), .B2(n6146), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9649 ( .A1(n5507), .A2(net76692), .B1(n6223), .B2(n6184), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9650 ( .A1(n8756), .A2(n6150), .B1(n6223), .B2(n6186), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9651 ( .A1(n8757), .A2(n6153), .B1(n6223), .B2(n6188), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9652 ( .A1(multOut[28]), .A2(net92392), .ZN(n8783) );
  INV_X4 U9653 ( .A(n10094), .ZN(n8759) );
  NAND2_X2 U9654 ( .A1(net77084), .A2(n10466), .ZN(n8763) );
  NAND2_X2 U9655 ( .A1(n8759), .A2(n8978), .ZN(n8762) );
  NAND2_X2 U9656 ( .A1(n6083), .A2(n8977), .ZN(n8761) );
  NAND2_X2 U9657 ( .A1(n6082), .A2(n8976), .ZN(n8760) );
  NAND4_X2 U9658 ( .A1(n8763), .A2(n8762), .A3(n8761), .A4(n8760), .ZN(n8890)
         );
  NAND2_X2 U9659 ( .A1(n8854), .A2(n8890), .ZN(n8764) );
  OAI22_X2 U9660 ( .A1(n4896), .A2(n9802), .B1(n4922), .B2(n9770), .ZN(n8769)
         );
  INV_X4 U9661 ( .A(n8772), .ZN(n8775) );
  INV_X4 U9662 ( .A(n8773), .ZN(n8774) );
  NAND2_X2 U9663 ( .A1(n8775), .A2(n8774), .ZN(n8779) );
  INV_X4 U9664 ( .A(n10441), .ZN(n10317) );
  NAND2_X2 U9665 ( .A1(net70701), .A2(n10317), .ZN(n8777) );
  NAND2_X2 U9666 ( .A1(n8777), .A2(n8776), .ZN(n8778) );
  AOI21_X4 U9667 ( .B1(n8780), .B2(n8779), .A(n8778), .ZN(n8781) );
  NAND3_X2 U9668 ( .A1(n8783), .A2(n8782), .A3(n8781), .ZN(dmem_addr_out[28])
         );
  INV_X4 U9669 ( .A(dmem_addr_out[28]), .ZN(n8791) );
  INV_X4 U9670 ( .A(dmem_read_in[12]), .ZN(n9108) );
  INV_X4 U9671 ( .A(dmem_read_in[4]), .ZN(n10083) );
  INV_X4 U9672 ( .A(dmem_read_in[28]), .ZN(n8786) );
  OAI211_X2 U9673 ( .C1(n8791), .C2(net76646), .A(n8790), .B(n8789), .ZN(n8792) );
  OAI22_X2 U9674 ( .A1(n5047), .A2(n6088), .B1(n6221), .B2(net76658), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9675 ( .A1(n5484), .A2(n6091), .B1(n6221), .B2(n6155), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9676 ( .A1(n5494), .A2(n6097), .B1(n6221), .B2(n6094), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9677 ( .A1(n5491), .A2(n6103), .B1(n6221), .B2(n6102), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9678 ( .A1(n5485), .A2(n6108), .B1(n6221), .B2(n6105), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9679 ( .A1(n5568), .A2(n6112), .B1(n6221), .B2(n6157), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9680 ( .A1(n5544), .A2(n6115), .B1(n6221), .B2(n6159), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9681 ( .A1(n5486), .A2(n6118), .B1(n6221), .B2(n6161), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9682 ( .A1(n5357), .A2(net76862), .B1(n6221), .B2(net76614), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9683 ( .A1(n5069), .A2(n6121), .B1(n6221), .B2(n6163), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9684 ( .A1(n5495), .A2(n6124), .B1(n6221), .B2(n6165), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9685 ( .A1(n5351), .A2(n6127), .B1(n6221), .B2(n6167), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9686 ( .A1(n5569), .A2(n6129), .B1(n6221), .B2(n6169), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9687 ( .A1(n5487), .A2(n6132), .B1(n6221), .B2(n6171), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9688 ( .A1(n5545), .A2(n6136), .B1(n6221), .B2(n6173), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9689 ( .A1(n6178), .A2(REGFILE_reg_out_29__28_), .ZN(n8793) );
  OAI22_X2 U9690 ( .A1(n5488), .A2(n6139), .B1(n6221), .B2(net76548), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9691 ( .A1(n6180), .A2(REGFILE_reg_out_30__28_), .ZN(n8794) );
  NAND2_X2 U9692 ( .A1(net76488), .A2(REGFILE_reg_out_31__28_), .ZN(n8795) );
  OAI22_X2 U9693 ( .A1(n5358), .A2(n6144), .B1(n6221), .B2(n6182), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9694 ( .A1(n5565), .A2(net76706), .B1(n6221), .B2(n6146), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9695 ( .A1(n5546), .A2(net76692), .B1(n6221), .B2(n6184), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9696 ( .A1(n5032), .A2(n6150), .B1(n6221), .B2(n6186), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9697 ( .A1(n5547), .A2(n6153), .B1(n6221), .B2(n6188), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9698 ( .A1(net73708), .A2(aluA[17]), .ZN(n8801) );
  OAI211_X2 U9699 ( .C1(n8360), .C2(n8798), .A(n8797), .B(n10649), .ZN(n8800)
         );
  NAND2_X2 U9700 ( .A1(n6190), .A2(n9041), .ZN(n8799) );
  NAND3_X4 U9701 ( .A1(n8801), .A2(n8800), .A3(n8799), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U9702 ( .A(n8803), .B(n8802), .ZN(n8807) );
  INV_X4 U9703 ( .A(n8804), .ZN(n8873) );
  NAND2_X2 U9704 ( .A1(n6190), .A2(n8873), .ZN(n8806) );
  NAND2_X2 U9705 ( .A1(net73708), .A2(aluA[18]), .ZN(n8805) );
  OAI211_X2 U9706 ( .C1(n8807), .C2(n6008), .A(n8806), .B(n8805), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9707 ( .A(n10053), .ZN(n8818) );
  OAI22_X2 U9708 ( .A1(n8810), .A2(net72312), .B1(n8809), .B2(n8808), .ZN(
        n9289) );
  XNOR2_X2 U9709 ( .A(n10931), .B(n4814), .ZN(n9290) );
  INV_X4 U9710 ( .A(n9290), .ZN(n8811) );
  AOI22_X2 U9711 ( .A1(n9289), .A2(n8811), .B1(n10931), .B2(n4814), .ZN(n8920)
         );
  INV_X4 U9712 ( .A(n8813), .ZN(n8812) );
  XNOR2_X2 U9713 ( .A(n10932), .B(n8812), .ZN(n8918) );
  OAI22_X2 U9714 ( .A1(n8813), .A2(n8967), .B1(n8920), .B2(n8918), .ZN(n9542)
         );
  INV_X4 U9715 ( .A(n9543), .ZN(n8814) );
  AOI22_X2 U9716 ( .A1(n9542), .A2(n8814), .B1(n10933), .B2(n4810), .ZN(n10054) );
  AOI22_X2 U9717 ( .A1(n9992), .A2(n9993), .B1(n8820), .B2(aluA[19]), .ZN(
        n9033) );
  XNOR2_X2 U9718 ( .A(n9033), .B(n9028), .ZN(n8835) );
  NAND2_X2 U9719 ( .A1(n8822), .A2(n8821), .ZN(n10241) );
  INV_X4 U9720 ( .A(n10241), .ZN(n8825) );
  INV_X4 U9721 ( .A(n8823), .ZN(n8937) );
  NAND2_X2 U9722 ( .A1(n8937), .A2(n10930), .ZN(n8824) );
  OAI21_X4 U9723 ( .B1(n6005), .B2(n8825), .A(n8824), .ZN(n10063) );
  INV_X4 U9724 ( .A(n10063), .ZN(n8832) );
  NAND2_X2 U9725 ( .A1(n8827), .A2(n8826), .ZN(n9018) );
  NAND2_X2 U9726 ( .A1(n6082), .A2(n9018), .ZN(n8831) );
  NAND2_X2 U9727 ( .A1(n9065), .A2(n5761), .ZN(n8829) );
  NAND2_X2 U9728 ( .A1(n8829), .A2(n8828), .ZN(n10240) );
  NAND2_X2 U9729 ( .A1(net77084), .A2(n10240), .ZN(n8830) );
  OAI211_X2 U9730 ( .C1(net71026), .C2(n8832), .A(n8831), .B(n8830), .ZN(n9986) );
  INV_X4 U9731 ( .A(n9986), .ZN(n8833) );
  NAND2_X2 U9732 ( .A1(multOut[18]), .A2(net81873), .ZN(n8868) );
  NAND2_X2 U9733 ( .A1(n8837), .A2(n8836), .ZN(n9397) );
  INV_X4 U9734 ( .A(n9397), .ZN(n8839) );
  NAND2_X2 U9735 ( .A1(n8937), .A2(net36391), .ZN(n8838) );
  OAI21_X4 U9736 ( .B1(n6005), .B2(n8839), .A(n8838), .ZN(n10065) );
  INV_X4 U9737 ( .A(n10065), .ZN(n8846) );
  NAND2_X2 U9738 ( .A1(n8841), .A2(n8840), .ZN(n9183) );
  NAND2_X2 U9739 ( .A1(n6082), .A2(n9183), .ZN(n8845) );
  NAND2_X2 U9740 ( .A1(n8843), .A2(n8842), .ZN(n9396) );
  NAND2_X2 U9741 ( .A1(net77084), .A2(n9396), .ZN(n8844) );
  OAI211_X2 U9742 ( .C1(net71026), .C2(n8846), .A(n8845), .B(n8844), .ZN(n9010) );
  INV_X4 U9743 ( .A(n9010), .ZN(n8848) );
  INV_X4 U9744 ( .A(n10445), .ZN(n10354) );
  NAND2_X2 U9745 ( .A1(net70701), .A2(n10354), .ZN(n8847) );
  INV_X4 U9746 ( .A(aluA[18]), .ZN(n8849) );
  NAND2_X2 U9747 ( .A1(net77084), .A2(n9975), .ZN(n8853) );
  NAND2_X2 U9748 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_11__MUX_N1), .A2(n6041), .ZN(
        n9341) );
  OAI211_X2 U9749 ( .C1(n9094), .C2(n10404), .A(n9093), .B(n9341), .ZN(n9408)
         );
  NAND2_X2 U9750 ( .A1(n6083), .A2(n9408), .ZN(n8852) );
  NAND2_X2 U9751 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_15__MUX_N1), .A2(n6041), .ZN(
        n9066) );
  NAND2_X2 U9752 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_7__MUX_N1), .A2(n9065), .ZN(
        n8850) );
  NAND2_X2 U9753 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_13__MUX_N1), .A2(n6041), .ZN(
        n9069) );
  OAI211_X2 U9754 ( .C1(n9094), .C2(n10396), .A(n9093), .B(n9069), .ZN(n9977)
         );
  AOI22_X2 U9755 ( .A1(n8728), .A2(n9978), .B1(n6081), .B2(n9977), .ZN(n8851)
         );
  NAND2_X2 U9756 ( .A1(n8854), .A2(n9011), .ZN(n8863) );
  NAND2_X2 U9757 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_14__MUX_N1), .A2(n6041), .ZN(
        n9077) );
  OAI211_X2 U9758 ( .C1(n9094), .C2(n9656), .A(n9093), .B(n9077), .ZN(n10233)
         );
  NAND2_X2 U9759 ( .A1(n6081), .A2(n10233), .ZN(n8860) );
  NAND2_X2 U9760 ( .A1(n6040), .A2(aluA[16]), .ZN(n9082) );
  NAND2_X2 U9761 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_8__MUX_N1), .A2(n9065), .ZN(
        net70717) );
  NAND2_X2 U9762 ( .A1(net70720), .A2(net70534), .ZN(n8856) );
  NAND4_X2 U9763 ( .A1(n9082), .A2(net70717), .A3(n8856), .A4(n8855), .ZN(
        n9548) );
  NAND2_X2 U9764 ( .A1(n8728), .A2(n9548), .ZN(n8859) );
  NAND2_X2 U9765 ( .A1(net77084), .A2(n9546), .ZN(n8858) );
  NAND2_X2 U9766 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_12__MUX_N1), .A2(n6040), .ZN(
        n9080) );
  OAI211_X2 U9767 ( .C1(n9094), .C2(n9954), .A(n9093), .B(n9080), .ZN(n10232)
         );
  NAND2_X2 U9768 ( .A1(n6083), .A2(n10232), .ZN(n8857) );
  NAND4_X2 U9769 ( .A1(n8860), .A2(n8859), .A3(n8858), .A4(n8857), .ZN(n9984)
         );
  NAND2_X2 U9770 ( .A1(n8861), .A2(n9984), .ZN(n8862) );
  NOR3_X4 U9771 ( .A1(n8866), .A2(n8865), .A3(n8864), .ZN(n8867) );
  NAND3_X2 U9772 ( .A1(n8869), .A2(n8868), .A3(n8867), .ZN(dmem_addr_out[18])
         );
  INV_X4 U9773 ( .A(dmem_addr_out[18]), .ZN(n8876) );
  INV_X4 U9774 ( .A(net70740), .ZN(net73167) );
  NAND2_X2 U9775 ( .A1(net73167), .A2(n8870), .ZN(n10079) );
  INV_X4 U9776 ( .A(n10079), .ZN(n10000) );
  INV_X4 U9777 ( .A(dmem_read_in[18]), .ZN(n8871) );
  OAI211_X2 U9778 ( .C1(n8876), .C2(net76646), .A(n8875), .B(n8874), .ZN(n8877) );
  NAND2_X2 U9779 ( .A1(net76270), .A2(n8877), .ZN(n8882) );
  OAI22_X2 U9780 ( .A1(n5088), .A2(n6088), .B1(net76660), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9781 ( .A1(n5886), .A2(n6091), .B1(n6156), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9782 ( .A1(n6192), .A2(n5115), .B1(n6195), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9783 ( .A1(n6196), .A2(n4980), .B1(n6199), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9784 ( .A1(n4925), .A2(n6097), .B1(n6095), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9785 ( .A1(n5089), .A2(n6103), .B1(n6102), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9786 ( .A1(n5878), .A2(n6108), .B1(n6106), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9787 ( .A1(n5138), .A2(n6112), .B1(n6158), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9788 ( .A1(n5139), .A2(n6115), .B1(n6160), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9789 ( .A1(n5262), .A2(n6118), .B1(n6162), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9790 ( .A1(n6200), .A2(n5365), .B1(n6204), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9791 ( .A1(n5263), .A2(net76862), .B1(net76616), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9792 ( .A1(n6205), .A2(n5401), .B1(n6208), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9793 ( .A1(n5140), .A2(n6121), .B1(n6164), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9794 ( .A1(n5071), .A2(n6124), .B1(n6166), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9795 ( .A1(n5090), .A2(n6127), .B1(n6168), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9796 ( .A1(n5141), .A2(n6129), .B1(n6170), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9797 ( .A1(n5857), .A2(n6132), .B1(n6172), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9798 ( .A1(n5142), .A2(n6136), .B1(n6174), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9799 ( .A1(n6209), .A2(n5913), .B1(n6212), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9800 ( .A1(REGFILE_reg_out_28__18_), .A2(n6177), .ZN(n8878) );
  NAND2_X2 U9801 ( .A1(n6178), .A2(REGFILE_reg_out_29__18_), .ZN(n8879) );
  OAI22_X2 U9802 ( .A1(n5785), .A2(n6139), .B1(net76550), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9803 ( .A1(n6180), .A2(REGFILE_reg_out_30__18_), .ZN(n8880) );
  NAND2_X2 U9804 ( .A1(net76488), .A2(REGFILE_reg_out_31__18_), .ZN(n8881) );
  OAI22_X2 U9805 ( .A1(n6215), .A2(n5685), .B1(net76320), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9806 ( .A1(n6217), .A2(n5366), .B1(n6220), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9807 ( .A1(n5030), .A2(n6144), .B1(n6183), .B2(n8882), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9808 ( .A1(n5264), .A2(net76706), .B1(n6147), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9809 ( .A1(n5143), .A2(net76692), .B1(n6185), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9810 ( .A1(n5072), .A2(n6150), .B1(n6187), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9811 ( .A1(n5091), .A2(n6153), .B1(n6189), .B2(n6023), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  XOR2_X2 U9812 ( .A(n8884), .B(n8883), .Z(n8889) );
  NAND2_X2 U9813 ( .A1(net70701), .A2(n10436), .ZN(n8887) );
  NAND2_X2 U9814 ( .A1(n8887), .A2(n8886), .ZN(n8888) );
  INV_X4 U9815 ( .A(n8890), .ZN(n8898) );
  NAND2_X2 U9816 ( .A1(n6083), .A2(n9547), .ZN(n8896) );
  NAND2_X2 U9817 ( .A1(net77084), .A2(n8891), .ZN(n8895) );
  NAND2_X2 U9818 ( .A1(n6082), .A2(n8928), .ZN(n8894) );
  NAND2_X2 U9819 ( .A1(n8759), .A2(n8892), .ZN(n8893) );
  NAND4_X2 U9820 ( .A1(n8896), .A2(n8895), .A3(n8894), .A4(n8893), .ZN(n8897)
         );
  INV_X4 U9821 ( .A(n8897), .ZN(n9768) );
  OAI22_X2 U9822 ( .A1(n10472), .A2(n8898), .B1(n9768), .B2(n10474), .ZN(n8900) );
  OAI22_X2 U9823 ( .A1(n4896), .A2(n9770), .B1(n9771), .B2(n9802), .ZN(n8899)
         );
  NAND2_X2 U9824 ( .A1(multOut[27]), .A2(net92392), .ZN(n8901) );
  NAND3_X4 U9825 ( .A1(n8903), .A2(n8902), .A3(n8901), .ZN(dmem_addr_out[27])
         );
  INV_X4 U9826 ( .A(dmem_addr_out[27]), .ZN(n8911) );
  INV_X4 U9827 ( .A(dmem_read_in[11]), .ZN(n9862) );
  INV_X4 U9828 ( .A(dmem_read_in[3]), .ZN(n10041) );
  INV_X4 U9829 ( .A(dmem_read_in[27]), .ZN(n8906) );
  OAI211_X2 U9830 ( .C1(n8911), .C2(net76646), .A(n8910), .B(n8909), .ZN(n8912) );
  NAND2_X2 U9831 ( .A1(net76270), .A2(n8912), .ZN(n8917) );
  OAI22_X2 U9832 ( .A1(n5548), .A2(n6088), .B1(net76660), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9833 ( .A1(n5489), .A2(n6091), .B1(n6156), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9834 ( .A1(n6192), .A2(n5562), .B1(n6195), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9835 ( .A1(n6196), .A2(n5567), .B1(n6199), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9836 ( .A1(n4955), .A2(n6097), .B1(n6095), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9837 ( .A1(n5492), .A2(n6103), .B1(n6102), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9838 ( .A1(n4949), .A2(n6108), .B1(n6106), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9839 ( .A1(n5493), .A2(n6112), .B1(n6158), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9840 ( .A1(n5549), .A2(n6115), .B1(n6160), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9841 ( .A1(n5490), .A2(n6118), .B1(n6162), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9842 ( .A1(n6200), .A2(n5432), .B1(n6204), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9843 ( .A1(n5359), .A2(net76862), .B1(net76616), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9844 ( .A1(n6205), .A2(n5434), .B1(n6208), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9845 ( .A1(n5352), .A2(n6121), .B1(n6164), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9846 ( .A1(n5496), .A2(n6124), .B1(n6166), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9847 ( .A1(n5353), .A2(n6127), .B1(n6168), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9848 ( .A1(n5354), .A2(n6129), .B1(n6170), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9849 ( .A1(n5360), .A2(n6132), .B1(n6172), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9850 ( .A1(n5355), .A2(n6136), .B1(n6174), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9851 ( .A1(n6209), .A2(n5435), .B1(n6212), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9852 ( .A1(REGFILE_reg_out_28__27_), .A2(n6177), .ZN(n8913) );
  NAND2_X2 U9853 ( .A1(n6178), .A2(REGFILE_reg_out_29__27_), .ZN(n8914) );
  OAI22_X2 U9854 ( .A1(n5361), .A2(n6139), .B1(net76550), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9855 ( .A1(n6180), .A2(REGFILE_reg_out_30__27_), .ZN(n8915) );
  NAND2_X2 U9856 ( .A1(net76488), .A2(REGFILE_reg_out_31__27_), .ZN(n8916) );
  OAI22_X2 U9857 ( .A1(n6215), .A2(n5436), .B1(net76320), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9858 ( .A1(n6217), .A2(n5542), .B1(n6220), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9859 ( .A1(n5497), .A2(n6144), .B1(n6183), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9860 ( .A1(n5566), .A2(net76706), .B1(n6147), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9861 ( .A1(n5550), .A2(net76692), .B1(n6185), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9862 ( .A1(n5362), .A2(n6150), .B1(n6187), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9863 ( .A1(n5356), .A2(n6153), .B1(n6189), .B2(n6025), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9864 ( .A(n8918), .ZN(n8919) );
  XNOR2_X2 U9865 ( .A(n8920), .B(n8919), .ZN(n8923) );
  XNOR2_X2 U9866 ( .A(n10932), .B(n10338), .ZN(n10432) );
  INV_X4 U9867 ( .A(n10432), .ZN(n8921) );
  NAND2_X2 U9868 ( .A1(multOut[22]), .A2(net92392), .ZN(n8947) );
  NAND2_X2 U9869 ( .A1(n10102), .A2(n9976), .ZN(n8927) );
  NAND2_X2 U9870 ( .A1(n9978), .A2(n4880), .ZN(n8926) );
  NAND2_X2 U9871 ( .A1(n6081), .A2(n9975), .ZN(n8925) );
  NAND2_X2 U9872 ( .A1(net77084), .A2(n8977), .ZN(n8924) );
  NAND4_X2 U9873 ( .A1(n8927), .A2(n8926), .A3(n8925), .A4(n8924), .ZN(n9552)
         );
  NAND2_X2 U9874 ( .A1(n10058), .A2(n9552), .ZN(n8934) );
  NAND2_X2 U9875 ( .A1(n8728), .A2(n9547), .ZN(n8932) );
  NAND2_X2 U9876 ( .A1(n4880), .A2(n9548), .ZN(n8931) );
  NAND2_X2 U9877 ( .A1(net77084), .A2(n8928), .ZN(n8930) );
  NAND2_X2 U9878 ( .A1(n6081), .A2(n9546), .ZN(n8929) );
  NAND4_X2 U9879 ( .A1(n8932), .A2(n8931), .A3(n8930), .A4(n8929), .ZN(n9293)
         );
  NAND2_X2 U9880 ( .A1(n10060), .A2(n9293), .ZN(n8933) );
  NAND2_X2 U9881 ( .A1(n8934), .A2(n8933), .ZN(n8945) );
  INV_X4 U9882 ( .A(n9018), .ZN(n8936) );
  NAND2_X2 U9883 ( .A1(n8937), .A2(n5761), .ZN(n8935) );
  NAND2_X2 U9884 ( .A1(n10064), .A2(n9302), .ZN(n8941) );
  INV_X4 U9885 ( .A(n9183), .ZN(n8939) );
  OAI21_X4 U9886 ( .B1(n6005), .B2(n8939), .A(n8938), .ZN(n9982) );
  NAND2_X2 U9887 ( .A1(n10066), .A2(n9982), .ZN(n8940) );
  NAND2_X2 U9888 ( .A1(n8941), .A2(n8940), .ZN(n10070) );
  MUX2_X2 U9889 ( .A(n8942), .B(n10070), .S(net71026), .Z(n8944) );
  NOR3_X4 U9890 ( .A1(n8945), .A2(n8944), .A3(n8943), .ZN(n8946) );
  NAND3_X2 U9891 ( .A1(n8948), .A2(n8947), .A3(n8946), .ZN(dmem_addr_out[22])
         );
  INV_X4 U9892 ( .A(dmem_addr_out[22]), .ZN(n8955) );
  INV_X4 U9893 ( .A(n8950), .ZN(n8964) );
  INV_X4 U9894 ( .A(dmem_read_in[22]), .ZN(n8951) );
  OAI211_X2 U9895 ( .C1(n8955), .C2(net76646), .A(n8954), .B(n8953), .ZN(n8956) );
  OAI22_X2 U9896 ( .A1(n5144), .A2(n6088), .B1(net76660), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9897 ( .A1(n4983), .A2(n6091), .B1(n6156), .B2(n8961), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9898 ( .A1(n6192), .A2(n5367), .B1(n6195), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9899 ( .A1(n6196), .A2(n5621), .B1(n6199), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9900 ( .A1(n5265), .A2(n6097), .B1(n6095), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9901 ( .A1(n5145), .A2(n6103), .B1(n6102), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9902 ( .A1(n5017), .A2(n6108), .B1(n6106), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9903 ( .A1(n5092), .A2(n6112), .B1(n6158), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9904 ( .A1(n5146), .A2(n6115), .B1(n6160), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9905 ( .A1(n5266), .A2(n6118), .B1(n6162), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9906 ( .A1(n6200), .A2(n5368), .B1(n6204), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9907 ( .A1(n5267), .A2(net76862), .B1(net76616), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9908 ( .A1(n6205), .A2(n5504), .B1(n6208), .B2(n8961), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9909 ( .A1(n5147), .A2(n6121), .B1(n6164), .B2(n8961), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9910 ( .A1(n5268), .A2(n6124), .B1(n6166), .B2(n8961), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9911 ( .A1(n5148), .A2(n6127), .B1(n6168), .B2(n8961), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9912 ( .A1(n5149), .A2(n6129), .B1(n6170), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9913 ( .A1(n5269), .A2(n6132), .B1(n6172), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9914 ( .A1(n5150), .A2(n6136), .B1(n6174), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9915 ( .A1(n6209), .A2(n5402), .B1(n6212), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9916 ( .A1(REGFILE_reg_out_28__22_), .A2(n6177), .ZN(n8957) );
  OAI21_X4 U9917 ( .B1(n6213), .B2(n6027), .A(n8957), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9918 ( .A1(n6178), .A2(REGFILE_reg_out_29__22_), .ZN(n8958) );
  OAI21_X4 U9919 ( .B1(n6138), .B2(n6027), .A(n8958), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9920 ( .A1(n5270), .A2(n6139), .B1(net76550), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9921 ( .A1(n6180), .A2(REGFILE_reg_out_30__22_), .ZN(n8959) );
  OAI21_X4 U9922 ( .B1(n6142), .B2(n6027), .A(n8959), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9923 ( .A1(net76488), .A2(REGFILE_reg_out_31__22_), .ZN(n8960) );
  OAI21_X4 U9924 ( .B1(net76480), .B2(n6027), .A(n8960), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9925 ( .A1(n6215), .A2(n5403), .B1(net76320), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9926 ( .A1(n6217), .A2(n5498), .B1(n6220), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9927 ( .A1(n5271), .A2(n6144), .B1(n6183), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9928 ( .A1(n5272), .A2(net76706), .B1(n6147), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9929 ( .A1(n5151), .A2(net76692), .B1(n6185), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9930 ( .A1(n5273), .A2(n6150), .B1(n6187), .B2(n6027), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9931 ( .A1(n5152), .A2(n6153), .B1(n6189), .B2(n8961), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U9932 ( .A(n8963), .B(n8962), .ZN(n8966) );
  NAND2_X2 U9933 ( .A1(n6190), .A2(n8964), .ZN(n8965) );
  OAI221_X2 U9934 ( .B1(n8967), .B2(n4962), .C1(n9533), .C2(n8966), .A(n8965), 
        .ZN(PCLOGIC_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9935 ( .A1(net73708), .A2(n10930), .ZN(n8973) );
  OAI211_X2 U9936 ( .C1(n8349), .C2(n8970), .A(n8969), .B(n10649), .ZN(n8972)
         );
  NAND2_X2 U9937 ( .A1(n6190), .A2(n9000), .ZN(n8971) );
  MUX2_X2 U9938 ( .A(n8974), .B(n9298), .S(net71026), .Z(n8986) );
  INV_X4 U9939 ( .A(n9802), .ZN(n8985) );
  INV_X4 U9940 ( .A(n8975), .ZN(n8982) );
  NAND2_X2 U9941 ( .A1(n8728), .A2(n8976), .ZN(n8981) );
  NAND2_X2 U9942 ( .A1(n6081), .A2(n8977), .ZN(n8980) );
  AOI22_X2 U9943 ( .A1(net77084), .A2(n8978), .B1(n6083), .B2(n9976), .ZN(
        n8979) );
  OAI22_X2 U9944 ( .A1(n10474), .A2(n8982), .B1(n5061), .B2(n10472), .ZN(n8984) );
  AOI211_X4 U9945 ( .C1(n8986), .C2(n8985), .A(n8984), .B(n8983), .ZN(n8996)
         );
  XNOR2_X2 U9946 ( .A(n8988), .B(n8987), .ZN(n8993) );
  NAND2_X2 U9947 ( .A1(n8991), .A2(n8990), .ZN(n8992) );
  NAND2_X2 U9948 ( .A1(multOut[25]), .A2(net92392), .ZN(n8994) );
  OAI211_X2 U9949 ( .C1(n8996), .C2(net72163), .A(n8995), .B(n8994), .ZN(
        dmem_addr_out[25]) );
  INV_X4 U9950 ( .A(dmem_addr_out[25]), .ZN(n9003) );
  INV_X4 U9951 ( .A(dmem_read_in[9]), .ZN(n9373) );
  INV_X4 U9952 ( .A(dmem_read_in[25]), .ZN(n8998) );
  OAI211_X2 U9953 ( .C1(n9003), .C2(net76646), .A(n9002), .B(n9001), .ZN(n9004) );
  NAND2_X2 U9954 ( .A1(net76270), .A2(n9004), .ZN(n9009) );
  OAI22_X2 U9955 ( .A1(n5153), .A2(n6088), .B1(net76660), .B2(n6029), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9956 ( .A1(n5274), .A2(n6091), .B1(n6156), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9957 ( .A1(n6192), .A2(n5551), .B1(n6195), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9958 ( .A1(n6196), .A2(n5501), .B1(n6199), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9959 ( .A1(n5275), .A2(n6097), .B1(n6095), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9960 ( .A1(n5154), .A2(n6103), .B1(n6102), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9961 ( .A1(n5276), .A2(n6108), .B1(n6106), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9962 ( .A1(n5155), .A2(n6112), .B1(n6158), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9963 ( .A1(n5508), .A2(n6115), .B1(n6160), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9964 ( .A1(n5441), .A2(n6118), .B1(n6162), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9965 ( .A1(n6200), .A2(n5552), .B1(n6204), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9966 ( .A1(n5442), .A2(net76862), .B1(net76616), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9967 ( .A1(n6205), .A2(n5404), .B1(n6208), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9968 ( .A1(n5156), .A2(n6121), .B1(n6164), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9969 ( .A1(n5277), .A2(n6124), .B1(n6166), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9970 ( .A1(n5157), .A2(n6127), .B1(n6168), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9971 ( .A1(n5158), .A2(n6129), .B1(n6170), .B2(n6029), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9972 ( .A1(n5278), .A2(n6132), .B1(n6172), .B2(n6029), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9973 ( .A1(n5159), .A2(n6136), .B1(n6174), .B2(n6029), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9974 ( .A1(n6209), .A2(n5405), .B1(n6212), .B2(n6029), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9975 ( .A1(REGFILE_reg_out_28__25_), .A2(n6177), .ZN(n9005) );
  OAI21_X4 U9976 ( .B1(n6213), .B2(n6029), .A(n9005), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9977 ( .A1(n6178), .A2(REGFILE_reg_out_29__25_), .ZN(n9006) );
  OAI21_X4 U9978 ( .B1(n6138), .B2(n6029), .A(n9006), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9979 ( .A1(n5443), .A2(n6139), .B1(net76550), .B2(n6029), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9980 ( .A1(n6180), .A2(REGFILE_reg_out_30__25_), .ZN(n9007) );
  OAI21_X4 U9981 ( .B1(n6142), .B2(n6029), .A(n9007), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9982 ( .A1(net76488), .A2(REGFILE_reg_out_31__25_), .ZN(n9008) );
  OAI21_X4 U9983 ( .B1(net76480), .B2(n6029), .A(n9008), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9984 ( .A1(n6215), .A2(n5406), .B1(net76320), .B2(n6029), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9985 ( .A1(n6217), .A2(n5369), .B1(n6220), .B2(n6029), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9986 ( .A1(n5279), .A2(n6144), .B1(n6183), .B2(n6029), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9987 ( .A1(n5444), .A2(net76706), .B1(n6147), .B2(n6029), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9988 ( .A1(n5509), .A2(net76692), .B1(n6185), .B2(n6029), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9989 ( .A1(n5445), .A2(n6150), .B1(n6187), .B2(n6029), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9990 ( .A1(n5510), .A2(n6153), .B1(n6189), .B2(n6030), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  AOI22_X2 U9991 ( .A1(net71092), .A2(n9011), .B1(net71094), .B2(n9010), .ZN(
        n9026) );
  NAND2_X2 U9992 ( .A1(net77084), .A2(n9548), .ZN(n9016) );
  NAND2_X2 U9993 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_10__MUX_N1), .A2(n6041), .ZN(
        n9361) );
  OAI211_X2 U9994 ( .C1(n9094), .C2(n10109), .A(n9093), .B(n9361), .ZN(n10230)
         );
  NAND2_X2 U9995 ( .A1(n6083), .A2(n10230), .ZN(n9015) );
  NAND2_X2 U9996 ( .A1(n6081), .A2(n10232), .ZN(n9014) );
  NAND2_X2 U9997 ( .A1(n8728), .A2(n10233), .ZN(n9013) );
  NAND4_X2 U9998 ( .A1(n9016), .A2(n9015), .A3(n9014), .A4(n9013), .ZN(n9194)
         );
  NAND2_X2 U9999 ( .A1(n10280), .A2(n9194), .ZN(n9025) );
  INV_X4 U10000 ( .A(n9606), .ZN(net71085) );
  NAND2_X2 U10001 ( .A1(n6081), .A2(n10241), .ZN(n9022) );
  NAND2_X2 U10002 ( .A1(net77086), .A2(n10238), .ZN(n9021) );
  NAND2_X2 U10003 ( .A1(n8728), .A2(n10240), .ZN(n9020) );
  NAND2_X2 U10004 ( .A1(n6083), .A2(n9018), .ZN(n9019) );
  NAND4_X2 U10005 ( .A1(n9022), .A2(n9021), .A3(n9020), .A4(n9019), .ZN(n9182)
         );
  NAND3_X2 U10006 ( .A1(n9026), .A2(n9025), .A3(n9024), .ZN(n9027) );
  MUX2_X2 U10007 ( .A(n9027), .B(multOut[17]), .S(net76452), .Z(n9038) );
  INV_X4 U10008 ( .A(n9028), .ZN(n9032) );
  NAND2_X2 U10009 ( .A1(n9030), .A2(aluA[18]), .ZN(n9031) );
  XNOR2_X2 U10010 ( .A(n9052), .B(n9053), .ZN(n9036) );
  NAND2_X2 U10011 ( .A1(net71078), .A2(aluA[17]), .ZN(n9034) );
  OAI22_X2 U10012 ( .A1(n9036), .A2(net70691), .B1(n9035), .B2(n9034), .ZN(
        n9037) );
  NOR2_X4 U10013 ( .A1(n9038), .A2(n9037), .ZN(n9044) );
  INV_X4 U10014 ( .A(n9044), .ZN(dmem_addr_out[17]) );
  INV_X4 U10015 ( .A(dmem_read_in[17]), .ZN(n9039) );
  OAI211_X2 U10016 ( .C1(n9044), .C2(net76646), .A(n9043), .B(n9042), .ZN(
        n9045) );
  OAI22_X2 U10017 ( .A1(n5093), .A2(n6088), .B1(net76660), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10018 ( .A1(n5073), .A2(n6091), .B1(n6156), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10019 ( .A1(n6192), .A2(n5370), .B1(n6194), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10020 ( .A1(n6196), .A2(n5620), .B1(n6198), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10021 ( .A1(n5280), .A2(n6097), .B1(n6095), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10022 ( .A1(n5160), .A2(n6103), .B1(n6102), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10023 ( .A1(n5018), .A2(n6108), .B1(n6106), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10024 ( .A1(n5094), .A2(n6112), .B1(n6158), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10025 ( .A1(n5095), .A2(n6115), .B1(n6160), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10026 ( .A1(n5074), .A2(n6118), .B1(n6162), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10027 ( .A1(n6200), .A2(n5116), .B1(n6203), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10028 ( .A1(n5075), .A2(net76862), .B1(net76616), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10029 ( .A1(n6205), .A2(n5407), .B1(n6207), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10030 ( .A1(n5161), .A2(n6121), .B1(n6164), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10031 ( .A1(n5281), .A2(n6124), .B1(n6166), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10032 ( .A1(n5162), .A2(n6127), .B1(n6168), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10033 ( .A1(n5096), .A2(n6129), .B1(n6170), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10034 ( .A1(n5019), .A2(n6132), .B1(n6172), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10035 ( .A1(n5097), .A2(n6136), .B1(n6174), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10036 ( .A1(n6209), .A2(n5027), .B1(n6211), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10037 ( .A1(REGFILE_reg_out_28__17_), .A2(n6177), .ZN(n9046) );
  NAND2_X2 U10038 ( .A1(n6178), .A2(REGFILE_reg_out_29__17_), .ZN(n9047) );
  OAI22_X2 U10039 ( .A1(n5020), .A2(n6139), .B1(net76550), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10040 ( .A1(n6180), .A2(REGFILE_reg_out_30__17_), .ZN(n9048) );
  NAND2_X2 U10041 ( .A1(net76488), .A2(REGFILE_reg_out_31__17_), .ZN(n9049) );
  OAI22_X2 U10042 ( .A1(n6215), .A2(n5111), .B1(net76318), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10043 ( .A1(n6217), .A2(n5117), .B1(n6219), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10044 ( .A1(n5076), .A2(n6144), .B1(n6183), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10045 ( .A1(n5077), .A2(net76706), .B1(n6147), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10046 ( .A1(n5098), .A2(net76692), .B1(n6185), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10047 ( .A1(n5078), .A2(n6150), .B1(n6187), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10048 ( .A1(n5099), .A2(n6153), .B1(n6189), .B2(n6032), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10049 ( .A1(multOut[12]), .A2(net92392), .ZN(n9106) );
  XNOR2_X2 U10050 ( .A(n9351), .B(n9075), .ZN(n9352) );
  INV_X4 U10051 ( .A(n9352), .ZN(n9063) );
  AOI22_X2 U10052 ( .A1(n9053), .A2(n9052), .B1(n9051), .B2(aluA[17]), .ZN(
        n9179) );
  INV_X4 U10053 ( .A(n9179), .ZN(n9056) );
  AOI22_X2 U10054 ( .A1(n9178), .A2(n9056), .B1(n9055), .B2(aluA[16]), .ZN(
        n10287) );
  OAI22_X2 U10055 ( .A1(n9058), .A2(n10463), .B1(n10287), .B2(n4807), .ZN(
        n10253) );
  XNOR2_X2 U10056 ( .A(n9059), .B(n10247), .ZN(n10254) );
  AOI22_X2 U10057 ( .A1(n10253), .A2(n10254), .B1(
        WIRE_ALU_A_MUX2TO1_32BIT_14__MUX_N1), .B2(n9059), .ZN(n9393) );
  XNOR2_X2 U10058 ( .A(n9060), .B(n10368), .ZN(n9392) );
  INV_X4 U10059 ( .A(n9392), .ZN(n9062) );
  NAND2_X2 U10060 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_13__MUX_N1), .A2(n9060), .ZN(
        n9061) );
  XNOR2_X2 U10061 ( .A(n9063), .B(n9353), .ZN(n9064) );
  NAND2_X2 U10062 ( .A1(net71271), .A2(n9064), .ZN(n9105) );
  NAND2_X2 U10063 ( .A1(net70720), .A2(net80189), .ZN(n9067) );
  NAND2_X2 U10064 ( .A1(n10931), .A2(n9065), .ZN(n10462) );
  NAND2_X2 U10065 ( .A1(n10102), .A2(n10239), .ZN(n9074) );
  NAND2_X2 U10066 ( .A1(net77086), .A2(n9838), .ZN(n9073) );
  NAND2_X2 U10067 ( .A1(n6083), .A2(n10240), .ZN(n9072) );
  NAND2_X2 U10068 ( .A1(n6081), .A2(n10238), .ZN(n9071) );
  NAND4_X2 U10069 ( .A1(n9074), .A2(n9073), .A3(n9072), .A4(n9071), .ZN(n9403)
         );
  INV_X4 U10070 ( .A(n10423), .ZN(n10373) );
  NAND2_X2 U10071 ( .A1(n8759), .A2(n9500), .ZN(n9086) );
  NAND2_X2 U10072 ( .A1(net77086), .A2(n9621), .ZN(n9085) );
  NAND2_X2 U10073 ( .A1(n6083), .A2(n9396), .ZN(n9084) );
  NAND2_X2 U10074 ( .A1(n6081), .A2(n9395), .ZN(n9083) );
  NAND4_X2 U10075 ( .A1(n9086), .A2(n9085), .A3(n9084), .A4(n9083), .ZN(n9837)
         );
  NAND2_X2 U10076 ( .A1(n10066), .A2(n9837), .ZN(n9092) );
  NAND2_X2 U10077 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_7__MUX_N1), .A2(n6040), .ZN(
        n9594) );
  NAND2_X2 U10078 ( .A1(net70696), .A2(n9581), .ZN(n9580) );
  NAND2_X2 U10079 ( .A1(n9594), .A2(n9580), .ZN(n9493) );
  NAND2_X2 U10080 ( .A1(n6081), .A2(n9493), .ZN(n9090) );
  NAND2_X2 U10081 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_9__MUX_N1), .A2(n6041), .ZN(
        n9342) );
  OAI211_X2 U10082 ( .C1(n9094), .C2(net71273), .A(n9093), .B(n9342), .ZN(
        n9407) );
  NAND2_X2 U10083 ( .A1(n8759), .A2(n9407), .ZN(n9089) );
  NAND2_X2 U10084 ( .A1(net77086), .A2(n9408), .ZN(n9088) );
  NAND2_X2 U10085 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_5__MUX_N1), .A2(n6041), .ZN(
        n9598) );
  NAND2_X2 U10086 ( .A1(n9598), .A2(n9580), .ZN(n9585) );
  NAND2_X2 U10087 ( .A1(n4880), .A2(n9585), .ZN(n9087) );
  NAND4_X2 U10088 ( .A1(n9090), .A2(n9089), .A3(n9088), .A4(n9087), .ZN(n9852)
         );
  NAND2_X2 U10089 ( .A1(n10058), .A2(n9852), .ZN(n9091) );
  NAND2_X2 U10090 ( .A1(n9092), .A2(n9091), .ZN(n9102) );
  NAND2_X2 U10091 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_6__MUX_N1), .A2(n6040), .ZN(
        n9618) );
  NAND2_X2 U10092 ( .A1(n9618), .A2(n9580), .ZN(n9845) );
  NAND2_X2 U10093 ( .A1(n4880), .A2(n9845), .ZN(n9098) );
  NAND2_X2 U10094 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_8__MUX_N1), .A2(n6040), .ZN(
        n9498) );
  OAI211_X2 U10095 ( .C1(net70535), .C2(n9094), .A(n9498), .B(n9093), .ZN(
        n10231) );
  NAND2_X2 U10096 ( .A1(n6081), .A2(n10231), .ZN(n9097) );
  NAND2_X2 U10097 ( .A1(net77086), .A2(n10232), .ZN(n9096) );
  NAND2_X2 U10098 ( .A1(n8728), .A2(n10230), .ZN(n9095) );
  NAND4_X2 U10099 ( .A1(n9098), .A2(n9097), .A3(n9096), .A4(n9095), .ZN(n9404)
         );
  INV_X4 U10100 ( .A(n9404), .ZN(n9100) );
  NOR2_X4 U10101 ( .A1(n9102), .A2(n9101), .ZN(n9103) );
  NAND4_X2 U10102 ( .A1(n9106), .A2(n9105), .A3(n9104), .A4(n9103), .ZN(
        dmem_addr_out[12]) );
  NAND2_X2 U10103 ( .A1(net76650), .A2(dmem_addr_out[12]), .ZN(n9112) );
  INV_X4 U10104 ( .A(n9107), .ZN(n9110) );
  AOI21_X4 U10105 ( .B1(n9110), .B2(net77030), .A(n9109), .ZN(n9111) );
  NAND3_X2 U10106 ( .A1(n9112), .A2(net70740), .A3(n9111), .ZN(n9113) );
  NAND2_X2 U10107 ( .A1(n6034), .A2(n4992), .ZN(n9115) );
  NAND2_X2 U10108 ( .A1(n4867), .A2(REGFILE_reg_out_0__12_), .ZN(n9114) );
  NAND2_X2 U10109 ( .A1(n9115), .A2(n9114), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10110 ( .A1(n6034), .A2(n4990), .ZN(n9117) );
  NAND2_X2 U10111 ( .A1(n6093), .A2(REGFILE_reg_out_10__12_), .ZN(n9116) );
  NAND2_X2 U10112 ( .A1(n9117), .A2(n9116), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10113 ( .A1(n6034), .A2(n4998), .ZN(n9119) );
  NAND2_X2 U10114 ( .A1(REGFILE_reg_out_11__12_), .A2(n4869), .ZN(n9118) );
  NAND2_X2 U10115 ( .A1(n9119), .A2(n9118), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10116 ( .A1(n6034), .A2(n4993), .ZN(n9121) );
  NAND2_X2 U10117 ( .A1(n9121), .A2(n9120), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10118 ( .A1(n6034), .A2(n6096), .ZN(n9123) );
  NAND2_X2 U10119 ( .A1(n9123), .A2(n9122), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10120 ( .A1(n6034), .A2(n6101), .ZN(n9125) );
  NAND2_X2 U10121 ( .A1(n4805), .A2(REGFILE_reg_out_14__12_), .ZN(n9124) );
  NAND2_X2 U10122 ( .A1(n9125), .A2(n9124), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10123 ( .A1(n6034), .A2(n6107), .ZN(n9127) );
  NAND2_X2 U10124 ( .A1(n9127), .A2(n9126), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10125 ( .A1(n6034), .A2(n4994), .ZN(n9129) );
  NAND2_X2 U10126 ( .A1(n4891), .A2(REGFILE_reg_out_16__12_), .ZN(n9128) );
  NAND2_X2 U10127 ( .A1(n9129), .A2(n9128), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10128 ( .A1(n6034), .A2(n4999), .ZN(n9131) );
  NAND2_X2 U10129 ( .A1(n4892), .A2(REGFILE_reg_out_17__12_), .ZN(n9130) );
  NAND2_X2 U10130 ( .A1(n9131), .A2(n9130), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10131 ( .A1(n6034), .A2(n5000), .ZN(n9133) );
  NAND2_X2 U10132 ( .A1(n4884), .A2(REGFILE_reg_out_18__12_), .ZN(n9132) );
  NAND2_X2 U10133 ( .A1(n9133), .A2(n9132), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10134 ( .A1(n6033), .A2(n5001), .ZN(n9135) );
  NAND2_X2 U10135 ( .A1(REGFILE_reg_out_19__12_), .A2(n4876), .ZN(n9134) );
  NAND2_X2 U10136 ( .A1(n9135), .A2(n9134), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10137 ( .A1(n6033), .A2(n4997), .ZN(n9137) );
  NAND2_X2 U10138 ( .A1(n4877), .A2(REGFILE_reg_out_1__12_), .ZN(n9136) );
  NAND2_X2 U10139 ( .A1(n9137), .A2(n9136), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10140 ( .A1(n6033), .A2(n4903), .ZN(n9139) );
  NAND2_X2 U10141 ( .A1(REGFILE_reg_out_20__12_), .A2(n4868), .ZN(n9138) );
  NAND2_X2 U10142 ( .A1(n9139), .A2(n9138), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10143 ( .A1(n6033), .A2(n4904), .ZN(n9141) );
  NAND2_X2 U10144 ( .A1(n4882), .A2(REGFILE_reg_out_21__12_), .ZN(n9140) );
  NAND2_X2 U10145 ( .A1(n9141), .A2(n9140), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10146 ( .A1(n6033), .A2(n4905), .ZN(n9143) );
  NAND2_X2 U10147 ( .A1(n4888), .A2(REGFILE_reg_out_22__12_), .ZN(n9142) );
  NAND2_X2 U10148 ( .A1(n9143), .A2(n9142), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10149 ( .A1(n6033), .A2(n4906), .ZN(n9145) );
  NAND2_X2 U10150 ( .A1(n4883), .A2(REGFILE_reg_out_23__12_), .ZN(n9144) );
  NAND2_X2 U10151 ( .A1(n9145), .A2(n9144), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10152 ( .A1(n6033), .A2(n4995), .ZN(n9147) );
  NAND2_X2 U10153 ( .A1(n4875), .A2(REGFILE_reg_out_24__12_), .ZN(n9146) );
  NAND2_X2 U10154 ( .A1(n9147), .A2(n9146), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10155 ( .A1(n6033), .A2(n5002), .ZN(n9149) );
  NAND2_X2 U10156 ( .A1(n4878), .A2(REGFILE_reg_out_25__12_), .ZN(n9148) );
  NAND2_X2 U10157 ( .A1(n9149), .A2(n9148), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10158 ( .A1(n6033), .A2(n5003), .ZN(n9151) );
  NAND2_X2 U10159 ( .A1(n4893), .A2(REGFILE_reg_out_26__12_), .ZN(n9150) );
  NAND2_X2 U10160 ( .A1(n9151), .A2(n9150), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10161 ( .A1(n6033), .A2(n5004), .ZN(n9153) );
  NAND2_X2 U10162 ( .A1(REGFILE_reg_out_27__12_), .A2(n4872), .ZN(n9152) );
  NAND2_X2 U10163 ( .A1(n9153), .A2(n9152), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10164 ( .A1(n6033), .A2(n4806), .ZN(n9155) );
  NAND2_X2 U10165 ( .A1(n9155), .A2(n9154), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10166 ( .A1(n6033), .A2(n10607), .ZN(n9157) );
  NAND2_X2 U10167 ( .A1(n6178), .A2(REGFILE_reg_out_29__12_), .ZN(n9156) );
  NAND2_X2 U10168 ( .A1(n9157), .A2(n9156), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10169 ( .A1(n6033), .A2(n5005), .ZN(n9159) );
  NAND2_X2 U10170 ( .A1(n4879), .A2(REGFILE_reg_out_2__12_), .ZN(n9158) );
  NAND2_X2 U10171 ( .A1(n9159), .A2(n9158), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10172 ( .A1(n6033), .A2(n10614), .ZN(n9161) );
  NAND2_X2 U10173 ( .A1(n6180), .A2(REGFILE_reg_out_30__12_), .ZN(n9160) );
  NAND2_X2 U10174 ( .A1(n9161), .A2(n9160), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10175 ( .A1(n6034), .A2(net70574), .ZN(n9163) );
  NAND2_X2 U10176 ( .A1(net76488), .A2(REGFILE_reg_out_31__12_), .ZN(n9162) );
  NAND2_X2 U10177 ( .A1(n9163), .A2(n9162), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10178 ( .A1(n6034), .A2(n5009), .ZN(n9165) );
  NAND2_X2 U10180 ( .A1(n9165), .A2(n9164), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10181 ( .A1(n6034), .A2(n4996), .ZN(n9167) );
  NAND2_X2 U10182 ( .A1(REGFILE_reg_out_4__12_), .A2(n4870), .ZN(n9166) );
  NAND2_X2 U10183 ( .A1(n9167), .A2(n9166), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10184 ( .A1(n6034), .A2(n5006), .ZN(n9169) );
  NAND2_X2 U10185 ( .A1(n4885), .A2(REGFILE_reg_out_5__12_), .ZN(n9168) );
  NAND2_X2 U10186 ( .A1(n9169), .A2(n9168), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10187 ( .A1(n6034), .A2(n6148), .ZN(n9171) );
  NAND2_X2 U10188 ( .A1(n4889), .A2(REGFILE_reg_out_6__12_), .ZN(n9170) );
  NAND2_X2 U10189 ( .A1(n9171), .A2(n9170), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10190 ( .A1(n6033), .A2(n5007), .ZN(n9173) );
  NAND2_X2 U10191 ( .A1(n4886), .A2(REGFILE_reg_out_7__12_), .ZN(n9172) );
  NAND2_X2 U10192 ( .A1(n9173), .A2(n9172), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10193 ( .A1(n6033), .A2(n4991), .ZN(n9175) );
  NAND2_X2 U10195 ( .A1(n9175), .A2(n9174), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10196 ( .A1(n6034), .A2(n5008), .ZN(n9177) );
  NAND2_X2 U10197 ( .A1(n4887), .A2(REGFILE_reg_out_9__12_), .ZN(n9176) );
  NAND2_X2 U10198 ( .A1(n9177), .A2(n9176), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10199 ( .A1(multOut[16]), .A2(net92392), .ZN(n9202) );
  XNOR2_X2 U10200 ( .A(n9179), .B(n9178), .ZN(n9180) );
  NAND2_X2 U10201 ( .A1(net71271), .A2(n9180), .ZN(n9201) );
  NAND2_X2 U10202 ( .A1(n6081), .A2(n9397), .ZN(n9187) );
  NAND2_X2 U10203 ( .A1(net77086), .A2(n9395), .ZN(n9186) );
  NAND2_X2 U10204 ( .A1(n8759), .A2(n9396), .ZN(n9185) );
  NAND2_X2 U10205 ( .A1(n6083), .A2(n9183), .ZN(n9184) );
  NAND4_X2 U10206 ( .A1(n9187), .A2(n9186), .A3(n9185), .A4(n9184), .ZN(n10277) );
  NAND2_X2 U10207 ( .A1(n10066), .A2(n10277), .ZN(n9193) );
  NAND2_X2 U10208 ( .A1(net77086), .A2(n9978), .ZN(n9191) );
  NAND2_X2 U10209 ( .A1(n6083), .A2(n9407), .ZN(n9190) );
  NAND2_X2 U10210 ( .A1(n6081), .A2(n9408), .ZN(n9189) );
  NAND2_X2 U10211 ( .A1(n8759), .A2(n9977), .ZN(n9188) );
  NAND4_X2 U10212 ( .A1(n9191), .A2(n9190), .A3(n9189), .A4(n9188), .ZN(n10278) );
  NAND2_X2 U10213 ( .A1(n10058), .A2(n10278), .ZN(n9192) );
  NAND2_X2 U10214 ( .A1(n9193), .A2(n9192), .ZN(n9198) );
  INV_X4 U10215 ( .A(n9194), .ZN(n9196) );
  NAND4_X2 U10216 ( .A1(n9202), .A2(n9201), .A3(n9200), .A4(n9199), .ZN(
        dmem_addr_out[16]) );
  AOI21_X4 U10217 ( .B1(n9205), .B2(n9204), .A(net76278), .ZN(n9268) );
  NAND2_X2 U10218 ( .A1(n6036), .A2(n4992), .ZN(n9207) );
  NAND2_X2 U10219 ( .A1(n4867), .A2(REGFILE_reg_out_0__16_), .ZN(n9206) );
  NAND2_X2 U10220 ( .A1(n9207), .A2(n9206), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10221 ( .A1(n6036), .A2(n4990), .ZN(n9209) );
  NAND2_X2 U10222 ( .A1(n6093), .A2(REGFILE_reg_out_10__16_), .ZN(n9208) );
  NAND2_X2 U10223 ( .A1(n9209), .A2(n9208), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10224 ( .A1(n6036), .A2(n4998), .ZN(n9211) );
  NAND2_X2 U10225 ( .A1(REGFILE_reg_out_11__16_), .A2(n4869), .ZN(n9210) );
  NAND2_X2 U10226 ( .A1(n9211), .A2(n9210), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10227 ( .A1(n6036), .A2(n4993), .ZN(n9213) );
  NAND2_X2 U10228 ( .A1(n9213), .A2(n9212), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10229 ( .A1(n6036), .A2(n6096), .ZN(n9215) );
  NAND2_X2 U10230 ( .A1(n6100), .A2(REGFILE_reg_out_13__16_), .ZN(n9214) );
  NAND2_X2 U10231 ( .A1(n9215), .A2(n9214), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10232 ( .A1(n6036), .A2(n6101), .ZN(n9217) );
  NAND2_X2 U10233 ( .A1(n4805), .A2(REGFILE_reg_out_14__16_), .ZN(n9216) );
  NAND2_X2 U10234 ( .A1(n9217), .A2(n9216), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10235 ( .A1(n6036), .A2(n6107), .ZN(n9219) );
  NAND2_X2 U10236 ( .A1(n9219), .A2(n9218), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10237 ( .A1(n6036), .A2(n4994), .ZN(n9221) );
  NAND2_X2 U10238 ( .A1(n4891), .A2(REGFILE_reg_out_16__16_), .ZN(n9220) );
  NAND2_X2 U10239 ( .A1(n9221), .A2(n9220), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10240 ( .A1(n6036), .A2(n4999), .ZN(n9223) );
  NAND2_X2 U10241 ( .A1(n4892), .A2(REGFILE_reg_out_17__16_), .ZN(n9222) );
  NAND2_X2 U10242 ( .A1(n9223), .A2(n9222), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10243 ( .A1(n6036), .A2(n5000), .ZN(n9225) );
  NAND2_X2 U10244 ( .A1(n9225), .A2(n9224), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10245 ( .A1(n6035), .A2(n5001), .ZN(n9227) );
  NAND2_X2 U10246 ( .A1(REGFILE_reg_out_19__16_), .A2(n4876), .ZN(n9226) );
  NAND2_X2 U10247 ( .A1(n9227), .A2(n9226), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10248 ( .A1(n6035), .A2(n4997), .ZN(n9229) );
  NAND2_X2 U10249 ( .A1(n4877), .A2(REGFILE_reg_out_1__16_), .ZN(n9228) );
  NAND2_X2 U10250 ( .A1(n9229), .A2(n9228), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10251 ( .A1(n6035), .A2(n4903), .ZN(n9231) );
  NAND2_X2 U10252 ( .A1(REGFILE_reg_out_20__16_), .A2(n4868), .ZN(n9230) );
  NAND2_X2 U10253 ( .A1(n9231), .A2(n9230), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10254 ( .A1(n6035), .A2(n4904), .ZN(n9233) );
  NAND2_X2 U10255 ( .A1(n4882), .A2(REGFILE_reg_out_21__16_), .ZN(n9232) );
  NAND2_X2 U10256 ( .A1(n9233), .A2(n9232), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10257 ( .A1(n6035), .A2(n4905), .ZN(n9235) );
  NAND2_X2 U10258 ( .A1(n9235), .A2(n9234), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10259 ( .A1(n6035), .A2(n4906), .ZN(n9237) );
  NAND2_X2 U10260 ( .A1(n4883), .A2(REGFILE_reg_out_23__16_), .ZN(n9236) );
  NAND2_X2 U10261 ( .A1(n9237), .A2(n9236), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10262 ( .A1(n6035), .A2(n4995), .ZN(n9239) );
  NAND2_X2 U10263 ( .A1(n4875), .A2(REGFILE_reg_out_24__16_), .ZN(n9238) );
  NAND2_X2 U10264 ( .A1(n9239), .A2(n9238), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10265 ( .A1(n6035), .A2(n5002), .ZN(n9241) );
  NAND2_X2 U10266 ( .A1(n9241), .A2(n9240), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10267 ( .A1(n6035), .A2(n5003), .ZN(n9243) );
  NAND2_X2 U10268 ( .A1(n4893), .A2(REGFILE_reg_out_26__16_), .ZN(n9242) );
  NAND2_X2 U10269 ( .A1(n9243), .A2(n9242), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10270 ( .A1(n6035), .A2(n5004), .ZN(n9245) );
  NAND2_X2 U10271 ( .A1(n9245), .A2(n9244), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10272 ( .A1(n6035), .A2(n4806), .ZN(n9247) );
  NAND2_X2 U10273 ( .A1(REGFILE_reg_out_28__16_), .A2(n6177), .ZN(n9246) );
  NAND2_X2 U10274 ( .A1(n9247), .A2(n9246), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10275 ( .A1(n6035), .A2(n10607), .ZN(n9249) );
  NAND2_X2 U10276 ( .A1(n6178), .A2(REGFILE_reg_out_29__16_), .ZN(n9248) );
  NAND2_X2 U10277 ( .A1(n9249), .A2(n9248), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10278 ( .A1(n6035), .A2(n5005), .ZN(n9251) );
  NAND2_X2 U10279 ( .A1(n4879), .A2(REGFILE_reg_out_2__16_), .ZN(n9250) );
  NAND2_X2 U10280 ( .A1(n9251), .A2(n9250), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10281 ( .A1(n6035), .A2(n10614), .ZN(n9253) );
  NAND2_X2 U10282 ( .A1(n6180), .A2(REGFILE_reg_out_30__16_), .ZN(n9252) );
  NAND2_X2 U10283 ( .A1(n9253), .A2(n9252), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10284 ( .A1(n6036), .A2(net70574), .ZN(n9255) );
  NAND2_X2 U10285 ( .A1(net76488), .A2(REGFILE_reg_out_31__16_), .ZN(n9254) );
  NAND2_X2 U10286 ( .A1(n9255), .A2(n9254), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10287 ( .A1(n6036), .A2(n5009), .ZN(n9257) );
  NAND2_X2 U10288 ( .A1(n9257), .A2(n9256), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10289 ( .A1(n6036), .A2(n4996), .ZN(n9259) );
  NAND2_X2 U10290 ( .A1(REGFILE_reg_out_4__16_), .A2(n4870), .ZN(n9258) );
  NAND2_X2 U10291 ( .A1(n9259), .A2(n9258), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10292 ( .A1(n6036), .A2(n5006), .ZN(n9261) );
  NAND2_X2 U10293 ( .A1(n4885), .A2(REGFILE_reg_out_5__16_), .ZN(n9260) );
  NAND2_X2 U10294 ( .A1(n9261), .A2(n9260), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10295 ( .A1(n6036), .A2(n6148), .ZN(n9263) );
  NAND2_X2 U10296 ( .A1(n9263), .A2(n9262), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10297 ( .A1(n6036), .A2(n5007), .ZN(n9265) );
  NAND2_X2 U10298 ( .A1(n4886), .A2(REGFILE_reg_out_7__16_), .ZN(n9264) );
  NAND2_X2 U10299 ( .A1(n9265), .A2(n9264), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10300 ( .A1(n6035), .A2(n4991), .ZN(n9267) );
  NAND2_X2 U10301 ( .A1(n4890), .A2(REGFILE_reg_out_8__16_), .ZN(n9266) );
  NAND2_X2 U10302 ( .A1(n9267), .A2(n9266), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10303 ( .A1(n6035), .A2(n5008), .ZN(n9270) );
  NAND2_X2 U10304 ( .A1(n4887), .A2(REGFILE_reg_out_9__16_), .ZN(n9269) );
  NAND2_X2 U10305 ( .A1(n9270), .A2(n9269), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10306 ( .A1(n10649), .A2(n9272), .ZN(n9275) );
  NAND2_X2 U10307 ( .A1(n6190), .A2(n10003), .ZN(n9274) );
  NAND2_X2 U10308 ( .A1(net73708), .A2(aluA[19]), .ZN(n9273) );
  OAI211_X2 U10309 ( .C1(n9276), .C2(n9275), .A(n9274), .B(n9273), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U10310 ( .A(n9278), .B(n9277), .ZN(n9282) );
  INV_X4 U10311 ( .A(n9279), .ZN(n10080) );
  NAND2_X2 U10312 ( .A1(n6190), .A2(n10080), .ZN(n9281) );
  NAND2_X2 U10313 ( .A1(net73708), .A2(aluA[20]), .ZN(n9280) );
  OAI211_X2 U10314 ( .C1(n9282), .C2(n9533), .A(n9281), .B(n9280), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10315 ( .A1(net73708), .A2(n10931), .ZN(n9288) );
  OAI211_X2 U10316 ( .C1(n8353), .C2(n9285), .A(n9284), .B(n10649), .ZN(n9287)
         );
  NAND2_X2 U10317 ( .A1(n6190), .A2(n9316), .ZN(n9286) );
  XNOR2_X2 U10318 ( .A(n9290), .B(n9289), .ZN(n9292) );
  XNOR2_X2 U10319 ( .A(n10931), .B(n9306), .ZN(n10429) );
  INV_X4 U10320 ( .A(n10429), .ZN(n10336) );
  NAND2_X2 U10321 ( .A1(multOut[23]), .A2(net92392), .ZN(n9311) );
  NAND2_X2 U10322 ( .A1(n10058), .A2(n9293), .ZN(n9296) );
  NAND2_X2 U10323 ( .A1(n10060), .A2(n9294), .ZN(n9295) );
  NAND2_X2 U10324 ( .A1(n9296), .A2(n9295), .ZN(n9309) );
  NAND2_X2 U10325 ( .A1(n10064), .A2(n9297), .ZN(n9300) );
  NAND2_X2 U10326 ( .A1(n10066), .A2(n9298), .ZN(n9299) );
  NAND2_X2 U10327 ( .A1(n9300), .A2(n9299), .ZN(n9305) );
  NAND2_X2 U10328 ( .A1(n10064), .A2(n9301), .ZN(n9304) );
  NAND2_X2 U10329 ( .A1(n10066), .A2(n9302), .ZN(n9303) );
  NAND2_X2 U10330 ( .A1(n9304), .A2(n9303), .ZN(n9558) );
  MUX2_X2 U10331 ( .A(n9305), .B(n9558), .S(net71026), .Z(n9308) );
  NOR3_X4 U10332 ( .A1(n9309), .A2(n9308), .A3(n9307), .ZN(n9310) );
  NAND3_X2 U10333 ( .A1(n9312), .A2(n9311), .A3(n9310), .ZN(dmem_addr_out[23])
         );
  INV_X4 U10334 ( .A(dmem_addr_out[23]), .ZN(n9319) );
  INV_X4 U10335 ( .A(dmem_read_in[7]), .ZN(n10505) );
  INV_X4 U10336 ( .A(dmem_read_in[23]), .ZN(n9314) );
  OAI211_X2 U10337 ( .C1(n9319), .C2(net76646), .A(n9318), .B(n9317), .ZN(
        n9320) );
  OAI22_X2 U10338 ( .A1(n5511), .A2(n6088), .B1(net76660), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10339 ( .A1(n5446), .A2(n6091), .B1(n6156), .B2(n9325), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10340 ( .A1(n6192), .A2(n5553), .B1(n6195), .B2(n9325), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10341 ( .A1(n6196), .A2(n5502), .B1(n6199), .B2(n9325), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10342 ( .A1(n5282), .A2(n6097), .B1(n6095), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10343 ( .A1(n5163), .A2(n6103), .B1(n6102), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10344 ( .A1(n5283), .A2(n6108), .B1(n6106), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10345 ( .A1(n5164), .A2(n6112), .B1(n6158), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10346 ( .A1(n5512), .A2(n6115), .B1(n6160), .B2(n9325), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10347 ( .A1(n5447), .A2(n6118), .B1(n6162), .B2(n9325), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10348 ( .A1(n6200), .A2(n5371), .B1(n6204), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10349 ( .A1(n5284), .A2(net76862), .B1(net76616), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10350 ( .A1(n6206), .A2(n5408), .B1(n6208), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10351 ( .A1(n5165), .A2(n6121), .B1(n6164), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10352 ( .A1(n5285), .A2(n6124), .B1(n6166), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10353 ( .A1(n5166), .A2(n6127), .B1(n6168), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10354 ( .A1(n5513), .A2(n6129), .B1(n6170), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10355 ( .A1(n5448), .A2(n6132), .B1(n6172), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10356 ( .A1(n5167), .A2(n6136), .B1(n6174), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10357 ( .A1(n6209), .A2(n5409), .B1(n6212), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10358 ( .A1(REGFILE_reg_out_28__23_), .A2(n6177), .ZN(n9321) );
  OAI21_X4 U10359 ( .B1(n6213), .B2(n6038), .A(n9321), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10360 ( .A1(n6178), .A2(REGFILE_reg_out_29__23_), .ZN(n9322) );
  OAI21_X4 U10361 ( .B1(n6138), .B2(n6038), .A(n9322), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10362 ( .A1(n5449), .A2(n6139), .B1(net76550), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10363 ( .A1(n6180), .A2(REGFILE_reg_out_30__23_), .ZN(n9323) );
  OAI21_X4 U10364 ( .B1(n6142), .B2(n6038), .A(n9323), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10365 ( .A1(net76488), .A2(REGFILE_reg_out_31__23_), .ZN(n9324) );
  OAI21_X4 U10366 ( .B1(net76480), .B2(n6038), .A(n9324), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10367 ( .A1(n6215), .A2(n5410), .B1(net76320), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10368 ( .A1(n6218), .A2(n5372), .B1(n6220), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10369 ( .A1(n5286), .A2(n6144), .B1(n6183), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10370 ( .A1(n5450), .A2(net76706), .B1(n6147), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10371 ( .A1(n5514), .A2(net76692), .B1(n6185), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10372 ( .A1(n5287), .A2(n6150), .B1(n6187), .B2(n6038), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10373 ( .A1(n5168), .A2(n6153), .B1(n6189), .B2(n9325), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10374 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_2__MUX_N1), .A2(n6040), .ZN(
        n10096) );
  NAND2_X2 U10375 ( .A1(n10096), .A2(n9580), .ZN(n10013) );
  NAND2_X2 U10376 ( .A1(n4880), .A2(n10013), .ZN(n9329) );
  NAND2_X2 U10377 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_4__MUX_N1), .A2(n6040), .ZN(
        n9939) );
  NAND2_X2 U10378 ( .A1(n9939), .A2(n9580), .ZN(n9844) );
  NAND2_X2 U10379 ( .A1(n9844), .A2(n6082), .ZN(n9328) );
  NAND2_X2 U10380 ( .A1(net77086), .A2(n10231), .ZN(n9327) );
  NAND2_X2 U10381 ( .A1(n8759), .A2(n9845), .ZN(n9326) );
  NAND4_X2 U10382 ( .A1(n9329), .A2(n9328), .A3(n9327), .A4(n9326), .ZN(n9492)
         );
  INV_X4 U10383 ( .A(n9492), .ZN(n9336) );
  NAND2_X2 U10384 ( .A1(net77086), .A2(n9407), .ZN(n9334) );
  NAND2_X2 U10385 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_3__MUX_N1), .A2(n6041), .ZN(
        n10019) );
  NAND2_X2 U10386 ( .A1(n10019), .A2(n9580), .ZN(n9935) );
  NAND2_X2 U10387 ( .A1(n4880), .A2(n9935), .ZN(n9333) );
  NAND2_X2 U10388 ( .A1(n6082), .A2(n9585), .ZN(n9332) );
  NAND2_X2 U10389 ( .A1(n10102), .A2(n9493), .ZN(n9331) );
  NAND4_X2 U10390 ( .A1(n9334), .A2(n9333), .A3(n9332), .A4(n9331), .ZN(n10124) );
  INV_X4 U10391 ( .A(n10124), .ZN(n9335) );
  OAI22_X2 U10392 ( .A1(n10474), .A2(n9336), .B1(n10472), .B2(n9335), .ZN(
        n9338) );
  NAND2_X2 U10393 ( .A1(net70720), .A2(n5761), .ZN(n9339) );
  NAND2_X2 U10394 ( .A1(n10102), .A2(n9839), .ZN(n9347) );
  OAI211_X2 U10395 ( .C1(net70868), .C2(n10327), .A(n9343), .B(n9342), .ZN(
        n10024) );
  NAND2_X2 U10396 ( .A1(net77086), .A2(n10024), .ZN(n9346) );
  NAND2_X2 U10397 ( .A1(n6083), .A2(n10239), .ZN(n9345) );
  NAND2_X2 U10398 ( .A1(n6082), .A2(n9838), .ZN(n9344) );
  NAND4_X2 U10399 ( .A1(n9347), .A2(n9346), .A3(n9345), .A4(n9344), .ZN(n9491)
         );
  INV_X4 U10400 ( .A(n9491), .ZN(n9348) );
  NOR2_X4 U10401 ( .A1(n9350), .A2(n9349), .ZN(n9371) );
  AOI22_X2 U10402 ( .A1(n9353), .A2(n9352), .B1(
        WIRE_ALU_A_MUX2TO1_32BIT_12__MUX_N1), .B2(n9351), .ZN(n9833) );
  XNOR2_X2 U10403 ( .A(n9354), .B(n10375), .ZN(n9832) );
  INV_X4 U10404 ( .A(n9832), .ZN(n9356) );
  XNOR2_X2 U10405 ( .A(n9357), .B(n10125), .ZN(n10132) );
  AOI22_X2 U10406 ( .A1(n10131), .A2(n10132), .B1(
        WIRE_ALU_A_MUX2TO1_32BIT_10__MUX_N1), .B2(n9357), .ZN(n9511) );
  XNOR2_X2 U10407 ( .A(n9508), .B(n10382), .ZN(n9507) );
  XNOR2_X2 U10408 ( .A(n9511), .B(n9507), .ZN(n9368) );
  NAND2_X2 U10409 ( .A1(n8759), .A2(n9621), .ZN(n9365) );
  NAND2_X2 U10410 ( .A1(net77086), .A2(n9945), .ZN(n9364) );
  NAND2_X2 U10411 ( .A1(n6083), .A2(n9395), .ZN(n9363) );
  NAND2_X2 U10412 ( .A1(n6082), .A2(n9500), .ZN(n9362) );
  NAND4_X2 U10413 ( .A1(n9365), .A2(n9364), .A3(n9363), .A4(n9362), .ZN(n10126) );
  INV_X4 U10414 ( .A(n10126), .ZN(n9366) );
  INV_X4 U10415 ( .A(dmem_addr_out[9]), .ZN(n9377) );
  OAI22_X2 U10416 ( .A1(n5169), .A2(n6088), .B1(net76660), .B2(n6043), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10417 ( .A1(n5616), .A2(n6091), .B1(n6156), .B2(n6044), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10418 ( .A1(n6193), .A2(n5373), .B1(n6195), .B2(n6044), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10419 ( .A1(n6196), .A2(n5653), .B1(n6199), .B2(n6044), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10420 ( .A1(n5288), .A2(n6097), .B1(n6095), .B2(n6044), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10421 ( .A1(n5170), .A2(n6103), .B1(n6102), .B2(n6044), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10422 ( .A1(n4976), .A2(n6108), .B1(n6106), .B2(n6044), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10423 ( .A1(n5171), .A2(n6112), .B1(n6044), .B2(n6158), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10424 ( .A1(n5172), .A2(n6115), .B1(n6160), .B2(n6044), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10425 ( .A1(n5289), .A2(n6118), .B1(n6162), .B2(n6044), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10426 ( .A1(n6200), .A2(n5374), .B1(n6204), .B2(n6044), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10427 ( .A1(n5290), .A2(net76862), .B1(net76616), .B2(n6044), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10428 ( .A1(n6206), .A2(n5411), .B1(n6208), .B2(n6044), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10429 ( .A1(n5173), .A2(n6121), .B1(n6164), .B2(n6044), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10430 ( .A1(n5291), .A2(n6124), .B1(n6166), .B2(n6044), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10431 ( .A1(n5174), .A2(n6127), .B1(n6168), .B2(n6044), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10432 ( .A1(n5100), .A2(n6129), .B1(n6170), .B2(n6043), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10433 ( .A1(n5021), .A2(n6132), .B1(n6172), .B2(n6043), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10434 ( .A1(n5175), .A2(n6136), .B1(n6174), .B2(n6043), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10435 ( .A1(n6210), .A2(n5412), .B1(n6212), .B2(n6043), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10436 ( .A1(REGFILE_reg_out_28__9_), .A2(n6177), .ZN(n9379) );
  NAND2_X2 U10437 ( .A1(n6178), .A2(REGFILE_reg_out_29__9_), .ZN(n9380) );
  OAI22_X2 U10438 ( .A1(n5022), .A2(n6139), .B1(net76550), .B2(n6043), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10439 ( .A1(n6180), .A2(REGFILE_reg_out_30__9_), .ZN(n9381) );
  NAND2_X2 U10440 ( .A1(n5688), .A2(REGFILE_reg_out_31__9_), .ZN(n9382) );
  OAI22_X2 U10441 ( .A1(n6216), .A2(n5112), .B1(net76320), .B2(n6043), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10442 ( .A1(n6218), .A2(n5375), .B1(n6220), .B2(n6043), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10443 ( .A1(n5292), .A2(n6144), .B1(n6183), .B2(n6043), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10444 ( .A1(n5293), .A2(net76706), .B1(n6147), .B2(n6043), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10445 ( .A1(n5176), .A2(net76692), .B1(n6185), .B2(n6043), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10446 ( .A1(n5294), .A2(n6150), .B1(n6187), .B2(n6043), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10447 ( .A1(n5177), .A2(n6153), .B1(n6189), .B2(n6044), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U10448 ( .A(n9385), .B(n9384), .ZN(n9387) );
  NAND2_X2 U10449 ( .A1(n6190), .A2(n10139), .ZN(n9386) );
  OAI221_X2 U10450 ( .B1(n10125), .B2(n4962), .C1(n6008), .C2(n9387), .A(n9386), .ZN(PCLOGIC_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  XOR2_X2 U10451 ( .A(n9389), .B(n9388), .Z(n9391) );
  NAND2_X2 U10452 ( .A1(n6190), .A2(n9422), .ZN(n9390) );
  OAI221_X2 U10453 ( .B1(n10368), .B2(n4962), .C1(n9391), .C2(n9533), .A(n9390), .ZN(PCLOGIC_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10454 ( .A1(multOut[13]), .A2(net92392), .ZN(n9420) );
  XNOR2_X2 U10455 ( .A(n9393), .B(n9392), .ZN(n9394) );
  NAND2_X2 U10456 ( .A1(net71271), .A2(n9394), .ZN(n9419) );
  NAND2_X2 U10457 ( .A1(n10102), .A2(n9395), .ZN(n9401) );
  NAND2_X2 U10458 ( .A1(net77086), .A2(n9500), .ZN(n9400) );
  NAND2_X2 U10459 ( .A1(n6082), .A2(n9396), .ZN(n9399) );
  NAND2_X2 U10460 ( .A1(n6083), .A2(n9397), .ZN(n9398) );
  NAND4_X2 U10461 ( .A1(n9401), .A2(n9400), .A3(n9399), .A4(n9398), .ZN(n10248) );
  NAND2_X2 U10462 ( .A1(n10066), .A2(n9403), .ZN(n9406) );
  NAND2_X2 U10463 ( .A1(n10058), .A2(n9404), .ZN(n9405) );
  NAND2_X2 U10464 ( .A1(n9406), .A2(n9405), .ZN(n9416) );
  NAND2_X2 U10465 ( .A1(n4880), .A2(n9493), .ZN(n9412) );
  NAND2_X2 U10466 ( .A1(n6082), .A2(n9407), .ZN(n9411) );
  NAND2_X2 U10467 ( .A1(n8759), .A2(n9408), .ZN(n9410) );
  NAND2_X2 U10468 ( .A1(net77086), .A2(n9977), .ZN(n9409) );
  NAND4_X2 U10469 ( .A1(n9412), .A2(n9411), .A3(n9410), .A4(n9409), .ZN(n10246) );
  INV_X4 U10470 ( .A(n10246), .ZN(n9414) );
  NOR2_X4 U10471 ( .A1(n9416), .A2(n9415), .ZN(n9417) );
  NAND4_X2 U10472 ( .A1(n9420), .A2(n9419), .A3(n9418), .A4(n9417), .ZN(
        dmem_addr_out[13]) );
  NAND2_X2 U10473 ( .A1(net76650), .A2(dmem_addr_out[13]), .ZN(n9424) );
  INV_X4 U10474 ( .A(dmem_read_in[13]), .ZN(n9816) );
  NAND3_X2 U10475 ( .A1(n9424), .A2(net70740), .A3(n9423), .ZN(n9425) );
  NAND2_X2 U10476 ( .A1(n6047), .A2(n4992), .ZN(n9428) );
  NAND2_X2 U10477 ( .A1(n4867), .A2(REGFILE_reg_out_0__13_), .ZN(n9427) );
  NAND2_X2 U10478 ( .A1(n9428), .A2(n9427), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10479 ( .A1(n6047), .A2(n4990), .ZN(n9430) );
  NAND2_X2 U10480 ( .A1(n9430), .A2(n9429), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10481 ( .A1(n6047), .A2(n4998), .ZN(n9432) );
  NAND2_X2 U10482 ( .A1(net148736), .A2(n4869), .ZN(n9431) );
  NAND2_X2 U10483 ( .A1(n9432), .A2(n9431), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10484 ( .A1(n6047), .A2(n4993), .ZN(n9434) );
  NAND2_X2 U10485 ( .A1(n9434), .A2(n9433), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10486 ( .A1(n6047), .A2(n6096), .ZN(n9436) );
  NAND2_X2 U10487 ( .A1(n6100), .A2(REGFILE_reg_out_13__13_), .ZN(n9435) );
  NAND2_X2 U10488 ( .A1(n9436), .A2(n9435), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10489 ( .A1(n6047), .A2(n6101), .ZN(n9438) );
  NAND2_X2 U10490 ( .A1(n9438), .A2(n9437), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10491 ( .A1(n6047), .A2(n6107), .ZN(n9440) );
  NAND2_X2 U10492 ( .A1(n4804), .A2(REGFILE_reg_out_15__13_), .ZN(n9439) );
  NAND2_X2 U10493 ( .A1(n9440), .A2(n9439), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10494 ( .A1(n6047), .A2(n4994), .ZN(n9442) );
  NAND2_X2 U10495 ( .A1(n9442), .A2(n9441), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10496 ( .A1(n6047), .A2(n4999), .ZN(n9444) );
  NAND2_X2 U10497 ( .A1(n4892), .A2(REGFILE_reg_out_17__13_), .ZN(n9443) );
  NAND2_X2 U10498 ( .A1(n9444), .A2(n9443), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10499 ( .A1(n6047), .A2(n5000), .ZN(n9446) );
  NAND2_X2 U10500 ( .A1(n4884), .A2(REGFILE_reg_out_18__13_), .ZN(n9445) );
  NAND2_X2 U10501 ( .A1(n9446), .A2(n9445), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10502 ( .A1(n6046), .A2(n5001), .ZN(n9448) );
  NAND2_X2 U10503 ( .A1(REGFILE_reg_out_19__13_), .A2(n4876), .ZN(n9447) );
  NAND2_X2 U10504 ( .A1(n9448), .A2(n9447), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10505 ( .A1(n6046), .A2(n4997), .ZN(n9450) );
  NAND2_X2 U10506 ( .A1(n9450), .A2(n9449), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10507 ( .A1(n6046), .A2(n4903), .ZN(n9452) );
  NAND2_X2 U10508 ( .A1(REGFILE_reg_out_20__13_), .A2(n4868), .ZN(n9451) );
  NAND2_X2 U10509 ( .A1(n9452), .A2(n9451), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10510 ( .A1(n6046), .A2(n4904), .ZN(n9454) );
  NAND2_X2 U10511 ( .A1(n4882), .A2(REGFILE_reg_out_21__13_), .ZN(n9453) );
  NAND2_X2 U10512 ( .A1(n9454), .A2(n9453), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10513 ( .A1(n6046), .A2(n4905), .ZN(n9456) );
  NAND2_X2 U10514 ( .A1(n4888), .A2(REGFILE_reg_out_22__13_), .ZN(n9455) );
  NAND2_X2 U10515 ( .A1(n9456), .A2(n9455), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10516 ( .A1(n6046), .A2(n4906), .ZN(n9458) );
  NAND2_X2 U10517 ( .A1(n4883), .A2(REGFILE_reg_out_23__13_), .ZN(n9457) );
  NAND2_X2 U10518 ( .A1(n9458), .A2(n9457), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10519 ( .A1(n6046), .A2(n4995), .ZN(n9460) );
  NAND2_X2 U10520 ( .A1(n9460), .A2(n9459), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10521 ( .A1(n6046), .A2(n5002), .ZN(n9462) );
  NAND2_X2 U10522 ( .A1(n4878), .A2(REGFILE_reg_out_25__13_), .ZN(n9461) );
  NAND2_X2 U10523 ( .A1(n9462), .A2(n9461), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10524 ( .A1(n6046), .A2(n5003), .ZN(n9464) );
  NAND2_X2 U10525 ( .A1(n9464), .A2(n9463), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10526 ( .A1(n6046), .A2(n5004), .ZN(n9466) );
  NAND2_X2 U10527 ( .A1(REGFILE_reg_out_27__13_), .A2(n4872), .ZN(n9465) );
  NAND2_X2 U10528 ( .A1(n9466), .A2(n9465), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10529 ( .A1(n6046), .A2(n4806), .ZN(n9468) );
  NAND2_X2 U10530 ( .A1(n9468), .A2(n9467), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10531 ( .A1(n6046), .A2(n10607), .ZN(n9470) );
  NAND2_X2 U10532 ( .A1(n6178), .A2(REGFILE_reg_out_29__13_), .ZN(n9469) );
  NAND2_X2 U10533 ( .A1(n9470), .A2(n9469), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10534 ( .A1(n6047), .A2(n5005), .ZN(n9472) );
  NAND2_X2 U10535 ( .A1(n9472), .A2(n9471), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10536 ( .A1(n6046), .A2(n10614), .ZN(n9474) );
  NAND2_X2 U10537 ( .A1(n9474), .A2(n9473), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10538 ( .A1(n6047), .A2(net70574), .ZN(n9476) );
  NAND2_X2 U10539 ( .A1(n5688), .A2(REGFILE_reg_out_31__13_), .ZN(n9475) );
  NAND2_X2 U10540 ( .A1(n9476), .A2(n9475), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10541 ( .A1(n6047), .A2(n5009), .ZN(n9478) );
  NAND2_X2 U10542 ( .A1(REGFILE_reg_out_3__13_), .A2(n4871), .ZN(n9477) );
  NAND2_X2 U10543 ( .A1(n9478), .A2(n9477), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10544 ( .A1(n6046), .A2(n4996), .ZN(n9480) );
  NAND2_X2 U10545 ( .A1(REGFILE_reg_out_4__13_), .A2(n4870), .ZN(n9479) );
  NAND2_X2 U10546 ( .A1(n9480), .A2(n9479), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10547 ( .A1(n6046), .A2(n5006), .ZN(n9482) );
  NAND2_X2 U10548 ( .A1(n4885), .A2(REGFILE_reg_out_5__13_), .ZN(n9481) );
  NAND2_X2 U10549 ( .A1(n9482), .A2(n9481), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10550 ( .A1(n6047), .A2(n6148), .ZN(n9484) );
  NAND2_X2 U10551 ( .A1(n4889), .A2(REGFILE_reg_out_6__13_), .ZN(n9483) );
  NAND2_X2 U10552 ( .A1(n9484), .A2(n9483), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10553 ( .A1(n6046), .A2(n5007), .ZN(n9486) );
  NAND2_X2 U10554 ( .A1(n4886), .A2(REGFILE_reg_out_7__13_), .ZN(n9485) );
  NAND2_X2 U10555 ( .A1(n9486), .A2(n9485), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10556 ( .A1(n6047), .A2(n4991), .ZN(n9488) );
  NAND2_X2 U10557 ( .A1(n9488), .A2(n9487), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10558 ( .A1(n6047), .A2(n5008), .ZN(n9490) );
  NAND2_X2 U10559 ( .A1(n4887), .A2(REGFILE_reg_out_9__13_), .ZN(n9489) );
  NAND2_X2 U10560 ( .A1(n9490), .A2(n9489), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  AOI22_X2 U10561 ( .A1(net71092), .A2(n9492), .B1(net71094), .B2(n9491), .ZN(
        n9505) );
  NAND2_X2 U10562 ( .A1(n6082), .A2(n9935), .ZN(n9497) );
  NAND2_X2 U10563 ( .A1(n4880), .A2(n10091), .ZN(n9496) );
  NAND2_X2 U10564 ( .A1(n10102), .A2(n9585), .ZN(n9495) );
  NAND2_X2 U10565 ( .A1(net77086), .A2(n9493), .ZN(n9494) );
  NAND4_X2 U10566 ( .A1(n9497), .A2(n9496), .A3(n9495), .A4(n9494), .ZN(n9690)
         );
  NAND2_X2 U10567 ( .A1(n10280), .A2(n9690), .ZN(n9504) );
  OAI211_X2 U10568 ( .C1(net72312), .C2(net70868), .A(n9499), .B(n9498), .ZN(
        n10103) );
  AOI22_X2 U10569 ( .A1(net77084), .A2(n10103), .B1(n8728), .B2(n9945), .ZN(
        n9502) );
  AOI22_X2 U10570 ( .A1(n6082), .A2(n9621), .B1(n6083), .B2(n9500), .ZN(n9501)
         );
  NAND2_X2 U10571 ( .A1(n9502), .A2(n9501), .ZN(n9685) );
  INV_X4 U10572 ( .A(n10419), .ZN(n10387) );
  NAND3_X2 U10573 ( .A1(n9505), .A2(n9504), .A3(n9503), .ZN(n9506) );
  INV_X4 U10575 ( .A(n9507), .ZN(n9510) );
  NAND2_X2 U10576 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_9__MUX_N1), .A2(n9508), .ZN(
        n9509) );
  XNOR2_X2 U10577 ( .A(n9610), .B(n9611), .ZN(n9513) );
  NAND2_X2 U10578 ( .A1(net71078), .A2(WIRE_ALU_A_MUX2TO1_32BIT_8__MUX_N1), 
        .ZN(n9512) );
  NOR2_X4 U10579 ( .A1(n9515), .A2(n9514), .ZN(n9519) );
  OAI22_X2 U10581 ( .A1(n5977), .A2(n6091), .B1(n6156), .B2(n6049), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10582 ( .A1(n6193), .A2(n5376), .B1(n6195), .B2(n6049), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  INV_X4 U10583 ( .A(REGFILE_reg_out_12__8_), .ZN(n9521) );
  OAI22_X2 U10584 ( .A1(n6196), .A2(n9521), .B1(n6199), .B2(n6049), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10585 ( .A1(n5295), .A2(n6097), .B1(n6095), .B2(n6049), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10586 ( .A1(n5178), .A2(n6103), .B1(n6102), .B2(n6049), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10587 ( .A1(n5910), .A2(n6108), .B1(n6106), .B2(n6049), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10588 ( .A1(n5179), .A2(n6112), .B1(n6158), .B2(n6048), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10589 ( .A1(n5180), .A2(n6115), .B1(n6160), .B2(n4801), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10590 ( .A1(n5296), .A2(n6118), .B1(n6162), .B2(n6048), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10591 ( .A1(n6200), .A2(n5377), .B1(n6204), .B2(n6049), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10592 ( .A1(n5297), .A2(net76862), .B1(net76616), .B2(n4801), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10593 ( .A1(n6206), .A2(n5413), .B1(n6208), .B2(n6049), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10594 ( .A1(n5181), .A2(n6121), .B1(n6164), .B2(n6048), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10595 ( .A1(n5298), .A2(n6124), .B1(n6166), .B2(n4801), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10596 ( .A1(n5182), .A2(n6127), .B1(n6168), .B2(n6049), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10597 ( .A1(n5183), .A2(n6129), .B1(n6170), .B2(n6048), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10598 ( .A1(n5869), .A2(n6132), .B1(n6172), .B2(n6048), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10599 ( .A1(n5184), .A2(n6136), .B1(n6174), .B2(n6048), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10600 ( .A1(n6210), .A2(n5978), .B1(n6212), .B2(n4801), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10601 ( .A1(REGFILE_reg_out_28__8_), .A2(n6175), .ZN(n9522) );
  NAND2_X2 U10602 ( .A1(n6178), .A2(REGFILE_reg_out_29__8_), .ZN(n9523) );
  OAI22_X2 U10603 ( .A1(n9524), .A2(n6139), .B1(net76550), .B2(n4801), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10604 ( .A1(n6180), .A2(REGFILE_reg_out_30__8_), .ZN(n9525) );
  NAND2_X2 U10605 ( .A1(n5688), .A2(REGFILE_reg_out_31__8_), .ZN(n9526) );
  OAI22_X2 U10606 ( .A1(n6216), .A2(n5028), .B1(net76320), .B2(n4801), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10607 ( .A1(n6218), .A2(n5378), .B1(n6220), .B2(n6048), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  INV_X4 U10608 ( .A(REGFILE_reg_out_5__8_), .ZN(n9527) );
  OAI22_X2 U10609 ( .A1(n9527), .A2(n6144), .B1(n6183), .B2(n6048), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10610 ( .A1(n5079), .A2(net76706), .B1(n6147), .B2(n4801), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10611 ( .A1(n5101), .A2(net76692), .B1(n6185), .B2(n4801), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10612 ( .A1(n4972), .A2(n6150), .B1(n6187), .B2(n4801), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10613 ( .A1(n5102), .A2(n6153), .B1(n6189), .B2(n6049), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  XOR2_X2 U10614 ( .A(n9530), .B(n9529), .Z(n9534) );
  NAND2_X2 U10615 ( .A1(n6190), .A2(n9531), .ZN(n9532) );
  OAI221_X2 U10616 ( .B1(n9535), .B2(n4962), .C1(n9534), .C2(n6008), .A(n9532), 
        .ZN(PCLOGIC_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10617 ( .A1(net73708), .A2(n10933), .ZN(n9541) );
  OAI211_X2 U10618 ( .C1(n8357), .C2(n9538), .A(n9537), .B(n10649), .ZN(n9540)
         );
  NAND2_X2 U10619 ( .A1(n6190), .A2(n9569), .ZN(n9539) );
  XNOR2_X2 U10620 ( .A(n9543), .B(n9542), .ZN(n9545) );
  INV_X4 U10621 ( .A(n10431), .ZN(n10343) );
  NAND2_X2 U10622 ( .A1(multOut[21]), .A2(net92392), .ZN(n9564) );
  NAND2_X2 U10623 ( .A1(n10102), .A2(n9546), .ZN(n9551) );
  NAND2_X2 U10624 ( .A1(net77086), .A2(n9547), .ZN(n9550) );
  AOI22_X2 U10625 ( .A1(n6082), .A2(n9548), .B1(n6083), .B2(n10233), .ZN(n9549) );
  NAND2_X2 U10626 ( .A1(n10058), .A2(n10059), .ZN(n9554) );
  NAND2_X2 U10627 ( .A1(n10060), .A2(n9552), .ZN(n9553) );
  NAND2_X2 U10628 ( .A1(n9554), .A2(n9553), .ZN(n9562) );
  NAND2_X2 U10629 ( .A1(n10064), .A2(n9982), .ZN(n9556) );
  NAND2_X2 U10630 ( .A1(n10066), .A2(n10063), .ZN(n9555) );
  NAND2_X2 U10631 ( .A1(n9556), .A2(n9555), .ZN(n9557) );
  MUX2_X2 U10632 ( .A(n9558), .B(n9557), .S(net71026), .Z(n9561) );
  NAND3_X2 U10633 ( .A1(n9565), .A2(n9564), .A3(n9563), .ZN(dmem_addr_out[21])
         );
  INV_X4 U10634 ( .A(dmem_addr_out[21]), .ZN(n9572) );
  INV_X4 U10635 ( .A(dmem_read_in[5]), .ZN(n9817) );
  INV_X4 U10636 ( .A(dmem_read_in[21]), .ZN(n9567) );
  OAI211_X2 U10637 ( .C1(n9572), .C2(net76646), .A(n9571), .B(n9570), .ZN(
        n9573) );
  OAI22_X2 U10638 ( .A1(n5185), .A2(n6089), .B1(net76658), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  INV_X4 U10639 ( .A(REGFILE_reg_out_10__21_), .ZN(n9574) );
  OAI22_X2 U10640 ( .A1(n9574), .A2(n6092), .B1(n6155), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10641 ( .A1(n6192), .A2(n5379), .B1(n6195), .B2(n9579), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10642 ( .A1(n6196), .A2(n5810), .B1(n6199), .B2(n9579), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10643 ( .A1(n5299), .A2(n6098), .B1(n6095), .B2(n9579), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10644 ( .A1(n5186), .A2(n6104), .B1(n6102), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10645 ( .A1(n5300), .A2(n6109), .B1(n6106), .B2(n9579), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10646 ( .A1(n5187), .A2(n6113), .B1(n6157), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10647 ( .A1(n5188), .A2(n6116), .B1(n6159), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10648 ( .A1(n5301), .A2(n6119), .B1(n6161), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10649 ( .A1(n6200), .A2(n5380), .B1(n6204), .B2(n9579), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10650 ( .A1(n5302), .A2(net76864), .B1(net76614), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10651 ( .A1(n6205), .A2(n5505), .B1(n6208), .B2(n9579), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10652 ( .A1(n5189), .A2(n6122), .B1(n6163), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10653 ( .A1(n5303), .A2(n6125), .B1(n6165), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10654 ( .A1(n5190), .A2(n6128), .B1(n6167), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10655 ( .A1(n5191), .A2(n6130), .B1(n6169), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10656 ( .A1(n5807), .A2(n6133), .B1(n6171), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10657 ( .A1(n5192), .A2(n6137), .B1(n6173), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10658 ( .A1(n6209), .A2(n5034), .B1(n6212), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10659 ( .A1(REGFILE_reg_out_28__21_), .A2(n6175), .ZN(n9575) );
  OAI21_X4 U10660 ( .B1(n6213), .B2(n6051), .A(n9575), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10661 ( .A1(n6178), .A2(REGFILE_reg_out_29__21_), .ZN(n9576) );
  OAI21_X4 U10662 ( .B1(n6138), .B2(n6051), .A(n9576), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10663 ( .A1(n5304), .A2(n6140), .B1(net76548), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10664 ( .A1(n6180), .A2(REGFILE_reg_out_30__21_), .ZN(n9577) );
  OAI21_X4 U10665 ( .B1(n6142), .B2(n6051), .A(n9577), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10666 ( .A1(n5688), .A2(REGFILE_reg_out_31__21_), .ZN(n9578) );
  OAI21_X4 U10667 ( .B1(net76480), .B2(n6051), .A(n9578), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10668 ( .A1(n6215), .A2(n5414), .B1(net76320), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10669 ( .A1(n6217), .A2(n5499), .B1(n6220), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10670 ( .A1(n5305), .A2(n6145), .B1(n6182), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10671 ( .A1(n5306), .A2(net76708), .B1(n6147), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10672 ( .A1(n5193), .A2(net76694), .B1(n6184), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10673 ( .A1(n5307), .A2(n6151), .B1(n6186), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10674 ( .A1(n5194), .A2(n6154), .B1(n6188), .B2(n6051), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10675 ( .A1(net77086), .A2(n9844), .ZN(n9584) );
  NAND2_X2 U10676 ( .A1(n6082), .A2(net70727), .ZN(n9583) );
  INV_X4 U10677 ( .A(n9934), .ZN(n9590) );
  NAND2_X2 U10678 ( .A1(n8759), .A2(n9935), .ZN(n9588) );
  NAND2_X2 U10679 ( .A1(n6082), .A2(n10091), .ZN(n9587) );
  INV_X4 U10680 ( .A(n9655), .ZN(n9589) );
  OAI22_X2 U10681 ( .A1(n10474), .A2(n9590), .B1(n10472), .B2(n9589), .ZN(
        n9592) );
  NAND2_X2 U10682 ( .A1(n10931), .A2(net70720), .ZN(n9596) );
  NAND2_X2 U10683 ( .A1(net70719), .A2(net80189), .ZN(n9595) );
  NAND4_X2 U10684 ( .A1(n9596), .A2(n9595), .A3(n9594), .A4(n9593), .ZN(n10023) );
  NAND2_X2 U10685 ( .A1(n10102), .A2(n10023), .ZN(n9604) );
  NAND2_X2 U10686 ( .A1(n10933), .A2(net70720), .ZN(n9600) );
  NAND4_X2 U10687 ( .A1(n9600), .A2(n9599), .A3(n9598), .A4(n9597), .ZN(n10158) );
  NAND2_X2 U10688 ( .A1(net77086), .A2(n10158), .ZN(n9603) );
  NAND2_X2 U10689 ( .A1(n6083), .A2(n9839), .ZN(n9602) );
  NAND2_X2 U10690 ( .A1(n6082), .A2(n10024), .ZN(n9601) );
  NAND4_X2 U10691 ( .A1(n9604), .A2(n9603), .A3(n9602), .A4(n9601), .ZN(n9933)
         );
  INV_X4 U10692 ( .A(n9933), .ZN(n9605) );
  NOR2_X4 U10693 ( .A1(n9608), .A2(n9607), .ZN(n9631) );
  AOI22_X2 U10695 ( .A1(n9611), .A2(n9610), .B1(
        WIRE_ALU_A_MUX2TO1_32BIT_8__MUX_N1), .B2(n9609), .ZN(n9683) );
  XNOR2_X2 U10696 ( .A(n9612), .B(n10464), .ZN(n9682) );
  INV_X4 U10697 ( .A(n9682), .ZN(n9614) );
  NAND2_X2 U10698 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_7__MUX_N1), .A2(n9612), .ZN(
        n9613) );
  AOI22_X2 U10699 ( .A1(n9663), .A2(n9664), .B1(
        WIRE_ALU_A_MUX2TO1_32BIT_6__MUX_N1), .B2(n9615), .ZN(n9959) );
  XNOR2_X2 U10700 ( .A(n9956), .B(n10396), .ZN(n9955) );
  XNOR2_X2 U10701 ( .A(n9959), .B(n9955), .ZN(n9628) );
  NAND2_X2 U10702 ( .A1(n8759), .A2(n10103), .ZN(n9625) );
  NAND2_X2 U10703 ( .A1(n10932), .A2(net70720), .ZN(n9620) );
  NAND4_X2 U10704 ( .A1(n9620), .A2(n9619), .A3(n9618), .A4(n9617), .ZN(n10101) );
  NAND2_X2 U10705 ( .A1(net77086), .A2(n10101), .ZN(n9624) );
  NAND2_X2 U10706 ( .A1(n4880), .A2(n9621), .ZN(n9623) );
  NAND2_X2 U10707 ( .A1(n6082), .A2(n9945), .ZN(n9622) );
  NAND4_X2 U10708 ( .A1(n9625), .A2(n9624), .A3(n9623), .A4(n9622), .ZN(n9658)
         );
  INV_X4 U10709 ( .A(n9658), .ZN(n9626) );
  OAI22_X2 U10712 ( .A1(n5515), .A2(n6089), .B1(n6053), .B2(net76658), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10713 ( .A1(n5043), .A2(n6092), .B1(n6054), .B2(n6155), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10716 ( .A1(n6196), .A2(n5660), .B1(n6054), .B2(n6199), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10717 ( .A1(n5308), .A2(n6098), .B1(n6054), .B2(n6095), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10720 ( .A1(n5309), .A2(n6109), .B1(n6054), .B2(n6106), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10722 ( .A1(n5196), .A2(n6116), .B1(n6054), .B2(n6159), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10723 ( .A1(n5310), .A2(n6119), .B1(n6054), .B2(n6161), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10724 ( .A1(n6200), .A2(n5381), .B1(n6054), .B2(n6204), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10725 ( .A1(n5311), .A2(net76864), .B1(n6054), .B2(net76614), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10726 ( .A1(n6205), .A2(n5415), .B1(n6054), .B2(n6208), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10727 ( .A1(n5197), .A2(n6122), .B1(n6054), .B2(n6163), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10728 ( .A1(n5312), .A2(n6125), .B1(n6054), .B2(n6165), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10729 ( .A1(n5198), .A2(n6128), .B1(n6054), .B2(n6167), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10732 ( .A1(n5313), .A2(n6133), .B1(n6053), .B2(n6171), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10734 ( .A1(n9641), .A2(n6137), .B1(n6053), .B2(n6173), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10735 ( .A1(n6210), .A2(n5416), .B1(n6053), .B2(n6212), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10736 ( .A1(REGFILE_reg_out_28__5_), .A2(n6175), .ZN(n9642) );
  NAND2_X2 U10737 ( .A1(n6178), .A2(REGFILE_reg_out_29__5_), .ZN(n9643) );
  OAI22_X2 U10738 ( .A1(n4984), .A2(n6140), .B1(n6053), .B2(net76548), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10739 ( .A1(n6180), .A2(REGFILE_reg_out_30__5_), .ZN(n9644) );
  NAND2_X2 U10740 ( .A1(n5688), .A2(REGFILE_reg_out_31__5_), .ZN(n9645) );
  OAI22_X2 U10741 ( .A1(n6216), .A2(n4985), .B1(n6053), .B2(net76320), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10742 ( .A1(n6217), .A2(n5554), .B1(n6053), .B2(n6220), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10743 ( .A1(n5044), .A2(n6145), .B1(n6053), .B2(n6182), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10744 ( .A1(n5451), .A2(net76708), .B1(n6053), .B2(n6147), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10745 ( .A1(n5516), .A2(net76694), .B1(n6053), .B2(n6184), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10746 ( .A1(n5314), .A2(n6151), .B1(n6053), .B2(n6186), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10747 ( .A1(n5199), .A2(n6154), .B1(n6054), .B2(n6188), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10748 ( .A1(n10102), .A2(n9844), .ZN(n9650) );
  NAND2_X2 U10749 ( .A1(n4880), .A2(net70727), .ZN(n9649) );
  NAND2_X2 U10750 ( .A1(net77086), .A2(n9845), .ZN(n9648) );
  NAND2_X2 U10751 ( .A1(n6082), .A2(n10013), .ZN(n9647) );
  NAND4_X2 U10752 ( .A1(n9650), .A2(n9649), .A3(n9648), .A4(n9647), .ZN(n9687)
         );
  NAND2_X2 U10753 ( .A1(n8759), .A2(n10024), .ZN(n9654) );
  NAND2_X2 U10754 ( .A1(net77086), .A2(n10023), .ZN(n9653) );
  NAND2_X2 U10755 ( .A1(n6083), .A2(n9838), .ZN(n9652) );
  NAND2_X2 U10756 ( .A1(n6082), .A2(n9839), .ZN(n9651) );
  NAND4_X2 U10757 ( .A1(n9654), .A2(n9653), .A3(n9652), .A4(n9651), .ZN(n9686)
         );
  AOI22_X2 U10758 ( .A1(net71092), .A2(n9687), .B1(net71094), .B2(n9686), .ZN(
        n9661) );
  NAND2_X2 U10759 ( .A1(n10280), .A2(n9655), .ZN(n9660) );
  INV_X4 U10760 ( .A(n9657), .ZN(n10394) );
  AOI21_X4 U10761 ( .B1(net71085), .B2(n9658), .A(n5052), .ZN(n9659) );
  NAND3_X2 U10762 ( .A1(n9661), .A2(n9660), .A3(n9659), .ZN(n9662) );
  XNOR2_X2 U10763 ( .A(n9664), .B(n9663), .ZN(n9666) );
  NAND2_X2 U10764 ( .A1(net71078), .A2(WIRE_ALU_A_MUX2TO1_32BIT_6__MUX_N1), 
        .ZN(n9665) );
  NOR2_X4 U10765 ( .A1(n9668), .A2(n9667), .ZN(n9673) );
  OAI22_X2 U10766 ( .A1(n5437), .A2(n6089), .B1(n4802), .B2(net76658), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10768 ( .A1(n9675), .A2(n6092), .B1(n4802), .B2(n6155), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10769 ( .A1(n6193), .A2(n5382), .B1(n4802), .B2(n6194), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10770 ( .A1(n6197), .A2(n5417), .B1(n6057), .B2(n6198), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10771 ( .A1(n5315), .A2(n6098), .B1(n6056), .B2(n6095), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10772 ( .A1(n5200), .A2(n6104), .B1(n6102), .B2(n6057), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10773 ( .A1(n4982), .A2(n6109), .B1(n6057), .B2(n6106), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10774 ( .A1(n5517), .A2(n6113), .B1(n6057), .B2(n6157), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10775 ( .A1(n5201), .A2(n6116), .B1(n6057), .B2(n6159), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10776 ( .A1(n5316), .A2(n6119), .B1(n6056), .B2(n6161), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10777 ( .A1(n6201), .A2(n5383), .B1(n6056), .B2(n6203), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10778 ( .A1(n5317), .A2(net76864), .B1(n4802), .B2(net76614), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10779 ( .A1(n6206), .A2(n5418), .B1(n4802), .B2(n6207), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10780 ( .A1(n5202), .A2(n6122), .B1(n6057), .B2(n6163), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10781 ( .A1(n5318), .A2(n6125), .B1(n6056), .B2(n6165), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10782 ( .A1(n5203), .A2(n6128), .B1(n6056), .B2(n6167), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10783 ( .A1(n5204), .A2(n6130), .B1(n6057), .B2(n6169), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  INV_X4 U10784 ( .A(n5764), .ZN(n9676) );
  OAI22_X2 U10785 ( .A1(n9676), .A2(n6133), .B1(n6056), .B2(n6171), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10786 ( .A1(n5103), .A2(n6137), .B1(n6056), .B2(n6173), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10787 ( .A1(n6210), .A2(n5113), .B1(n4802), .B2(n6211), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10788 ( .A1(REGFILE_reg_out_28__6_), .A2(n6175), .ZN(n9677) );
  NAND2_X2 U10789 ( .A1(n6178), .A2(REGFILE_reg_out_29__6_), .ZN(n9678) );
  OAI22_X2 U10790 ( .A1(n5319), .A2(n6140), .B1(n4802), .B2(net76548), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10791 ( .A1(n6180), .A2(REGFILE_reg_out_30__6_), .ZN(n9679) );
  NAND2_X2 U10792 ( .A1(n5688), .A2(REGFILE_reg_out_31__6_), .ZN(n9680) );
  OAI22_X2 U10793 ( .A1(n6216), .A2(n5419), .B1(n6056), .B2(net76318), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10794 ( .A1(n6218), .A2(n5384), .B1(n6057), .B2(n6219), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10795 ( .A1(n5320), .A2(n6145), .B1(n6057), .B2(n6182), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10796 ( .A1(n5321), .A2(net76708), .B1(n4802), .B2(n6147), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10797 ( .A1(n5205), .A2(net76694), .B1(n6056), .B2(n6184), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10798 ( .A1(n5322), .A2(n6151), .B1(n4802), .B2(n6186), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10799 ( .A1(n5206), .A2(n6154), .B1(n6057), .B2(n6188), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U10801 ( .A(n9683), .B(n9682), .ZN(n9684) );
  NAND2_X2 U10802 ( .A1(net71271), .A2(n9684), .ZN(n9697) );
  INV_X4 U10803 ( .A(n10391), .ZN(n10307) );
  NAND2_X2 U10804 ( .A1(n10066), .A2(n9686), .ZN(n9689) );
  NAND2_X2 U10805 ( .A1(n10058), .A2(n9687), .ZN(n9688) );
  NAND2_X2 U10806 ( .A1(n9689), .A2(n9688), .ZN(n9694) );
  INV_X4 U10807 ( .A(n9690), .ZN(n9692) );
  NAND2_X2 U10808 ( .A1(n6060), .A2(n4992), .ZN(n9706) );
  NAND2_X2 U10809 ( .A1(n4867), .A2(REGFILE_reg_out_0__7_), .ZN(n9705) );
  NAND2_X2 U10810 ( .A1(n9706), .A2(n9705), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10811 ( .A1(n6060), .A2(n4990), .ZN(n9708) );
  NAND2_X2 U10812 ( .A1(n9708), .A2(n9707), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10813 ( .A1(n6059), .A2(n4998), .ZN(n9710) );
  NAND2_X2 U10814 ( .A1(REGFILE_reg_out_11__7_), .A2(n4869), .ZN(n9709) );
  NAND2_X2 U10815 ( .A1(n9710), .A2(n9709), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10816 ( .A1(n6060), .A2(n4993), .ZN(n9712) );
  NAND2_X2 U10817 ( .A1(REGFILE_reg_out_12__7_), .A2(n4873), .ZN(n9711) );
  NAND2_X2 U10818 ( .A1(n9712), .A2(n9711), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10819 ( .A1(n6060), .A2(n6096), .ZN(n9714) );
  NAND2_X2 U10820 ( .A1(n6100), .A2(REGFILE_reg_out_13__7_), .ZN(n9713) );
  NAND2_X2 U10821 ( .A1(n9714), .A2(n9713), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10822 ( .A1(n9765), .A2(n6101), .ZN(n9716) );
  NAND2_X2 U10823 ( .A1(n4805), .A2(REGFILE_reg_out_14__7_), .ZN(n9715) );
  NAND2_X2 U10824 ( .A1(n9716), .A2(n9715), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10825 ( .A1(n6059), .A2(n6107), .ZN(n9718) );
  NAND2_X2 U10826 ( .A1(n4804), .A2(REGFILE_reg_out_15__7_), .ZN(n9717) );
  NAND2_X2 U10827 ( .A1(n9718), .A2(n9717), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10828 ( .A1(n6060), .A2(n4994), .ZN(n9720) );
  NAND2_X2 U10829 ( .A1(n4891), .A2(REGFILE_reg_out_16__7_), .ZN(n9719) );
  NAND2_X2 U10830 ( .A1(n9720), .A2(n9719), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10831 ( .A1(n6060), .A2(n4999), .ZN(n9722) );
  NAND2_X2 U10832 ( .A1(n4892), .A2(REGFILE_reg_out_17__7_), .ZN(n9721) );
  NAND2_X2 U10833 ( .A1(n9722), .A2(n9721), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10834 ( .A1(n6060), .A2(n5000), .ZN(n9724) );
  NAND2_X2 U10835 ( .A1(n4884), .A2(REGFILE_reg_out_18__7_), .ZN(n9723) );
  NAND2_X2 U10836 ( .A1(n9724), .A2(n9723), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10837 ( .A1(n6060), .A2(n5001), .ZN(n9726) );
  NAND2_X2 U10838 ( .A1(REGFILE_reg_out_19__7_), .A2(n4876), .ZN(n9725) );
  NAND2_X2 U10839 ( .A1(n9726), .A2(n9725), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10840 ( .A1(n6060), .A2(n4997), .ZN(n9728) );
  NAND2_X2 U10841 ( .A1(n4877), .A2(REGFILE_reg_out_1__7_), .ZN(n9727) );
  NAND2_X2 U10842 ( .A1(n9728), .A2(n9727), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10843 ( .A1(n6060), .A2(n4903), .ZN(n9730) );
  NAND2_X2 U10844 ( .A1(REGFILE_reg_out_20__7_), .A2(n4868), .ZN(n9729) );
  NAND2_X2 U10845 ( .A1(n9730), .A2(n9729), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10846 ( .A1(n6060), .A2(n4904), .ZN(n9732) );
  NAND2_X2 U10847 ( .A1(n4882), .A2(REGFILE_reg_out_21__7_), .ZN(n9731) );
  NAND2_X2 U10848 ( .A1(n9732), .A2(n9731), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10849 ( .A1(n6060), .A2(n4905), .ZN(n9734) );
  NAND2_X2 U10850 ( .A1(n4888), .A2(REGFILE_reg_out_22__7_), .ZN(n9733) );
  NAND2_X2 U10851 ( .A1(n9734), .A2(n9733), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10852 ( .A1(n6060), .A2(n4906), .ZN(n9736) );
  NAND2_X2 U10853 ( .A1(n4883), .A2(REGFILE_reg_out_23__7_), .ZN(n9735) );
  NAND2_X2 U10854 ( .A1(n9736), .A2(n9735), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10855 ( .A1(n6060), .A2(n4995), .ZN(n9738) );
  NAND2_X2 U10856 ( .A1(n4875), .A2(REGFILE_reg_out_24__7_), .ZN(n9737) );
  NAND2_X2 U10857 ( .A1(n9738), .A2(n9737), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10858 ( .A1(n6060), .A2(n5002), .ZN(n9740) );
  NAND2_X2 U10859 ( .A1(n9740), .A2(n9739), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10860 ( .A1(n6060), .A2(n5003), .ZN(n9742) );
  NAND2_X2 U10861 ( .A1(n4893), .A2(REGFILE_reg_out_26__7_), .ZN(n9741) );
  NAND2_X2 U10862 ( .A1(n9742), .A2(n9741), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10863 ( .A1(n6060), .A2(n5004), .ZN(n9744) );
  NAND2_X2 U10864 ( .A1(n9744), .A2(n9743), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10865 ( .A1(n6060), .A2(n4806), .ZN(n9746) );
  NAND2_X2 U10866 ( .A1(REGFILE_reg_out_28__7_), .A2(n10604), .ZN(n9745) );
  NAND2_X2 U10867 ( .A1(n9746), .A2(n9745), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10868 ( .A1(n6059), .A2(n10607), .ZN(n9748) );
  NAND2_X2 U10869 ( .A1(n6178), .A2(REGFILE_reg_out_29__7_), .ZN(n9747) );
  NAND2_X2 U10870 ( .A1(n9748), .A2(n9747), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10871 ( .A1(n6059), .A2(n5005), .ZN(n9750) );
  NAND2_X2 U10872 ( .A1(n9750), .A2(n9749), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10873 ( .A1(n6059), .A2(n10614), .ZN(n9752) );
  NAND2_X2 U10874 ( .A1(n6180), .A2(REGFILE_reg_out_30__7_), .ZN(n9751) );
  NAND2_X2 U10875 ( .A1(n9752), .A2(n9751), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10876 ( .A1(n6059), .A2(net70574), .ZN(n9754) );
  NAND2_X2 U10877 ( .A1(n5688), .A2(REGFILE_reg_out_31__7_), .ZN(n9753) );
  NAND2_X2 U10878 ( .A1(n9754), .A2(n9753), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10879 ( .A1(n6059), .A2(n5009), .ZN(n9756) );
  NAND2_X2 U10880 ( .A1(REGFILE_reg_out_3__7_), .A2(n4871), .ZN(n9755) );
  NAND2_X2 U10881 ( .A1(n9756), .A2(n9755), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10882 ( .A1(n6059), .A2(n4996), .ZN(n9758) );
  NAND2_X2 U10883 ( .A1(REGFILE_reg_out_4__7_), .A2(n4870), .ZN(n9757) );
  NAND2_X2 U10884 ( .A1(n9758), .A2(n9757), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10885 ( .A1(n6059), .A2(n5006), .ZN(n9760) );
  NAND2_X2 U10886 ( .A1(n4885), .A2(REGFILE_reg_out_5__7_), .ZN(n9759) );
  NAND2_X2 U10887 ( .A1(n9760), .A2(n9759), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10888 ( .A1(n6059), .A2(n6148), .ZN(n9761) );
  NAND2_X2 U10889 ( .A1(n9761), .A2(net71936), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10890 ( .A1(n6059), .A2(n5007), .ZN(n9762) );
  NAND2_X2 U10891 ( .A1(n9762), .A2(net71934), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10892 ( .A1(n6059), .A2(n4991), .ZN(n9764) );
  NAND2_X2 U10893 ( .A1(n4890), .A2(REGFILE_reg_out_8__7_), .ZN(n9763) );
  NAND2_X2 U10894 ( .A1(n9764), .A2(n9763), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10895 ( .A1(n6059), .A2(n5008), .ZN(n9767) );
  NAND2_X2 U10896 ( .A1(n4887), .A2(REGFILE_reg_out_9__7_), .ZN(n9766) );
  NAND2_X2 U10897 ( .A1(n9767), .A2(n9766), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10898 ( .A1(multOut[26]), .A2(net92392), .ZN(n9787) );
  OAI22_X2 U10899 ( .A1(n9768), .A2(n10472), .B1(n5061), .B2(n10474), .ZN(
        n9773) );
  INV_X4 U10900 ( .A(n9774), .ZN(n9775) );
  NOR2_X4 U10901 ( .A1(n9775), .A2(net70691), .ZN(n9784) );
  INV_X4 U10902 ( .A(n9776), .ZN(n9779) );
  INV_X4 U10903 ( .A(n9777), .ZN(n9778) );
  NAND2_X2 U10904 ( .A1(n9779), .A2(n9778), .ZN(n9783) );
  INV_X4 U10905 ( .A(n10444), .ZN(n10325) );
  NAND2_X2 U10906 ( .A1(net70701), .A2(n10325), .ZN(n9781) );
  NAND2_X2 U10907 ( .A1(n9781), .A2(n9780), .ZN(n9782) );
  NAND3_X2 U10908 ( .A1(n9787), .A2(n9786), .A3(n9785), .ZN(dmem_addr_out[26])
         );
  INV_X4 U10909 ( .A(dmem_addr_out[26]), .ZN(n9794) );
  INV_X4 U10910 ( .A(dmem_read_in[10]), .ZN(n10137) );
  INV_X4 U10911 ( .A(dmem_read_in[26]), .ZN(n9789) );
  OAI211_X2 U10912 ( .C1(n9794), .C2(net76646), .A(n9793), .B(n9792), .ZN(
        n9795) );
  NAND2_X2 U10913 ( .A1(net76270), .A2(n9795), .ZN(n9800) );
  OAI22_X2 U10914 ( .A1(n5518), .A2(n6089), .B1(net76658), .B2(n6062), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10915 ( .A1(n5452), .A2(n6092), .B1(n6155), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10916 ( .A1(n6193), .A2(n5555), .B1(n6194), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10917 ( .A1(n6197), .A2(n5503), .B1(n6198), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10918 ( .A1(n5323), .A2(n6098), .B1(n6095), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10919 ( .A1(n5207), .A2(n6104), .B1(n6102), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10920 ( .A1(n5324), .A2(n6109), .B1(n6106), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10921 ( .A1(n5208), .A2(n6113), .B1(n6157), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10922 ( .A1(n5519), .A2(n6116), .B1(n6159), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10923 ( .A1(n5453), .A2(n6119), .B1(n6161), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10924 ( .A1(n6201), .A2(n5385), .B1(n6203), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10925 ( .A1(n5325), .A2(net76864), .B1(net76614), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10926 ( .A1(n6206), .A2(n5420), .B1(n6207), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10927 ( .A1(n5209), .A2(n6122), .B1(n6163), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10928 ( .A1(n5326), .A2(n6125), .B1(n6165), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10929 ( .A1(n5210), .A2(n6128), .B1(n6167), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10930 ( .A1(n5211), .A2(n6130), .B1(n6169), .B2(n6062), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10931 ( .A1(n5327), .A2(n6133), .B1(n6171), .B2(n6062), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10932 ( .A1(n5212), .A2(n6137), .B1(n6173), .B2(n6062), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10933 ( .A1(n6210), .A2(n5421), .B1(n6211), .B2(n6062), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10934 ( .A1(REGFILE_reg_out_28__26_), .A2(n6175), .ZN(n9796) );
  OAI21_X4 U10935 ( .B1(n6214), .B2(n6062), .A(n9796), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10936 ( .A1(n6178), .A2(REGFILE_reg_out_29__26_), .ZN(n9797) );
  OAI21_X4 U10937 ( .B1(n10532), .B2(n6062), .A(n9797), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10938 ( .A1(n5454), .A2(n6140), .B1(net76548), .B2(n6062), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10939 ( .A1(n6180), .A2(REGFILE_reg_out_30__26_), .ZN(n9798) );
  OAI21_X4 U10940 ( .B1(n10534), .B2(n6062), .A(n9798), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10941 ( .A1(n5688), .A2(REGFILE_reg_out_31__26_), .ZN(n9799) );
  OAI21_X4 U10942 ( .B1(net70509), .B2(n6062), .A(n9799), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10943 ( .A1(n6216), .A2(n5422), .B1(net76318), .B2(n6062), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10944 ( .A1(n6218), .A2(n5556), .B1(n6219), .B2(n6062), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10945 ( .A1(n5455), .A2(n6145), .B1(n6182), .B2(n6062), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10946 ( .A1(n5456), .A2(net76708), .B1(n6147), .B2(n6062), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10947 ( .A1(n5520), .A2(net76694), .B1(n6184), .B2(n6062), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10948 ( .A1(n5457), .A2(n6151), .B1(n6186), .B2(n6062), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10949 ( .A1(n5521), .A2(n6154), .B1(n6188), .B2(n6063), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10950 ( .A1(n4922), .A2(n9802), .B1(n9801), .B2(n10472), .ZN(n9808) );
  OAI22_X2 U10951 ( .A1(net70710), .A2(n9805), .B1(n9804), .B2(n9803), .ZN(
        n9807) );
  AOI211_X4 U10952 ( .C1(n9808), .C2(net70697), .A(n9807), .B(n9806), .ZN(
        n9815) );
  NAND2_X2 U10953 ( .A1(multOut[29]), .A2(net92392), .ZN(n9814) );
  XNOR2_X2 U10954 ( .A(n9810), .B(n9809), .ZN(n9812) );
  INV_X4 U10955 ( .A(dmem_addr_out[29]), .ZN(n9825) );
  INV_X4 U10956 ( .A(dmem_read_in[29]), .ZN(n9820) );
  OAI211_X2 U10957 ( .C1(n9825), .C2(net76646), .A(n9824), .B(n9823), .ZN(
        n9826) );
  OAI22_X2 U10958 ( .A1(n5522), .A2(n6089), .B1(n6222), .B2(net76658), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10959 ( .A1(n5458), .A2(n6092), .B1(n6222), .B2(n6155), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10960 ( .A1(n5328), .A2(n6098), .B1(n6222), .B2(n6094), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  INV_X4 U10961 ( .A(REGFILE_reg_out_14__29_), .ZN(n9827) );
  OAI22_X2 U10962 ( .A1(n9827), .A2(n6104), .B1(n6222), .B2(n6102), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10963 ( .A1(n9828), .A2(n6109), .B1(n6222), .B2(n6105), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10964 ( .A1(n5213), .A2(n6113), .B1(n6222), .B2(n6157), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10965 ( .A1(n5126), .A2(n6116), .B1(n6222), .B2(n6159), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10966 ( .A1(n5459), .A2(n6119), .B1(n6222), .B2(n6161), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10967 ( .A1(n4977), .A2(net76864), .B1(n6222), .B2(net76614), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10968 ( .A1(n4988), .A2(n6122), .B1(n6222), .B2(n6163), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10969 ( .A1(n5460), .A2(n6125), .B1(n6222), .B2(n6165), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10970 ( .A1(net71824), .A2(n6128), .B1(n6222), .B2(n6167), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10971 ( .A1(n5123), .A2(n6130), .B1(n6222), .B2(n6169), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10972 ( .A1(n4974), .A2(n6133), .B1(n6222), .B2(n6171), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10973 ( .A1(n5214), .A2(n6137), .B1(n6222), .B2(n6173), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10974 ( .A1(n6178), .A2(REGFILE_reg_out_29__29_), .ZN(n9829) );
  OAI22_X2 U10975 ( .A1(n5461), .A2(n6140), .B1(n6222), .B2(net76548), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10976 ( .A1(n6180), .A2(REGFILE_reg_out_30__29_), .ZN(n9830) );
  OAI22_X2 U10977 ( .A1(n5125), .A2(n6145), .B1(n6222), .B2(n6182), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10978 ( .A1(n5462), .A2(net76708), .B1(n6222), .B2(n6146), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10979 ( .A1(n5523), .A2(net76694), .B1(n6222), .B2(n6184), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10980 ( .A1(n5463), .A2(n6151), .B1(n6222), .B2(n6186), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10981 ( .A1(n5987), .A2(n6154), .B1(n6222), .B2(n6188), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U10982 ( .A1(multOut[11]), .A2(net92392), .ZN(n9861) );
  XNOR2_X2 U10983 ( .A(n9833), .B(n9832), .ZN(n9834) );
  NAND2_X2 U10984 ( .A1(net71271), .A2(n9834), .ZN(n9860) );
  NAND2_X2 U10985 ( .A1(n8759), .A2(n9838), .ZN(n9843) );
  NAND2_X2 U10986 ( .A1(net105360), .A2(n9839), .ZN(n9842) );
  NAND2_X2 U10987 ( .A1(n6083), .A2(n10238), .ZN(n9841) );
  NAND2_X2 U10988 ( .A1(n6082), .A2(n10239), .ZN(n9840) );
  NAND4_X2 U10989 ( .A1(n9843), .A2(n9842), .A3(n9841), .A4(n9840), .ZN(n10122) );
  NAND2_X2 U10990 ( .A1(n10066), .A2(n10122), .ZN(n9851) );
  NAND2_X2 U10991 ( .A1(n8759), .A2(n10231), .ZN(n9849) );
  NAND2_X2 U10992 ( .A1(n6083), .A2(n9844), .ZN(n9848) );
  NAND2_X2 U10993 ( .A1(net105360), .A2(n10230), .ZN(n9847) );
  NAND2_X2 U10994 ( .A1(n6082), .A2(n9845), .ZN(n9846) );
  NAND4_X2 U10995 ( .A1(n9849), .A2(n9848), .A3(n9847), .A4(n9846), .ZN(n10123) );
  NAND2_X2 U10996 ( .A1(n10058), .A2(n10123), .ZN(n9850) );
  NAND2_X2 U10997 ( .A1(n9851), .A2(n9850), .ZN(n9857) );
  INV_X4 U10998 ( .A(n9852), .ZN(n9855) );
  NAND4_X2 U10999 ( .A1(n9861), .A2(n9860), .A3(n9859), .A4(n9858), .ZN(
        dmem_addr_out[11]) );
  NAND2_X2 U11000 ( .A1(net76650), .A2(dmem_addr_out[11]), .ZN(n9866) );
  NAND3_X2 U11001 ( .A1(n9866), .A2(net70740), .A3(n9865), .ZN(n9867) );
  NAND2_X2 U11002 ( .A1(n6066), .A2(n4992), .ZN(n9870) );
  NAND2_X2 U11003 ( .A1(n4867), .A2(REGFILE_reg_out_0__11_), .ZN(n9869) );
  NAND2_X2 U11004 ( .A1(n9870), .A2(n9869), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11005 ( .A1(n6066), .A2(n4990), .ZN(n9872) );
  NAND2_X2 U11006 ( .A1(n6093), .A2(n5907), .ZN(n9871) );
  NAND2_X2 U11007 ( .A1(n9872), .A2(n9871), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11008 ( .A1(n6066), .A2(n4998), .ZN(n9874) );
  NAND2_X2 U11009 ( .A1(REGFILE_reg_out_11__11_), .A2(n4869), .ZN(n9873) );
  NAND2_X2 U11010 ( .A1(n9874), .A2(n9873), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11011 ( .A1(n6066), .A2(n4993), .ZN(n9876) );
  NAND2_X2 U11012 ( .A1(n9876), .A2(n9875), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11013 ( .A1(n6066), .A2(n6096), .ZN(n9878) );
  NAND2_X2 U11014 ( .A1(n9878), .A2(n9877), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11015 ( .A1(n6066), .A2(n6101), .ZN(n9880) );
  NAND2_X2 U11016 ( .A1(n4805), .A2(REGFILE_reg_out_14__11_), .ZN(n9879) );
  NAND2_X2 U11017 ( .A1(n9880), .A2(n9879), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11018 ( .A1(n6066), .A2(n6107), .ZN(n9882) );
  NAND2_X2 U11019 ( .A1(n4804), .A2(REGFILE_reg_out_15__11_), .ZN(n9881) );
  NAND2_X2 U11020 ( .A1(n9882), .A2(n9881), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11021 ( .A1(n6066), .A2(n4994), .ZN(n9884) );
  NAND2_X2 U11022 ( .A1(n4891), .A2(REGFILE_reg_out_16__11_), .ZN(n9883) );
  NAND2_X2 U11023 ( .A1(n9884), .A2(n9883), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11024 ( .A1(n6066), .A2(n4999), .ZN(n9886) );
  NAND2_X2 U11025 ( .A1(n4892), .A2(REGFILE_reg_out_17__11_), .ZN(n9885) );
  NAND2_X2 U11026 ( .A1(n9886), .A2(n9885), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11027 ( .A1(n6066), .A2(n5000), .ZN(n9888) );
  NAND2_X2 U11028 ( .A1(n4884), .A2(REGFILE_reg_out_18__11_), .ZN(n9887) );
  NAND2_X2 U11029 ( .A1(n9888), .A2(n9887), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11030 ( .A1(n6065), .A2(n5001), .ZN(n9890) );
  NAND2_X2 U11031 ( .A1(REGFILE_reg_out_19__11_), .A2(n4876), .ZN(n9889) );
  NAND2_X2 U11032 ( .A1(n9890), .A2(n9889), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11033 ( .A1(n6065), .A2(n4997), .ZN(n9892) );
  NAND2_X2 U11034 ( .A1(n4877), .A2(REGFILE_reg_out_1__11_), .ZN(n9891) );
  NAND2_X2 U11035 ( .A1(n9892), .A2(n9891), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11036 ( .A1(n6065), .A2(n4903), .ZN(n9894) );
  NAND2_X2 U11037 ( .A1(REGFILE_reg_out_20__11_), .A2(n4868), .ZN(n9893) );
  NAND2_X2 U11038 ( .A1(n9894), .A2(n9893), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11039 ( .A1(n6065), .A2(n4904), .ZN(n9896) );
  NAND2_X2 U11040 ( .A1(n4882), .A2(REGFILE_reg_out_21__11_), .ZN(n9895) );
  NAND2_X2 U11041 ( .A1(n9896), .A2(n9895), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11042 ( .A1(n6065), .A2(n4905), .ZN(n9898) );
  NAND2_X2 U11043 ( .A1(n4888), .A2(REGFILE_reg_out_22__11_), .ZN(n9897) );
  NAND2_X2 U11044 ( .A1(n9898), .A2(n9897), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11045 ( .A1(n6065), .A2(n4906), .ZN(n9900) );
  NAND2_X2 U11046 ( .A1(n4883), .A2(REGFILE_reg_out_23__11_), .ZN(n9899) );
  NAND2_X2 U11047 ( .A1(n9900), .A2(n9899), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11048 ( .A1(n6065), .A2(n4995), .ZN(n9902) );
  NAND2_X2 U11049 ( .A1(n4875), .A2(REGFILE_reg_out_24__11_), .ZN(n9901) );
  NAND2_X2 U11050 ( .A1(n9902), .A2(n9901), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11051 ( .A1(n6065), .A2(n5002), .ZN(n9904) );
  NAND2_X2 U11052 ( .A1(n4878), .A2(REGFILE_reg_out_25__11_), .ZN(n9903) );
  NAND2_X2 U11053 ( .A1(n9904), .A2(n9903), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11054 ( .A1(n6065), .A2(n5003), .ZN(n9906) );
  NAND2_X2 U11055 ( .A1(n4893), .A2(REGFILE_reg_out_26__11_), .ZN(n9905) );
  NAND2_X2 U11056 ( .A1(n9906), .A2(n9905), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11057 ( .A1(n6065), .A2(n5004), .ZN(n9908) );
  NAND2_X2 U11058 ( .A1(n9908), .A2(n9907), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11059 ( .A1(n6065), .A2(n4806), .ZN(n9910) );
  NAND2_X2 U11060 ( .A1(n9910), .A2(n9909), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11061 ( .A1(n6065), .A2(n10607), .ZN(n9912) );
  NAND2_X2 U11062 ( .A1(n6178), .A2(REGFILE_reg_out_29__11_), .ZN(n9911) );
  NAND2_X2 U11063 ( .A1(n9912), .A2(n9911), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11064 ( .A1(n6065), .A2(n5005), .ZN(n9914) );
  NAND2_X2 U11065 ( .A1(n4879), .A2(REGFILE_reg_out_2__11_), .ZN(n9913) );
  NAND2_X2 U11066 ( .A1(n9914), .A2(n9913), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11067 ( .A1(n6066), .A2(n10614), .ZN(n9916) );
  NAND2_X2 U11068 ( .A1(n6180), .A2(REGFILE_reg_out_30__11_), .ZN(n9915) );
  NAND2_X2 U11069 ( .A1(n9916), .A2(n9915), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11070 ( .A1(n6065), .A2(net70574), .ZN(n9918) );
  NAND2_X2 U11071 ( .A1(n5688), .A2(REGFILE_reg_out_31__11_), .ZN(n9917) );
  NAND2_X2 U11072 ( .A1(n9918), .A2(n9917), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11073 ( .A1(n6066), .A2(n5009), .ZN(n9920) );
  NAND2_X2 U11074 ( .A1(REGFILE_reg_out_3__11_), .A2(n4871), .ZN(n9919) );
  NAND2_X2 U11075 ( .A1(n9920), .A2(n9919), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11076 ( .A1(n6066), .A2(n4996), .ZN(n9922) );
  NAND2_X2 U11077 ( .A1(REGFILE_reg_out_4__11_), .A2(n4870), .ZN(n9921) );
  NAND2_X2 U11078 ( .A1(n9922), .A2(n9921), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11079 ( .A1(n6066), .A2(n5006), .ZN(n9924) );
  NAND2_X2 U11080 ( .A1(n4885), .A2(REGFILE_reg_out_5__11_), .ZN(n9923) );
  NAND2_X2 U11081 ( .A1(n9924), .A2(n9923), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11082 ( .A1(n6066), .A2(n6148), .ZN(n9926) );
  NAND2_X2 U11083 ( .A1(n4889), .A2(REGFILE_reg_out_6__11_), .ZN(n9925) );
  NAND2_X2 U11084 ( .A1(n9926), .A2(n9925), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11085 ( .A1(n6065), .A2(n5007), .ZN(n9928) );
  NAND2_X2 U11086 ( .A1(n4886), .A2(REGFILE_reg_out_7__11_), .ZN(n9927) );
  NAND2_X2 U11087 ( .A1(n9928), .A2(n9927), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11088 ( .A1(n6065), .A2(n4991), .ZN(n9930) );
  NAND2_X2 U11089 ( .A1(n4890), .A2(REGFILE_reg_out_8__11_), .ZN(n9929) );
  NAND2_X2 U11090 ( .A1(n9930), .A2(n9929), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11091 ( .A1(n6066), .A2(n5008), .ZN(n9932) );
  NAND2_X2 U11092 ( .A1(n4887), .A2(REGFILE_reg_out_9__11_), .ZN(n9931) );
  NAND2_X2 U11093 ( .A1(n9932), .A2(n9931), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  AOI22_X2 U11094 ( .A1(net71092), .A2(n9934), .B1(net71094), .B2(n9933), .ZN(
        n9952) );
  INV_X4 U11095 ( .A(n10091), .ZN(n9937) );
  INV_X4 U11096 ( .A(n9935), .ZN(n9936) );
  NAND2_X2 U11097 ( .A1(net70696), .A2(n6005), .ZN(n10014) );
  OAI221_X2 U11098 ( .B1(n9937), .B2(n10094), .C1(n9936), .C2(net70718), .A(
        n10014), .ZN(n10017) );
  NAND2_X2 U11099 ( .A1(n10280), .A2(n10017), .ZN(n9951) );
  NAND2_X2 U11100 ( .A1(n10102), .A2(n10101), .ZN(n9949) );
  NAND2_X2 U11101 ( .A1(net70720), .A2(aluA[20]), .ZN(n9944) );
  INV_X4 U11102 ( .A(n9938), .ZN(n9941) );
  INV_X4 U11103 ( .A(n9939), .ZN(n9940) );
  NAND2_X2 U11104 ( .A1(net105360), .A2(n10541), .ZN(n9948) );
  NAND2_X2 U11105 ( .A1(n4880), .A2(n9945), .ZN(n9947) );
  NAND2_X2 U11106 ( .A1(n6082), .A2(n10103), .ZN(n9946) );
  NAND4_X2 U11107 ( .A1(n9949), .A2(n9948), .A3(n9947), .A4(n9946), .ZN(n10016) );
  INV_X4 U11108 ( .A(n10306), .ZN(n10402) );
  NAND3_X2 U11109 ( .A1(n9952), .A2(n9951), .A3(n9950), .ZN(n9953) );
  MUX2_X2 U11110 ( .A(n9953), .B(multOut[4]), .S(net76452), .Z(n9963) );
  XNOR2_X2 U11111 ( .A(n10033), .B(n9954), .ZN(n10034) );
  INV_X4 U11112 ( .A(n9955), .ZN(n9958) );
  XNOR2_X2 U11113 ( .A(n10034), .B(n10035), .ZN(n9961) );
  NAND2_X2 U11114 ( .A1(net71078), .A2(WIRE_ALU_A_MUX2TO1_32BIT_4__MUX_N1), 
        .ZN(n9960) );
  OAI22_X2 U11115 ( .A1(n5524), .A2(n6089), .B1(net76658), .B2(n4803), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11116 ( .A1(n5464), .A2(n6092), .B1(n6155), .B2(n6068), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11117 ( .A1(n6193), .A2(n5557), .B1(n6194), .B2(n4803), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11118 ( .A1(n6197), .A2(n5033), .B1(n6198), .B2(n6067), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11119 ( .A1(n5465), .A2(n6098), .B1(n6094), .B2(n6067), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11120 ( .A1(n5525), .A2(n6104), .B1(n10519), .B2(n6067), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11121 ( .A1(n5329), .A2(n6109), .B1(n6105), .B2(n6067), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11122 ( .A1(n5215), .A2(n6113), .B1(n6157), .B2(n6067), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11123 ( .A1(n5526), .A2(n6116), .B1(n6159), .B2(n6067), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11124 ( .A1(n5466), .A2(n6119), .B1(n6161), .B2(n4803), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11125 ( .A1(n6201), .A2(n5438), .B1(n6203), .B2(n6068), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11126 ( .A1(n5048), .A2(net76864), .B1(net76614), .B2(n4803), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11127 ( .A1(n6206), .A2(n5423), .B1(n6207), .B2(n4803), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11128 ( .A1(n5216), .A2(n6122), .B1(n6163), .B2(n6067), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11129 ( .A1(n5467), .A2(n6125), .B1(n6165), .B2(n6068), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11130 ( .A1(n5527), .A2(n6128), .B1(n6167), .B2(n6068), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11131 ( .A1(n5528), .A2(n6130), .B1(n6169), .B2(n6068), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11132 ( .A1(n5468), .A2(n6133), .B1(n6171), .B2(n4803), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11133 ( .A1(n5217), .A2(n6137), .B1(n6067), .B2(n6173), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11134 ( .A1(n6210), .A2(n5424), .B1(n6211), .B2(n6068), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11135 ( .A1(REGFILE_reg_out_28__4_), .A2(n10604), .ZN(n9969) );
  NAND2_X2 U11136 ( .A1(n10608), .A2(REGFILE_reg_out_29__4_), .ZN(n9970) );
  OAI22_X2 U11137 ( .A1(n5770), .A2(n6140), .B1(net76548), .B2(n6068), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11138 ( .A1(n10615), .A2(REGFILE_reg_out_30__4_), .ZN(n9971) );
  NAND2_X2 U11139 ( .A1(net76488), .A2(REGFILE_reg_out_31__4_), .ZN(n9972) );
  OAI22_X2 U11141 ( .A1(n6216), .A2(n9973), .B1(net76318), .B2(n4803), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11142 ( .A1(n6218), .A2(n5386), .B1(n6219), .B2(n6067), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11143 ( .A1(n5330), .A2(n6145), .B1(n6182), .B2(n4803), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11144 ( .A1(n5469), .A2(net76708), .B1(n6146), .B2(n6068), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11145 ( .A1(n5529), .A2(net76694), .B1(n6184), .B2(n4803), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11146 ( .A1(n5331), .A2(n6151), .B1(n6186), .B2(n6068), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11147 ( .A1(n5218), .A2(n6154), .B1(n6188), .B2(n6067), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11148 ( .A1(n8759), .A2(n9975), .ZN(n9981) );
  NAND2_X2 U11149 ( .A1(net77086), .A2(n9976), .ZN(n9980) );
  AOI22_X2 U11150 ( .A1(n6082), .A2(n9978), .B1(n6083), .B2(n9977), .ZN(n9979)
         );
  NAND2_X2 U11151 ( .A1(net71092), .A2(n10057), .ZN(n9990) );
  MUX2_X2 U11152 ( .A(n9982), .B(n10065), .S(net71026), .Z(n9983) );
  NAND2_X2 U11153 ( .A1(net71094), .A2(n9983), .ZN(n9989) );
  NAND2_X2 U11154 ( .A1(n10280), .A2(n9984), .ZN(n9988) );
  AOI21_X4 U11155 ( .B1(net71085), .B2(n9986), .A(n9985), .ZN(n9987) );
  NAND4_X2 U11156 ( .A1(n9990), .A2(n9989), .A3(n9988), .A4(n9987), .ZN(n9991)
         );
  MUX2_X2 U11157 ( .A(n9991), .B(multOut[19]), .S(net76452), .Z(n9998) );
  XNOR2_X2 U11158 ( .A(n9993), .B(n9992), .ZN(n9996) );
  NAND2_X2 U11159 ( .A1(net71078), .A2(aluA[19]), .ZN(n9994) );
  OAI22_X2 U11160 ( .A1(n9996), .A2(net70691), .B1(n9995), .B2(n9994), .ZN(
        n9997) );
  NOR2_X4 U11161 ( .A1(n9998), .A2(n9997), .ZN(n10006) );
  INV_X4 U11162 ( .A(n10006), .ZN(dmem_addr_out[19]) );
  INV_X4 U11163 ( .A(dmem_read_in[19]), .ZN(n10001) );
  OAI211_X2 U11164 ( .C1(n10006), .C2(net76646), .A(n10005), .B(n10004), .ZN(
        n10007) );
  NAND2_X2 U11165 ( .A1(net76270), .A2(n10007), .ZN(n10012) );
  OAI22_X2 U11166 ( .A1(n5219), .A2(n6089), .B1(net76658), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11167 ( .A1(n5031), .A2(n6092), .B1(n6155), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11168 ( .A1(n6193), .A2(n5387), .B1(n6194), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11169 ( .A1(n6197), .A2(n5035), .B1(n6198), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11170 ( .A1(n5332), .A2(n6098), .B1(n6094), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11171 ( .A1(n5220), .A2(n6104), .B1(n6102), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11172 ( .A1(n4978), .A2(n6109), .B1(n6105), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11173 ( .A1(n5221), .A2(n6113), .B1(n6157), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11174 ( .A1(n5222), .A2(n6116), .B1(n6159), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11175 ( .A1(n5333), .A2(n6119), .B1(n6161), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11176 ( .A1(n6201), .A2(n5118), .B1(n6203), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11177 ( .A1(n5080), .A2(net76864), .B1(net76614), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11178 ( .A1(n6206), .A2(n5425), .B1(n6207), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11179 ( .A1(n5223), .A2(n6122), .B1(n6163), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11180 ( .A1(n5334), .A2(n6125), .B1(n6165), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11181 ( .A1(n5224), .A2(n6128), .B1(n6167), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11182 ( .A1(n5104), .A2(n6130), .B1(n6169), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11183 ( .A1(n4973), .A2(n6133), .B1(n6171), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11184 ( .A1(n5225), .A2(n6137), .B1(n6173), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11185 ( .A1(n6210), .A2(n5036), .B1(n6211), .B2(n10012), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11186 ( .A1(REGFILE_reg_out_28__19_), .A2(n10604), .ZN(n10008) );
  NAND2_X2 U11187 ( .A1(n10608), .A2(REGFILE_reg_out_29__19_), .ZN(n10009) );
  OAI22_X2 U11188 ( .A1(n5651), .A2(n6140), .B1(net76548), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11189 ( .A1(n10615), .A2(REGFILE_reg_out_30__19_), .ZN(n10010) );
  NAND2_X2 U11190 ( .A1(net76488), .A2(REGFILE_reg_out_31__19_), .ZN(n10011)
         );
  OAI22_X2 U11191 ( .A1(n6216), .A2(n5426), .B1(net76318), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11192 ( .A1(n6218), .A2(n5388), .B1(n6219), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11193 ( .A1(n5335), .A2(n6145), .B1(n6182), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11194 ( .A1(n5336), .A2(net76708), .B1(n6146), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11195 ( .A1(n5226), .A2(net76694), .B1(n6184), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11196 ( .A1(n5337), .A2(n6151), .B1(n6186), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11197 ( .A1(n5227), .A2(n6154), .B1(n6188), .B2(n6070), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11198 ( .A(net70727), .ZN(net71299) );
  INV_X4 U11199 ( .A(n10013), .ZN(n10015) );
  OAI221_X2 U11200 ( .B1(net71299), .B2(n10094), .C1(n10015), .C2(net70718), 
        .A(n10014), .ZN(n10092) );
  AOI222_X2 U11201 ( .A1(n10280), .A2(n10092), .B1(net71092), .B2(n10017), 
        .C1(net71094), .C2(n10016), .ZN(n10031) );
  NAND2_X2 U11202 ( .A1(net70720), .A2(aluA[19]), .ZN(n10021) );
  NAND2_X2 U11203 ( .A1(net70719), .A2(n5761), .ZN(n10020) );
  NAND4_X2 U11204 ( .A1(n10021), .A2(n10020), .A3(n10019), .A4(n10018), .ZN(
        n10022) );
  MUX2_X2 U11205 ( .A(n10023), .B(n10022), .S(n10099), .Z(n10156) );
  INV_X4 U11206 ( .A(n10156), .ZN(n10027) );
  NAND2_X2 U11207 ( .A1(n8759), .A2(n10158), .ZN(n10026) );
  NAND2_X2 U11208 ( .A1(n6083), .A2(n10024), .ZN(n10025) );
  OAI211_X2 U11209 ( .C1(net78051), .C2(n10027), .A(n10026), .B(n10025), .ZN(
        n10028) );
  INV_X4 U11210 ( .A(n10028), .ZN(n10093) );
  INV_X4 U11211 ( .A(n10407), .ZN(n10415) );
  NOR2_X4 U11212 ( .A1(n10029), .A2(n5040), .ZN(n10030) );
  NAND2_X2 U11213 ( .A1(n10031), .A2(n10030), .ZN(n10032) );
  AOI22_X2 U11214 ( .A1(n10035), .A2(n10034), .B1(
        WIRE_ALU_A_MUX2TO1_32BIT_4__MUX_N1), .B2(n10033), .ZN(n10111) );
  XNOR2_X2 U11215 ( .A(n10111), .B(n4813), .ZN(n10038) );
  NAND2_X2 U11216 ( .A1(net71078), .A2(WIRE_ALU_A_MUX2TO1_32BIT_3__MUX_N1), 
        .ZN(n10037) );
  OAI22_X2 U11217 ( .A1(n5530), .A2(n6089), .B1(net76658), .B2(n6072), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11218 ( .A1(n5470), .A2(n6092), .B1(n6073), .B2(n6155), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11219 ( .A1(n6193), .A2(n5389), .B1(n6194), .B2(n6073), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11220 ( .A1(n6197), .A2(n5427), .B1(n6073), .B2(n6198), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11221 ( .A1(n5471), .A2(n6098), .B1(n6095), .B2(n6072), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11222 ( .A1(n5531), .A2(n6104), .B1(n6073), .B2(n6102), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11223 ( .A1(n5338), .A2(n6109), .B1(n6073), .B2(n6106), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11224 ( .A1(n5228), .A2(n6113), .B1(n6073), .B2(n6157), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11225 ( .A1(n5532), .A2(n6116), .B1(n6073), .B2(n6159), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11226 ( .A1(n5472), .A2(n6119), .B1(n6073), .B2(n6161), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11227 ( .A1(n6201), .A2(n5558), .B1(n6073), .B2(n6203), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11228 ( .A1(n5473), .A2(net76864), .B1(n6073), .B2(net76614), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11229 ( .A1(n6206), .A2(n5428), .B1(n6073), .B2(n6207), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11230 ( .A1(n5229), .A2(n6122), .B1(n6073), .B2(n6163), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11231 ( .A1(n5339), .A2(n6125), .B1(n6073), .B2(n6165), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11232 ( .A1(n5230), .A2(n6128), .B1(n6073), .B2(n6167), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11233 ( .A1(n5533), .A2(n6130), .B1(n6169), .B2(n6072), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11234 ( .A(n5957), .ZN(n10047) );
  OAI22_X2 U11235 ( .A1(n10047), .A2(n6133), .B1(n6171), .B2(n6072), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11236 ( .A1(n5231), .A2(n6137), .B1(n6173), .B2(n6072), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11237 ( .A1(n6210), .A2(n5429), .B1(n6211), .B2(n6072), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11238 ( .A1(REGFILE_reg_out_28__3_), .A2(n6175), .ZN(n10048) );
  OAI22_X2 U11239 ( .A1(n5045), .A2(n6140), .B1(net76548), .B2(n6072), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11240 ( .A1(n10615), .A2(REGFILE_reg_out_30__3_), .ZN(n10050) );
  NAND2_X2 U11241 ( .A1(net76488), .A2(REGFILE_reg_out_31__3_), .ZN(n10051) );
  OAI22_X2 U11242 ( .A1(n6216), .A2(n5046), .B1(net76318), .B2(n6072), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11243 ( .A1(n6218), .A2(n5559), .B1(n6219), .B2(n6072), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11244 ( .A1(n5474), .A2(n6145), .B1(n6182), .B2(n6072), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11245 ( .A1(n5475), .A2(net76708), .B1(n6147), .B2(n6072), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11246 ( .A1(n5534), .A2(net76694), .B1(n6184), .B2(n6072), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11247 ( .A1(n5476), .A2(n6151), .B1(n6186), .B2(n6072), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11248 ( .A1(n5535), .A2(n6154), .B1(n6073), .B2(n6188), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U11249 ( .A(n10054), .B(n10053), .ZN(n10056) );
  NAND2_X2 U11250 ( .A1(multOut[20]), .A2(net92392), .ZN(n10076) );
  NAND2_X2 U11251 ( .A1(n10058), .A2(n10057), .ZN(n10062) );
  NAND2_X2 U11252 ( .A1(n10060), .A2(n10059), .ZN(n10061) );
  NAND2_X2 U11253 ( .A1(n10062), .A2(n10061), .ZN(n10074) );
  NAND2_X2 U11254 ( .A1(n10064), .A2(n10063), .ZN(n10068) );
  NAND2_X2 U11255 ( .A1(n10066), .A2(n10065), .ZN(n10067) );
  NAND2_X2 U11256 ( .A1(n10068), .A2(n10067), .ZN(n10069) );
  MUX2_X2 U11257 ( .A(n10070), .B(n10069), .S(net71026), .Z(n10073) );
  INV_X4 U11258 ( .A(aluA[20]), .ZN(n10071) );
  NAND3_X2 U11259 ( .A1(n10077), .A2(n10076), .A3(n10075), .ZN(
        dmem_addr_out[20]) );
  INV_X4 U11260 ( .A(dmem_read_in[20]), .ZN(n10078) );
  NAND2_X2 U11261 ( .A1(n5573), .A2(n10079), .ZN(n10085) );
  INV_X4 U11262 ( .A(dmem_addr_out[20]), .ZN(n10082) );
  NAND2_X2 U11263 ( .A1(n10080), .A2(net77030), .ZN(n10081) );
  OAI221_X2 U11264 ( .B1(net77999), .B2(n10083), .C1(n10082), .C2(net76646), 
        .A(n10081), .ZN(n10084) );
  OAI21_X4 U11265 ( .B1(n10085), .B2(n10084), .A(reset), .ZN(n10090) );
  OAI22_X2 U11266 ( .A1(n5232), .A2(n6089), .B1(net76658), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11267 ( .A1(n5821), .A2(n6092), .B1(n6155), .B2(n6075), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11268 ( .A1(n6193), .A2(n5390), .B1(n6194), .B2(n6075), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11269 ( .A1(n6197), .A2(n5682), .B1(n6198), .B2(n6075), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11270 ( .A1(n5340), .A2(n6098), .B1(n6094), .B2(n6075), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11271 ( .A1(n5233), .A2(n6104), .B1(n6102), .B2(n6075), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11272 ( .A1(n5081), .A2(n6109), .B1(n6105), .B2(n6075), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11273 ( .A1(n5105), .A2(n6113), .B1(n6157), .B2(n6075), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11274 ( .A1(n5234), .A2(n6116), .B1(n6159), .B2(n6075), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11275 ( .A1(n5341), .A2(n6119), .B1(n6161), .B2(n6075), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11276 ( .A1(n6201), .A2(n5391), .B1(n6203), .B2(n6075), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11277 ( .A1(n5342), .A2(net76864), .B1(net76614), .B2(n6075), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11278 ( .A1(n6206), .A2(n5506), .B1(n6207), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11279 ( .A1(n5235), .A2(n6122), .B1(n6163), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11280 ( .A1(n5343), .A2(n6125), .B1(n6165), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11281 ( .A1(n5236), .A2(n6128), .B1(n6167), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11282 ( .A1(n5237), .A2(n6130), .B1(n6169), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11283 ( .A1(n5661), .A2(n6133), .B1(n6171), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11284 ( .A1(n5238), .A2(n6137), .B1(n6173), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11285 ( .A1(n6210), .A2(n5681), .B1(n6211), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11286 ( .A1(REGFILE_reg_out_28__20_), .A2(n10604), .ZN(n10086) );
  OAI21_X4 U11287 ( .B1(n6214), .B2(n6075), .A(n10086), .ZN(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11288 ( .A1(n10608), .A2(REGFILE_reg_out_29__20_), .ZN(n10087) );
  OAI21_X4 U11289 ( .B1(n10532), .B2(n6075), .A(n10087), .ZN(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11290 ( .A1(n5023), .A2(n6140), .B1(net76548), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11291 ( .A1(n10615), .A2(REGFILE_reg_out_30__20_), .ZN(n10088) );
  OAI21_X4 U11292 ( .B1(n10534), .B2(n6075), .A(n10088), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11293 ( .A1(net76488), .A2(REGFILE_reg_out_31__20_), .ZN(n10089)
         );
  OAI21_X4 U11294 ( .B1(net70509), .B2(n6075), .A(n10089), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11295 ( .A1(n6216), .A2(n5037), .B1(net76318), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11296 ( .A1(n6218), .A2(n5500), .B1(n6219), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11297 ( .A1(n5344), .A2(n6145), .B1(n6182), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11298 ( .A1(n5345), .A2(net76708), .B1(n6146), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11299 ( .A1(n5239), .A2(net76694), .B1(n6184), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11300 ( .A1(n5346), .A2(n6151), .B1(n6186), .B2(n6076), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11301 ( .A1(n5240), .A2(n6154), .B1(n6188), .B2(n6075), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  MUX2_X2 U11302 ( .A(net70696), .B(n10091), .S(net77084), .Z(n10150) );
  AOI22_X2 U11303 ( .A1(n10280), .A2(n10150), .B1(net71092), .B2(n10092), .ZN(
        n10107) );
  INV_X4 U11304 ( .A(n10094), .ZN(n10102) );
  NAND2_X2 U11305 ( .A1(net70720), .A2(aluA[18]), .ZN(n10098) );
  NAND4_X2 U11306 ( .A1(n10098), .A2(n10097), .A3(n10096), .A4(n10095), .ZN(
        n10100) );
  MUX2_X2 U11307 ( .A(n10101), .B(n10100), .S(n10099), .Z(net70713) );
  INV_X4 U11308 ( .A(n10104), .ZN(n10414) );
  NOR2_X4 U11309 ( .A1(n10105), .A2(n5041), .ZN(n10106) );
  XNOR2_X2 U11310 ( .A(n10165), .B(n10109), .ZN(n10166) );
  INV_X4 U11311 ( .A(n10110), .ZN(n10112) );
  OAI22_X2 U11312 ( .A1(n10112), .A2(n10404), .B1(n10111), .B2(n4813), .ZN(
        n10167) );
  XNOR2_X2 U11313 ( .A(n10166), .B(n10167), .ZN(n10114) );
  NAND2_X2 U11314 ( .A1(net71078), .A2(WIRE_ALU_A_MUX2TO1_32BIT_2__MUX_N1), 
        .ZN(n10113) );
  OAI22_X2 U11315 ( .A1(n5536), .A2(n6089), .B1(net76658), .B2(net77116), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11316 ( .A1(n5477), .A2(n6092), .B1(n6155), .B2(net77114), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11317 ( .A1(n6193), .A2(n5560), .B1(n6194), .B2(net77116), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11318 ( .A1(n6197), .A2(n4989), .B1(net77116), .B2(n6198), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11319 ( .A1(n5478), .A2(n6098), .B1(n6094), .B2(net77116), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11320 ( .A1(n5537), .A2(n6104), .B1(n10519), .B2(net77114), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11321 ( .A1(n5347), .A2(n6109), .B1(n6105), .B2(net77114), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11322 ( .A1(n5241), .A2(n6113), .B1(n6157), .B2(net77116), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11323 ( .A1(n5538), .A2(n6116), .B1(n6159), .B2(net77114), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11324 ( .A1(n5479), .A2(n6119), .B1(n6161), .B2(net77114), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11325 ( .A1(n6201), .A2(n5392), .B1(n6203), .B2(net77116), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11327 ( .A1(n10116), .A2(net76864), .B1(net76614), .B2(net77114), 
        .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11328 ( .A1(n6206), .A2(n4986), .B1(net77116), .B2(n6207), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11329 ( .A1(n5242), .A2(n6122), .B1(n6163), .B2(net77114), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11330 ( .A1(n5348), .A2(n6125), .B1(n6165), .B2(net77114), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11331 ( .A1(n5243), .A2(n6128), .B1(n6167), .B2(net77116), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11332 ( .A1(n5539), .A2(n6130), .B1(n6169), .B2(net77114), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11334 ( .A1(n10117), .A2(n6133), .B1(n6171), .B2(net77116), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11335 ( .A1(n5244), .A2(n6137), .B1(n6173), .B2(net77114), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11336 ( .A1(n6210), .A2(n4987), .B1(n6211), .B2(net77116), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11337 ( .A1(REGFILE_reg_out_28__2_), .A2(n6175), .ZN(n10118) );
  NAND2_X2 U11338 ( .A1(n10608), .A2(REGFILE_reg_out_29__2_), .ZN(n10119) );
  OAI22_X2 U11339 ( .A1(n5480), .A2(n6140), .B1(net76548), .B2(net77116), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11340 ( .A1(n6180), .A2(REGFILE_reg_out_30__2_), .ZN(n10120) );
  OAI22_X2 U11342 ( .A1(n6216), .A2(n10121), .B1(net76318), .B2(net77114), 
        .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11343 ( .A1(n6218), .A2(n5561), .B1(n6219), .B2(net77116), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11344 ( .A1(n5481), .A2(n6145), .B1(n6182), .B2(net77114), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11345 ( .A1(n5482), .A2(net76708), .B1(n6146), .B2(net77114), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11346 ( .A1(n5540), .A2(net76694), .B1(n6184), .B2(net77116), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11347 ( .A1(n5483), .A2(n6151), .B1(n6186), .B2(net77114), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11348 ( .A1(n5541), .A2(n6154), .B1(n6188), .B2(net77116), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  AOI22_X2 U11349 ( .A1(net71092), .A2(n10123), .B1(net71094), .B2(n10122), 
        .ZN(n10129) );
  NAND2_X2 U11350 ( .A1(n10280), .A2(n10124), .ZN(n10128) );
  INV_X4 U11351 ( .A(n10421), .ZN(n10380) );
  NAND3_X2 U11352 ( .A1(n10129), .A2(n10128), .A3(n10127), .ZN(n10130) );
  XNOR2_X2 U11353 ( .A(n10132), .B(n10131), .ZN(n10134) );
  NAND2_X2 U11354 ( .A1(net71078), .A2(WIRE_ALU_A_MUX2TO1_32BIT_10__MUX_N1), 
        .ZN(n10133) );
  NOR2_X4 U11355 ( .A1(n10136), .A2(n10135), .ZN(n10141) );
  OAI22_X2 U11356 ( .A1(n5106), .A2(n6089), .B1(net76658), .B2(n6078), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11357 ( .A(REGFILE_reg_out_10__10_), .ZN(n10143) );
  OAI22_X2 U11358 ( .A1(n10143), .A2(n6092), .B1(n6155), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11359 ( .A1(n6193), .A2(n5119), .B1(n6194), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11360 ( .A1(n6197), .A2(n5775), .B1(n6198), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11361 ( .A1(n5024), .A2(n6098), .B1(n6094), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11362 ( .A1(n5107), .A2(n6104), .B1(n6102), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11363 ( .A1(n10144), .A2(n6109), .B1(n6105), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11364 ( .A1(n5245), .A2(n6113), .B1(n6157), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11365 ( .A1(n5108), .A2(n6116), .B1(n6159), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11366 ( .A1(n5774), .A2(n6119), .B1(n6161), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11367 ( .A1(n6201), .A2(n5393), .B1(n6203), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11368 ( .A1(n4979), .A2(net76864), .B1(net76614), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11369 ( .A1(n6206), .A2(n5430), .B1(n6207), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11370 ( .A1(n5246), .A2(n6122), .B1(n6163), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11371 ( .A1(n5082), .A2(n6125), .B1(n6165), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11372 ( .A1(n5109), .A2(n6128), .B1(n6167), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11373 ( .A1(n5110), .A2(n6130), .B1(n6169), .B2(n6078), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11374 ( .A1(n5025), .A2(n6133), .B1(n6171), .B2(n6078), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11375 ( .A1(n5247), .A2(n6137), .B1(n6173), .B2(n6078), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11376 ( .A1(n6210), .A2(n5877), .B1(n6211), .B2(n6078), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11377 ( .A1(REGFILE_reg_out_28__10_), .A2(n6177), .ZN(n10145) );
  NAND2_X2 U11378 ( .A1(n10608), .A2(REGFILE_reg_out_29__10_), .ZN(n10146) );
  OAI22_X2 U11379 ( .A1(n5773), .A2(n6140), .B1(net76548), .B2(n6078), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11380 ( .A1(n10615), .A2(REGFILE_reg_out_30__10_), .ZN(n10147) );
  NAND2_X2 U11381 ( .A1(net76488), .A2(REGFILE_reg_out_31__10_), .ZN(n10148)
         );
  OAI22_X2 U11382 ( .A1(n6216), .A2(n5114), .B1(net76318), .B2(n6078), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11383 ( .A1(n6218), .A2(n5120), .B1(n6219), .B2(n6078), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11384 ( .A1(n5083), .A2(n6145), .B1(n6182), .B2(n6078), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11385 ( .A1(n5349), .A2(net76708), .B1(n6146), .B2(n6078), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11386 ( .A1(n5248), .A2(net76694), .B1(n6184), .B2(n6078), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11387 ( .A1(n5350), .A2(n6151), .B1(n6186), .B2(n6078), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11388 ( .A1(n5249), .A2(n6154), .B1(n6188), .B2(n6079), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  AOI22_X2 U11389 ( .A1(n10280), .A2(n10151), .B1(net71092), .B2(n10150), .ZN(
        net71277) );
  NAND2_X2 U11390 ( .A1(n10930), .A2(net70719), .ZN(n10154) );
  NAND2_X2 U11391 ( .A1(net70720), .A2(aluA[17]), .ZN(n10153) );
  NAND3_X4 U11392 ( .A1(n10155), .A2(n10154), .A3(n10153), .ZN(n10163) );
  NAND2_X2 U11393 ( .A1(n10156), .A2(net78051), .ZN(n10157) );
  INV_X4 U11394 ( .A(n10157), .ZN(n10162) );
  INV_X4 U11395 ( .A(n10158), .ZN(n10160) );
  OAI22_X2 U11396 ( .A1(n10160), .A2(n10544), .B1(n10159), .B2(net71273), .ZN(
        n10161) );
  AOI211_X4 U11397 ( .C1(net77084), .C2(n10163), .A(n10162), .B(n10161), .ZN(
        net70709) );
  INV_X4 U11398 ( .A(n10164), .ZN(n10416) );
  AOI22_X2 U11399 ( .A1(n10167), .A2(n10166), .B1(
        WIRE_ALU_A_MUX2TO1_32BIT_2__MUX_N1), .B2(n10165), .ZN(net70731) );
  XNOR2_X2 U11400 ( .A(net70734), .B(net71273), .ZN(net70735) );
  NAND2_X2 U11401 ( .A1(net77104), .A2(n4992), .ZN(n10169) );
  NAND2_X2 U11402 ( .A1(n4867), .A2(REGFILE_reg_out_0__1_), .ZN(n10168) );
  NAND2_X2 U11403 ( .A1(n6093), .A2(REGFILE_reg_out_10__1_), .ZN(n10170) );
  NAND2_X2 U11404 ( .A1(net77102), .A2(n4998), .ZN(n10173) );
  NAND2_X2 U11405 ( .A1(REGFILE_reg_out_11__1_), .A2(n4869), .ZN(n10172) );
  NAND2_X2 U11406 ( .A1(n10173), .A2(n10172), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11407 ( .A1(net77102), .A2(n4993), .ZN(n10175) );
  NAND2_X2 U11408 ( .A1(REGFILE_reg_out_12__1_), .A2(n4873), .ZN(n10174) );
  NAND2_X2 U11409 ( .A1(n10175), .A2(n10174), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11410 ( .A1(net77104), .A2(n6096), .ZN(n10177) );
  NAND2_X2 U11411 ( .A1(n10177), .A2(n10176), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11412 ( .A1(net77104), .A2(n6101), .ZN(n10179) );
  NAND2_X2 U11413 ( .A1(n4805), .A2(REGFILE_reg_out_14__1_), .ZN(n10178) );
  NAND2_X2 U11414 ( .A1(n10179), .A2(n10178), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11415 ( .A1(net77100), .A2(n6107), .ZN(n10181) );
  NAND2_X2 U11416 ( .A1(n4804), .A2(REGFILE_reg_out_15__1_), .ZN(n10180) );
  NAND2_X2 U11417 ( .A1(n10181), .A2(n10180), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11418 ( .A1(net77104), .A2(n4994), .ZN(n10183) );
  NAND2_X2 U11419 ( .A1(n4891), .A2(REGFILE_reg_out_16__1_), .ZN(n10182) );
  NAND2_X2 U11420 ( .A1(n10183), .A2(n10182), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11421 ( .A1(net77102), .A2(n4999), .ZN(n10185) );
  NAND2_X2 U11422 ( .A1(n4892), .A2(REGFILE_reg_out_17__1_), .ZN(n10184) );
  NAND2_X2 U11423 ( .A1(net77104), .A2(n5000), .ZN(n10187) );
  NAND2_X2 U11424 ( .A1(n4884), .A2(REGFILE_reg_out_18__1_), .ZN(n10186) );
  NAND2_X2 U11425 ( .A1(net77100), .A2(n5001), .ZN(n10189) );
  NAND2_X2 U11426 ( .A1(REGFILE_reg_out_19__1_), .A2(n4876), .ZN(n10188) );
  NAND2_X2 U11427 ( .A1(n10189), .A2(n10188), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11428 ( .A1(net77100), .A2(n4903), .ZN(n10191) );
  NAND2_X2 U11429 ( .A1(REGFILE_reg_out_20__1_), .A2(n4868), .ZN(n10190) );
  NAND2_X2 U11430 ( .A1(net77100), .A2(n4904), .ZN(n10193) );
  NAND2_X2 U11431 ( .A1(n4882), .A2(REGFILE_reg_out_21__1_), .ZN(n10192) );
  NAND2_X2 U11432 ( .A1(n10193), .A2(n10192), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11433 ( .A1(n10947), .A2(n4905), .ZN(n10195) );
  NAND2_X2 U11435 ( .A1(n10195), .A2(n10194), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11436 ( .A1(net77102), .A2(n4906), .ZN(n10197) );
  NAND2_X2 U11437 ( .A1(n4883), .A2(REGFILE_reg_out_23__1_), .ZN(n10196) );
  NAND2_X2 U11438 ( .A1(net77102), .A2(n4995), .ZN(n10199) );
  NAND2_X2 U11439 ( .A1(n4875), .A2(REGFILE_reg_out_24__1_), .ZN(n10198) );
  NAND2_X2 U11440 ( .A1(n10199), .A2(n10198), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11441 ( .A1(net77100), .A2(n5002), .ZN(n10201) );
  NAND2_X2 U11442 ( .A1(n4878), .A2(REGFILE_reg_out_25__1_), .ZN(n10200) );
  NAND2_X2 U11443 ( .A1(n10201), .A2(n10200), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11444 ( .A1(net77100), .A2(n5003), .ZN(n10203) );
  NAND2_X2 U11445 ( .A1(n4893), .A2(REGFILE_reg_out_26__1_), .ZN(n10202) );
  NAND2_X2 U11446 ( .A1(net77104), .A2(n5004), .ZN(n10205) );
  NAND2_X2 U11447 ( .A1(REGFILE_reg_out_27__1_), .A2(n4872), .ZN(n10204) );
  NAND2_X2 U11448 ( .A1(REGFILE_reg_out_28__1_), .A2(n6175), .ZN(n10206) );
  NAND2_X2 U11449 ( .A1(n10608), .A2(REGFILE_reg_out_29__1_), .ZN(n10208) );
  NAND2_X2 U11450 ( .A1(net77102), .A2(n5005), .ZN(n10211) );
  NAND2_X2 U11451 ( .A1(n4879), .A2(REGFILE_reg_out_2__1_), .ZN(n10210) );
  NAND2_X2 U11452 ( .A1(n10211), .A2(n10210), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11453 ( .A1(n10615), .A2(REGFILE_reg_out_30__1_), .ZN(n10212) );
  NAND2_X2 U11454 ( .A1(net76488), .A2(REGFILE_reg_out_31__1_), .ZN(n10214) );
  NAND2_X2 U11455 ( .A1(REGFILE_reg_out_3__1_), .A2(n4871), .ZN(n10216) );
  NAND2_X2 U11456 ( .A1(n10217), .A2(n10216), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11457 ( .A1(net77100), .A2(n4996), .ZN(n10219) );
  NAND2_X2 U11458 ( .A1(REGFILE_reg_out_4__1_), .A2(n4870), .ZN(n10218) );
  NAND2_X2 U11459 ( .A1(net77102), .A2(n5006), .ZN(n10221) );
  NAND2_X2 U11460 ( .A1(n4885), .A2(REGFILE_reg_out_5__1_), .ZN(n10220) );
  NAND2_X2 U11461 ( .A1(net77102), .A2(n6148), .ZN(n10223) );
  NAND2_X2 U11462 ( .A1(n4889), .A2(REGFILE_reg_out_6__1_), .ZN(n10222) );
  NAND2_X2 U11463 ( .A1(n10223), .A2(n10222), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11464 ( .A1(net77100), .A2(n5007), .ZN(n10225) );
  NAND2_X2 U11465 ( .A1(n4886), .A2(REGFILE_reg_out_7__1_), .ZN(n10224) );
  NAND2_X2 U11466 ( .A1(n10225), .A2(n10224), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11467 ( .A1(net77104), .A2(n4991), .ZN(n10227) );
  NAND2_X2 U11468 ( .A1(n4890), .A2(REGFILE_reg_out_8__1_), .ZN(n10226) );
  NAND2_X2 U11469 ( .A1(n10227), .A2(n10226), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11470 ( .A1(net77102), .A2(n5008), .ZN(n10229) );
  NAND2_X2 U11471 ( .A1(n4887), .A2(REGFILE_reg_out_9__1_), .ZN(n10228) );
  NAND2_X2 U11472 ( .A1(n10229), .A2(n10228), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11473 ( .A1(n6082), .A2(n10230), .ZN(n10237) );
  NAND2_X2 U11474 ( .A1(n6083), .A2(n10231), .ZN(n10236) );
  NAND2_X2 U11475 ( .A1(n8759), .A2(n10232), .ZN(n10235) );
  NAND2_X2 U11476 ( .A1(net105360), .A2(n10233), .ZN(n10234) );
  NAND4_X2 U11477 ( .A1(n10237), .A2(n10236), .A3(n10235), .A4(n10234), .ZN(
        n10279) );
  NAND2_X2 U11478 ( .A1(n8728), .A2(n10238), .ZN(n10245) );
  NAND2_X2 U11479 ( .A1(net77084), .A2(n10239), .ZN(n10244) );
  NAND2_X2 U11480 ( .A1(n6082), .A2(n10240), .ZN(n10243) );
  NAND2_X2 U11481 ( .A1(n6083), .A2(n10241), .ZN(n10242) );
  NAND4_X2 U11482 ( .A1(n10245), .A2(n10244), .A3(n10243), .A4(n10242), .ZN(
        n10282) );
  AOI22_X2 U11483 ( .A1(net71092), .A2(n10279), .B1(net71094), .B2(n10282), 
        .ZN(n10251) );
  NAND2_X2 U11484 ( .A1(n10280), .A2(n10246), .ZN(n10250) );
  INV_X4 U11485 ( .A(n10425), .ZN(n10366) );
  NAND3_X2 U11486 ( .A1(n10251), .A2(n10250), .A3(n10249), .ZN(n10252) );
  MUX2_X2 U11487 ( .A(n10252), .B(multOut[14]), .S(net76452), .Z(n10258) );
  XNOR2_X2 U11488 ( .A(n10254), .B(n10253), .ZN(n10256) );
  NAND2_X2 U11489 ( .A1(net71078), .A2(WIRE_ALU_A_MUX2TO1_32BIT_14__MUX_N1), 
        .ZN(n10255) );
  NOR2_X4 U11490 ( .A1(n10258), .A2(n10257), .ZN(n10263) );
  INV_X4 U11491 ( .A(n10263), .ZN(dmem_addr_out[14]) );
  OAI211_X2 U11492 ( .C1(n10263), .C2(net76646), .A(net70740), .B(n10262), 
        .ZN(n10264) );
  NAND2_X2 U11493 ( .A1(reset), .A2(n10264), .ZN(n10276) );
  OAI22_X2 U11494 ( .A1(n5029), .A2(n6090), .B1(net76658), .B2(n10276), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11495 ( .A1(n5844), .A2(n10512), .B1(n6155), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11496 ( .A(n5777), .ZN(n10265) );
  OAI22_X2 U11497 ( .A1(n6193), .A2(n10265), .B1(n6194), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11498 ( .A1(n6197), .A2(n10266), .B1(n6198), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11499 ( .A1(n5843), .A2(n6099), .B1(n6094), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11500 ( .A1(n4928), .A2(n6104), .B1(n10519), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11501 ( .A(REGFILE_reg_out_15__14_), .ZN(n10267) );
  OAI22_X2 U11502 ( .A1(n10267), .A2(n6110), .B1(n6105), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11503 ( .A1(n5819), .A2(n6111), .B1(n6157), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11504 ( .A1(n4929), .A2(n6114), .B1(n6159), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11505 ( .A1(n5842), .A2(n6117), .B1(n6161), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11506 ( .A1(n6201), .A2(n5394), .B1(n6203), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11507 ( .A1(n5841), .A2(net76866), .B1(net76614), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11508 ( .A(n5781), .ZN(n10268) );
  OAI22_X2 U11509 ( .A1(n6206), .A2(n10268), .B1(n6207), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11510 ( .A1(n4930), .A2(n6120), .B1(n6163), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11511 ( .A1(n5837), .A2(n6123), .B1(n6165), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11512 ( .A1(n4931), .A2(n6126), .B1(n6167), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11513 ( .A1(n5662), .A2(n6131), .B1(n6169), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11514 ( .A1(n10269), .A2(n6134), .B1(n6171), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11515 ( .A1(n4936), .A2(n6135), .B1(n6173), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11516 ( .A1(n6210), .A2(n10270), .B1(n6211), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11517 ( .A1(n10608), .A2(REGFILE_reg_out_29__14_), .ZN(n10272) );
  OAI22_X2 U11518 ( .A1(n5838), .A2(n6141), .B1(net76548), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11519 ( .A1(n10615), .A2(REGFILE_reg_out_30__14_), .ZN(n10273) );
  NAND2_X2 U11520 ( .A1(net76488), .A2(REGFILE_reg_out_31__14_), .ZN(n10274)
         );
  OAI22_X2 U11521 ( .A1(n6216), .A2(n4981), .B1(net76318), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11522 ( .A1(n6218), .A2(n5395), .B1(n6219), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11523 ( .A(n5832), .ZN(n10275) );
  OAI22_X2 U11524 ( .A1(n10275), .A2(n6143), .B1(n6182), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11525 ( .A1(n4926), .A2(net76716), .B1(n6146), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11526 ( .A1(n4932), .A2(net76702), .B1(n6184), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11527 ( .A1(n4918), .A2(n6149), .B1(n6186), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11528 ( .A1(n4933), .A2(n6152), .B1(n6188), .B2(n6085), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  AOI22_X2 U11529 ( .A1(net71092), .A2(n10278), .B1(net71094), .B2(n10277), 
        .ZN(n10285) );
  NAND2_X2 U11530 ( .A1(n10280), .A2(n10279), .ZN(n10284) );
  NAND3_X2 U11531 ( .A1(n10285), .A2(n10284), .A3(n10283), .ZN(n10286) );
  MUX2_X2 U11532 ( .A(n10286), .B(multOut[15]), .S(net76452), .Z(n10292) );
  XNOR2_X2 U11533 ( .A(n10287), .B(n4807), .ZN(n10290) );
  NAND2_X2 U11534 ( .A1(net71078), .A2(WIRE_ALU_A_MUX2TO1_32BIT_15__MUX_N1), 
        .ZN(n10289) );
  NOR2_X4 U11535 ( .A1(n10292), .A2(n10291), .ZN(n10296) );
  INV_X4 U11536 ( .A(n10296), .ZN(dmem_addr_out[15]) );
  INV_X4 U11537 ( .A(dmem_read_in[15]), .ZN(n10504) );
  OAI211_X2 U11538 ( .C1(n10296), .C2(net76646), .A(net70740), .B(n10295), 
        .ZN(n10297) );
  OAI22_X2 U11539 ( .A1(n5250), .A2(n6090), .B1(net76658), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11540 ( .A1(n10298), .A2(n10512), .B1(n6155), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11541 ( .A1(n6193), .A2(n5121), .B1(n6194), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11542 ( .A1(n6197), .A2(n5856), .B1(n6198), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11543 ( .A1(n5714), .A2(n6099), .B1(n6094), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11544 ( .A1(n4941), .A2(n6103), .B1(n10519), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11545 ( .A1(n5866), .A2(n6110), .B1(n6105), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11546 ( .A1(n4954), .A2(n6111), .B1(n6157), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11547 ( .A1(n4942), .A2(n6114), .B1(n6159), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11548 ( .A1(n4901), .A2(n6117), .B1(n6161), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11549 ( .A1(n6201), .A2(n5122), .B1(n6203), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11550 ( .A1(n5656), .A2(net76866), .B1(net76614), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11551 ( .A1(n6206), .A2(n5431), .B1(n6207), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11552 ( .A1(n4943), .A2(n6120), .B1(n6163), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11553 ( .A1(n4919), .A2(n6123), .B1(n6165), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11554 ( .A1(n4934), .A2(n6126), .B1(n6167), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11555 ( .A1(n5251), .A2(n6131), .B1(n6169), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11556 ( .A1(n5784), .A2(n6134), .B1(n6171), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11557 ( .A1(n4944), .A2(n6135), .B1(n6173), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11558 ( .A1(n6210), .A2(n5683), .B1(n6211), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11559 ( .A1(n10608), .A2(REGFILE_reg_out_29__15_), .ZN(n10300) );
  OAI22_X2 U11560 ( .A1(n5917), .A2(n6141), .B1(net76548), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11561 ( .A1(n10615), .A2(REGFILE_reg_out_30__15_), .ZN(n10301) );
  NAND2_X2 U11562 ( .A1(net76488), .A2(REGFILE_reg_out_31__15_), .ZN(n10302)
         );
  OAI22_X2 U11563 ( .A1(n6216), .A2(n5038), .B1(net76318), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11564 ( .A1(n6218), .A2(n5396), .B1(n6219), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11565 ( .A1(n4902), .A2(n6143), .B1(n6182), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11566 ( .A1(n4948), .A2(net76716), .B1(n6146), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11567 ( .A1(n4945), .A2(net76702), .B1(n6184), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11568 ( .A1(n4927), .A2(n6149), .B1(n6186), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11569 ( .A1(n4935), .A2(n6152), .B1(n6188), .B2(n6087), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11570 ( .A1(n10303), .A2(net77040), .ZN(n10305) );
  XNOR2_X2 U11571 ( .A(net80189), .B(n10928), .ZN(n10434) );
  INV_X4 U11572 ( .A(n10434), .ZN(n10459) );
  NAND2_X2 U11573 ( .A1(n10306), .A2(n10399), .ZN(n10308) );
  XNOR2_X2 U11574 ( .A(net71027), .B(net70535), .ZN(net70703) );
  NOR2_X4 U11575 ( .A1(n10470), .A2(n10434), .ZN(n10311) );
  OAI21_X4 U11576 ( .B1(n10311), .B2(n10310), .A(n10309), .ZN(n10314) );
  AOI21_X4 U11577 ( .B1(n10442), .B2(n10314), .A(n10313), .ZN(n10318) );
  OAI21_X4 U11578 ( .B1(n10318), .B2(n10317), .A(n10316), .ZN(n10322) );
  INV_X4 U11579 ( .A(n10436), .ZN(n10321) );
  AOI21_X4 U11580 ( .B1(n10322), .B2(n10321), .A(n10320), .ZN(n10326) );
  NAND2_X2 U11581 ( .A1(aluA[26]), .A2(n10323), .ZN(n10324) );
  OAI21_X4 U11582 ( .B1(n10326), .B2(n10325), .A(n10324), .ZN(n10330) );
  INV_X4 U11583 ( .A(n10435), .ZN(n10329) );
  AOI21_X4 U11584 ( .B1(n10330), .B2(n10329), .A(n10328), .ZN(n10333) );
  OAI21_X4 U11585 ( .B1(n10430), .B2(n10333), .A(n10332), .ZN(n10337) );
  AOI21_X4 U11586 ( .B1(n10337), .B2(n10336), .A(n10335), .ZN(n10340) );
  NAND2_X2 U11587 ( .A1(n10932), .A2(n10338), .ZN(n10339) );
  OAI21_X4 U11588 ( .B1(n10432), .B2(n10340), .A(n10339), .ZN(n10344) );
  INV_X4 U11589 ( .A(n10443), .ZN(n10347) );
  INV_X4 U11590 ( .A(aluA[19]), .ZN(n10349) );
  INV_X4 U11591 ( .A(aluA[17]), .ZN(n10356) );
  INV_X4 U11592 ( .A(n10447), .ZN(n10360) );
  OAI21_X4 U11593 ( .B1(n10361), .B2(n10360), .A(n10359), .ZN(n10363) );
  OAI21_X4 U11594 ( .B1(n10374), .B2(n10373), .A(n10372), .ZN(n10377) );
  INV_X4 U11595 ( .A(n10411), .ZN(n10413) );
  OAI21_X4 U11596 ( .B1(n10413), .B2(n10416), .A(n10412), .ZN(n10486) );
  NAND2_X2 U11597 ( .A1(net70703), .A2(n10486), .ZN(net70838) );
  OAI21_X4 U11598 ( .B1(net70703), .B2(n10486), .A(net70838), .ZN(n10485) );
  INV_X4 U11599 ( .A(n10485), .ZN(n10417) );
  NOR4_X2 U11600 ( .A1(n10417), .A2(n10416), .A3(n10415), .A4(n10414), .ZN(
        n10454) );
  NAND2_X2 U11601 ( .A1(n10425), .A2(n10424), .ZN(n10426) );
  NOR3_X4 U11602 ( .A1(n10428), .A2(n10427), .A3(n10426), .ZN(n10453) );
  NAND2_X2 U11603 ( .A1(n10434), .A2(n10433), .ZN(n10437) );
  NAND4_X2 U11604 ( .A1(n10455), .A2(n10454), .A3(n10453), .A4(n10452), .ZN(
        n10456) );
  INV_X4 U11605 ( .A(n10456), .ZN(n10484) );
  MUX2_X2 U11606 ( .A(n10459), .B(n10458), .S(n10457), .Z(n10460) );
  NOR2_X4 U11607 ( .A1(n10461), .A2(n10460), .ZN(n10477) );
  OAI221_X2 U11608 ( .B1(net70866), .B2(n10464), .C1(net70868), .C2(n10463), 
        .A(n10462), .ZN(n10469) );
  INV_X4 U11609 ( .A(n10466), .ZN(n10467) );
  NOR2_X4 U11610 ( .A1(n10467), .A2(n10544), .ZN(n10468) );
  AOI211_X4 U11611 ( .C1(n10469), .C2(net105360), .A(n4811), .B(n10468), .ZN(
        n10473) );
  OAI221_X2 U11612 ( .B1(n4812), .B2(n10474), .C1(n10473), .C2(n10472), .A(
        n10471), .ZN(n10480) );
  NAND2_X2 U11613 ( .A1(n10480), .A2(n10475), .ZN(n10476) );
  MUX2_X2 U11614 ( .A(n10477), .B(n10476), .S(net70826), .Z(n10478) );
  NAND4_X2 U11615 ( .A1(net77040), .A2(n10494), .A3(net70826), .A4(n10484), 
        .ZN(n10479) );
  NAND2_X2 U11616 ( .A1(n10478), .A2(n10479), .ZN(n10501) );
  INV_X4 U11617 ( .A(n10479), .ZN(n10483) );
  INV_X4 U11618 ( .A(n10480), .ZN(n10481) );
  NOR2_X4 U11619 ( .A1(n10481), .A2(net70845), .ZN(n10482) );
  NOR2_X4 U11620 ( .A1(n10483), .A2(n10482), .ZN(n10499) );
  XNOR2_X2 U11621 ( .A(n10486), .B(n10485), .ZN(n10487) );
  XNOR2_X2 U11622 ( .A(n10487), .B(net70837), .ZN(n10489) );
  NAND2_X2 U11623 ( .A1(n10488), .A2(n10489), .ZN(n10497) );
  INV_X4 U11624 ( .A(n10489), .ZN(n10495) );
  MUX2_X2 U11625 ( .A(n10492), .B(n10491), .S(n10490), .Z(n10493) );
  MUX2_X2 U11626 ( .A(n10497), .B(n10496), .S(net70826), .Z(n10498) );
  NAND2_X2 U11627 ( .A1(n10499), .A2(n10498), .ZN(n10500) );
  MUX2_X2 U11628 ( .A(n10501), .B(n10500), .S(net70821), .Z(n10502) );
  MUX2_X2 U11629 ( .A(n10502), .B(multOut[31]), .S(net76452), .Z(
        dmem_addr_out[31]) );
  AOI22_X2 U11630 ( .A1(dmem_read_in[31]), .A2(dmem_dsize[0]), .B1(
        instructionAddr_out[31]), .B2(net77030), .ZN(n10510) );
  INV_X4 U11631 ( .A(dmem_addr_out[31]), .ZN(n10503) );
  NOR3_X4 U11632 ( .A1(n10508), .A2(n10507), .A3(n10506), .ZN(n10509) );
  AOI21_X4 U11633 ( .B1(n10510), .B2(n10509), .A(net76278), .ZN(n10511) );
  OAI22_X2 U11634 ( .A1(n10513), .A2(n10512), .B1(n6191), .B2(n6155), .ZN(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11635 ( .A(REGFILE_reg_out_11__31_), .ZN(n10514) );
  OAI22_X2 U11636 ( .A1(n6193), .A2(n10514), .B1(n6194), .B2(n6191), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11637 ( .A1(n6197), .A2(n10515), .B1(n6198), .B2(n6191), .ZN(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11638 ( .A1(n10518), .A2(n6099), .B1(n6191), .B2(n6094), .ZN(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11639 ( .A1(n10520), .A2(n6103), .B1(n6191), .B2(n6102), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11640 ( .A1(n10522), .A2(n6110), .B1(n6191), .B2(n6105), .ZN(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11641 ( .A1(n10523), .A2(n6111), .B1(n6191), .B2(n6157), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11642 ( .A1(n4917), .A2(n6114), .B1(n6191), .B2(n6159), .ZN(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11643 ( .A1(n10524), .A2(n6117), .B1(n6191), .B2(n6161), .ZN(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11644 ( .A1(n6201), .A2(n5026), .B1(n6203), .B2(n6191), .ZN(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11645 ( .A1(net70780), .A2(net76866), .B1(n6191), .B2(net76614), 
        .ZN(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11646 ( .A1(n6206), .A2(n10525), .B1(n6207), .B2(n6191), .ZN(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11647 ( .A1(n4939), .A2(n6120), .B1(n6191), .B2(n6163), .ZN(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11648 ( .A(REGFILE_reg_out_22__31_), .ZN(n10526) );
  OAI22_X2 U11649 ( .A1(n10526), .A2(n6123), .B1(n6191), .B2(n6165), .ZN(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11650 ( .A1(n4953), .A2(n6126), .B1(n6191), .B2(n6167), .ZN(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11651 ( .A1(n5999), .A2(n6131), .B1(n6191), .B2(n6169), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11652 ( .A(REGFILE_reg_out_25__31_), .ZN(n10527) );
  OAI22_X2 U11653 ( .A1(n10527), .A2(n6134), .B1(n6191), .B2(n6171), .ZN(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11654 ( .A(REGFILE_reg_out_26__31_), .ZN(n10528) );
  OAI22_X2 U11655 ( .A1(n10528), .A2(n6135), .B1(n6191), .B2(n6173), .ZN(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11656 ( .A(REGFILE_reg_out_27__31_), .ZN(n10529) );
  OAI22_X2 U11657 ( .A1(n6210), .A2(n10529), .B1(n6211), .B2(n6191), .ZN(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11658 ( .A1(REGFILE_reg_out_28__31_), .A2(n6175), .ZN(n10530) );
  NAND2_X2 U11659 ( .A1(n6178), .A2(REGFILE_reg_out_29__31_), .ZN(n10531) );
  OAI22_X2 U11660 ( .A1(net70761), .A2(n6141), .B1(n6191), .B2(net76548), .ZN(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11661 ( .A1(n6180), .A2(REGFILE_reg_out_30__31_), .ZN(n10533) );
  INV_X4 U11662 ( .A(REGFILE_reg_out_3__31_), .ZN(net70758) );
  OAI22_X2 U11663 ( .A1(n6216), .A2(net70758), .B1(net76318), .B2(n6191), .ZN(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11664 ( .A1(n6218), .A2(net70757), .B1(n6219), .B2(n6191), .ZN(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11665 ( .A(REGFILE_reg_out_5__31_), .ZN(net70755) );
  OAI22_X2 U11666 ( .A1(net70755), .A2(n6143), .B1(n6191), .B2(n6182), .ZN(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11667 ( .A(REGFILE_reg_out_6__31_), .ZN(net70752) );
  OAI22_X2 U11668 ( .A1(net70752), .A2(net76716), .B1(n6191), .B2(n6146), .ZN(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11669 ( .A(REGFILE_reg_out_7__31_), .ZN(net70750) );
  OAI22_X2 U11670 ( .A1(net70750), .A2(net76702), .B1(n6191), .B2(n6184), .ZN(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  INV_X4 U11671 ( .A(REGFILE_reg_out_8__31_), .ZN(n10536) );
  OAI22_X2 U11672 ( .A1(n10536), .A2(n6149), .B1(n6191), .B2(n6186), .ZN(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U11673 ( .A1(n10537), .A2(n6152), .B1(n6191), .B2(n6188), .ZN(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11674 ( .A1(instructionAddr_out[1]), .A2(n10538), .ZN(n10539) );
  XNOR2_X2 U11675 ( .A(n10539), .B(n5439), .ZN(n10644) );
  OAI211_X2 U11676 ( .C1(net70738), .C2(n10644), .A(n5572), .B(net70740), .ZN(
        net70737) );
  INV_X4 U11677 ( .A(net70737), .ZN(net70685) );
  INV_X4 U11678 ( .A(n10541), .ZN(n10545) );
  NAND2_X2 U11679 ( .A1(n10542), .A2(net70534), .ZN(n10543) );
  OAI21_X4 U11680 ( .B1(n10545), .B2(n10544), .A(n10543), .ZN(net70714) );
  INV_X4 U11681 ( .A(net70687), .ZN(net70684) );
  NAND2_X2 U11682 ( .A1(n10546), .A2(net76510), .ZN(n10548) );
  NAND2_X2 U11683 ( .A1(n10549), .A2(net76510), .ZN(n10551) );
  NAND2_X2 U11684 ( .A1(n6093), .A2(REGFILE_reg_out_10__0_), .ZN(n10550) );
  NAND2_X2 U11685 ( .A1(n10552), .A2(net76510), .ZN(n10554) );
  NAND2_X2 U11686 ( .A1(REGFILE_reg_out_11__0_), .A2(n4869), .ZN(n10553) );
  NAND2_X2 U11687 ( .A1(n10555), .A2(net76510), .ZN(n10557) );
  NAND2_X2 U11688 ( .A1(REGFILE_reg_out_12__0_), .A2(n4873), .ZN(n10556) );
  NAND2_X2 U11690 ( .A1(n4805), .A2(REGFILE_reg_out_14__0_), .ZN(n10560) );
  NAND2_X2 U11691 ( .A1(n4804), .A2(REGFILE_reg_out_15__0_), .ZN(n10562) );
  NAND2_X2 U11692 ( .A1(n10564), .A2(net76510), .ZN(n10566) );
  NAND2_X2 U11693 ( .A1(n4891), .A2(REGFILE_reg_out_16__0_), .ZN(n10565) );
  NAND2_X2 U11694 ( .A1(n10567), .A2(net76510), .ZN(n10569) );
  NAND2_X2 U11695 ( .A1(n10570), .A2(net76510), .ZN(n10572) );
  NAND2_X2 U11696 ( .A1(n4884), .A2(REGFILE_reg_out_18__0_), .ZN(n10571) );
  NAND2_X2 U11697 ( .A1(n10573), .A2(net76510), .ZN(n10575) );
  NAND2_X2 U11698 ( .A1(REGFILE_reg_out_19__0_), .A2(n4876), .ZN(n10574) );
  NAND2_X2 U11699 ( .A1(n10576), .A2(net76510), .ZN(n10578) );
  NAND2_X2 U11700 ( .A1(n4877), .A2(REGFILE_reg_out_1__0_), .ZN(n10577) );
  NAND2_X2 U11701 ( .A1(n10579), .A2(net76510), .ZN(n10581) );
  NAND2_X2 U11703 ( .A1(n10582), .A2(net76510), .ZN(n10584) );
  NAND2_X2 U11704 ( .A1(n4882), .A2(REGFILE_reg_out_21__0_), .ZN(n10583) );
  NAND2_X2 U11705 ( .A1(n10585), .A2(net76510), .ZN(n10587) );
  NAND2_X2 U11706 ( .A1(n4888), .A2(REGFILE_reg_out_22__0_), .ZN(n10586) );
  NAND2_X2 U11707 ( .A1(n10588), .A2(net76510), .ZN(n10590) );
  NAND2_X2 U11709 ( .A1(n10591), .A2(net76510), .ZN(n10593) );
  NAND2_X2 U11710 ( .A1(n4875), .A2(REGFILE_reg_out_24__0_), .ZN(n10592) );
  NAND2_X2 U11711 ( .A1(n10594), .A2(net76510), .ZN(n10596) );
  NAND2_X2 U11712 ( .A1(n4878), .A2(REGFILE_reg_out_25__0_), .ZN(n10595) );
  NAND2_X2 U11713 ( .A1(n10597), .A2(net76510), .ZN(n10599) );
  NAND2_X2 U11714 ( .A1(n4893), .A2(REGFILE_reg_out_26__0_), .ZN(n10598) );
  NAND2_X2 U11715 ( .A1(n10600), .A2(net76510), .ZN(n10602) );
  NAND2_X2 U11716 ( .A1(REGFILE_reg_out_27__0_), .A2(n4872), .ZN(n10601) );
  NAND2_X2 U11717 ( .A1(n10603), .A2(net76510), .ZN(n10606) );
  NAND2_X2 U11718 ( .A1(REGFILE_reg_out_28__0_), .A2(n6175), .ZN(n10605) );
  NAND2_X2 U11719 ( .A1(n10608), .A2(REGFILE_reg_out_29__0_), .ZN(n10609) );
  NAND2_X2 U11720 ( .A1(n10611), .A2(net76510), .ZN(n10613) );
  NAND2_X2 U11722 ( .A1(n10615), .A2(REGFILE_reg_out_30__0_), .ZN(n10616) );
  NAND2_X2 U11724 ( .A1(n10620), .A2(net76510), .ZN(n10622) );
  NAND2_X2 U11725 ( .A1(REGFILE_reg_out_3__0_), .A2(n4871), .ZN(n10621) );
  NAND2_X2 U11726 ( .A1(n10623), .A2(net76510), .ZN(n10625) );
  NAND2_X2 U11727 ( .A1(REGFILE_reg_out_4__0_), .A2(n4870), .ZN(n10624) );
  NAND2_X2 U11728 ( .A1(n10626), .A2(net76510), .ZN(n10628) );
  NAND2_X2 U11729 ( .A1(n4885), .A2(REGFILE_reg_out_5__0_), .ZN(n10627) );
  NAND2_X2 U11731 ( .A1(n10631), .A2(net76510), .ZN(n10633) );
  NAND2_X2 U11733 ( .A1(n10634), .A2(net76510), .ZN(n10636) );
  NAND2_X2 U11735 ( .A1(net76510), .A2(n10637), .ZN(n10639) );
  INV_X4 U11737 ( .A(net70535), .ZN(net70534) );
  NAND2_X2 U11738 ( .A1(net73708), .A2(net70534), .ZN(n10648) );
  INV_X4 U11739 ( .A(n10640), .ZN(n10641) );
  XNOR2_X2 U11740 ( .A(n10641), .B(net70529), .ZN(n10642) );
  INV_X4 U11741 ( .A(n10642), .ZN(n10643) );
  NAND2_X2 U11742 ( .A1(n10649), .A2(n10643), .ZN(n10645) );
  MUX2_X2 U11743 ( .A(n10646), .B(n10645), .S(n10644), .Z(n10647) );
  NAND2_X2 U11744 ( .A1(n10648), .A2(n10647), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11745 ( .A1(n10649), .A2(instruction[31]), .ZN(n10653) );
  MUX2_X2 U11746 ( .A(n10653), .B(n10652), .S(instructionAddr_out[31]), .Z(
        n10654) );
  NAND2_X2 U11747 ( .A1(n10655), .A2(n10654), .ZN(
        PCLOGIC_PC_REG_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U11748 ( .A1(net76488), .A2(REGFILE_reg_out_31__31_), .ZN(n10656)
         );
  INV_X4 U11749 ( .A(net70506), .ZN(dmem_writeEnable_out) );
  INV_X4 U11750 ( .A(REGFILE_reg_out_20__29_), .ZN(n10935) );
  INV_X4 U11751 ( .A(REGFILE_reg_out_28__30_), .ZN(n10937) );
  INV_X4 U11752 ( .A(REGFILE_reg_out_27__30_), .ZN(n10938) );
  INV_X4 U11753 ( .A(REGFILE_reg_out_20__30_), .ZN(n10939) );
  INV_X4 U11754 ( .A(REGFILE_reg_out_12__30_), .ZN(n10940) );
  INV_X4 U11755 ( .A(REGFILE_reg_out_11__30_), .ZN(n10941) );
  DFF_X1 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__0_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__0_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__5_), .QN(n5415) );
  DFF_X1 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__5_), .QN(n5312) );
  DFF_X1 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__5_), .QN(n5311) );
  DFF_X1 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__4_), .QN(n5465) );
  DFF_X1 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__4_), .QN(n5329) );
  DFF_X1 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__4_), .QN(n5526) );
  DFF_X1 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__4_), .QN(n5525) );
  DFF_X1 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__4_), .QN(n5438) );
  DFF_X1 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__4_), .QN(n5524) );
  DFF_X1 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__4_), .QN(n5528) );
  DFF_X1 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__4_), .QN(n5467) );
  DFF_X1 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__4_), .QN(n5466) );
  DFF_X1 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__4_), .QN(n5331) );
  DFF_X1 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__4_), .QN(n5469) );
  DFF_X1 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__4_), .QN(n5048) );
  DFF_X1 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__4_), .QN(n5527) );
  DFF_X1 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__4_), .QN(n5529) );
  DFF_X1 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__4_), .QN(n5330) );
  DFF_X1 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__4_), .QN(n5424) );
  DFF_X1 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__4_), .QN(n5423) );
  DFF_X1 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__4_), .QN(n5557) );
  DFF_X1 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__2_), .QN(n4989) );
  DFF_X1 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__2_), .QN(n5347) );
  DFF_X1 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__2_), .QN(n5482) );
  DFF_X1 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__2_), .QN(n5537) );
  DFF_X1 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__2_), .QN(n5539) );
  DFF_X1 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__2_), .QN(n5348) );
  DFF_X1 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__2_), .QN(n5479) );
  DFF_X1 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__2_), .QN(n5538) );
  DFF_X1 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__2_), .QN(n5477) );
  DFF_X1 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__2_), .QN(n5483) );
  DFF_X1 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__2_), .QN(n5481) );
  DFF_X1 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__2_), .QN(n5478) );
  DFF_X1 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__2_), .QN(n5560) );
  DFF_X1 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__2_), .QN(n5561) );
  DFF_X1 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__2_), .QN(n5541) );
  DFF_X1 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__2_), .QN(n5540) );
  DFF_X1 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__2_), .QN(n5480) );
  DFF_X1 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__2_), .QN(n5536) );
  DFF_X1 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__3_), .QN(n5338) );
  DFF_X1 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__3_), .QN(n5558) );
  DFF_X1 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__3_), .QN(n5427) );
  DFF_X1 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__3_), .QN(n5230) );
  DFF_X1 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__3_), .QN(n5339) );
  DFF_X1 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__3_), .QN(n5229) );
  DFF_X1 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__3_), .QN(n5472) );
  DFF_X1 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__3_), .QN(n5532) );
  DFF_X1 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__3_), .QN(n5228) );
  DFF_X1 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__3_), .QN(n5470) );
  DFF_X1 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__3_), .QN(n5535) );
  DFF_X1 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__3_), .QN(n5473) );
  DFF_X1 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__3_), .QN(n5531) );
  DFF_X1 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__3_), .QN(n5471) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[30]), .QN(n5014) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[29]), .QN(n5016) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[27]), .QN(n4969) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__27_), .QN(n5492) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__26_), .QN(n5519) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__26_), .QN(n5520) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[15]), .QN(n5064) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[12]), .QN(n4908) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__25_), .QN(n5510) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__25_), .QN(n5552) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__25_), .QN(n5509) );
  DFF_X2 PCLOGIC_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( .D(
        PCLOGIC_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        instructionAddr_out[11]), .QN(n5060) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__23_), .QN(n5512) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__23_), .QN(n5511) );
  DFF_X1 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__27_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__26_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__25_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__25_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__23_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(n5902), .QN(n9675) );
  DFF_X1 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__2_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__2_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__3_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__3_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__2_), .QN(n10121) );
  DFF_X1 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__2_), .QN(n10116) );
  DFF_X1 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__2_), .QN(n10117) );
  DFF_X1 REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_13__0_) );
  DFF_X1 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(n5982), .QN(n9973) );
  DFF_X1 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__5_), .QN(n9641) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(n5764) );
  DFF_X2 REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_15__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_0__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_27__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_26__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_25__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_22__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_21__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_19__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_18__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_16__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_12__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_4__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_3__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_1__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_10__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_6__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_17__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_2__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_23__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_20__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_9__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_8__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_7__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_5__0_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__2_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__3_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__2_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_28__4_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_31__4_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_30__4_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__4_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__5_), .QN(n9639) );
  DFF_X2 REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_11__5_), .QN(n9638) );
  DFF_X2 REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_24__5_), .QN(n9640) );
  DFF_X2 REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_29__5_) );
  DFF_X2 REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REGFILE_reg_out_14__0_) );
  INV_X8 U4890 ( .A(n4881), .ZN(n10945) );
  INV_X8 U4892 ( .A(n4881), .ZN(net78042) );
  AOI22_X2 U4900 ( .A1(REGFILE_reg_out_26__18_), .A2(net75439), .B1(n4818), 
        .B2(net75440), .ZN(n6545) );
  AOI22_X2 U4901 ( .A1(REGFILE_reg_out_30__20_), .A2(net84761), .B1(
        REGFILE_reg_out_2__20_), .B2(net82613), .ZN(n6498) );
  AOI22_X1 U4914 ( .A1(REGFILE_reg_out_30__27_), .A2(net77638), .B1(
        REGFILE_reg_out_2__27_), .B2(net75442), .ZN(n6337) );
  INV_X8 U4917 ( .A(n10947), .ZN(n10946) );
  AOI21_X4 U4929 ( .B1(net81874), .B2(n4970), .A(net76274), .ZN(n10947) );
  NAND2_X2 U4930 ( .A1(net73838), .A2(net77272), .ZN(n4830) );
  INV_X8 U4934 ( .A(net77856), .ZN(net77854) );
  INV_X1 U5036 ( .A(net73837), .ZN(n10948) );
  INV_X4 U5043 ( .A(n10948), .ZN(n10949) );
  INV_X2 U5049 ( .A(n10950), .ZN(n10951) );
  NAND2_X1 U5060 ( .A1(REGFILE_reg_out_28__0_), .A2(net77388), .ZN(n8237) );
  NAND2_X1 U5066 ( .A1(REGFILE_reg_out_28__22_), .A2(net77388), .ZN(n7267) );
  NAND2_X1 U5083 ( .A1(REGFILE_reg_out_28__23_), .A2(net77388), .ZN(n7222) );
  NAND2_X1 U5094 ( .A1(REGFILE_reg_out_4__23_), .A2(net77388), .ZN(n7232) );
  NAND2_X1 U5168 ( .A1(REGFILE_reg_out_12__23_), .A2(net77388), .ZN(n7242) );
  NAND2_X1 U5171 ( .A1(REGFILE_reg_out_20__23_), .A2(net77388), .ZN(n7252) );
  NAND2_X1 U5175 ( .A1(REGFILE_reg_out_28__24_), .A2(net77388), .ZN(n7177) );
  NAND2_X1 U5185 ( .A1(REGFILE_reg_out_4__24_), .A2(net77388), .ZN(n7187) );
  NAND2_X1 U5291 ( .A1(REGFILE_reg_out_12__24_), .A2(net77388), .ZN(n7197) );
  NAND2_X1 U5919 ( .A1(REGFILE_reg_out_20__24_), .A2(net77388), .ZN(n7207) );
  NAND2_X1 U6111 ( .A1(REGFILE_reg_out_4__25_), .A2(net77388), .ZN(n7142) );
  NAND2_X1 U6117 ( .A1(REGFILE_reg_out_12__25_), .A2(net77388), .ZN(n7152) );
  NAND2_X1 U6118 ( .A1(REGFILE_reg_out_20__25_), .A2(net77388), .ZN(n7162) );
  NAND2_X1 U6380 ( .A1(net77388), .A2(REGFILE_reg_out_20__27_), .ZN(n7058) );
  AOI22_X2 U6493 ( .A1(REGFILE_reg_out_21__31_), .A2(net77458), .B1(n5766), 
        .B2(net77388), .ZN(n6923) );
  NAND2_X1 U6537 ( .A1(net77298), .A2(REGFILE_reg_out_0__28_), .ZN(n7032) );
  NAND2_X1 U6546 ( .A1(net77298), .A2(REGFILE_reg_out_16__28_), .ZN(n7012) );
  NAND2_X1 U6547 ( .A1(REGFILE_reg_out_16__1_), .A2(net77300), .ZN(n8201) );
  NAND2_X1 U6679 ( .A1(net77300), .A2(REGFILE_reg_out_0__27_), .ZN(n7076) );
  NAND2_X1 U6756 ( .A1(REGFILE_reg_out_0__1_), .A2(net77300), .ZN(n8221) );
  NAND2_X1 U6833 ( .A1(REGFILE_reg_out_8__0_), .A2(net77300), .ZN(n8255) );
  NAND2_X1 U6834 ( .A1(REGFILE_reg_out_24__1_), .A2(net77300), .ZN(n8191) );
  NAND2_X1 U6895 ( .A1(REGFILE_reg_out_8__1_), .A2(net77300), .ZN(n8211) );
  NAND4_X2 U6947 ( .A1(net75417), .A2(net75416), .A3(net75415), .A4(net75414), 
        .ZN(net73849) );
  NAND4_X2 U6962 ( .A1(n6927), .A2(n6928), .A3(n6926), .A4(n6925), .ZN(n8401)
         );
  INV_X16 U6984 ( .A(instruction[11]), .ZN(n5574) );
  OAI22_X2 U7135 ( .A1(n9640), .A2(n6130), .B1(n6053), .B2(n6169), .ZN(
        REGFILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7213 ( .A1(n9639), .A2(n6104), .B1(n6054), .B2(n6102), .ZN(
        REGFILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7363 ( .A1(n6193), .A2(n9638), .B1(n6054), .B2(n6195), .ZN(
        REGFILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI211_X2 U7428 ( .C1(n9967), .C2(net76646), .A(net70740), .B(n9966), .ZN(
        n9968) );
  NOR2_X2 U7492 ( .A1(n4815), .A2(n5571), .ZN(n4898) );
  NAND2_X1 U7494 ( .A1(n4890), .A2(REGFILE_reg_out_8__12_), .ZN(n9174) );
  NAND2_X1 U7495 ( .A1(REGFILE_reg_out_8__12_), .A2(net77308), .ZN(n7729) );
  INV_X32 U7626 ( .A(instruction[8]), .ZN(net73879) );
  AOI22_X2 U8002 ( .A1(REGFILE_reg_out_1__30_), .A2(net77514), .B1(
        REGFILE_reg_out_0__30_), .B2(net77298), .ZN(n6938) );
  INV_X4 U8019 ( .A(n5842), .ZN(n10953) );
  NAND2_X2 U8072 ( .A1(net77346), .A2(REGFILE_reg_out_18__14_), .ZN(n7632) );
  INV_X4 U8082 ( .A(net76260), .ZN(net75481) );
  INV_X8 U8092 ( .A(n6050), .ZN(n6048) );
  INV_X8 U8106 ( .A(n6050), .ZN(n6049) );
  INV_X8 U8116 ( .A(n6050), .ZN(n4801) );
  OAI211_X4 U8126 ( .C1(n9519), .C2(net76646), .A(net70740), .B(n9518), .ZN(
        n9520) );
  OAI22_X2 U8136 ( .A1(n5195), .A2(n6113), .B1(n6054), .B2(n6157), .ZN(
        REGFILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  INV_X8 U8151 ( .A(dmem_addr_out[5]), .ZN(n9636) );
  OAI21_X2 U8161 ( .B1(net70509), .B2(n6072), .A(n10051), .ZN(
        REGFILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  AOI21_X2 U8171 ( .B1(net73878), .B2(net81974), .A(net73997), .ZN(n8374) );
  OAI21_X2 U8181 ( .B1(net77114), .B2(n10534), .A(n10120), .ZN(
        REGFILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  BUF_X4 U8196 ( .A(n10924), .Z(n5762) );
  MUX2_X2 U8574 ( .A(multOut[8]), .B(n9506), .S(net73585), .Z(n9515) );
  NAND2_X4 U8581 ( .A1(multOut[7]), .A2(net92392), .ZN(n9698) );
  NAND4_X4 U8996 ( .A1(n9630), .A2(n9631), .A3(n9632), .A4(n9629), .ZN(
        dmem_addr_out[5]) );
  NAND2_X4 U9003 ( .A1(multOut[5]), .A2(net92392), .ZN(n9630) );
  NAND2_X1 U9011 ( .A1(n4886), .A2(REGFILE_reg_out_7__0_), .ZN(n10632) );
  NAND2_X1 U9019 ( .A1(n4890), .A2(REGFILE_reg_out_8__0_), .ZN(n10635) );
  NAND2_X1 U9027 ( .A1(n4883), .A2(REGFILE_reg_out_23__0_), .ZN(n10589) );
  NAND2_X1 U9044 ( .A1(n4887), .A2(REGFILE_reg_out_9__0_), .ZN(n10638) );
  NAND2_X1 U9334 ( .A1(n4879), .A2(REGFILE_reg_out_2__0_), .ZN(n10612) );
  NAND2_X1 U9577 ( .A1(REGFILE_reg_out_20__0_), .A2(n4868), .ZN(n10580) );
  NAND2_X1 U10179 ( .A1(n4889), .A2(REGFILE_reg_out_6__0_), .ZN(n10629) );
  NAND2_X1 U10194 ( .A1(net76488), .A2(REGFILE_reg_out_31__0_), .ZN(n10618) );
  NAND2_X1 U10574 ( .A1(n6100), .A2(REGFILE_reg_out_13__0_), .ZN(n10558) );
  INV_X16 U10580 ( .A(net76508), .ZN(net76502) );
  NAND2_X1 U10694 ( .A1(n4888), .A2(REGFILE_reg_out_22__1_), .ZN(n10194) );
  NAND2_X1 U10710 ( .A1(REGFILE_reg_out_3__12_), .A2(n4871), .ZN(n9164) );
  NAND2_X1 U10711 ( .A1(REGFILE_reg_out_3__12_), .A2(net77416), .ZN(n7742) );
  AOI22_X4 U10714 ( .A1(REGFILE_reg_out_14__16_), .A2(net77780), .B1(n5611), 
        .B2(n5664), .ZN(n6569) );
  AOI22_X4 U10715 ( .A1(REGFILE_reg_out_14__18_), .A2(net77780), .B1(
        REGFILE_reg_out_13__18_), .B2(n6009), .ZN(n6537) );
  AOI22_X4 U10718 ( .A1(REGFILE_reg_out_0__18_), .A2(net120684), .B1(
        REGFILE_reg_out_10__18_), .B2(net83203), .ZN(n6534) );
  INV_X8 U10719 ( .A(instruction[11]), .ZN(net81974) );
  INV_X32 U10721 ( .A(instruction[11]), .ZN(net82618) );
  INV_X16 U10730 ( .A(instruction[11]), .ZN(n4820) );
  INV_X2 U10731 ( .A(net77328), .ZN(net77324) );
  INV_X4 U10733 ( .A(net77328), .ZN(net77320) );
  NAND2_X1 U10767 ( .A1(net82613), .A2(n5836), .ZN(n5942) );
  AOI21_X4 U10800 ( .B1(dmem_write_out[16]), .B2(net73509), .A(n5933), .ZN(
        n11001) );
  INV_X8 U11140 ( .A(n11001), .ZN(n10917) );
  INV_X8 U11326 ( .A(net78056), .ZN(net73509) );
  NAND3_X2 MULT_mult_6_U4863 ( .A1(MULT_mult_6_net119921), .A2(
        MULT_mult_6_n490), .A3(MULT_mult_6_net82029), .ZN(MULT_mult_6_n123) );
  CLKBUF_X3 MULT_mult_6_U4862 ( .A(MULT_mult_6_SUMB_9__10_), .Z(
        MULT_mult_6_net91419) );
  NAND2_X4 MULT_mult_6_U4861 ( .A1(MULT_mult_6_ab_23__2_), .A2(
        MULT_mult_6_n394), .ZN(MULT_mult_6_n2295) );
  NAND2_X4 MULT_mult_6_U4860 ( .A1(MULT_mult_6_CARRYB_13__6_), .A2(
        MULT_mult_6_SUMB_13__7_), .ZN(MULT_mult_6_n1976) );
  XNOR2_X2 MULT_mult_6_U4859 ( .A(MULT_mult_6_n173), .B(MULT_mult_6_ab_11__7_), 
        .ZN(MULT_mult_6_n1717) );
  NOR2_X1 MULT_mult_6_U4858 ( .A1(MULT_mult_6_net123000), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__17_) );
  NAND2_X4 MULT_mult_6_U4503 ( .A1(MULT_mult_6_net83919), .A2(
        MULT_mult_6_ab_5__14_), .ZN(MULT_mult_6_n479) );
  NAND2_X4 MULT_mult_6_U4466 ( .A1(MULT_mult_6_CARRYB_4__14_), .A2(
        MULT_mult_6_ab_5__14_), .ZN(MULT_mult_6_n480) );
  NAND2_X4 MULT_mult_6_U4373 ( .A1(MULT_mult_6_n805), .A2(MULT_mult_6_n660), 
        .ZN(MULT_mult_6_net81992) );
  INV_X2 MULT_mult_6_U4338 ( .A(MULT_mult_6_net123000), .ZN(
        MULT_mult_6_net123072) );
  NAND2_X2 MULT_mult_6_U3936 ( .A1(MULT_mult_6_CARRYB_18__1_), .A2(
        MULT_mult_6_SUMB_18__2_), .ZN(MULT_mult_6_net81097) );
  BUF_X8 MULT_mult_6_U3738 ( .A(MULT_mult_6_SUMB_18__2_), .Z(MULT_mult_6_n359)
         );
  NAND3_X2 MULT_mult_6_U3730 ( .A1(MULT_mult_6_net81216), .A2(MULT_mult_6_n461), .A3(MULT_mult_6_net81215), .ZN(MULT_mult_6_n2378) );
  NAND3_X2 MULT_mult_6_U3678 ( .A1(MULT_mult_6_n1964), .A2(MULT_mult_6_n1966), 
        .A3(MULT_mult_6_n1965), .ZN(MULT_mult_6_n2377) );
  BUF_X4 MULT_mult_6_U3672 ( .A(MULT_mult_6_SUMB_5__9_), .Z(MULT_mult_6_n1214)
         );
  CLKBUF_X2 MULT_mult_6_U3625 ( .A(MULT_mult_6_n2010), .Z(MULT_mult_6_n2376)
         );
  NAND2_X1 MULT_mult_6_U3603 ( .A1(MULT_mult_6_ab_10__16_), .A2(
        MULT_mult_6_CARRYB_9__16_), .ZN(MULT_mult_6_n2164) );
  NAND2_X2 MULT_mult_6_U3602 ( .A1(MULT_mult_6_n1730), .A2(MULT_mult_6_n1191), 
        .ZN(MULT_mult_6_n1629) );
  CLKBUF_X3 MULT_mult_6_U3585 ( .A(MULT_mult_6_n152), .Z(MULT_mult_6_n290) );
  NAND2_X2 MULT_mult_6_U3549 ( .A1(MULT_mult_6_net82548), .A2(
        MULT_mult_6_net149580), .ZN(MULT_mult_6_n1124) );
  INV_X8 MULT_mult_6_U3548 ( .A(MULT_mult_6_n1277), .ZN(MULT_mult_6_n1278) );
  INV_X4 MULT_mult_6_U3537 ( .A(MULT_mult_6_SUMB_12__8_), .ZN(MULT_mult_6_n313) );
  NAND2_X2 MULT_mult_6_U3536 ( .A1(MULT_mult_6_CARRYB_6__7_), .A2(
        MULT_mult_6_n1499), .ZN(MULT_mult_6_n1443) );
  NAND2_X4 MULT_mult_6_U3520 ( .A1(MULT_mult_6_ab_6__7_), .A2(MULT_mult_6_n853), .ZN(MULT_mult_6_n1331) );
  XNOR2_X2 MULT_mult_6_U3396 ( .A(MULT_mult_6_n1309), .B(MULT_mult_6_n1208), 
        .ZN(MULT_mult_6_n2375) );
  NAND2_X2 MULT_mult_6_U3395 ( .A1(MULT_mult_6_net88303), .A2(
        MULT_mult_6_CARRYB_11__10_), .ZN(MULT_mult_6_net92552) );
  INV_X16 MULT_mult_6_U3386 ( .A(MULT_mult_6_n90), .ZN(MULT_mult_6_net81424)
         );
  OR2_X2 MULT_mult_6_U3381 ( .A1(MULT_mult_6_net81424), .A2(
        MULT_mult_6_net77964), .ZN(MULT_mult_6_n353) );
  INV_X4 MULT_mult_6_U3379 ( .A(MULT_mult_6_CARRYB_21__4_), .ZN(
        MULT_mult_6_n73) );
  INV_X2 MULT_mult_6_U3233 ( .A(MULT_mult_6_net88887), .ZN(
        MULT_mult_6_net88800) );
  NAND2_X4 MULT_mult_6_U3232 ( .A1(MULT_mult_6_n1582), .A2(
        MULT_mult_6_net84708), .ZN(MULT_mult_6_net92542) );
  INV_X2 MULT_mult_6_U3114 ( .A(MULT_mult_6_CARRYB_23__2_), .ZN(
        MULT_mult_6_net147938) );
  INV_X2 MULT_mult_6_U3056 ( .A(MULT_mult_6_n585), .ZN(MULT_mult_6_n289) );
  INV_X2 MULT_mult_6_U2811 ( .A(MULT_mult_6_n1456), .ZN(
        MULT_mult_6_SUMB_5__11_) );
  INV_X4 MULT_mult_6_U2772 ( .A(MULT_mult_6_n1456), .ZN(MULT_mult_6_n2374) );
  NAND2_X2 MULT_mult_6_U2734 ( .A1(MULT_mult_6_SUMB_8__13_), .A2(
        MULT_mult_6_net89149), .ZN(MULT_mult_6_net81375) );
  NAND2_X4 MULT_mult_6_U2648 ( .A1(MULT_mult_6_n1383), .A2(MULT_mult_6_n1382), 
        .ZN(MULT_mult_6_n11) );
  CLKBUF_X3 MULT_mult_6_U2579 ( .A(MULT_mult_6_SUMB_21__1_), .Z(
        MULT_mult_6_n1280) );
  NAND2_X2 MULT_mult_6_U2526 ( .A1(MULT_mult_6_ab_21__1_), .A2(
        MULT_mult_6_SUMB_20__2_), .ZN(MULT_mult_6_n2161) );
  NAND2_X4 MULT_mult_6_U2452 ( .A1(MULT_mult_6_ab_22__1_), .A2(
        MULT_mult_6_CARRYB_21__1_), .ZN(MULT_mult_6_net82542) );
  CLKBUF_X3 MULT_mult_6_U2379 ( .A(MULT_mult_6_SUMB_15__4_), .Z(
        MULT_mult_6_n871) );
  NAND3_X2 MULT_mult_6_U2338 ( .A1(MULT_mult_6_net81110), .A2(
        MULT_mult_6_net81111), .A3(MULT_mult_6_net81112), .ZN(
        MULT_mult_6_n2373) );
  XNOR2_X2 MULT_mult_6_U2335 ( .A(MULT_mult_6_n2372), .B(
        MULT_mult_6_CARRYB_23__0_), .ZN(multOut[7]) );
  XNOR2_X2 MULT_mult_6_U2254 ( .A(MULT_mult_6_n23), .B(MULT_mult_6_ab_24__0_), 
        .ZN(MULT_mult_6_n2372) );
  NAND2_X2 MULT_mult_6_U2252 ( .A1(MULT_mult_6_SUMB_9__5_), .A2(
        MULT_mult_6_ab_10__4_), .ZN(MULT_mult_6_n1924) );
  NAND2_X2 MULT_mult_6_U2194 ( .A1(MULT_mult_6_ab_14__3_), .A2(
        MULT_mult_6_CARRYB_13__3_), .ZN(MULT_mult_6_n1967) );
  XNOR2_X2 MULT_mult_6_U2193 ( .A(MULT_mult_6_ab_4__5_), .B(
        MULT_mult_6_CARRYB_3__5_), .ZN(MULT_mult_6_n2371) );
  XNOR2_X2 MULT_mult_6_U2160 ( .A(MULT_mult_6_n2371), .B(
        MULT_mult_6_SUMB_3__6_), .ZN(MULT_mult_6_SUMB_4__5_) );
  NAND3_X2 MULT_mult_6_U2159 ( .A1(MULT_mult_6_n1926), .A2(MULT_mult_6_n1925), 
        .A3(MULT_mult_6_n1924), .ZN(MULT_mult_6_n2370) );
  INV_X32 MULT_mult_6_U2093 ( .A(MULT_mult_6_ab_3__7_), .ZN(MULT_mult_6_n2369)
         );
  XNOR2_X2 MULT_mult_6_U2086 ( .A(MULT_mult_6_n566), .B(MULT_mult_6_n2369), 
        .ZN(MULT_mult_6_net85734) );
  XNOR2_X2 MULT_mult_6_U2002 ( .A(MULT_mult_6_n396), .B(
        MULT_mult_6_CARRYB_17__1_), .ZN(MULT_mult_6_SUMB_18__1_) );
  XOR2_X2 MULT_mult_6_U1995 ( .A(MULT_mult_6_ab_19__0_), .B(
        MULT_mult_6_SUMB_18__1_), .Z(MULT_mult_6_n1812) );
  XNOR2_X1 MULT_mult_6_U1973 ( .A(MULT_mult_6_CARRYB_14__1_), .B(
        MULT_mult_6_ab_15__1_), .ZN(MULT_mult_6_n2368) );
  XNOR2_X2 MULT_mult_6_U1869 ( .A(MULT_mult_6_SUMB_14__2_), .B(
        MULT_mult_6_n2368), .ZN(MULT_mult_6_SUMB_15__1_) );
  XOR2_X2 MULT_mult_6_U1774 ( .A(MULT_mult_6_CARRYB_9__1_), .B(
        MULT_mult_6_ab_10__1_), .Z(MULT_mult_6_n1470) );
  NAND2_X4 MULT_mult_6_U1772 ( .A1(MULT_mult_6_SUMB_1__16_), .A2(
        MULT_mult_6_ab_2__15_), .ZN(MULT_mult_6_n1985) );
  XNOR2_X2 MULT_mult_6_U1767 ( .A(MULT_mult_6_ab_4__20_), .B(
        MULT_mult_6_CARRYB_3__20_), .ZN(MULT_mult_6_n2367) );
  NAND2_X4 MULT_mult_6_U1738 ( .A1(MULT_mult_6_net84070), .A2(
        MULT_mult_6_net81256), .ZN(MULT_mult_6_net84071) );
  INV_X2 MULT_mult_6_U1629 ( .A(MULT_mult_6_SUMB_14__9_), .ZN(
        MULT_mult_6_net88934) );
  NAND2_X4 MULT_mult_6_U1527 ( .A1(MULT_mult_6_n877), .A2(MULT_mult_6_n878), 
        .ZN(MULT_mult_6_n1626) );
  NAND2_X2 MULT_mult_6_U1275 ( .A1(MULT_mult_6_n1554), .A2(MULT_mult_6_n1555), 
        .ZN(MULT_mult_6_n150) );
  NAND2_X4 MULT_mult_6_U1215 ( .A1(MULT_mult_6_SUMB_6__17_), .A2(
        MULT_mult_6_ab_7__16_), .ZN(MULT_mult_6_n2250) );
  NAND2_X2 MULT_mult_6_U1214 ( .A1(MULT_mult_6_n372), .A2(
        MULT_mult_6_ab_22__2_), .ZN(MULT_mult_6_net80926) );
  BUF_X4 MULT_mult_6_U1181 ( .A(MULT_mult_6_CARRYB_21__6_), .Z(
        MULT_mult_6_net89008) );
  INV_X4 MULT_mult_6_U1178 ( .A(MULT_mult_6_n1274), .ZN(MULT_mult_6_n1275) );
  NAND2_X2 MULT_mult_6_U1165 ( .A1(MULT_mult_6_n224), .A2(MULT_mult_6_n225), 
        .ZN(MULT_mult_6_n227) );
  INV_X4 MULT_mult_6_U1156 ( .A(MULT_mult_6_n541), .ZN(MULT_mult_6_n542) );
  NAND2_X4 MULT_mult_6_U1153 ( .A1(MULT_mult_6_n597), .A2(
        MULT_mult_6_ab_25__0_), .ZN(MULT_mult_6_net81531) );
  NAND2_X2 MULT_mult_6_U1126 ( .A1(MULT_mult_6_CARRYB_24__2_), .A2(
        MULT_mult_6_ab_25__2_), .ZN(MULT_mult_6_n131) );
  XOR2_X2 MULT_mult_6_U997 ( .A(MULT_mult_6_CARRYB_2__13_), .B(
        MULT_mult_6_ab_3__13_), .Z(MULT_mult_6_n2366) );
  INV_X4 MULT_mult_6_U995 ( .A(MULT_mult_6_CARRYB_24__2_), .ZN(
        MULT_mult_6_n129) );
  NAND2_X2 MULT_mult_6_U961 ( .A1(MULT_mult_6_n1033), .A2(MULT_mult_6_n1034), 
        .ZN(MULT_mult_6_net81070) );
  NAND2_X4 MULT_mult_6_U938 ( .A1(MULT_mult_6_n2363), .A2(MULT_mult_6_n334), 
        .ZN(MULT_mult_6_net147939) );
  INV_X32 MULT_mult_6_U899 ( .A(MULT_mult_6_net121380), .ZN(MULT_mult_6_n2365)
         );
  XNOR2_X2 MULT_mult_6_U886 ( .A(MULT_mult_6_net86519), .B(MULT_mult_6_n2365), 
        .ZN(MULT_mult_6_n2364) );
  XNOR2_X2 MULT_mult_6_U884 ( .A(MULT_mult_6_net86519), .B(
        MULT_mult_6_net121380), .ZN(MULT_mult_6_n2363) );
  INV_X4 MULT_mult_6_U837 ( .A(MULT_mult_6_n1718), .ZN(MULT_mult_6_n634) );
  INV_X2 MULT_mult_6_U832 ( .A(MULT_mult_6_net86662), .ZN(
        MULT_mult_6_net148235) );
  INV_X2 MULT_mult_6_U828 ( .A(MULT_mult_6_SUMB_11__6_), .ZN(MULT_mult_6_n1274) );
  INV_X16 MULT_mult_6_U808 ( .A(MULT_mult_6_net70491), .ZN(MULT_mult_6_n26) );
  NAND2_X4 MULT_mult_6_U804 ( .A1(MULT_mult_6_n1029), .A2(MULT_mult_6_n1030), 
        .ZN(MULT_mult_6_n1032) );
  NAND2_X4 MULT_mult_6_U716 ( .A1(MULT_mult_6_n2370), .A2(MULT_mult_6_n563), 
        .ZN(MULT_mult_6_n1832) );
  NAND2_X2 MULT_mult_6_U704 ( .A1(MULT_mult_6_ab_15__1_), .A2(
        MULT_mult_6_CARRYB_14__1_), .ZN(MULT_mult_6_n653) );
  NAND2_X2 MULT_mult_6_U703 ( .A1(MULT_mult_6_ab_16__1_), .A2(
        MULT_mult_6_CARRYB_15__1_), .ZN(MULT_mult_6_n648) );
  BUF_X2 MULT_mult_6_U693 ( .A(MULT_mult_6_SUMB_6__7_), .Z(MULT_mult_6_n1208)
         );
  NAND2_X2 MULT_mult_6_U684 ( .A1(MULT_mult_6_SUMB_2__13_), .A2(
        MULT_mult_6_n1324), .ZN(MULT_mult_6_n2007) );
  NAND2_X2 MULT_mult_6_U682 ( .A1(MULT_mult_6_SUMB_2__13_), .A2(
        MULT_mult_6_ab_3__12_), .ZN(MULT_mult_6_n2008) );
  NAND2_X1 MULT_mult_6_U672 ( .A1(MULT_mult_6_ab_3__17_), .A2(
        MULT_mult_6_CARRYB_2__17_), .ZN(MULT_mult_6_n1714) );
  NAND3_X4 MULT_mult_6_U658 ( .A1(MULT_mult_6_net80941), .A2(
        MULT_mult_6_net80942), .A3(MULT_mult_6_net80940), .ZN(
        MULT_mult_6_CARRYB_22__6_) );
  NAND2_X4 MULT_mult_6_U639 ( .A1(MULT_mult_6_net79863), .A2(MULT_mult_6_n1090), .ZN(MULT_mult_6_net80110) );
  NAND2_X4 MULT_mult_6_U637 ( .A1(MULT_mult_6_n58), .A2(MULT_mult_6_n59), .ZN(
        MULT_mult_6_n61) );
  NAND2_X4 MULT_mult_6_U633 ( .A1(MULT_mult_6_n1431), .A2(MULT_mult_6_n1432), 
        .ZN(MULT_mult_6_n1434) );
  NAND2_X4 MULT_mult_6_U628 ( .A1(MULT_mult_6_n60), .A2(MULT_mult_6_n61), .ZN(
        MULT_mult_6_n933) );
  INV_X2 MULT_mult_6_U617 ( .A(MULT_mult_6_n544), .ZN(MULT_mult_6_n547) );
  NAND3_X2 MULT_mult_6_U579 ( .A1(MULT_mult_6_n892), .A2(MULT_mult_6_n893), 
        .A3(MULT_mult_6_n894), .ZN(MULT_mult_6_CARRYB_17__12_) );
  XNOR2_X2 MULT_mult_6_U569 ( .A(MULT_mult_6_CARRYB_7__9_), .B(
        MULT_mult_6_ab_8__9_), .ZN(MULT_mult_6_n2362) );
  NAND2_X2 MULT_mult_6_U505 ( .A1(MULT_mult_6_CARRYB_5__6_), .A2(
        MULT_mult_6_SUMB_5__7_), .ZN(MULT_mult_6_n1949) );
  NAND2_X2 MULT_mult_6_U485 ( .A1(MULT_mult_6_CARRYB_5__6_), .A2(
        MULT_mult_6_ab_6__6_), .ZN(MULT_mult_6_n1951) );
  INV_X4 MULT_mult_6_U467 ( .A(MULT_mult_6_ab_2__16_), .ZN(MULT_mult_6_n280)
         );
  INV_X2 MULT_mult_6_U465 ( .A(MULT_mult_6_n280), .ZN(MULT_mult_6_n2361) );
  NAND2_X4 MULT_mult_6_U455 ( .A1(MULT_mult_6_CARRYB_21__3_), .A2(
        MULT_mult_6_ab_22__3_), .ZN(MULT_mult_6_n502) );
  NAND2_X4 MULT_mult_6_U448 ( .A1(MULT_mult_6_n817), .A2(MULT_mult_6_net87363), 
        .ZN(MULT_mult_6_net82029) );
  NAND2_X2 MULT_mult_6_U446 ( .A1(MULT_mult_6_n9), .A2(MULT_mult_6_net92568), 
        .ZN(MULT_mult_6_n499) );
  INV_X2 MULT_mult_6_U444 ( .A(MULT_mult_6_net92790), .ZN(MULT_mult_6_net92568) );
  NAND2_X2 MULT_mult_6_U443 ( .A1(MULT_mult_6_net85461), .A2(MULT_mult_6_n517), 
        .ZN(MULT_mult_6_SUMB_8__13_) );
  NAND2_X4 MULT_mult_6_U430 ( .A1(MULT_mult_6_net85461), .A2(MULT_mult_6_n517), 
        .ZN(MULT_mult_6_n2360) );
  NAND2_X2 MULT_mult_6_U428 ( .A1(MULT_mult_6_CARRYB_8__12_), .A2(
        MULT_mult_6_ab_9__12_), .ZN(MULT_mult_6_net81373) );
  INV_X4 MULT_mult_6_U402 ( .A(MULT_mult_6_CARRYB_8__12_), .ZN(
        MULT_mult_6_net84868) );
  NAND2_X2 MULT_mult_6_U350 ( .A1(MULT_mult_6_net81070), .A2(MULT_mult_6_n193), 
        .ZN(MULT_mult_6_n486) );
  NAND2_X2 MULT_mult_6_U330 ( .A1(MULT_mult_6_net85044), .A2(
        MULT_mult_6_net88455), .ZN(MULT_mult_6_n2117) );
  INV_X2 MULT_mult_6_U309 ( .A(MULT_mult_6_n2358), .ZN(MULT_mult_6_n2359) );
  INV_X1 MULT_mult_6_U290 ( .A(MULT_mult_6_CARRYB_1__16_), .ZN(
        MULT_mult_6_n2358) );
  INV_X2 MULT_mult_6_U287 ( .A(MULT_mult_6_n565), .ZN(MULT_mult_6_net85399) );
  NAND2_X2 MULT_mult_6_U262 ( .A1(MULT_mult_6_net121452), .A2(
        MULT_mult_6_net121451), .ZN(MULT_mult_6_n193) );
  XOR2_X2 MULT_mult_6_U253 ( .A(MULT_mult_6_ab_1__24_), .B(
        MULT_mult_6_ab_0__25_), .Z(MULT_mult_6_n2357) );
  NAND2_X2 MULT_mult_6_U236 ( .A1(MULT_mult_6_CARRYB_27__2_), .A2(
        MULT_mult_6_ab_28__2_), .ZN(MULT_mult_6_n115) );
  INV_X8 MULT_mult_6_U217 ( .A(MULT_mult_6_CARRYB_26__2_), .ZN(
        MULT_mult_6_net83054) );
  NAND2_X2 MULT_mult_6_U178 ( .A1(MULT_mult_6_CARRYB_3__13_), .A2(
        MULT_mult_6_n212), .ZN(MULT_mult_6_n213) );
  NAND2_X4 MULT_mult_6_U177 ( .A1(MULT_mult_6_n214), .A2(MULT_mult_6_n213), 
        .ZN(MULT_mult_6_n857) );
  INV_X2 MULT_mult_6_U160 ( .A(MULT_mult_6_SUMB_3__14_), .ZN(MULT_mult_6_n910)
         );
  INV_X4 MULT_mult_6_U148 ( .A(MULT_mult_6_n939), .ZN(MULT_mult_6_n221) );
  XNOR2_X2 MULT_mult_6_U140 ( .A(MULT_mult_6_n2001), .B(MULT_mult_6_n221), 
        .ZN(MULT_mult_6_n1261) );
  INV_X2 MULT_mult_6_U105 ( .A(MULT_mult_6_net89104), .ZN(MULT_mult_6_n582) );
  INV_X4 MULT_mult_6_U67 ( .A(MULT_mult_6_n476), .ZN(MULT_mult_6_n12) );
  NAND2_X2 MULT_mult_6_U65 ( .A1(MULT_mult_6_net123363), .A2(
        MULT_mult_6_ab_28__1_), .ZN(MULT_mult_6_net79880) );
  INV_X2 MULT_mult_6_U40 ( .A(MULT_mult_6_net83054), .ZN(MULT_mult_6_n2356) );
  NAND2_X2 MULT_mult_6_U35 ( .A1(MULT_mult_6_net91001), .A2(
        MULT_mult_6_net88699), .ZN(MULT_mult_6_net80673) );
  NAND3_X4 MULT_mult_6_U30 ( .A1(MULT_mult_6_net80673), .A2(
        MULT_mult_6_net80672), .A3(MULT_mult_6_net80671), .ZN(
        MULT_mult_6_CARRYB_20__7_) );
  NAND2_X2 MULT_mult_6_U29 ( .A1(MULT_mult_6_net119817), .A2(
        MULT_mult_6_CARRYB_3__14_), .ZN(MULT_mult_6_n529) );
  NAND2_X2 MULT_mult_6_U17 ( .A1(MULT_mult_6_n581), .A2(MULT_mult_6_n582), 
        .ZN(MULT_mult_6_n584) );
  NOR2_X1 MULT_mult_6_U15 ( .A1(MULT_mult_6_n348), .A2(MULT_mult_6_net92311), 
        .ZN(MULT_mult_6_n1181) );
  INV_X4 MULT_mult_6_U4857 ( .A(MULT_mult_6_net70435), .ZN(multOut[31]) );
  NOR2_X4 MULT_mult_6_U4856 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70443), .ZN(MULT_mult_6_ab_26__3_) );
  NOR2_X4 MULT_mult_6_U4855 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70447), .ZN(MULT_mult_6_ab_24__2_) );
  NOR2_X4 MULT_mult_6_U4854 ( .A1(MULT_mult_6_net77906), .A2(
        MULT_mult_6_net70447), .ZN(MULT_mult_6_ab_24__6_) );
  NOR2_X4 MULT_mult_6_U4853 ( .A1(MULT_mult_6_net77858), .A2(
        MULT_mult_6_net70449), .ZN(MULT_mult_6_ab_23__0_) );
  NOR2_X4 MULT_mult_6_U4852 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70449), .ZN(MULT_mult_6_ab_23__2_) );
  NOR2_X4 MULT_mult_6_U4851 ( .A1(MULT_mult_6_net77900), .A2(
        MULT_mult_6_net70449), .ZN(MULT_mult_6_ab_23__5_) );
  NOR2_X4 MULT_mult_6_U4850 ( .A1(MULT_mult_6_net77908), .A2(
        MULT_mult_6_net70449), .ZN(MULT_mult_6_ab_23__6_) );
  NOR2_X4 MULT_mult_6_U4849 ( .A1(MULT_mult_6_net77858), .A2(
        MULT_mult_6_net70451), .ZN(MULT_mult_6_ab_22__0_) );
  NOR2_X4 MULT_mult_6_U4848 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70451), .ZN(MULT_mult_6_ab_22__4_) );
  NOR2_X4 MULT_mult_6_U4847 ( .A1(MULT_mult_6_net77908), .A2(
        MULT_mult_6_net70451), .ZN(MULT_mult_6_ab_22__6_) );
  NOR2_X4 MULT_mult_6_U4846 ( .A1(MULT_mult_6_net77868), .A2(
        MULT_mult_6_net70453), .ZN(MULT_mult_6_ab_21__1_) );
  NOR2_X4 MULT_mult_6_U4845 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70453), .ZN(MULT_mult_6_ab_21__3_) );
  NOR2_X4 MULT_mult_6_U4844 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70453), .ZN(MULT_mult_6_ab_21__4_) );
  NOR2_X4 MULT_mult_6_U4843 ( .A1(MULT_mult_6_net77858), .A2(
        MULT_mult_6_net70455), .ZN(MULT_mult_6_ab_20__0_) );
  NOR2_X4 MULT_mult_6_U4842 ( .A1(MULT_mult_6_net77868), .A2(
        MULT_mult_6_net70455), .ZN(MULT_mult_6_ab_20__1_) );
  NOR2_X4 MULT_mult_6_U4841 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70455), .ZN(MULT_mult_6_ab_20__2_) );
  NOR2_X4 MULT_mult_6_U4840 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70455), .ZN(MULT_mult_6_ab_20__4_) );
  NOR2_X4 MULT_mult_6_U4839 ( .A1(MULT_mult_6_net77914), .A2(
        MULT_mult_6_net70455), .ZN(MULT_mult_6_ab_20__7_) );
  NOR2_X4 MULT_mult_6_U4838 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net70455), .ZN(MULT_mult_6_ab_20__8_) );
  NOR2_X4 MULT_mult_6_U4837 ( .A1(MULT_mult_6_net77858), .A2(
        MULT_mult_6_net70457), .ZN(MULT_mult_6_ab_19__0_) );
  NOR2_X4 MULT_mult_6_U4836 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70457), .ZN(MULT_mult_6_ab_19__2_) );
  NOR2_X4 MULT_mult_6_U4835 ( .A1(MULT_mult_6_net77900), .A2(
        MULT_mult_6_net70457), .ZN(MULT_mult_6_ab_19__5_) );
  NOR2_X4 MULT_mult_6_U4834 ( .A1(MULT_mult_6_net77914), .A2(
        MULT_mult_6_net70457), .ZN(MULT_mult_6_ab_19__7_) );
  NOR2_X4 MULT_mult_6_U4833 ( .A1(MULT_mult_6_net77860), .A2(
        MULT_mult_6_net70459), .ZN(MULT_mult_6_ab_18__0_) );
  NOR2_X4 MULT_mult_6_U4832 ( .A1(MULT_mult_6_net77868), .A2(
        MULT_mult_6_net70459), .ZN(MULT_mult_6_ab_18__1_) );
  NOR2_X4 MULT_mult_6_U4831 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70459), .ZN(MULT_mult_6_ab_18__2_) );
  NOR2_X4 MULT_mult_6_U4830 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70459), .ZN(MULT_mult_6_ab_18__4_) );
  NOR2_X4 MULT_mult_6_U4829 ( .A1(MULT_mult_6_net77900), .A2(
        MULT_mult_6_net70459), .ZN(MULT_mult_6_ab_18__5_) );
  NOR2_X4 MULT_mult_6_U4828 ( .A1(MULT_mult_6_net77860), .A2(
        MULT_mult_6_net70461), .ZN(MULT_mult_6_ab_17__0_) );
  NOR2_X4 MULT_mult_6_U4827 ( .A1(MULT_mult_6_net77868), .A2(
        MULT_mult_6_net70461), .ZN(MULT_mult_6_ab_17__1_) );
  NOR2_X4 MULT_mult_6_U4826 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70461), .ZN(MULT_mult_6_ab_17__2_) );
  NOR2_X4 MULT_mult_6_U4825 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70461), .ZN(MULT_mult_6_ab_17__3_) );
  NOR2_X4 MULT_mult_6_U4824 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70461), .ZN(MULT_mult_6_ab_17__4_) );
  NOR2_X4 MULT_mult_6_U4823 ( .A1(MULT_mult_6_net77900), .A2(
        MULT_mult_6_net70461), .ZN(MULT_mult_6_ab_17__5_) );
  NOR2_X4 MULT_mult_6_U4822 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net70461), .ZN(MULT_mult_6_ab_17__8_) );
  NOR2_X4 MULT_mult_6_U4821 ( .A1(MULT_mult_6_net77860), .A2(
        MULT_mult_6_net70463), .ZN(MULT_mult_6_ab_16__0_) );
  NOR2_X4 MULT_mult_6_U4820 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70463), .ZN(MULT_mult_6_ab_16__2_) );
  NOR2_X4 MULT_mult_6_U4819 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70463), .ZN(MULT_mult_6_ab_16__3_) );
  NOR2_X4 MULT_mult_6_U4818 ( .A1(MULT_mult_6_net77900), .A2(
        MULT_mult_6_net70463), .ZN(MULT_mult_6_ab_16__5_) );
  NOR2_X4 MULT_mult_6_U4817 ( .A1(MULT_mult_6_net77908), .A2(
        MULT_mult_6_net70463), .ZN(MULT_mult_6_ab_16__6_) );
  NOR2_X4 MULT_mult_6_U4816 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net70463), .ZN(MULT_mult_6_ab_16__8_) );
  NOR2_X4 MULT_mult_6_U4815 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__2_) );
  NOR2_X4 MULT_mult_6_U4814 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__4_) );
  NOR2_X4 MULT_mult_6_U4813 ( .A1(MULT_mult_6_net77900), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__5_) );
  NOR2_X4 MULT_mult_6_U4812 ( .A1(MULT_mult_6_net77914), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__7_) );
  NOR2_X4 MULT_mult_6_U4811 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__8_) );
  NOR2_X4 MULT_mult_6_U4810 ( .A1(MULT_mult_6_net77868), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__1_) );
  NOR2_X4 MULT_mult_6_U4809 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__3_) );
  NOR2_X4 MULT_mult_6_U4808 ( .A1(MULT_mult_6_net77900), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__5_) );
  NOR2_X4 MULT_mult_6_U4807 ( .A1(MULT_mult_6_net77900), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__5_) );
  NOR2_X4 MULT_mult_6_U4806 ( .A1(MULT_mult_6_net77860), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__0_) );
  NOR2_X4 MULT_mult_6_U4805 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__3_) );
  NOR2_X4 MULT_mult_6_U4804 ( .A1(MULT_mult_6_net77900), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__5_) );
  NOR2_X4 MULT_mult_6_U4803 ( .A1(MULT_mult_6_net77908), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__6_) );
  NOR2_X4 MULT_mult_6_U4802 ( .A1(MULT_mult_6_net77860), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__0_) );
  NOR2_X4 MULT_mult_6_U4801 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__3_) );
  NOR2_X4 MULT_mult_6_U4800 ( .A1(MULT_mult_6_net77866), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__1_) );
  NOR2_X4 MULT_mult_6_U4799 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__3_) );
  NOR2_X4 MULT_mult_6_U4798 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__4_) );
  NOR2_X4 MULT_mult_6_U4797 ( .A1(MULT_mult_6_net81424), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__15_) );
  NOR2_X4 MULT_mult_6_U4796 ( .A1(MULT_mult_6_net80727), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__20_) );
  NOR2_X4 MULT_mult_6_U4795 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__2_) );
  NOR2_X4 MULT_mult_6_U4794 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__3_) );
  NOR2_X4 MULT_mult_6_U4793 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__4_) );
  NOR2_X4 MULT_mult_6_U4792 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__8_) );
  NOR2_X4 MULT_mult_6_U4791 ( .A1(MULT_mult_6_net80727), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__20_) );
  NOR2_X4 MULT_mult_6_U4790 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net77924), .ZN(MULT_mult_6_ab_8__8_) );
  NOR2_X4 MULT_mult_6_U4789 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net77926), .ZN(MULT_mult_6_ab_8__13_) );
  NOR2_X4 MULT_mult_6_U4788 ( .A1(MULT_mult_6_net80727), .A2(
        MULT_mult_6_net77926), .ZN(MULT_mult_6_ab_8__20_) );
  NOR2_X4 MULT_mult_6_U4787 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net77930), .ZN(MULT_mult_6_ab_7__3_) );
  NOR2_X4 MULT_mult_6_U4786 ( .A1(MULT_mult_6_net77906), .A2(
        MULT_mult_6_net77930), .ZN(MULT_mult_6_ab_7__6_) );
  NOR2_X4 MULT_mult_6_U4785 ( .A1(MULT_mult_6_net77912), .A2(
        MULT_mult_6_net77930), .ZN(MULT_mult_6_ab_7__7_) );
  NOR2_X4 MULT_mult_6_U4784 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net77930), .ZN(MULT_mult_6_ab_7__9_) );
  NOR2_X4 MULT_mult_6_U4783 ( .A1(MULT_mult_6_net123000), .A2(
        MULT_mult_6_net77932), .ZN(MULT_mult_6_ab_7__17_) );
  NOR2_X4 MULT_mult_6_U4782 ( .A1(MULT_mult_6_net77860), .A2(
        MULT_mult_6_net77938), .ZN(MULT_mult_6_ab_6__0_) );
  NOR2_X4 MULT_mult_6_U4781 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net77938), .ZN(MULT_mult_6_ab_6__2_) );
  NOR2_X4 MULT_mult_6_U4780 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net77938), .ZN(MULT_mult_6_ab_6__4_) );
  NOR2_X4 MULT_mult_6_U4779 ( .A1(MULT_mult_6_net77912), .A2(
        MULT_mult_6_net77938), .ZN(MULT_mult_6_ab_6__7_) );
  NOR2_X4 MULT_mult_6_U4778 ( .A1(MULT_mult_6_net81424), .A2(
        MULT_mult_6_net77940), .ZN(MULT_mult_6_ab_6__15_) );
  NOR2_X4 MULT_mult_6_U4777 ( .A1(MULT_mult_6_net77866), .A2(
        MULT_mult_6_net77946), .ZN(MULT_mult_6_ab_5__1_) );
  NOR2_X4 MULT_mult_6_U4776 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net77946), .ZN(MULT_mult_6_ab_5__8_) );
  NOR2_X4 MULT_mult_6_U4775 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net119855), .ZN(MULT_mult_6_ab_4__2_) );
  NOR2_X4 MULT_mult_6_U4774 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net77956), .ZN(MULT_mult_6_ab_4__3_) );
  NOR2_X4 MULT_mult_6_U4773 ( .A1(MULT_mult_6_net77906), .A2(
        MULT_mult_6_net119855), .ZN(MULT_mult_6_ab_4__6_) );
  NOR2_X4 MULT_mult_6_U4772 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net119855), .ZN(MULT_mult_6_ab_4__8_) );
  NOR2_X4 MULT_mult_6_U4771 ( .A1(MULT_mult_6_net77906), .A2(
        MULT_mult_6_net77966), .ZN(MULT_mult_6_ab_3__6_) );
  NOR2_X4 MULT_mult_6_U4770 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net77966), .ZN(MULT_mult_6_ab_3__8_) );
  NOR2_X4 MULT_mult_6_U4769 ( .A1(MULT_mult_6_net82890), .A2(
        MULT_mult_6_net77964), .ZN(MULT_mult_6_ab_3__17_) );
  NOR2_X4 MULT_mult_6_U4768 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net77970), .ZN(MULT_mult_6_ab_2__8_) );
  NOR2_X4 MULT_mult_6_U4767 ( .A1(MULT_mult_6_net81673), .A2(
        MULT_mult_6_net77878), .ZN(MULT_mult_6_ab_0__2_) );
  NOR2_X4 MULT_mult_6_U4766 ( .A1(MULT_mult_6_net77882), .A2(
        MULT_mult_6_net83263), .ZN(MULT_mult_6_ab_1__3_) );
  NOR2_X4 MULT_mult_6_U4765 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net83263), .ZN(MULT_mult_6_ab_1__4_) );
  NOR2_X4 MULT_mult_6_U4764 ( .A1(MULT_mult_6_net81673), .A2(
        MULT_mult_6_net77898), .ZN(MULT_mult_6_ab_0__5_) );
  NOR2_X4 MULT_mult_6_U4763 ( .A1(MULT_mult_6_net70476), .A2(
        MULT_mult_6_net82149), .ZN(MULT_mult_6_ab_0__21_) );
  AND2_X2 MULT_mult_6_U4762 ( .A1(net36488), .A2(MULT_mult_6_net80392), .ZN(
        MULT_mult_6_ab_0__31_) );
  INV_X4 MULT_mult_6_U4761 ( .A(MULT_mult_6_n2352), .ZN(
        MULT_mult_6_SUMB_1__29_) );
  XNOR2_X2 MULT_mult_6_U4760 ( .A(MULT_mult_6_ab_1__29_), .B(
        MULT_mult_6_ab_0__30_), .ZN(MULT_mult_6_n2352) );
  INV_X4 MULT_mult_6_U4759 ( .A(MULT_mult_6_n2351), .ZN(
        MULT_mult_6_SUMB_1__28_) );
  XNOR2_X2 MULT_mult_6_U4758 ( .A(MULT_mult_6_ab_1__28_), .B(
        MULT_mult_6_ab_0__29_), .ZN(MULT_mult_6_n2351) );
  INV_X4 MULT_mult_6_U4757 ( .A(MULT_mult_6_n2350), .ZN(
        MULT_mult_6_SUMB_1__27_) );
  INV_X4 MULT_mult_6_U4756 ( .A(MULT_mult_6_n2349), .ZN(
        MULT_mult_6_SUMB_1__26_) );
  XNOR2_X2 MULT_mult_6_U4755 ( .A(MULT_mult_6_ab_1__26_), .B(
        MULT_mult_6_ab_0__27_), .ZN(MULT_mult_6_n2349) );
  INV_X4 MULT_mult_6_U4754 ( .A(MULT_mult_6_n2348), .ZN(
        MULT_mult_6_CARRYB_1__26_) );
  NAND2_X2 MULT_mult_6_U4753 ( .A1(MULT_mult_6_ab_0__27_), .A2(
        MULT_mult_6_ab_1__26_), .ZN(MULT_mult_6_n2348) );
  INV_X4 MULT_mult_6_U4752 ( .A(MULT_mult_6_n2347), .ZN(
        MULT_mult_6_SUMB_1__23_) );
  XNOR2_X2 MULT_mult_6_U4751 ( .A(MULT_mult_6_n2196), .B(MULT_mult_6_ab_0__23_), .ZN(MULT_mult_6_n2346) );
  XNOR2_X2 MULT_mult_6_U4750 ( .A(MULT_mult_6_ab_0__22_), .B(
        MULT_mult_6_ab_1__21_), .ZN(MULT_mult_6_n2344) );
  XNOR2_X2 MULT_mult_6_U4749 ( .A(MULT_mult_6_ab_1__20_), .B(
        MULT_mult_6_ab_0__21_), .ZN(MULT_mult_6_n2342) );
  XNOR2_X2 MULT_mult_6_U4748 ( .A(MULT_mult_6_ab_1__19_), .B(
        MULT_mult_6_ab_0__20_), .ZN(MULT_mult_6_n2340) );
  XNOR2_X2 MULT_mult_6_U4747 ( .A(MULT_mult_6_n237), .B(MULT_mult_6_ab_0__13_), 
        .ZN(MULT_mult_6_n2337) );
  INV_X4 MULT_mult_6_U4746 ( .A(MULT_mult_6_n2336), .ZN(
        MULT_mult_6_CARRYB_1__12_) );
  INV_X4 MULT_mult_6_U4745 ( .A(MULT_mult_6_n2333), .ZN(
        MULT_mult_6_SUMB_1__10_) );
  XNOR2_X2 MULT_mult_6_U4744 ( .A(MULT_mult_6_ab_1__10_), .B(
        MULT_mult_6_ab_0__11_), .ZN(MULT_mult_6_n2333) );
  INV_X4 MULT_mult_6_U4743 ( .A(MULT_mult_6_n2331), .ZN(MULT_mult_6_SUMB_1__9_) );
  INV_X4 MULT_mult_6_U4742 ( .A(MULT_mult_6_n1517), .ZN(
        MULT_mult_6_CARRYB_1__9_) );
  INV_X4 MULT_mult_6_U4741 ( .A(MULT_mult_6__UDW__112739_net78703), .ZN(
        MULT_mult_6_SUMB_1__6_) );
  INV_X4 MULT_mult_6_U4740 ( .A(MULT_mult_6_n2330), .ZN(MULT_mult_6_SUMB_1__5_) );
  XNOR2_X2 MULT_mult_6_U4739 ( .A(MULT_mult_6_ab_1__5_), .B(
        MULT_mult_6_ab_0__6_), .ZN(MULT_mult_6_n2330) );
  INV_X4 MULT_mult_6_U4738 ( .A(MULT_mult_6_n2328), .ZN(MULT_mult_6_SUMB_1__4_) );
  INV_X4 MULT_mult_6_U4737 ( .A(MULT_mult_6_n2326), .ZN(MULT_mult_6_SUMB_1__3_) );
  XNOR2_X2 MULT_mult_6_U4736 ( .A(MULT_mult_6_ab_1__3_), .B(MULT_mult_6_n870), 
        .ZN(MULT_mult_6_n2326) );
  NAND2_X2 MULT_mult_6_U4735 ( .A1(MULT_mult_6_n870), .A2(MULT_mult_6_ab_1__3_), .ZN(MULT_mult_6_n2325) );
  INV_X4 MULT_mult_6_U4734 ( .A(MULT_mult_6_n2324), .ZN(MULT_mult_6_SUMB_1__2_) );
  INV_X4 MULT_mult_6_U4733 ( .A(MULT_mult_6_n2323), .ZN(
        MULT_mult_6_CARRYB_1__2_) );
  NAND2_X2 MULT_mult_6_U4732 ( .A1(MULT_mult_6_ab_0__3_), .A2(
        MULT_mult_6_ab_1__2_), .ZN(MULT_mult_6_n2323) );
  INV_X4 MULT_mult_6_U4731 ( .A(MULT_mult_6_n2322), .ZN(
        MULT_mult_6_CARRYB_1__0_) );
  NAND2_X2 MULT_mult_6_U4730 ( .A1(MULT_mult_6_ab_0__1_), .A2(
        MULT_mult_6_ab_1__0_), .ZN(MULT_mult_6_n2322) );
  NOR2_X1 MULT_mult_6_U4729 ( .A1(MULT_mult_6_net70475), .A2(
        MULT_mult_6_net80643), .ZN(MULT_mult_6_ab_10__21_) );
  NOR2_X1 MULT_mult_6_U4728 ( .A1(MULT_mult_6_net77956), .A2(MULT_mult_6_n2355), .ZN(MULT_mult_6_ab_4__27_) );
  NOR2_X1 MULT_mult_6_U4727 ( .A1(MULT_mult_6_net70463), .A2(
        MULT_mult_6_net81424), .ZN(MULT_mult_6_ab_16__15_) );
  NOR2_X1 MULT_mult_6_U4726 ( .A1(MULT_mult_6_net70473), .A2(
        MULT_mult_6_net80727), .ZN(MULT_mult_6_ab_11__20_) );
  XOR2_X2 MULT_mult_6_U4725 ( .A(MULT_mult_6_CARRYB_9__21_), .B(
        MULT_mult_6_ab_10__21_), .Z(MULT_mult_6_n2321) );
  XOR2_X2 MULT_mult_6_U4724 ( .A(MULT_mult_6_SUMB_3__28_), .B(
        MULT_mult_6_n2320), .Z(MULT_mult_6_SUMB_4__27_) );
  XOR2_X2 MULT_mult_6_U4723 ( .A(MULT_mult_6_CARRYB_3__27_), .B(
        MULT_mult_6_ab_4__27_), .Z(MULT_mult_6_n2320) );
  XOR2_X2 MULT_mult_6_U4722 ( .A(MULT_mult_6_SUMB_10__21_), .B(
        MULT_mult_6_n2319), .Z(MULT_mult_6_SUMB_11__20_) );
  XOR2_X2 MULT_mult_6_U4721 ( .A(MULT_mult_6_CARRYB_10__20_), .B(
        MULT_mult_6_ab_11__20_), .Z(MULT_mult_6_n2319) );
  NOR2_X1 MULT_mult_6_U4720 ( .A1(MULT_mult_6_net124723), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__16_) );
  NAND3_X2 MULT_mult_6_U4719 ( .A1(MULT_mult_6_n2316), .A2(MULT_mult_6_n2317), 
        .A3(MULT_mult_6_n2318), .ZN(MULT_mult_6_CARRYB_13__16_) );
  NAND2_X1 MULT_mult_6_U4718 ( .A1(MULT_mult_6_ab_13__16_), .A2(
        MULT_mult_6_CARRYB_12__16_), .ZN(MULT_mult_6_n2318) );
  NAND2_X1 MULT_mult_6_U4717 ( .A1(MULT_mult_6_CARRYB_12__16_), .A2(
        MULT_mult_6_SUMB_12__17_), .ZN(MULT_mult_6_n2316) );
  NAND3_X2 MULT_mult_6_U4716 ( .A1(MULT_mult_6_n2313), .A2(MULT_mult_6_n2314), 
        .A3(MULT_mult_6_n2315), .ZN(MULT_mult_6_CARRYB_4__24_) );
  NAND2_X1 MULT_mult_6_U4715 ( .A1(MULT_mult_6_CARRYB_3__24_), .A2(
        MULT_mult_6_SUMB_3__25_), .ZN(MULT_mult_6_n2315) );
  NAND2_X1 MULT_mult_6_U4714 ( .A1(MULT_mult_6_ab_4__24_), .A2(
        MULT_mult_6_SUMB_3__25_), .ZN(MULT_mult_6_n2314) );
  NAND2_X1 MULT_mult_6_U4713 ( .A1(MULT_mult_6_ab_4__24_), .A2(
        MULT_mult_6_CARRYB_3__24_), .ZN(MULT_mult_6_n2313) );
  NAND3_X2 MULT_mult_6_U4712 ( .A1(MULT_mult_6_n2310), .A2(MULT_mult_6_n2311), 
        .A3(MULT_mult_6_n2312), .ZN(MULT_mult_6_CARRYB_3__25_) );
  NAND2_X2 MULT_mult_6_U4711 ( .A1(MULT_mult_6_n1219), .A2(
        MULT_mult_6_CARRYB_2__25_), .ZN(MULT_mult_6_n2312) );
  NAND2_X2 MULT_mult_6_U4710 ( .A1(MULT_mult_6_n1219), .A2(
        MULT_mult_6_ab_3__25_), .ZN(MULT_mult_6_n2311) );
  NAND2_X1 MULT_mult_6_U4709 ( .A1(MULT_mult_6_ab_3__25_), .A2(
        MULT_mult_6_CARRYB_2__25_), .ZN(MULT_mult_6_n2310) );
  NAND2_X1 MULT_mult_6_U4708 ( .A1(MULT_mult_6_ab_12__16_), .A2(
        MULT_mult_6_CARRYB_11__16_), .ZN(MULT_mult_6_n2307) );
  NOR2_X1 MULT_mult_6_U4707 ( .A1(MULT_mult_6_net80727), .A2(
        MULT_mult_6_net77940), .ZN(MULT_mult_6_ab_6__20_) );
  NOR2_X1 MULT_mult_6_U4706 ( .A1(MULT_mult_6_net80727), .A2(
        MULT_mult_6_net77932), .ZN(MULT_mult_6_ab_7__20_) );
  NAND3_X2 MULT_mult_6_U4705 ( .A1(MULT_mult_6_net79959), .A2(
        MULT_mult_6_net79960), .A3(MULT_mult_6_net79961), .ZN(
        MULT_mult_6_CARRYB_7__20_) );
  NAND3_X2 MULT_mult_6_U4704 ( .A1(MULT_mult_6_net79955), .A2(
        MULT_mult_6_net79956), .A3(MULT_mult_6_net79957), .ZN(
        MULT_mult_6_CARRYB_8__19_) );
  NAND3_X2 MULT_mult_6_U4703 ( .A1(MULT_mult_6_net79951), .A2(
        MULT_mult_6_net79952), .A3(MULT_mult_6_net79953), .ZN(
        MULT_mult_6_CARRYB_9__18_) );
  NAND2_X1 MULT_mult_6_U4702 ( .A1(MULT_mult_6_ab_9__16_), .A2(
        MULT_mult_6_CARRYB_8__16_), .ZN(MULT_mult_6_n2306) );
  NOR2_X1 MULT_mult_6_U4701 ( .A1(MULT_mult_6_n175), .A2(MULT_mult_6_net70492), 
        .ZN(MULT_mult_6_ab_2__29_) );
  XNOR2_X2 MULT_mult_6_U4700 ( .A(MULT_mult_6_ab_1__27_), .B(
        MULT_mult_6_ab_0__28_), .ZN(MULT_mult_6_n2350) );
  NOR2_X1 MULT_mult_6_U4699 ( .A1(MULT_mult_6_net84698), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__14_) );
  NAND2_X2 MULT_mult_6_U4698 ( .A1(MULT_mult_6_CARRYB_8__19_), .A2(
        MULT_mult_6_SUMB_8__20_), .ZN(MULT_mult_6_n2291) );
  NAND2_X1 MULT_mult_6_U4697 ( .A1(MULT_mult_6_ab_9__19_), .A2(
        MULT_mult_6_CARRYB_8__19_), .ZN(MULT_mult_6_n2289) );
  NAND2_X2 MULT_mult_6_U4696 ( .A1(MULT_mult_6_n851), .A2(
        MULT_mult_6_CARRYB_7__20_), .ZN(MULT_mult_6_n2288) );
  NAND2_X2 MULT_mult_6_U4695 ( .A1(MULT_mult_6_n851), .A2(
        MULT_mult_6_ab_8__20_), .ZN(MULT_mult_6_n2287) );
  NAND2_X1 MULT_mult_6_U4694 ( .A1(MULT_mult_6_ab_8__20_), .A2(
        MULT_mult_6_CARRYB_7__20_), .ZN(MULT_mult_6_n2286) );
  NAND3_X2 MULT_mult_6_U4693 ( .A1(MULT_mult_6_net80273), .A2(
        MULT_mult_6_net80274), .A3(MULT_mult_6_net80275), .ZN(
        MULT_mult_6_CARRYB_16__13_) );
  NAND2_X1 MULT_mult_6_U4692 ( .A1(MULT_mult_6_ab_23__6_), .A2(
        MULT_mult_6_n351), .ZN(MULT_mult_6_n2283) );
  NOR2_X1 MULT_mult_6_U4691 ( .A1(MULT_mult_6_n955), .A2(MULT_mult_6_net77956), 
        .ZN(MULT_mult_6_ab_4__21_) );
  NAND2_X1 MULT_mult_6_U4690 ( .A1(MULT_mult_6_ab_6__19_), .A2(MULT_mult_6_n56), .ZN(MULT_mult_6_n2279) );
  NAND2_X1 MULT_mult_6_U4689 ( .A1(MULT_mult_6_ab_4__21_), .A2(
        MULT_mult_6_CARRYB_3__21_), .ZN(MULT_mult_6_n2278) );
  INV_X8 MULT_mult_6_U4688 ( .A(n10907), .ZN(MULT_mult_6_net70492) );
  NOR2_X2 MULT_mult_6_U4687 ( .A1(MULT_mult_6_net77966), .A2(MULT_mult_6_n2354), .ZN(MULT_mult_6_ab_3__28_) );
  NOR2_X1 MULT_mult_6_U4686 ( .A1(MULT_mult_6_n2355), .A2(MULT_mult_6_net77966), .ZN(MULT_mult_6_ab_3__27_) );
  NOR2_X1 MULT_mult_6_U4685 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70457), .ZN(MULT_mult_6_ab_19__3_) );
  NAND3_X2 MULT_mult_6_U4684 ( .A1(MULT_mult_6_n2273), .A2(MULT_mult_6_n2274), 
        .A3(MULT_mult_6_n2275), .ZN(MULT_mult_6_CARRYB_19__3_) );
  NAND2_X2 MULT_mult_6_U4683 ( .A1(MULT_mult_6_SUMB_18__4_), .A2(
        MULT_mult_6_ab_19__3_), .ZN(MULT_mult_6_n2274) );
  NAND3_X2 MULT_mult_6_U4682 ( .A1(MULT_mult_6_n2272), .A2(
        MULT_mult_6_net80356), .A3(MULT_mult_6_net80355), .ZN(
        MULT_mult_6_CARRYB_8__14_) );
  INV_X8 MULT_mult_6_U4681 ( .A(n10908), .ZN(MULT_mult_6_n2354) );
  NOR2_X1 MULT_mult_6_U4680 ( .A1(MULT_mult_6_n242), .A2(MULT_mult_6_n2353), 
        .ZN(MULT_mult_6_ab_1__30_) );
  NAND3_X2 MULT_mult_6_U4679 ( .A1(MULT_mult_6_n2269), .A2(MULT_mult_6_n2270), 
        .A3(MULT_mult_6_n2271), .ZN(MULT_mult_6_CARRYB_8__22_) );
  NAND2_X1 MULT_mult_6_U4678 ( .A1(MULT_mult_6_CARRYB_7__22_), .A2(
        MULT_mult_6_SUMB_7__23_), .ZN(MULT_mult_6_n2271) );
  NAND2_X1 MULT_mult_6_U4677 ( .A1(MULT_mult_6_ab_8__22_), .A2(
        MULT_mult_6_SUMB_7__23_), .ZN(MULT_mult_6_n2270) );
  NAND2_X1 MULT_mult_6_U4676 ( .A1(MULT_mult_6_ab_8__22_), .A2(
        MULT_mult_6_CARRYB_7__22_), .ZN(MULT_mult_6_n2269) );
  NAND2_X1 MULT_mult_6_U4675 ( .A1(MULT_mult_6_ab_7__23_), .A2(
        MULT_mult_6_CARRYB_6__23_), .ZN(MULT_mult_6_n2266) );
  NAND3_X2 MULT_mult_6_U4674 ( .A1(MULT_mult_6_n2263), .A2(MULT_mult_6_n2264), 
        .A3(MULT_mult_6_n2265), .ZN(MULT_mult_6_CARRYB_3__27_) );
  NAND2_X1 MULT_mult_6_U4673 ( .A1(MULT_mult_6_CARRYB_2__27_), .A2(
        MULT_mult_6_SUMB_2__28_), .ZN(MULT_mult_6_n2265) );
  NAND2_X1 MULT_mult_6_U4672 ( .A1(MULT_mult_6_ab_3__27_), .A2(
        MULT_mult_6_SUMB_2__28_), .ZN(MULT_mult_6_n2264) );
  NAND2_X1 MULT_mult_6_U4671 ( .A1(MULT_mult_6_ab_3__27_), .A2(
        MULT_mult_6_CARRYB_2__27_), .ZN(MULT_mult_6_n2263) );
  NAND2_X2 MULT_mult_6_U4670 ( .A1(MULT_mult_6_n347), .A2(
        MULT_mult_6_SUMB_1__29_), .ZN(MULT_mult_6_n2262) );
  NAND2_X2 MULT_mult_6_U4669 ( .A1(MULT_mult_6_ab_2__28_), .A2(
        MULT_mult_6_SUMB_1__29_), .ZN(MULT_mult_6_n2261) );
  NAND2_X2 MULT_mult_6_U4668 ( .A1(MULT_mult_6_ab_2__28_), .A2(
        MULT_mult_6_n347), .ZN(MULT_mult_6_n2260) );
  XOR2_X2 MULT_mult_6_U4667 ( .A(MULT_mult_6_n2259), .B(
        MULT_mult_6_SUMB_1__29_), .Z(MULT_mult_6_SUMB_2__28_) );
  XOR2_X2 MULT_mult_6_U4666 ( .A(MULT_mult_6_ab_2__28_), .B(MULT_mult_6_n347), 
        .Z(MULT_mult_6_n2259) );
  NAND2_X1 MULT_mult_6_U4665 ( .A1(MULT_mult_6_ab_19__11_), .A2(
        MULT_mult_6_CARRYB_18__11_), .ZN(MULT_mult_6_n2256) );
  NAND3_X2 MULT_mult_6_U4664 ( .A1(MULT_mult_6_net80449), .A2(
        MULT_mult_6_n2255), .A3(MULT_mult_6_net80451), .ZN(
        MULT_mult_6_CARRYB_18__12_) );
  NAND2_X2 MULT_mult_6_U4663 ( .A1(MULT_mult_6_ab_8__15_), .A2(
        MULT_mult_6_SUMB_7__16_), .ZN(MULT_mult_6_n2253) );
  NAND3_X4 MULT_mult_6_U4662 ( .A1(MULT_mult_6_n2251), .A2(MULT_mult_6_n2250), 
        .A3(MULT_mult_6_n2249), .ZN(MULT_mult_6_CARRYB_7__16_) );
  NAND2_X1 MULT_mult_6_U4661 ( .A1(MULT_mult_6_ab_5__19_), .A2(
        MULT_mult_6_CARRYB_4__19_), .ZN(MULT_mult_6_n2240) );
  NAND2_X1 MULT_mult_6_U4660 ( .A1(MULT_mult_6_ab_4__20_), .A2(
        MULT_mult_6_CARRYB_3__20_), .ZN(MULT_mult_6_n2237) );
  NAND3_X2 MULT_mult_6_U4659 ( .A1(MULT_mult_6_net80521), .A2(
        MULT_mult_6_net80522), .A3(MULT_mult_6_net80523), .ZN(
        MULT_mult_6_CARRYB_11__16_) );
  NAND3_X2 MULT_mult_6_U4658 ( .A1(MULT_mult_6_net80518), .A2(
        MULT_mult_6_net80519), .A3(MULT_mult_6_net80520), .ZN(
        MULT_mult_6_CARRYB_10__17_) );
  NAND3_X2 MULT_mult_6_U4657 ( .A1(MULT_mult_6_n2225), .A2(MULT_mult_6_n2226), 
        .A3(MULT_mult_6_n2227), .ZN(MULT_mult_6_CARRYB_14__16_) );
  NAND2_X1 MULT_mult_6_U4656 ( .A1(MULT_mult_6_ab_14__16_), .A2(
        MULT_mult_6_n1250), .ZN(MULT_mult_6_n2226) );
  NAND2_X1 MULT_mult_6_U4655 ( .A1(MULT_mult_6_ab_14__16_), .A2(
        MULT_mult_6_CARRYB_13__16_), .ZN(MULT_mult_6_n2225) );
  NAND3_X2 MULT_mult_6_U4654 ( .A1(MULT_mult_6_n2222), .A2(MULT_mult_6_n2223), 
        .A3(MULT_mult_6_n2224), .ZN(MULT_mult_6_CARRYB_13__17_) );
  NAND2_X2 MULT_mult_6_U4653 ( .A1(MULT_mult_6_ab_13__17_), .A2(
        MULT_mult_6_CARRYB_12__17_), .ZN(MULT_mult_6_n2222) );
  NAND2_X2 MULT_mult_6_U4652 ( .A1(MULT_mult_6_ab_10__19_), .A2(
        MULT_mult_6_CARRYB_9__19_), .ZN(MULT_mult_6_n2219) );
  NAND2_X2 MULT_mult_6_U4651 ( .A1(MULT_mult_6_ab_9__20_), .A2(
        MULT_mult_6_n1278), .ZN(MULT_mult_6_n2217) );
  NAND2_X1 MULT_mult_6_U4650 ( .A1(MULT_mult_6_ab_9__20_), .A2(
        MULT_mult_6_CARRYB_8__20_), .ZN(MULT_mult_6_n2216) );
  XOR2_X2 MULT_mult_6_U4649 ( .A(MULT_mult_6_n2214), .B(MULT_mult_6_n1278), 
        .Z(MULT_mult_6_SUMB_9__20_) );
  NOR2_X1 MULT_mult_6_U4648 ( .A1(MULT_mult_6_net77908), .A2(
        MULT_mult_6_net70455), .ZN(MULT_mult_6_ab_20__6_) );
  NOR2_X2 MULT_mult_6_U4647 ( .A1(MULT_mult_6_net123000), .A2(
        MULT_mult_6_net77948), .ZN(MULT_mult_6_ab_5__17_) );
  NAND2_X2 MULT_mult_6_U4646 ( .A1(MULT_mult_6_ab_6__16_), .A2(
        MULT_mult_6_SUMB_5__17_), .ZN(MULT_mult_6_n2206) );
  XNOR2_X2 MULT_mult_6_U4645 ( .A(MULT_mult_6_ab_5__19_), .B(
        MULT_mult_6_CARRYB_4__19_), .ZN(MULT_mult_6_n2197) );
  NOR2_X1 MULT_mult_6_U4644 ( .A1(MULT_mult_6_net80643), .A2(
        MULT_mult_6_net77932), .ZN(MULT_mult_6_ab_7__21_) );
  NOR2_X1 MULT_mult_6_U4643 ( .A1(MULT_mult_6_net80643), .A2(
        MULT_mult_6_net77926), .ZN(MULT_mult_6_ab_8__21_) );
  NOR2_X1 MULT_mult_6_U4642 ( .A1(MULT_mult_6_net80643), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__21_) );
  NOR2_X1 MULT_mult_6_U4641 ( .A1(MULT_mult_6_net70470), .A2(
        MULT_mult_6_net77932), .ZN(MULT_mult_6_ab_7__18_) );
  NAND3_X4 MULT_mult_6_U4640 ( .A1(MULT_mult_6_n2193), .A2(MULT_mult_6_n2194), 
        .A3(MULT_mult_6_n2192), .ZN(MULT_mult_6_CARRYB_3__20_) );
  NAND2_X2 MULT_mult_6_U4639 ( .A1(MULT_mult_6_CARRYB_1__21_), .A2(
        MULT_mult_6_n1692), .ZN(MULT_mult_6_n2191) );
  NAND2_X2 MULT_mult_6_U4638 ( .A1(MULT_mult_6_SUMB_15__9_), .A2(
        MULT_mult_6_CARRYB_15__8_), .ZN(MULT_mult_6_n2301) );
  XNOR2_X2 MULT_mult_6_U4637 ( .A(MULT_mult_6_ab_14__16_), .B(
        MULT_mult_6_CARRYB_13__16_), .ZN(MULT_mult_6_n2188) );
  NOR2_X2 MULT_mult_6_U4636 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70453), .ZN(MULT_mult_6_ab_21__2_) );
  NAND3_X2 MULT_mult_6_U4635 ( .A1(MULT_mult_6_n2185), .A2(MULT_mult_6_n2186), 
        .A3(MULT_mult_6_n2187), .ZN(MULT_mult_6_CARRYB_21__2_) );
  NAND2_X2 MULT_mult_6_U4634 ( .A1(MULT_mult_6_SUMB_20__3_), .A2(
        MULT_mult_6_ab_21__2_), .ZN(MULT_mult_6_n2186) );
  NAND3_X4 MULT_mult_6_U4633 ( .A1(MULT_mult_6_n2301), .A2(MULT_mult_6_n2300), 
        .A3(MULT_mult_6_n2299), .ZN(MULT_mult_6_CARRYB_16__8_) );
  NOR2_X1 MULT_mult_6_U4632 ( .A1(MULT_mult_6_net123000), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__17_) );
  NOR2_X1 MULT_mult_6_U4631 ( .A1(MULT_mult_6_net123000), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__17_) );
  XNOR2_X2 MULT_mult_6_U4630 ( .A(MULT_mult_6_ab_8__22_), .B(
        MULT_mult_6_CARRYB_7__22_), .ZN(MULT_mult_6_n2184) );
  XNOR2_X2 MULT_mult_6_U4629 ( .A(MULT_mult_6_n2184), .B(
        MULT_mult_6_SUMB_7__23_), .ZN(MULT_mult_6_SUMB_8__22_) );
  NAND3_X2 MULT_mult_6_U4628 ( .A1(MULT_mult_6_n877), .A2(MULT_mult_6_n2182), 
        .A3(MULT_mult_6_n2183), .ZN(MULT_mult_6_CARRYB_7__22_) );
  NAND2_X1 MULT_mult_6_U4627 ( .A1(MULT_mult_6_CARRYB_6__22_), .A2(
        MULT_mult_6_SUMB_6__23_), .ZN(MULT_mult_6_n2183) );
  NAND2_X1 MULT_mult_6_U4626 ( .A1(MULT_mult_6_ab_7__22_), .A2(
        MULT_mult_6_SUMB_6__23_), .ZN(MULT_mult_6_n2182) );
  NAND3_X2 MULT_mult_6_U4625 ( .A1(MULT_mult_6_n2179), .A2(MULT_mult_6_n2180), 
        .A3(MULT_mult_6_n2181), .ZN(MULT_mult_6_CARRYB_6__23_) );
  NAND3_X2 MULT_mult_6_U4624 ( .A1(MULT_mult_6_n2176), .A2(MULT_mult_6_n2177), 
        .A3(MULT_mult_6_n2178), .ZN(MULT_mult_6_CARRYB_4__25_) );
  NAND2_X1 MULT_mult_6_U4623 ( .A1(MULT_mult_6_CARRYB_3__25_), .A2(
        MULT_mult_6_SUMB_3__26_), .ZN(MULT_mult_6_n2178) );
  NAND2_X1 MULT_mult_6_U4622 ( .A1(MULT_mult_6_ab_4__25_), .A2(
        MULT_mult_6_SUMB_3__26_), .ZN(MULT_mult_6_n2177) );
  NAND2_X1 MULT_mult_6_U4621 ( .A1(MULT_mult_6_ab_4__25_), .A2(
        MULT_mult_6_CARRYB_3__25_), .ZN(MULT_mult_6_n2176) );
  NAND3_X2 MULT_mult_6_U4620 ( .A1(MULT_mult_6_n2173), .A2(MULT_mult_6_n2174), 
        .A3(MULT_mult_6_n2175), .ZN(MULT_mult_6_CARRYB_3__26_) );
  NAND2_X2 MULT_mult_6_U4619 ( .A1(MULT_mult_6_CARRYB_2__26_), .A2(
        MULT_mult_6_n1197), .ZN(MULT_mult_6_n2175) );
  NAND2_X2 MULT_mult_6_U4618 ( .A1(MULT_mult_6_ab_3__26_), .A2(
        MULT_mult_6_n1197), .ZN(MULT_mult_6_n2174) );
  NAND2_X1 MULT_mult_6_U4617 ( .A1(MULT_mult_6_ab_3__26_), .A2(
        MULT_mult_6_CARRYB_2__26_), .ZN(MULT_mult_6_n2173) );
  XOR2_X2 MULT_mult_6_U4616 ( .A(MULT_mult_6_n2172), .B(MULT_mult_6_n1197), 
        .Z(MULT_mult_6_SUMB_3__26_) );
  XOR2_X2 MULT_mult_6_U4615 ( .A(MULT_mult_6_ab_3__26_), .B(
        MULT_mult_6_CARRYB_2__26_), .Z(MULT_mult_6_n2172) );
  NAND2_X2 MULT_mult_6_U4614 ( .A1(MULT_mult_6_n349), .A2(
        MULT_mult_6_SUMB_1__26_), .ZN(MULT_mult_6_n2167) );
  NAND2_X2 MULT_mult_6_U4613 ( .A1(MULT_mult_6_ab_20__1_), .A2(
        MULT_mult_6_SUMB_19__2_), .ZN(MULT_mult_6_n2160) );
  NAND2_X1 MULT_mult_6_U4612 ( .A1(MULT_mult_6_ab_7__13_), .A2(
        MULT_mult_6_CARRYB_6__13_), .ZN(MULT_mult_6_n2159) );
  NOR2_X1 MULT_mult_6_U4611 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net70459), .ZN(MULT_mult_6_ab_18__9_) );
  NOR2_X1 MULT_mult_6_U4610 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70451), .ZN(MULT_mult_6_ab_22__2_) );
  INV_X4 MULT_mult_6_U4609 ( .A(MULT_mult_6_n896), .ZN(MULT_mult_6_n2148) );
  NAND3_X4 MULT_mult_6_U4608 ( .A1(MULT_mult_6_n2143), .A2(MULT_mult_6_n2144), 
        .A3(MULT_mult_6_n2145), .ZN(MULT_mult_6_CARRYB_2__19_) );
  NAND2_X2 MULT_mult_6_U4607 ( .A1(MULT_mult_6_CARRYB_1__19_), .A2(
        MULT_mult_6_ab_2__19_), .ZN(MULT_mult_6_n2145) );
  NOR2_X1 MULT_mult_6_U4606 ( .A1(MULT_mult_6_net70453), .A2(
        MULT_mult_6_net91660), .ZN(MULT_mult_6_ab_21__10_) );
  NAND3_X2 MULT_mult_6_U4605 ( .A1(MULT_mult_6_n2256), .A2(MULT_mult_6_n2257), 
        .A3(MULT_mult_6_n2258), .ZN(MULT_mult_6_CARRYB_19__11_) );
  NAND3_X4 MULT_mult_6_U4604 ( .A1(MULT_mult_6_n2138), .A2(MULT_mult_6_n2137), 
        .A3(MULT_mult_6_n2136), .ZN(MULT_mult_6_CARRYB_4__19_) );
  NAND2_X2 MULT_mult_6_U4603 ( .A1(MULT_mult_6_ab_4__19_), .A2(
        MULT_mult_6_CARRYB_3__19_), .ZN(MULT_mult_6_n2136) );
  NAND3_X2 MULT_mult_6_U4602 ( .A1(MULT_mult_6_n2132), .A2(MULT_mult_6_n2133), 
        .A3(MULT_mult_6_n2134), .ZN(MULT_mult_6_CARRYB_21__9_) );
  NAND2_X1 MULT_mult_6_U4601 ( .A1(MULT_mult_6_SUMB_20__10_), .A2(
        MULT_mult_6_n370), .ZN(MULT_mult_6_n2134) );
  NAND2_X1 MULT_mult_6_U4600 ( .A1(MULT_mult_6_ab_21__9_), .A2(
        MULT_mult_6_n568), .ZN(MULT_mult_6_n2133) );
  NAND2_X1 MULT_mult_6_U4599 ( .A1(MULT_mult_6_ab_21__9_), .A2(
        MULT_mult_6_n370), .ZN(MULT_mult_6_n2132) );
  NAND3_X2 MULT_mult_6_U4598 ( .A1(MULT_mult_6_n2129), .A2(MULT_mult_6_n2130), 
        .A3(MULT_mult_6_n2131), .ZN(MULT_mult_6_CARRYB_20__10_) );
  NAND2_X1 MULT_mult_6_U4597 ( .A1(MULT_mult_6_ab_20__10_), .A2(
        MULT_mult_6_CARRYB_19__10_), .ZN(MULT_mult_6_n2129) );
  NOR2_X1 MULT_mult_6_U4596 ( .A1(MULT_mult_6_net70456), .A2(
        MULT_mult_6_net77924), .ZN(MULT_mult_6_ab_8__11_) );
  NAND2_X2 MULT_mult_6_U4595 ( .A1(MULT_mult_6_ab_13__12_), .A2(
        MULT_mult_6_SUMB_12__13_), .ZN(MULT_mult_6_n2124) );
  NAND2_X2 MULT_mult_6_U4594 ( .A1(MULT_mult_6_ab_14__12_), .A2(
        MULT_mult_6_SUMB_13__13_), .ZN(MULT_mult_6_n2121) );
  XNOR2_X2 MULT_mult_6_U4593 ( .A(MULT_mult_6_SUMB_20__11_), .B(
        MULT_mult_6_ab_21__10_), .ZN(MULT_mult_6_n2119) );
  XNOR2_X2 MULT_mult_6_U4592 ( .A(MULT_mult_6_n2119), .B(
        MULT_mult_6_CARRYB_20__10_), .ZN(MULT_mult_6_SUMB_21__10_) );
  XNOR2_X2 MULT_mult_6_U4591 ( .A(MULT_mult_6_n2112), .B(
        MULT_mult_6_SUMB_5__18_), .ZN(MULT_mult_6_SUMB_6__17_) );
  XNOR2_X2 MULT_mult_6_U4590 ( .A(MULT_mult_6_n2111), .B(
        MULT_mult_6_SUMB_2__19_), .ZN(MULT_mult_6_SUMB_3__18_) );
  XNOR2_X2 MULT_mult_6_U4589 ( .A(MULT_mult_6_n2110), .B(MULT_mult_6_n1209), 
        .ZN(MULT_mult_6_SUMB_19__3_) );
  NOR2_X1 MULT_mult_6_U4588 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70463), .ZN(MULT_mult_6_ab_16__4_) );
  NAND3_X2 MULT_mult_6_U4587 ( .A1(MULT_mult_6_n2101), .A2(MULT_mult_6_n2102), 
        .A3(MULT_mult_6_n2100), .ZN(MULT_mult_6_CARRYB_20__0_) );
  NAND2_X2 MULT_mult_6_U4586 ( .A1(MULT_mult_6_ab_20__0_), .A2(
        MULT_mult_6_SUMB_19__1_), .ZN(MULT_mult_6_n2101) );
  NOR2_X1 MULT_mult_6_U4585 ( .A1(MULT_mult_6_net70486), .A2(MULT_mult_6_n331), 
        .ZN(MULT_mult_6_ab_2__26_) );
  NOR2_X1 MULT_mult_6_U4584 ( .A1(MULT_mult_6_net85716), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__11_) );
  NAND3_X2 MULT_mult_6_U4583 ( .A1(MULT_mult_6_net81178), .A2(
        MULT_mult_6_net81179), .A3(MULT_mult_6_net81180), .ZN(
        MULT_mult_6_CARRYB_22__8_) );
  NAND3_X2 MULT_mult_6_U4582 ( .A1(MULT_mult_6_n2096), .A2(MULT_mult_6_n2098), 
        .A3(MULT_mult_6_n2097), .ZN(MULT_mult_6_CARRYB_16__11_) );
  NAND2_X1 MULT_mult_6_U4581 ( .A1(MULT_mult_6_ab_16__11_), .A2(
        MULT_mult_6_n1187), .ZN(MULT_mult_6_n2096) );
  NAND3_X2 MULT_mult_6_U4580 ( .A1(MULT_mult_6_n2092), .A2(MULT_mult_6_n2093), 
        .A3(MULT_mult_6_n2094), .ZN(MULT_mult_6_CARRYB_15__11_) );
  NAND2_X1 MULT_mult_6_U4579 ( .A1(MULT_mult_6_n1545), .A2(
        MULT_mult_6_net125062), .ZN(MULT_mult_6_n2094) );
  NAND2_X1 MULT_mult_6_U4578 ( .A1(MULT_mult_6_ab_15__11_), .A2(
        MULT_mult_6_n1545), .ZN(MULT_mult_6_n2092) );
  NAND2_X2 MULT_mult_6_U4577 ( .A1(MULT_mult_6_ab_3__24_), .A2(
        MULT_mult_6_SUMB_2__25_), .ZN(MULT_mult_6_n2169) );
  NAND3_X4 MULT_mult_6_U4576 ( .A1(MULT_mult_6_n2168), .A2(MULT_mult_6_n2169), 
        .A3(MULT_mult_6_n2170), .ZN(MULT_mult_6_CARRYB_3__24_) );
  NOR2_X1 MULT_mult_6_U4575 ( .A1(MULT_mult_6_net91660), .A2(
        MULT_mult_6_net77930), .ZN(MULT_mult_6_ab_7__10_) );
  NAND3_X2 MULT_mult_6_U4574 ( .A1(MULT_mult_6_net81205), .A2(
        MULT_mult_6_net81204), .A3(MULT_mult_6_net81206), .ZN(
        MULT_mult_6_CARRYB_5__12_) );
  NAND2_X2 MULT_mult_6_U4573 ( .A1(MULT_mult_6_SUMB_7__10_), .A2(
        MULT_mult_6_CARRYB_7__9_), .ZN(MULT_mult_6_n2085) );
  NAND3_X4 MULT_mult_6_U4572 ( .A1(MULT_mult_6_net81212), .A2(
        MULT_mult_6_net81213), .A3(MULT_mult_6_net81211), .ZN(
        MULT_mult_6_CARRYB_7__11_) );
  NAND2_X2 MULT_mult_6_U4571 ( .A1(MULT_mult_6_SUMB_5__9_), .A2(
        MULT_mult_6_ab_6__8_), .ZN(MULT_mult_6_n2078) );
  NAND2_X1 MULT_mult_6_U4570 ( .A1(MULT_mult_6_ab_6__13_), .A2(
        MULT_mult_6_CARRYB_5__13_), .ZN(MULT_mult_6_n2068) );
  NAND3_X4 MULT_mult_6_U4569 ( .A1(MULT_mult_6_net81262), .A2(
        MULT_mult_6_net81261), .A3(MULT_mult_6_net81260), .ZN(
        MULT_mult_6_CARRYB_10__10_) );
  NAND3_X4 MULT_mult_6_U4568 ( .A1(MULT_mult_6_net81258), .A2(
        MULT_mult_6_net81259), .A3(MULT_mult_6_n2067), .ZN(
        MULT_mult_6_CARRYB_9__11_) );
  NAND2_X1 MULT_mult_6_U4567 ( .A1(MULT_mult_6_CARRYB_8__11_), .A2(
        MULT_mult_6_ab_9__11_), .ZN(MULT_mult_6_n2067) );
  NOR2_X1 MULT_mult_6_U4566 ( .A1(MULT_mult_6_net70470), .A2(
        MULT_mult_6_net77926), .ZN(MULT_mult_6_ab_8__18_) );
  NOR2_X1 MULT_mult_6_U4565 ( .A1(MULT_mult_6_n182), .A2(MULT_mult_6_net70475), 
        .ZN(MULT_mult_6_ab_10__18_) );
  NOR2_X1 MULT_mult_6_U4564 ( .A1(MULT_mult_6_n182), .A2(MULT_mult_6_net70473), 
        .ZN(MULT_mult_6_ab_11__18_) );
  NOR2_X1 MULT_mult_6_U4563 ( .A1(MULT_mult_6_n182), .A2(MULT_mult_6_net70471), 
        .ZN(MULT_mult_6_ab_12__18_) );
  NOR2_X1 MULT_mult_6_U4562 ( .A1(MULT_mult_6_net70469), .A2(MULT_mult_6_n182), 
        .ZN(MULT_mult_6_ab_13__18_) );
  NAND2_X1 MULT_mult_6_U4561 ( .A1(MULT_mult_6_CARRYB_19__10_), .A2(
        MULT_mult_6_SUMB_19__11_), .ZN(MULT_mult_6_n2131) );
  NOR2_X1 MULT_mult_6_U4560 ( .A1(MULT_mult_6_net70465), .A2(
        MULT_mult_6_net124723), .ZN(MULT_mult_6_ab_15__16_) );
  XOR2_X2 MULT_mult_6_U4559 ( .A(MULT_mult_6_CARRYB_14__16_), .B(
        MULT_mult_6_ab_15__16_), .Z(MULT_mult_6_n2066) );
  XNOR2_X2 MULT_mult_6_U4558 ( .A(MULT_mult_6_n2065), .B(
        MULT_mult_6_SUMB_14__13_), .ZN(MULT_mult_6_SUMB_15__12_) );
  NOR2_X1 MULT_mult_6_U4557 ( .A1(MULT_mult_6_net77898), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__5_) );
  NOR2_X1 MULT_mult_6_U4556 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net77930), .ZN(MULT_mult_6_ab_7__8_) );
  NAND2_X1 MULT_mult_6_U4555 ( .A1(MULT_mult_6_ab_11__5_), .A2(
        MULT_mult_6_CARRYB_10__5_), .ZN(MULT_mult_6_n2063) );
  NAND2_X1 MULT_mult_6_U4554 ( .A1(MULT_mult_6_ab_9__15_), .A2(
        MULT_mult_6_CARRYB_8__15_), .ZN(MULT_mult_6_n2050) );
  INV_X4 MULT_mult_6_U4553 ( .A(MULT_mult_6_CARRYB_5__17_), .ZN(
        MULT_mult_6_n2044) );
  NAND2_X1 MULT_mult_6_U4552 ( .A1(MULT_mult_6_ab_19__11_), .A2(
        MULT_mult_6_SUMB_18__12_), .ZN(MULT_mult_6_n2257) );
  NAND2_X1 MULT_mult_6_U4551 ( .A1(MULT_mult_6_SUMB_9__20_), .A2(
        MULT_mult_6_CARRYB_9__19_), .ZN(MULT_mult_6_n2221) );
  NAND2_X1 MULT_mult_6_U4550 ( .A1(MULT_mult_6_SUMB_9__20_), .A2(
        MULT_mult_6_ab_10__19_), .ZN(MULT_mult_6_n2220) );
  NAND2_X2 MULT_mult_6_U4549 ( .A1(MULT_mult_6_ab_24__5_), .A2(
        MULT_mult_6_SUMB_23__6_), .ZN(MULT_mult_6_net79969) );
  NAND2_X2 MULT_mult_6_U4548 ( .A1(MULT_mult_6_SUMB_16__6_), .A2(
        MULT_mult_6_CARRYB_16__5_), .ZN(MULT_mult_6_n2039) );
  NAND2_X2 MULT_mult_6_U4547 ( .A1(MULT_mult_6_ab_17__5_), .A2(
        MULT_mult_6_SUMB_16__6_), .ZN(MULT_mult_6_n2038) );
  XNOR2_X2 MULT_mult_6_U4546 ( .A(MULT_mult_6_ab_8__20_), .B(
        MULT_mult_6_CARRYB_7__20_), .ZN(MULT_mult_6_n2036) );
  XNOR2_X2 MULT_mult_6_U4545 ( .A(MULT_mult_6_n851), .B(MULT_mult_6_n2036), 
        .ZN(MULT_mult_6_SUMB_8__20_) );
  NOR2_X1 MULT_mult_6_U4544 ( .A1(MULT_mult_6_net70457), .A2(
        MULT_mult_6_net83784), .ZN(MULT_mult_6_ab_19__12_) );
  NAND2_X2 MULT_mult_6_U4543 ( .A1(MULT_mult_6_ab_7__14_), .A2(
        MULT_mult_6_SUMB_6__15_), .ZN(MULT_mult_6_n2035) );
  NAND3_X4 MULT_mult_6_U4542 ( .A1(MULT_mult_6_n2033), .A2(MULT_mult_6_n2034), 
        .A3(MULT_mult_6_n2032), .ZN(MULT_mult_6_CARRYB_6__15_) );
  NAND2_X2 MULT_mult_6_U4541 ( .A1(MULT_mult_6_SUMB_5__16_), .A2(
        MULT_mult_6_n847), .ZN(MULT_mult_6_n2034) );
  NAND2_X2 MULT_mult_6_U4540 ( .A1(MULT_mult_6_ab_6__15_), .A2(
        MULT_mult_6_SUMB_5__16_), .ZN(MULT_mult_6_n2033) );
  NOR2_X2 MULT_mult_6_U4539 ( .A1(MULT_mult_6_net70471), .A2(
        MULT_mult_6_net86565), .ZN(MULT_mult_6_ab_12__19_) );
  NOR2_X2 MULT_mult_6_U4538 ( .A1(MULT_mult_6_net86565), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__19_) );
  NOR2_X2 MULT_mult_6_U4537 ( .A1(MULT_mult_6_net86565), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__19_) );
  NOR2_X2 MULT_mult_6_U4536 ( .A1(MULT_mult_6_net86565), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__19_) );
  NOR2_X2 MULT_mult_6_U4535 ( .A1(MULT_mult_6_net86565), .A2(
        MULT_mult_6_net77932), .ZN(MULT_mult_6_ab_7__19_) );
  NOR2_X2 MULT_mult_6_U4534 ( .A1(MULT_mult_6_net86565), .A2(
        MULT_mult_6_net119855), .ZN(MULT_mult_6_ab_4__19_) );
  XNOR2_X2 MULT_mult_6_U4533 ( .A(MULT_mult_6_n2031), .B(
        MULT_mult_6_SUMB_8__16_), .ZN(MULT_mult_6_SUMB_9__15_) );
  XNOR2_X2 MULT_mult_6_U4532 ( .A(MULT_mult_6_net81493), .B(
        MULT_mult_6_net88868), .ZN(MULT_mult_6_SUMB_22__3_) );
  NOR2_X1 MULT_mult_6_U4531 ( .A1(MULT_mult_6_net77912), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__7_) );
  NAND2_X2 MULT_mult_6_U4530 ( .A1(MULT_mult_6_CARRYB_24__0_), .A2(
        MULT_mult_6_ab_25__0_), .ZN(MULT_mult_6_n2025) );
  NAND2_X2 MULT_mult_6_U4529 ( .A1(MULT_mult_6_ab_12__7_), .A2(
        MULT_mult_6_SUMB_11__8_), .ZN(MULT_mult_6_n2020) );
  NAND3_X2 MULT_mult_6_U4528 ( .A1(MULT_mult_6_n2016), .A2(MULT_mult_6_n2017), 
        .A3(MULT_mult_6_n2018), .ZN(MULT_mult_6_CARRYB_9__7_) );
  NAND2_X2 MULT_mult_6_U4527 ( .A1(MULT_mult_6_ab_3__20_), .A2(
        MULT_mult_6_SUMB_2__21_), .ZN(MULT_mult_6_n2193) );
  NAND2_X2 MULT_mult_6_U4526 ( .A1(MULT_mult_6_SUMB_2__21_), .A2(
        MULT_mult_6_CARRYB_2__20_), .ZN(MULT_mult_6_n2194) );
  NOR2_X1 MULT_mult_6_U4525 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70443), .ZN(MULT_mult_6_ab_26__4_) );
  NAND3_X4 MULT_mult_6_U4524 ( .A1(MULT_mult_6_n2069), .A2(MULT_mult_6_n2070), 
        .A3(MULT_mult_6_n2068), .ZN(MULT_mult_6_CARRYB_6__13_) );
  XNOR2_X2 MULT_mult_6_U4523 ( .A(MULT_mult_6_n1425), .B(MULT_mult_6_ab_7__8_), 
        .ZN(MULT_mult_6_n2014) );
  NAND2_X2 MULT_mult_6_U4522 ( .A1(MULT_mult_6_net88702), .A2(
        MULT_mult_6_ab_19__7_), .ZN(MULT_mult_6_n2011) );
  NAND2_X2 MULT_mult_6_U4521 ( .A1(MULT_mult_6_n938), .A2(
        MULT_mult_6_CARRYB_7__8_), .ZN(MULT_mult_6_n2006) );
  XNOR2_X2 MULT_mult_6_U4520 ( .A(MULT_mult_6_net149004), .B(
        MULT_mult_6_net81586), .ZN(MULT_mult_6_SUMB_7__10_) );
  NOR2_X1 MULT_mult_6_U4519 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net70459), .ZN(MULT_mult_6_ab_18__12_) );
  NOR2_X1 MULT_mult_6_U4518 ( .A1(MULT_mult_6_net85716), .A2(
        MULT_mult_6_net70463), .ZN(MULT_mult_6_ab_16__11_) );
  NOR2_X1 MULT_mult_6_U4517 ( .A1(MULT_mult_6_net85716), .A2(
        MULT_mult_6_net70461), .ZN(MULT_mult_6_ab_17__11_) );
  NOR2_X1 MULT_mult_6_U4516 ( .A1(MULT_mult_6_net85716), .A2(
        MULT_mult_6_net70457), .ZN(MULT_mult_6_ab_19__11_) );
  NOR2_X1 MULT_mult_6_U4515 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__2_) );
  NAND3_X2 MULT_mult_6_U4514 ( .A1(MULT_mult_6_n1995), .A2(MULT_mult_6_n1996), 
        .A3(MULT_mult_6_n1997), .ZN(MULT_mult_6_CARRYB_12__2_) );
  NAND2_X2 MULT_mult_6_U4513 ( .A1(MULT_mult_6_ab_12__2_), .A2(
        MULT_mult_6_SUMB_11__3_), .ZN(MULT_mult_6_n1996) );
  XNOR2_X2 MULT_mult_6_U4512 ( .A(MULT_mult_6_n1993), .B(MULT_mult_6_n1253), 
        .ZN(MULT_mult_6_SUMB_14__4_) );
  NAND2_X2 MULT_mult_6_U4511 ( .A1(MULT_mult_6_ab_25__4_), .A2(
        MULT_mult_6_SUMB_24__5_), .ZN(MULT_mult_6_n2114) );
  NAND2_X2 MULT_mult_6_U4510 ( .A1(MULT_mult_6_SUMB_8__9_), .A2(
        MULT_mult_6_ab_9__8_), .ZN(MULT_mult_6_n2087) );
  NAND2_X2 MULT_mult_6_U4509 ( .A1(MULT_mult_6_CARRYB_8__8_), .A2(
        MULT_mult_6_SUMB_8__9_), .ZN(MULT_mult_6_n2088) );
  NOR2_X1 MULT_mult_6_U4508 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__3_) );
  NAND2_X2 MULT_mult_6_U4507 ( .A1(MULT_mult_6_n17), .A2(MULT_mult_6_ab_15__3_), .ZN(MULT_mult_6_n1991) );
  NAND3_X2 MULT_mult_6_U4506 ( .A1(MULT_mult_6_n1986), .A2(MULT_mult_6_n1985), 
        .A3(MULT_mult_6_n1984), .ZN(MULT_mult_6_CARRYB_2__15_) );
  NAND3_X4 MULT_mult_6_U4505 ( .A1(MULT_mult_6_net81713), .A2(
        MULT_mult_6_net81714), .A3(MULT_mult_6_n1983), .ZN(
        MULT_mult_6_CARRYB_6__12_) );
  NAND2_X2 MULT_mult_6_U4504 ( .A1(MULT_mult_6_SUMB_4__14_), .A2(
        MULT_mult_6_n1255), .ZN(MULT_mult_6_n1982) );
  NAND2_X2 MULT_mult_6_U4502 ( .A1(MULT_mult_6_ab_14__6_), .A2(
        MULT_mult_6_SUMB_13__7_), .ZN(MULT_mult_6_n1975) );
  NAND3_X4 MULT_mult_6_U4501 ( .A1(MULT_mult_6_net80845), .A2(
        MULT_mult_6_net80844), .A3(MULT_mult_6_n2159), .ZN(
        MULT_mult_6_CARRYB_7__13_) );
  NAND2_X1 MULT_mult_6_U4500 ( .A1(MULT_mult_6_ab_2__25_), .A2(
        MULT_mult_6_SUMB_1__26_), .ZN(MULT_mult_6_n2166) );
  NAND2_X1 MULT_mult_6_U4499 ( .A1(MULT_mult_6_ab_2__25_), .A2(
        MULT_mult_6_n349), .ZN(MULT_mult_6_n2165) );
  NAND2_X1 MULT_mult_6_U4498 ( .A1(MULT_mult_6_ab_20__10_), .A2(
        MULT_mult_6_SUMB_19__11_), .ZN(MULT_mult_6_n2130) );
  NOR2_X2 MULT_mult_6_U4497 ( .A1(MULT_mult_6_net91660), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__10_) );
  NAND2_X2 MULT_mult_6_U4496 ( .A1(MULT_mult_6_CARRYB_14__2_), .A2(
        MULT_mult_6_SUMB_14__3_), .ZN(MULT_mult_6_n1972) );
  NAND2_X2 MULT_mult_6_U4495 ( .A1(MULT_mult_6_ab_15__2_), .A2(
        MULT_mult_6_SUMB_14__3_), .ZN(MULT_mult_6_n1971) );
  NAND3_X2 MULT_mult_6_U4494 ( .A1(MULT_mult_6_n1962), .A2(MULT_mult_6_n1961), 
        .A3(MULT_mult_6_n1963), .ZN(MULT_mult_6_CARRYB_4__9_) );
  NAND2_X2 MULT_mult_6_U4493 ( .A1(MULT_mult_6_ab_6__23_), .A2(
        MULT_mult_6_CARRYB_5__23_), .ZN(MULT_mult_6_n2179) );
  NAND2_X1 MULT_mult_6_U4492 ( .A1(MULT_mult_6_CARRYB_5__23_), .A2(
        MULT_mult_6_n1231), .ZN(MULT_mult_6_n2181) );
  NAND3_X4 MULT_mult_6_U4491 ( .A1(MULT_mult_6_net80791), .A2(
        MULT_mult_6_net80792), .A3(MULT_mult_6_net80793), .ZN(
        MULT_mult_6_CARRYB_4__23_) );
  NOR2_X1 MULT_mult_6_U4490 ( .A1(MULT_mult_6_net84358), .A2(
        MULT_mult_6_net77948), .ZN(MULT_mult_6_ab_5__23_) );
  NAND2_X1 MULT_mult_6_U4489 ( .A1(MULT_mult_6_ab_5__23_), .A2(
        MULT_mult_6_CARRYB_4__23_), .ZN(MULT_mult_6_n1960) );
  NAND2_X1 MULT_mult_6_U4488 ( .A1(MULT_mult_6_CARRYB_4__23_), .A2(
        MULT_mult_6_SUMB_4__24_), .ZN(MULT_mult_6_n1958) );
  NAND3_X2 MULT_mult_6_U4487 ( .A1(MULT_mult_6_n1955), .A2(MULT_mult_6_n1956), 
        .A3(MULT_mult_6_n1957), .ZN(MULT_mult_6_CARRYB_17__13_) );
  NAND2_X1 MULT_mult_6_U4486 ( .A1(MULT_mult_6_CARRYB_16__13_), .A2(
        MULT_mult_6_SUMB_16__14_), .ZN(MULT_mult_6_n1957) );
  NAND2_X1 MULT_mult_6_U4485 ( .A1(MULT_mult_6_ab_17__13_), .A2(
        MULT_mult_6_SUMB_16__14_), .ZN(MULT_mult_6_n1956) );
  NAND2_X1 MULT_mult_6_U4484 ( .A1(MULT_mult_6_ab_17__13_), .A2(
        MULT_mult_6_CARRYB_16__13_), .ZN(MULT_mult_6_n1955) );
  NAND2_X2 MULT_mult_6_U4483 ( .A1(MULT_mult_6_CARRYB_15__14_), .A2(
        MULT_mult_6_n1269), .ZN(MULT_mult_6_n1954) );
  NAND2_X2 MULT_mult_6_U4482 ( .A1(MULT_mult_6_ab_16__14_), .A2(
        MULT_mult_6_n1269), .ZN(MULT_mult_6_n1953) );
  XNOR2_X2 MULT_mult_6_U4481 ( .A(MULT_mult_6_ab_10__16_), .B(
        MULT_mult_6_CARRYB_9__16_), .ZN(MULT_mult_6_net81945) );
  NAND2_X2 MULT_mult_6_U4480 ( .A1(MULT_mult_6_SUMB_19__9_), .A2(
        MULT_mult_6_ab_20__8_), .ZN(MULT_mult_6_net81956) );
  NOR2_X1 MULT_mult_6_U4479 ( .A1(MULT_mult_6_net77906), .A2(
        MULT_mult_6_net77938), .ZN(MULT_mult_6_ab_6__6_) );
  NAND3_X2 MULT_mult_6_U4478 ( .A1(MULT_mult_6_n1949), .A2(MULT_mult_6_n1950), 
        .A3(MULT_mult_6_n1951), .ZN(MULT_mult_6_CARRYB_6__6_) );
  NOR2_X1 MULT_mult_6_U4477 ( .A1(MULT_mult_6_net70470), .A2(
        MULT_mult_6_net119855), .ZN(MULT_mult_6_ab_4__18_) );
  NOR2_X1 MULT_mult_6_U4476 ( .A1(MULT_mult_6_net70470), .A2(
        MULT_mult_6_net77948), .ZN(MULT_mult_6_ab_5__18_) );
  NOR2_X1 MULT_mult_6_U4475 ( .A1(MULT_mult_6_net70470), .A2(
        MULT_mult_6_net77940), .ZN(MULT_mult_6_ab_6__18_) );
  XNOR2_X2 MULT_mult_6_U4474 ( .A(MULT_mult_6_n1256), .B(MULT_mult_6_n1942), 
        .ZN(MULT_mult_6_SUMB_6__13_) );
  NAND2_X2 MULT_mult_6_U4473 ( .A1(MULT_mult_6_ab_7__15_), .A2(
        MULT_mult_6_SUMB_6__16_), .ZN(MULT_mult_6_n2209) );
  NAND3_X4 MULT_mult_6_U4472 ( .A1(MULT_mult_6_n1940), .A2(MULT_mult_6_n1939), 
        .A3(MULT_mult_6_n1938), .ZN(MULT_mult_6_CARRYB_14__9_) );
  XNOR2_X2 MULT_mult_6_U4471 ( .A(MULT_mult_6_n176), .B(MULT_mult_6_ab_17__4_), 
        .ZN(MULT_mult_6_n1936) );
  NAND2_X1 MULT_mult_6_U4470 ( .A1(MULT_mult_6_ab_2__22_), .A2(
        MULT_mult_6_CARRYB_1__22_), .ZN(MULT_mult_6_n1930) );
  NAND2_X2 MULT_mult_6_U4469 ( .A1(MULT_mult_6_net82045), .A2(
        MULT_mult_6_net82046), .ZN(MULT_mult_6_n2347) );
  NAND3_X2 MULT_mult_6_U4468 ( .A1(MULT_mult_6_n1926), .A2(MULT_mult_6_n1925), 
        .A3(MULT_mult_6_n1924), .ZN(MULT_mult_6_CARRYB_10__4_) );
  NAND2_X2 MULT_mult_6_U4467 ( .A1(MULT_mult_6_CARRYB_9__4_), .A2(
        MULT_mult_6_ab_10__4_), .ZN(MULT_mult_6_n1925) );
  NAND2_X2 MULT_mult_6_U4465 ( .A1(MULT_mult_6_ab_9__4_), .A2(
        MULT_mult_6_SUMB_8__5_), .ZN(MULT_mult_6_n1923) );
  NAND3_X2 MULT_mult_6_U4464 ( .A1(MULT_mult_6_n1922), .A2(MULT_mult_6_n1921), 
        .A3(MULT_mult_6_n1920), .ZN(MULT_mult_6_CARRYB_13__5_) );
  NAND3_X2 MULT_mult_6_U4463 ( .A1(MULT_mult_6_n1946), .A2(MULT_mult_6_n1945), 
        .A3(MULT_mult_6_n1944), .ZN(MULT_mult_6_CARRYB_4__8_) );
  XNOR2_X2 MULT_mult_6_U4462 ( .A(MULT_mult_6_net82154), .B(
        MULT_mult_6_net90731), .ZN(MULT_mult_6_SUMB_6__11_) );
  NOR2_X1 MULT_mult_6_U4461 ( .A1(MULT_mult_6_net82239), .A2(
        MULT_mult_6_net77966), .ZN(MULT_mult_6_ab_3__25_) );
  NOR2_X2 MULT_mult_6_U4460 ( .A1(MULT_mult_6_net82239), .A2(
        MULT_mult_6_net77956), .ZN(MULT_mult_6_ab_4__25_) );
  NOR2_X2 MULT_mult_6_U4459 ( .A1(MULT_mult_6_net82239), .A2(
        MULT_mult_6_net77946), .ZN(MULT_mult_6_ab_5__25_) );
  NAND3_X2 MULT_mult_6_U4458 ( .A1(MULT_mult_6_n1914), .A2(MULT_mult_6_n1916), 
        .A3(MULT_mult_6_n1915), .ZN(MULT_mult_6_CARRYB_20__2_) );
  NAND3_X4 MULT_mult_6_U4457 ( .A1(MULT_mult_6_n1907), .A2(MULT_mult_6_n1906), 
        .A3(MULT_mult_6_n1905), .ZN(MULT_mult_6_CARRYB_3__8_) );
  XNOR2_X2 MULT_mult_6_U4456 ( .A(MULT_mult_6_CARRYB_3__21_), .B(
        MULT_mult_6_ab_4__21_), .ZN(MULT_mult_6_n1904) );
  XOR2_X1 MULT_mult_6_U4455 ( .A(MULT_mult_6_ab_20__0_), .B(
        MULT_mult_6_CARRYB_19__0_), .Z(MULT_mult_6_n2099) );
  NOR2_X1 MULT_mult_6_U4454 ( .A1(MULT_mult_6_net84698), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__14_) );
  NOR2_X1 MULT_mult_6_U4453 ( .A1(MULT_mult_6_net84698), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__14_) );
  NOR2_X1 MULT_mult_6_U4452 ( .A1(MULT_mult_6_net84698), .A2(
        MULT_mult_6_net70463), .ZN(MULT_mult_6_ab_16__14_) );
  NAND3_X2 MULT_mult_6_U4451 ( .A1(MULT_mult_6_n2245), .A2(MULT_mult_6_n2246), 
        .A3(MULT_mult_6_n2247), .ZN(MULT_mult_6_CARRYB_6__17_) );
  NAND2_X1 MULT_mult_6_U4450 ( .A1(MULT_mult_6_ab_3__24_), .A2(
        MULT_mult_6_CARRYB_2__24_), .ZN(MULT_mult_6_n2168) );
  NAND2_X2 MULT_mult_6_U4449 ( .A1(MULT_mult_6_CARRYB_16__3_), .A2(
        MULT_mult_6_ab_17__3_), .ZN(MULT_mult_6_n2106) );
  XNOR2_X2 MULT_mult_6_U4448 ( .A(MULT_mult_6_n1902), .B(MULT_mult_6_n1248), 
        .ZN(MULT_mult_6_SUMB_12__7_) );
  XNOR2_X2 MULT_mult_6_U4447 ( .A(MULT_mult_6_n1899), .B(MULT_mult_6_n1379), 
        .ZN(MULT_mult_6_SUMB_13__6_) );
  NAND2_X2 MULT_mult_6_U4446 ( .A1(MULT_mult_6_SUMB_3__20_), .A2(
        MULT_mult_6_CARRYB_3__19_), .ZN(MULT_mult_6_n2138) );
  INV_X4 MULT_mult_6_U4445 ( .A(MULT_mult_6_n2341), .ZN(
        MULT_mult_6_CARRYB_1__20_) );
  XNOR2_X2 MULT_mult_6_U4444 ( .A(MULT_mult_6_CARRYB_12__16_), .B(
        MULT_mult_6_ab_13__16_), .ZN(MULT_mult_6_n2296) );
  NAND3_X4 MULT_mult_6_U4443 ( .A1(MULT_mult_6_n1898), .A2(MULT_mult_6_n1897), 
        .A3(MULT_mult_6_n1896), .ZN(MULT_mult_6_CARRYB_5__16_) );
  NAND2_X2 MULT_mult_6_U4442 ( .A1(MULT_mult_6_n1242), .A2(
        MULT_mult_6_CARRYB_4__16_), .ZN(MULT_mult_6_n1898) );
  NAND2_X2 MULT_mult_6_U4441 ( .A1(MULT_mult_6_n861), .A2(
        MULT_mult_6_SUMB_3__18_), .ZN(MULT_mult_6_n1895) );
  NAND2_X2 MULT_mult_6_U4440 ( .A1(MULT_mult_6_SUMB_3__18_), .A2(
        MULT_mult_6_ab_4__17_), .ZN(MULT_mult_6_n1894) );
  INV_X1 MULT_mult_6_U4439 ( .A(MULT_mult_6_ab_6__16_), .ZN(MULT_mult_6_n1890)
         );
  XNOR2_X2 MULT_mult_6_U4438 ( .A(MULT_mult_6_n1889), .B(
        MULT_mult_6_CARRYB_8__20_), .ZN(MULT_mult_6_n2214) );
  XNOR2_X2 MULT_mult_6_U4437 ( .A(MULT_mult_6_CARRYB_2__19_), .B(
        MULT_mult_6_ab_3__19_), .ZN(MULT_mult_6_n1887) );
  XNOR2_X2 MULT_mult_6_U4436 ( .A(MULT_mult_6_n1887), .B(
        MULT_mult_6_SUMB_2__20_), .ZN(MULT_mult_6_SUMB_3__19_) );
  XNOR2_X2 MULT_mult_6_U4435 ( .A(MULT_mult_6_n1886), .B(
        MULT_mult_6_CARRYB_9__19_), .ZN(MULT_mult_6_n2215) );
  NAND2_X2 MULT_mult_6_U4434 ( .A1(MULT_mult_6_CARRYB_2__18_), .A2(
        MULT_mult_6_SUMB_2__19_), .ZN(MULT_mult_6_n2147) );
  NAND2_X2 MULT_mult_6_U4433 ( .A1(MULT_mult_6_ab_6__20_), .A2(
        MULT_mult_6_CARRYB_5__20_), .ZN(MULT_mult_6_net79937) );
  NAND3_X4 MULT_mult_6_U4432 ( .A1(MULT_mult_6_n2053), .A2(MULT_mult_6_n2052), 
        .A3(MULT_mult_6_n2051), .ZN(MULT_mult_6_CARRYB_2__20_) );
  XNOR2_X2 MULT_mult_6_U4431 ( .A(MULT_mult_6_n1880), .B(MULT_mult_6_n1217), 
        .ZN(MULT_mult_6_SUMB_5__8_) );
  NAND3_X4 MULT_mult_6_U4430 ( .A1(MULT_mult_6_n2286), .A2(MULT_mult_6_n2287), 
        .A3(MULT_mult_6_n2288), .ZN(MULT_mult_6_CARRYB_8__20_) );
  NOR2_X1 MULT_mult_6_U4429 ( .A1(MULT_mult_6_net70449), .A2(
        MULT_mult_6_net77920), .ZN(MULT_mult_6_ab_23__8_) );
  NOR2_X1 MULT_mult_6_U4428 ( .A1(MULT_mult_6_net81424), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__15_) );
  NAND3_X2 MULT_mult_6_U4427 ( .A1(MULT_mult_6_n1877), .A2(MULT_mult_6_n1878), 
        .A3(MULT_mult_6_n1879), .ZN(MULT_mult_6_CARRYB_11__17_) );
  NAND2_X1 MULT_mult_6_U4426 ( .A1(MULT_mult_6_CARRYB_10__17_), .A2(
        MULT_mult_6_SUMB_10__18_), .ZN(MULT_mult_6_n1879) );
  NAND2_X1 MULT_mult_6_U4425 ( .A1(MULT_mult_6_ab_11__17_), .A2(
        MULT_mult_6_SUMB_10__18_), .ZN(MULT_mult_6_n1878) );
  NAND2_X1 MULT_mult_6_U4424 ( .A1(MULT_mult_6_ab_11__17_), .A2(
        MULT_mult_6_CARRYB_10__17_), .ZN(MULT_mult_6_n1877) );
  NAND2_X1 MULT_mult_6_U4423 ( .A1(MULT_mult_6_ab_10__18_), .A2(
        MULT_mult_6_CARRYB_9__18_), .ZN(MULT_mult_6_n1874) );
  XOR2_X2 MULT_mult_6_U4422 ( .A(MULT_mult_6_n1873), .B(
        MULT_mult_6_SUMB_10__18_), .Z(MULT_mult_6_SUMB_11__17_) );
  XOR2_X2 MULT_mult_6_U4421 ( .A(MULT_mult_6_ab_11__17_), .B(
        MULT_mult_6_CARRYB_10__17_), .Z(MULT_mult_6_n1873) );
  NAND2_X1 MULT_mult_6_U4420 ( .A1(MULT_mult_6_ab_14__15_), .A2(
        MULT_mult_6_CARRYB_13__15_), .ZN(MULT_mult_6_n1872) );
  NAND2_X1 MULT_mult_6_U4419 ( .A1(MULT_mult_6_CARRYB_13__15_), .A2(
        MULT_mult_6_SUMB_13__16_), .ZN(MULT_mult_6_n1870) );
  NAND2_X2 MULT_mult_6_U4418 ( .A1(MULT_mult_6_ab_3__18_), .A2(
        MULT_mult_6_SUMB_2__19_), .ZN(MULT_mult_6_n2146) );
  NOR2_X1 MULT_mult_6_U4417 ( .A1(MULT_mult_6_net77898), .A2(
        MULT_mult_6_net77966), .ZN(MULT_mult_6_ab_3__5_) );
  NOR2_X2 MULT_mult_6_U4416 ( .A1(MULT_mult_6_net77898), .A2(
        MULT_mult_6_net77970), .ZN(MULT_mult_6_ab_2__5_) );
  NAND3_X2 MULT_mult_6_U4415 ( .A1(MULT_mult_6_n1866), .A2(MULT_mult_6_n1867), 
        .A3(MULT_mult_6_n1868), .ZN(MULT_mult_6_CARRYB_2__5_) );
  NAND2_X1 MULT_mult_6_U4414 ( .A1(MULT_mult_6_ab_2__5_), .A2(
        MULT_mult_6_CARRYB_1__5_), .ZN(MULT_mult_6_n1868) );
  NAND2_X2 MULT_mult_6_U4413 ( .A1(MULT_mult_6_ab_2__5_), .A2(
        MULT_mult_6_SUMB_1__6_), .ZN(MULT_mult_6_n1867) );
  XOR2_X2 MULT_mult_6_U4412 ( .A(MULT_mult_6_SUMB_1__6_), .B(MULT_mult_6_n1865), .Z(MULT_mult_6_SUMB_2__5_) );
  XOR2_X2 MULT_mult_6_U4411 ( .A(MULT_mult_6_CARRYB_1__5_), .B(
        MULT_mult_6_ab_2__5_), .Z(MULT_mult_6_n1865) );
  NOR2_X1 MULT_mult_6_U4410 ( .A1(MULT_mult_6_net77912), .A2(
        MULT_mult_6_net77924), .ZN(MULT_mult_6_ab_8__7_) );
  NAND2_X2 MULT_mult_6_U4409 ( .A1(MULT_mult_6_SUMB_5__17_), .A2(
        MULT_mult_6_CARRYB_5__16_), .ZN(MULT_mult_6_n2207) );
  NOR2_X1 MULT_mult_6_U4408 ( .A1(MULT_mult_6_net84698), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__14_) );
  NAND2_X2 MULT_mult_6_U4407 ( .A1(MULT_mult_6_n1251), .A2(MULT_mult_6_n2195), 
        .ZN(MULT_mult_6_n2156) );
  NOR2_X1 MULT_mult_6_U4406 ( .A1(MULT_mult_6_net91660), .A2(
        MULT_mult_6_net70459), .ZN(MULT_mult_6_ab_18__10_) );
  NOR2_X2 MULT_mult_6_U4405 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70457), .ZN(MULT_mult_6_ab_19__4_) );
  INV_X1 MULT_mult_6_U4404 ( .A(MULT_mult_6_ab_19__4_), .ZN(MULT_mult_6_n1857)
         );
  XNOR2_X2 MULT_mult_6_U4403 ( .A(MULT_mult_6_n1904), .B(
        MULT_mult_6_SUMB_3__22_), .ZN(MULT_mult_6_SUMB_4__21_) );
  NAND2_X2 MULT_mult_6_U4402 ( .A1(MULT_mult_6_SUMB_7__17_), .A2(
        MULT_mult_6_CARRYB_7__16_), .ZN(MULT_mult_6_n2298) );
  XNOR2_X2 MULT_mult_6_U4401 ( .A(MULT_mult_6_SUMB_12__17_), .B(
        MULT_mult_6_n2296), .ZN(MULT_mult_6_SUMB_13__16_) );
  NAND3_X4 MULT_mult_6_U4400 ( .A1(MULT_mult_6_n2161), .A2(MULT_mult_6_n2162), 
        .A3(MULT_mult_6_n2163), .ZN(MULT_mult_6_CARRYB_21__1_) );
  NOR2_X1 MULT_mult_6_U4399 ( .A1(MULT_mult_6_net77868), .A2(
        MULT_mult_6_net70451), .ZN(MULT_mult_6_ab_22__1_) );
  NAND2_X2 MULT_mult_6_U4398 ( .A1(MULT_mult_6_ab_17__1_), .A2(
        MULT_mult_6_SUMB_16__2_), .ZN(MULT_mult_6_net82534) );
  NAND2_X4 MULT_mult_6_U4397 ( .A1(MULT_mult_6_n1892), .A2(MULT_mult_6_n2205), 
        .ZN(MULT_mult_6_n2064) );
  NAND2_X1 MULT_mult_6_U4396 ( .A1(MULT_mult_6_ab_24__5_), .A2(
        MULT_mult_6_CARRYB_23__5_), .ZN(MULT_mult_6_net79970) );
  NAND3_X2 MULT_mult_6_U4395 ( .A1(MULT_mult_6_n2025), .A2(
        MULT_mult_6_net81530), .A3(MULT_mult_6_net81531), .ZN(
        MULT_mult_6_CARRYB_25__0_) );
  INV_X2 MULT_mult_6_U4394 ( .A(MULT_mult_6_ab_25__4_), .ZN(
        MULT_mult_6_net82550) );
  NAND2_X4 MULT_mult_6_U4393 ( .A1(MULT_mult_6_net82551), .A2(
        MULT_mult_6_net82550), .ZN(MULT_mult_6_n1855) );
  NOR2_X4 MULT_mult_6_U4392 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__12_) );
  INV_X1 MULT_mult_6_U4391 ( .A(MULT_mult_6_ab_16__11_), .ZN(MULT_mult_6_n1881) );
  INV_X1 MULT_mult_6_U4390 ( .A(MULT_mult_6_ab_15__12_), .ZN(MULT_mult_6_n1851) );
  INV_X4 MULT_mult_6_U4389 ( .A(MULT_mult_6_n1881), .ZN(MULT_mult_6_n1846) );
  XNOR2_X2 MULT_mult_6_U4388 ( .A(MULT_mult_6_net82601), .B(
        MULT_mult_6_net121926), .ZN(MULT_mult_6_SUMB_9__4_) );
  NAND2_X1 MULT_mult_6_U4387 ( .A1(MULT_mult_6_ab_11__14_), .A2(
        MULT_mult_6_CARRYB_10__14_), .ZN(MULT_mult_6_n1842) );
  NAND2_X1 MULT_mult_6_U4386 ( .A1(MULT_mult_6_ab_10__15_), .A2(
        MULT_mult_6_CARRYB_9__15_), .ZN(MULT_mult_6_n1839) );
  XNOR2_X2 MULT_mult_6_U4385 ( .A(MULT_mult_6_n11), .B(MULT_mult_6_n1270), 
        .ZN(MULT_mult_6_SUMB_17__5_) );
  XNOR2_X2 MULT_mult_6_U4384 ( .A(MULT_mult_6_n1836), .B(MULT_mult_6_n1325), 
        .ZN(MULT_mult_6_SUMB_8__9_) );
  NOR2_X1 MULT_mult_6_U4383 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__4_) );
  NAND2_X2 MULT_mult_6_U4382 ( .A1(MULT_mult_6_ab_11__5_), .A2(
        MULT_mult_6_SUMB_10__6_), .ZN(MULT_mult_6_n2062) );
  XNOR2_X2 MULT_mult_6_U4381 ( .A(MULT_mult_6_ab_2__21_), .B(
        MULT_mult_6_CARRYB_1__21_), .ZN(MULT_mult_6_n1828) );
  NAND3_X4 MULT_mult_6_U4380 ( .A1(MULT_mult_6_n2189), .A2(MULT_mult_6_n2190), 
        .A3(MULT_mult_6_n2191), .ZN(MULT_mult_6_CARRYB_2__21_) );
  XNOR2_X2 MULT_mult_6_U4379 ( .A(MULT_mult_6_n1820), .B(MULT_mult_6_n1264), 
        .ZN(MULT_mult_6_SUMB_7__9_) );
  INV_X8 MULT_mult_6_U4378 ( .A(MULT_mult_6_n1888), .ZN(MULT_mult_6_n1816) );
  NAND2_X1 MULT_mult_6_U4377 ( .A1(MULT_mult_6_ab_15__11_), .A2(
        MULT_mult_6_net125062), .ZN(MULT_mult_6_n2093) );
  NOR2_X1 MULT_mult_6_U4376 ( .A1(MULT_mult_6_net77858), .A2(
        MULT_mult_6_net70453), .ZN(MULT_mult_6_ab_21__0_) );
  NAND2_X2 MULT_mult_6_U4375 ( .A1(MULT_mult_6_ab_19__0_), .A2(
        MULT_mult_6_CARRYB_18__0_), .ZN(MULT_mult_6_n1814) );
  NAND2_X2 MULT_mult_6_U4374 ( .A1(MULT_mult_6_ab_19__0_), .A2(
        MULT_mult_6_SUMB_18__1_), .ZN(MULT_mult_6_n1813) );
  NAND3_X2 MULT_mult_6_U4372 ( .A1(MULT_mult_6_n1809), .A2(MULT_mult_6_n1810), 
        .A3(MULT_mult_6_n1811), .ZN(MULT_mult_6_CARRYB_18__0_) );
  NAND3_X4 MULT_mult_6_U4371 ( .A1(MULT_mult_6_n1805), .A2(MULT_mult_6_n1807), 
        .A3(MULT_mult_6_n1806), .ZN(MULT_mult_6_CARRYB_21__0_) );
  NAND3_X2 MULT_mult_6_U4370 ( .A1(MULT_mult_6_n1802), .A2(MULT_mult_6_n1803), 
        .A3(MULT_mult_6_n1804), .ZN(MULT_mult_6_CARRYB_10__3_) );
  NAND3_X2 MULT_mult_6_U4369 ( .A1(MULT_mult_6_net82848), .A2(
        MULT_mult_6_net82849), .A3(MULT_mult_6_net82850), .ZN(
        MULT_mult_6_CARRYB_9__3_) );
  NAND2_X2 MULT_mult_6_U4368 ( .A1(MULT_mult_6_n36), .A2(
        MULT_mult_6_SUMB_22__1_), .ZN(MULT_mult_6_n1801) );
  NAND2_X2 MULT_mult_6_U4367 ( .A1(MULT_mult_6_ab_23__0_), .A2(
        MULT_mult_6_CARRYB_22__0_), .ZN(MULT_mult_6_n1800) );
  NAND2_X2 MULT_mult_6_U4366 ( .A1(MULT_mult_6_ab_12__13_), .A2(
        MULT_mult_6_SUMB_11__14_), .ZN(MULT_mult_6_n1794) );
  INV_X4 MULT_mult_6_U4365 ( .A(MULT_mult_6_CARRYB_5__16_), .ZN(
        MULT_mult_6_n1891) );
  NAND2_X2 MULT_mult_6_U4364 ( .A1(MULT_mult_6_n2373), .A2(MULT_mult_6_n868), 
        .ZN(MULT_mult_6_n1913) );
  NOR2_X1 MULT_mult_6_U4363 ( .A1(MULT_mult_6_net77898), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__5_) );
  INV_X1 MULT_mult_6_U4362 ( .A(MULT_mult_6_ab_11__5_), .ZN(MULT_mult_6_n1835)
         );
  NAND3_X2 MULT_mult_6_U4361 ( .A1(MULT_mult_6_n1786), .A2(MULT_mult_6_n1785), 
        .A3(MULT_mult_6_n1787), .ZN(MULT_mult_6_CARRYB_9__5_) );
  INV_X4 MULT_mult_6_U4360 ( .A(MULT_mult_6_n1835), .ZN(MULT_mult_6_n1782) );
  NAND2_X2 MULT_mult_6_U4359 ( .A1(MULT_mult_6_n1891), .A2(MULT_mult_6_n1890), 
        .ZN(MULT_mult_6_n1892) );
  NOR2_X2 MULT_mult_6_U4358 ( .A1(MULT_mult_6_net80643), .A2(
        MULT_mult_6_net77964), .ZN(MULT_mult_6_ab_3__21_) );
  NOR2_X1 MULT_mult_6_U4357 ( .A1(MULT_mult_6_net70478), .A2(
        MULT_mult_6_net77940), .ZN(MULT_mult_6_ab_6__22_) );
  NOR2_X1 MULT_mult_6_U4356 ( .A1(MULT_mult_6_net70478), .A2(
        MULT_mult_6_net77932), .ZN(MULT_mult_6_ab_7__22_) );
  NOR2_X1 MULT_mult_6_U4355 ( .A1(MULT_mult_6_net70478), .A2(
        MULT_mult_6_net77926), .ZN(MULT_mult_6_ab_8__22_) );
  NOR2_X1 MULT_mult_6_U4354 ( .A1(MULT_mult_6_net70477), .A2(
        MULT_mult_6_net70478), .ZN(MULT_mult_6_ab_9__22_) );
  NAND2_X4 MULT_mult_6_U4353 ( .A1(MULT_mult_6_n1121), .A2(MULT_mult_6_n2149), 
        .ZN(MULT_mult_6_SUMB_24__5_) );
  NAND2_X2 MULT_mult_6_U4352 ( .A1(MULT_mult_6_n173), .A2(
        MULT_mult_6_SUMB_10__8_), .ZN(MULT_mult_6_n1779) );
  NAND3_X2 MULT_mult_6_U4351 ( .A1(MULT_mult_6_n1776), .A2(MULT_mult_6_n1775), 
        .A3(MULT_mult_6_n1774), .ZN(MULT_mult_6_CARRYB_10__8_) );
  XNOR2_X2 MULT_mult_6_U4350 ( .A(MULT_mult_6_CARRYB_15__6_), .B(
        MULT_mult_6_ab_16__6_), .ZN(MULT_mult_6_n1856) );
  NAND2_X2 MULT_mult_6_U4349 ( .A1(MULT_mult_6_SUMB_18__5_), .A2(
        MULT_mult_6_CARRYB_18__4_), .ZN(MULT_mult_6_n2236) );
  NOR2_X2 MULT_mult_6_U4348 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__13_) );
  INV_X1 MULT_mult_6_U4347 ( .A(MULT_mult_6_ab_15__11_), .ZN(MULT_mult_6_n1769) );
  NAND2_X4 MULT_mult_6_U4346 ( .A1(MULT_mult_6_n1770), .A2(
        MULT_mult_6_ab_15__11_), .ZN(MULT_mult_6_n1771) );
  NAND3_X4 MULT_mult_6_U4345 ( .A1(MULT_mult_6_net80561), .A2(
        MULT_mult_6_net80562), .A3(MULT_mult_6_net80563), .ZN(
        MULT_mult_6_CARRYB_15__8_) );
  NAND3_X2 MULT_mult_6_U4344 ( .A1(MULT_mult_6_net80879), .A2(
        MULT_mult_6_net80880), .A3(MULT_mult_6_n2154), .ZN(
        MULT_mult_6_CARRYB_18__9_) );
  XNOR2_X2 MULT_mult_6_U4343 ( .A(MULT_mult_6_CARRYB_6__17_), .B(
        MULT_mult_6_ab_7__17_), .ZN(MULT_mult_6_n1766) );
  NAND2_X4 MULT_mult_6_U4342 ( .A1(MULT_mult_6_n1850), .A2(MULT_mult_6_n1851), 
        .ZN(MULT_mult_6_n1853) );
  INV_X4 MULT_mult_6_U4341 ( .A(MULT_mult_6_ab_8__8_), .ZN(MULT_mult_6_n1830)
         );
  NAND2_X4 MULT_mult_6_U4340 ( .A1(MULT_mult_6_n1761), .A2(MULT_mult_6_n1760), 
        .ZN(MULT_mult_6_n1763) );
  NAND2_X2 MULT_mult_6_U4339 ( .A1(MULT_mult_6_n621), .A2(MULT_mult_6_n1830), 
        .ZN(MULT_mult_6_n1762) );
  NAND3_X2 MULT_mult_6_U4337 ( .A1(MULT_mult_6_n2283), .A2(MULT_mult_6_n2284), 
        .A3(MULT_mult_6_n2285), .ZN(MULT_mult_6_CARRYB_23__6_) );
  XNOR2_X2 MULT_mult_6_U4336 ( .A(MULT_mult_6_n2171), .B(MULT_mult_6_net122087), .ZN(MULT_mult_6_SUMB_21__2_) );
  NAND2_X2 MULT_mult_6_U4335 ( .A1(MULT_mult_6_CARRYB_11__7_), .A2(
        MULT_mult_6_SUMB_11__8_), .ZN(MULT_mult_6_n2021) );
  NAND3_X4 MULT_mult_6_U4334 ( .A1(MULT_mult_6_n2006), .A2(MULT_mult_6_n2004), 
        .A3(MULT_mult_6_n2005), .ZN(MULT_mult_6_CARRYB_8__8_) );
  NAND2_X4 MULT_mult_6_U4333 ( .A1(MULT_mult_6_n1853), .A2(MULT_mult_6_n1852), 
        .ZN(MULT_mult_6_n2065) );
  INV_X4 MULT_mult_6_U4332 ( .A(MULT_mult_6_net82834), .ZN(
        MULT_mult_6_net83172) );
  XNOR2_X2 MULT_mult_6_U4331 ( .A(MULT_mult_6_CARRYB_19__8_), .B(
        MULT_mult_6_ab_20__8_), .ZN(MULT_mult_6_n1754) );
  XNOR2_X2 MULT_mult_6_U4330 ( .A(MULT_mult_6_n1754), .B(MULT_mult_6_net89289), 
        .ZN(MULT_mult_6_SUMB_20__8_) );
  XNOR2_X2 MULT_mult_6_U4329 ( .A(MULT_mult_6_CARRYB_2__14_), .B(
        MULT_mult_6_ab_3__14_), .ZN(MULT_mult_6_n1792) );
  XNOR2_X2 MULT_mult_6_U4328 ( .A(MULT_mult_6_SUMB_11__14_), .B(
        MULT_mult_6_n1753), .ZN(MULT_mult_6_SUMB_12__13_) );
  NAND3_X2 MULT_mult_6_U4327 ( .A1(MULT_mult_6_n2003), .A2(MULT_mult_6_n2002), 
        .A3(MULT_mult_6_n1700), .ZN(MULT_mult_6_CARRYB_7__9_) );
  INV_X1 MULT_mult_6_U4326 ( .A(MULT_mult_6_ab_7__15_), .ZN(MULT_mult_6_n2043)
         );
  INV_X8 MULT_mult_6_U4325 ( .A(MULT_mult_6_CARRYB_6__15_), .ZN(
        MULT_mult_6_n1750) );
  NAND2_X4 MULT_mult_6_U4324 ( .A1(MULT_mult_6_n1751), .A2(MULT_mult_6_n1752), 
        .ZN(MULT_mult_6_n2204) );
  NAND2_X4 MULT_mult_6_U4323 ( .A1(MULT_mult_6_n1750), .A2(MULT_mult_6_n1749), 
        .ZN(MULT_mult_6_n1752) );
  NAND2_X2 MULT_mult_6_U4322 ( .A1(MULT_mult_6_n2043), .A2(
        MULT_mult_6_CARRYB_6__15_), .ZN(MULT_mult_6_n1751) );
  NOR2_X1 MULT_mult_6_U4321 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__13_) );
  NOR2_X1 MULT_mult_6_U4320 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__13_) );
  NOR2_X1 MULT_mult_6_U4319 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net70461), .ZN(MULT_mult_6_ab_17__13_) );
  NOR2_X1 MULT_mult_6_U4318 ( .A1(MULT_mult_6_net70459), .A2(
        MULT_mult_6_net70460), .ZN(MULT_mult_6_ab_18__13_) );
  NAND2_X2 MULT_mult_6_U4317 ( .A1(MULT_mult_6_ab_6__10_), .A2(
        MULT_mult_6_CARRYB_5__10_), .ZN(MULT_mult_6_n1747) );
  NAND2_X1 MULT_mult_6_U4316 ( .A1(MULT_mult_6_ab_5__10_), .A2(
        MULT_mult_6_CARRYB_4__10_), .ZN(MULT_mult_6_n1744) );
  NAND2_X2 MULT_mult_6_U4315 ( .A1(MULT_mult_6_ab_9__14_), .A2(
        MULT_mult_6_n1235), .ZN(MULT_mult_6_n2294) );
  XNOR2_X2 MULT_mult_6_U4314 ( .A(MULT_mult_6_n1743), .B(MULT_mult_6_net89255), 
        .ZN(MULT_mult_6_SUMB_15__9_) );
  XNOR2_X2 MULT_mult_6_U4313 ( .A(MULT_mult_6_n1741), .B(
        MULT_mult_6_SUMB_4__17_), .ZN(MULT_mult_6_SUMB_5__16_) );
  NAND2_X1 MULT_mult_6_U4312 ( .A1(MULT_mult_6_ab_3__21_), .A2(
        MULT_mult_6_CARRYB_2__21_), .ZN(MULT_mult_6_n1933) );
  INV_X2 MULT_mult_6_U4311 ( .A(MULT_mult_6_net83357), .ZN(
        MULT_mult_6_net83358) );
  NOR2_X2 MULT_mult_6_U4310 ( .A1(MULT_mult_6_net80727), .A2(
        MULT_mult_6_net77964), .ZN(MULT_mult_6_ab_3__20_) );
  INV_X4 MULT_mult_6_U4309 ( .A(MULT_mult_6_CARRYB_2__20_), .ZN(
        MULT_mult_6_n1739) );
  INV_X4 MULT_mult_6_U4308 ( .A(MULT_mult_6_ab_3__20_), .ZN(MULT_mult_6_n1738)
         );
  XNOR2_X2 MULT_mult_6_U4307 ( .A(MULT_mult_6_ab_4__20_), .B(
        MULT_mult_6_CARRYB_3__20_), .ZN(MULT_mult_6_n1737) );
  XNOR2_X2 MULT_mult_6_U4306 ( .A(MULT_mult_6_n1737), .B(
        MULT_mult_6_SUMB_3__21_), .ZN(MULT_mult_6_SUMB_4__20_) );
  XNOR2_X2 MULT_mult_6_U4305 ( .A(MULT_mult_6_n1736), .B(
        MULT_mult_6_SUMB_7__16_), .ZN(MULT_mult_6_SUMB_8__15_) );
  NAND2_X4 MULT_mult_6_U4304 ( .A1(MULT_mult_6_ab_6__16_), .A2(
        MULT_mult_6_CARRYB_5__16_), .ZN(MULT_mult_6_n2205) );
  INV_X4 MULT_mult_6_U4303 ( .A(MULT_mult_6_CARRYB_3__19_), .ZN(
        MULT_mult_6_n1817) );
  NAND3_X4 MULT_mult_6_U4302 ( .A1(MULT_mult_6_n1913), .A2(MULT_mult_6_n1912), 
        .A3(MULT_mult_6_n1911), .ZN(MULT_mult_6_CARRYB_19__2_) );
  INV_X4 MULT_mult_6_U4301 ( .A(MULT_mult_6_n1734), .ZN(MULT_mult_6_n1735) );
  NAND2_X4 MULT_mult_6_U4300 ( .A1(MULT_mult_6_n1735), .A2(
        MULT_mult_6_net82760), .ZN(MULT_mult_6_CARRYB_4__12_) );
  XNOR2_X2 MULT_mult_6_U4299 ( .A(MULT_mult_6_n288), .B(MULT_mult_6_n2014), 
        .ZN(MULT_mult_6_SUMB_7__8_) );
  XNOR2_X2 MULT_mult_6_U4298 ( .A(MULT_mult_6_n1193), .B(MULT_mult_6_ab_12__6_), .ZN(MULT_mult_6_n1764) );
  NAND2_X1 MULT_mult_6_U4297 ( .A1(MULT_mult_6_ab_7__16_), .A2(
        MULT_mult_6_CARRYB_6__16_), .ZN(MULT_mult_6_n2249) );
  NAND2_X2 MULT_mult_6_U4296 ( .A1(MULT_mult_6_ab_7__9_), .A2(
        MULT_mult_6_SUMB_6__10_), .ZN(MULT_mult_6_n2002) );
  NAND2_X2 MULT_mult_6_U4295 ( .A1(MULT_mult_6_SUMB_12__6_), .A2(
        MULT_mult_6_CARRYB_12__5_), .ZN(MULT_mult_6_n1922) );
  NAND2_X2 MULT_mult_6_U4294 ( .A1(MULT_mult_6_SUMB_12__8_), .A2(
        MULT_mult_6_CARRYB_12__7_), .ZN(MULT_mult_6_n2024) );
  XNOR2_X2 MULT_mult_6_U4293 ( .A(MULT_mult_6_SUMB_13__13_), .B(
        MULT_mult_6_net83535), .ZN(MULT_mult_6_SUMB_14__12_) );
  XNOR2_X2 MULT_mult_6_U4292 ( .A(MULT_mult_6_CARRYB_4__17_), .B(
        MULT_mult_6_ab_5__17_), .ZN(MULT_mult_6_n1729) );
  XNOR2_X2 MULT_mult_6_U4291 ( .A(MULT_mult_6_SUMB_4__18_), .B(
        MULT_mult_6_n1729), .ZN(MULT_mult_6_SUMB_5__17_) );
  NAND2_X2 MULT_mult_6_U4290 ( .A1(MULT_mult_6_ab_17__5_), .A2(
        MULT_mult_6_n1201), .ZN(MULT_mult_6_n2037) );
  NAND2_X4 MULT_mult_6_U4289 ( .A1(MULT_mult_6_n1848), .A2(MULT_mult_6_n1849), 
        .ZN(MULT_mult_6_n2095) );
  INV_X2 MULT_mult_6_U4288 ( .A(MULT_mult_6_n1733), .ZN(MULT_mult_6_n1726) );
  NAND2_X4 MULT_mult_6_U4287 ( .A1(MULT_mult_6_n1725), .A2(MULT_mult_6_n1726), 
        .ZN(MULT_mult_6_n1728) );
  NAND3_X2 MULT_mult_6_U4286 ( .A1(MULT_mult_6_n1722), .A2(MULT_mult_6_n1723), 
        .A3(MULT_mult_6_n1724), .ZN(MULT_mult_6_CARRYB_4__18_) );
  NAND2_X2 MULT_mult_6_U4285 ( .A1(MULT_mult_6_ab_4__18_), .A2(
        MULT_mult_6_CARRYB_3__18_), .ZN(MULT_mult_6_n1723) );
  NAND2_X2 MULT_mult_6_U4284 ( .A1(MULT_mult_6_CARRYB_18__4_), .A2(
        MULT_mult_6_ab_19__4_), .ZN(MULT_mult_6_n1859) );
  INV_X2 MULT_mult_6_U4283 ( .A(MULT_mult_6_ab_4__19_), .ZN(MULT_mult_6_n1888)
         );
  NAND2_X2 MULT_mult_6_U4282 ( .A1(MULT_mult_6_n1888), .A2(
        MULT_mult_6_CARRYB_3__19_), .ZN(MULT_mult_6_n1818) );
  NOR2_X1 MULT_mult_6_U4281 ( .A1(MULT_mult_6_net84358), .A2(
        MULT_mult_6_net77956), .ZN(MULT_mult_6_ab_4__23_) );
  NOR2_X1 MULT_mult_6_U4280 ( .A1(MULT_mult_6_net84358), .A2(
        MULT_mult_6_net77932), .ZN(MULT_mult_6_ab_7__23_) );
  NOR2_X1 MULT_mult_6_U4279 ( .A1(MULT_mult_6_net77926), .A2(
        MULT_mult_6_net84358), .ZN(MULT_mult_6_ab_8__23_) );
  XNOR2_X2 MULT_mult_6_U4278 ( .A(MULT_mult_6_n1717), .B(MULT_mult_6_n1249), 
        .ZN(MULT_mult_6_SUMB_11__7_) );
  NAND2_X2 MULT_mult_6_U4277 ( .A1(MULT_mult_6_ab_3__17_), .A2(
        MULT_mult_6_SUMB_2__18_), .ZN(MULT_mult_6_n1715) );
  INV_X1 MULT_mult_6_U4276 ( .A(MULT_mult_6_ab_9__15_), .ZN(MULT_mult_6_n1708)
         );
  NAND2_X2 MULT_mult_6_U4275 ( .A1(MULT_mult_6_ab_5__18_), .A2(
        MULT_mult_6_n1768), .ZN(MULT_mult_6_n2139) );
  NAND2_X1 MULT_mult_6_U4274 ( .A1(MULT_mult_6_ab_10__18_), .A2(
        MULT_mult_6_SUMB_9__19_), .ZN(MULT_mult_6_n1875) );
  NOR2_X1 MULT_mult_6_U4273 ( .A1(MULT_mult_6_net81424), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__15_) );
  NAND2_X2 MULT_mult_6_U4272 ( .A1(MULT_mult_6_CARRYB_4__17_), .A2(
        MULT_mult_6_SUMB_4__18_), .ZN(MULT_mult_6_n2201) );
  NAND2_X2 MULT_mult_6_U4271 ( .A1(MULT_mult_6_ab_13__6_), .A2(
        MULT_mult_6_n553), .ZN(MULT_mult_6_n2000) );
  NAND2_X2 MULT_mult_6_U4270 ( .A1(MULT_mult_6_CARRYB_17__4_), .A2(
        MULT_mult_6_SUMB_17__5_), .ZN(MULT_mult_6_n2042) );
  XNOR2_X2 MULT_mult_6_U4269 ( .A(MULT_mult_6_CARRYB_14__5_), .B(
        MULT_mult_6_ab_15__5_), .ZN(MULT_mult_6_n1721) );
  XNOR2_X2 MULT_mult_6_U4268 ( .A(MULT_mult_6_n1500), .B(MULT_mult_6_ab_16__4_), .ZN(MULT_mult_6_n1731) );
  NAND2_X2 MULT_mult_6_U4267 ( .A1(MULT_mult_6_SUMB_8__6_), .A2(
        MULT_mult_6_ab_9__5_), .ZN(MULT_mult_6_n1787) );
  NAND2_X2 MULT_mult_6_U4266 ( .A1(MULT_mult_6_SUMB_17__5_), .A2(
        MULT_mult_6_ab_18__4_), .ZN(MULT_mult_6_n2041) );
  NAND2_X2 MULT_mult_6_U4265 ( .A1(MULT_mult_6_ab_14__5_), .A2(
        MULT_mult_6_SUMB_13__6_), .ZN(MULT_mult_6_n1703) );
  INV_X1 MULT_mult_6_U4264 ( .A(MULT_mult_6_ab_7__9_), .ZN(MULT_mult_6_n1698)
         );
  NAND2_X1 MULT_mult_6_U4263 ( .A1(MULT_mult_6_ab_27__3_), .A2(
        MULT_mult_6_SUMB_26__4_), .ZN(MULT_mult_6_net80817) );
  NAND3_X4 MULT_mult_6_U4262 ( .A1(MULT_mult_6_n1977), .A2(MULT_mult_6_n1979), 
        .A3(MULT_mult_6_n1978), .ZN(MULT_mult_6_CARRYB_15__5_) );
  NAND2_X2 MULT_mult_6_U4261 ( .A1(MULT_mult_6_n1222), .A2(
        MULT_mult_6_CARRYB_14__3_), .ZN(MULT_mult_6_n1990) );
  NAND3_X4 MULT_mult_6_U4260 ( .A1(MULT_mult_6_n2088), .A2(MULT_mult_6_n2087), 
        .A3(MULT_mult_6_n2086), .ZN(MULT_mult_6_CARRYB_9__8_) );
  NAND2_X1 MULT_mult_6_U4259 ( .A1(MULT_mult_6_CARRYB_18__11_), .A2(
        MULT_mult_6_SUMB_18__12_), .ZN(MULT_mult_6_n2258) );
  XNOR2_X2 MULT_mult_6_U4258 ( .A(MULT_mult_6_CARRYB_13__15_), .B(
        MULT_mult_6_ab_14__15_), .ZN(MULT_mult_6_n1697) );
  XNOR2_X2 MULT_mult_6_U4257 ( .A(MULT_mult_6_SUMB_13__16_), .B(
        MULT_mult_6_n1697), .ZN(MULT_mult_6_SUMB_14__15_) );
  INV_X1 MULT_mult_6_U4256 ( .A(MULT_mult_6_ab_26__3_), .ZN(
        MULT_mult_6_net83797) );
  XNOR2_X2 MULT_mult_6_U4255 ( .A(MULT_mult_6_n1695), .B(MULT_mult_6_n1119), 
        .ZN(MULT_mult_6_SUMB_6__15_) );
  NAND2_X1 MULT_mult_6_U4254 ( .A1(MULT_mult_6_ab_6__23_), .A2(
        MULT_mult_6_n1231), .ZN(MULT_mult_6_n2180) );
  NOR2_X2 MULT_mult_6_U4253 ( .A1(MULT_mult_6_net84358), .A2(
        MULT_mult_6_net77940), .ZN(MULT_mult_6_ab_6__23_) );
  NAND3_X2 MULT_mult_6_U4252 ( .A1(MULT_mult_6_n1689), .A2(MULT_mult_6_n1690), 
        .A3(MULT_mult_6_n1691), .ZN(MULT_mult_6_CARRYB_10__20_) );
  NAND2_X1 MULT_mult_6_U4251 ( .A1(MULT_mult_6_CARRYB_9__20_), .A2(
        MULT_mult_6_SUMB_9__21_), .ZN(MULT_mult_6_n1691) );
  NAND2_X1 MULT_mult_6_U4250 ( .A1(MULT_mult_6_ab_10__20_), .A2(
        MULT_mult_6_SUMB_9__21_), .ZN(MULT_mult_6_n1690) );
  NAND2_X1 MULT_mult_6_U4249 ( .A1(MULT_mult_6_ab_10__20_), .A2(
        MULT_mult_6_CARRYB_9__20_), .ZN(MULT_mult_6_n1689) );
  NAND3_X2 MULT_mult_6_U4248 ( .A1(MULT_mult_6_n1686), .A2(MULT_mult_6_n1687), 
        .A3(MULT_mult_6_n1688), .ZN(MULT_mult_6_CARRYB_9__21_) );
  NAND2_X1 MULT_mult_6_U4247 ( .A1(MULT_mult_6_ab_9__21_), .A2(
        MULT_mult_6_CARRYB_8__21_), .ZN(MULT_mult_6_n1686) );
  NAND3_X4 MULT_mult_6_U4246 ( .A1(MULT_mult_6_n2140), .A2(MULT_mult_6_n2141), 
        .A3(MULT_mult_6_n2139), .ZN(MULT_mult_6_CARRYB_5__18_) );
  NAND3_X4 MULT_mult_6_U4245 ( .A1(MULT_mult_6_n1680), .A2(MULT_mult_6_n1681), 
        .A3(MULT_mult_6_n1682), .ZN(MULT_mult_6_CARRYB_6__18_) );
  NAND2_X2 MULT_mult_6_U4244 ( .A1(MULT_mult_6_ab_6__18_), .A2(
        MULT_mult_6_CARRYB_5__18_), .ZN(MULT_mult_6_n1682) );
  NAND2_X2 MULT_mult_6_U4243 ( .A1(MULT_mult_6_CARRYB_5__18_), .A2(
        MULT_mult_6_SUMB_5__19_), .ZN(MULT_mult_6_n1680) );
  NAND3_X4 MULT_mult_6_U4242 ( .A1(MULT_mult_6_n2121), .A2(MULT_mult_6_n2120), 
        .A3(MULT_mult_6_n2122), .ZN(MULT_mult_6_CARRYB_14__12_) );
  NAND3_X2 MULT_mult_6_U4241 ( .A1(MULT_mult_6_n1919), .A2(MULT_mult_6_n1918), 
        .A3(MULT_mult_6_n1917), .ZN(MULT_mult_6_CARRYB_12__6_) );
  NAND2_X2 MULT_mult_6_U4240 ( .A1(MULT_mult_6_n854), .A2(
        MULT_mult_6_ab_13__6_), .ZN(MULT_mult_6_n1999) );
  NAND2_X2 MULT_mult_6_U4239 ( .A1(MULT_mult_6_CARRYB_12__6_), .A2(
        MULT_mult_6_SUMB_12__7_), .ZN(MULT_mult_6_n1998) );
  NAND2_X2 MULT_mult_6_U4238 ( .A1(MULT_mult_6_CARRYB_6__9_), .A2(
        MULT_mult_6_ab_7__9_), .ZN(MULT_mult_6_n1700) );
  NOR2_X1 MULT_mult_6_U4237 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__3_) );
  NOR2_X2 MULT_mult_6_U4236 ( .A1(MULT_mult_6_net77866), .A2(
        MULT_mult_6_net70443), .ZN(MULT_mult_6_ab_26__1_) );
  NAND2_X2 MULT_mult_6_U4235 ( .A1(MULT_mult_6_ab_13__3_), .A2(
        MULT_mult_6_SUMB_12__4_), .ZN(MULT_mult_6_n1677) );
  NAND2_X2 MULT_mult_6_U4234 ( .A1(MULT_mult_6_CARRYB_12__3_), .A2(
        MULT_mult_6_SUMB_12__4_), .ZN(MULT_mult_6_n1676) );
  NAND2_X2 MULT_mult_6_U4233 ( .A1(MULT_mult_6_ab_11__3_), .A2(
        MULT_mult_6_SUMB_10__4_), .ZN(MULT_mult_6_n1671) );
  NAND2_X1 MULT_mult_6_U4232 ( .A1(MULT_mult_6_ab_11__3_), .A2(
        MULT_mult_6_CARRYB_10__3_), .ZN(MULT_mult_6_n1670) );
  NAND3_X4 MULT_mult_6_U4231 ( .A1(MULT_mult_6_n1668), .A2(MULT_mult_6_n1669), 
        .A3(MULT_mult_6_n1667), .ZN(MULT_mult_6_CARRYB_17__2_) );
  NAND2_X2 MULT_mult_6_U4230 ( .A1(MULT_mult_6_ab_17__2_), .A2(
        MULT_mult_6_SUMB_16__3_), .ZN(MULT_mult_6_n1667) );
  NAND3_X4 MULT_mult_6_U4229 ( .A1(MULT_mult_6_n1666), .A2(MULT_mult_6_n1665), 
        .A3(MULT_mult_6_n1664), .ZN(MULT_mult_6_CARRYB_16__2_) );
  NAND2_X2 MULT_mult_6_U4228 ( .A1(MULT_mult_6_CARRYB_15__2_), .A2(
        MULT_mult_6_SUMB_15__3_), .ZN(MULT_mult_6_n1666) );
  NAND2_X2 MULT_mult_6_U4227 ( .A1(MULT_mult_6_ab_16__2_), .A2(
        MULT_mult_6_SUMB_15__3_), .ZN(MULT_mult_6_n1665) );
  NAND2_X2 MULT_mult_6_U4226 ( .A1(MULT_mult_6_ab_16__2_), .A2(
        MULT_mult_6_CARRYB_15__2_), .ZN(MULT_mult_6_n1664) );
  XNOR2_X2 MULT_mult_6_U4225 ( .A(MULT_mult_6_SUMB_3__19_), .B(
        MULT_mult_6_ab_4__18_), .ZN(MULT_mult_6_n1693) );
  XNOR2_X2 MULT_mult_6_U4224 ( .A(MULT_mult_6_CARRYB_20__9_), .B(
        MULT_mult_6_ab_21__9_), .ZN(MULT_mult_6_n1663) );
  XNOR2_X2 MULT_mult_6_U4223 ( .A(MULT_mult_6_n1663), .B(MULT_mult_6_n568), 
        .ZN(MULT_mult_6_SUMB_21__9_) );
  NAND3_X4 MULT_mult_6_U4222 ( .A1(MULT_mult_6_n1895), .A2(MULT_mult_6_n1894), 
        .A3(MULT_mult_6_n1893), .ZN(MULT_mult_6_CARRYB_4__17_) );
  INV_X4 MULT_mult_6_U4221 ( .A(MULT_mult_6_ab_8__11_), .ZN(MULT_mult_6_n1838)
         );
  INV_X4 MULT_mult_6_U4220 ( .A(MULT_mult_6_n1838), .ZN(MULT_mult_6_n1660) );
  NAND2_X4 MULT_mult_6_U4219 ( .A1(MULT_mult_6_n1659), .A2(MULT_mult_6_n1660), 
        .ZN(MULT_mult_6_n1662) );
  NAND2_X2 MULT_mult_6_U4218 ( .A1(MULT_mult_6_CARRYB_7__11_), .A2(
        MULT_mult_6_n1838), .ZN(MULT_mult_6_n1661) );
  NAND3_X4 MULT_mult_6_U4217 ( .A1(MULT_mult_6_n1657), .A2(MULT_mult_6_n1656), 
        .A3(MULT_mult_6_n1655), .ZN(MULT_mult_6_CARRYB_3__9_) );
  NAND2_X2 MULT_mult_6_U4216 ( .A1(MULT_mult_6_ab_3__9_), .A2(
        MULT_mult_6_SUMB_2__10_), .ZN(MULT_mult_6_n1657) );
  NAND2_X2 MULT_mult_6_U4215 ( .A1(MULT_mult_6_n1246), .A2(
        MULT_mult_6_SUMB_2__10_), .ZN(MULT_mult_6_n1656) );
  NAND3_X2 MULT_mult_6_U4214 ( .A1(MULT_mult_6_n1652), .A2(MULT_mult_6_n1653), 
        .A3(MULT_mult_6_n1654), .ZN(MULT_mult_6_CARRYB_2__10_) );
  XOR2_X2 MULT_mult_6_U4213 ( .A(MULT_mult_6_n1651), .B(
        MULT_mult_6_SUMB_1__11_), .Z(MULT_mult_6_SUMB_2__10_) );
  NOR2_X4 MULT_mult_6_U4212 ( .A1(MULT_mult_6_n392), .A2(MULT_mult_6_net70452), 
        .ZN(MULT_mult_6_ab_0__9_) );
  XNOR2_X2 MULT_mult_6_U4211 ( .A(MULT_mult_6_ab_4__7_), .B(
        MULT_mult_6_CARRYB_3__7_), .ZN(MULT_mult_6_n1649) );
  NAND2_X4 MULT_mult_6_U4210 ( .A1(MULT_mult_6_n1700), .A2(MULT_mult_6_n1701), 
        .ZN(MULT_mult_6_n1820) );
  NOR2_X2 MULT_mult_6_U4209 ( .A1(MULT_mult_6_net77912), .A2(
        MULT_mult_6_net77966), .ZN(MULT_mult_6_ab_3__7_) );
  INV_X4 MULT_mult_6_U4208 ( .A(MULT_mult_6_CARRYB_25__3_), .ZN(
        MULT_mult_6_net83796) );
  NOR2_X4 MULT_mult_6_U4207 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__4_) );
  NAND3_X4 MULT_mult_6_U4206 ( .A1(MULT_mult_6_n1647), .A2(MULT_mult_6_n1646), 
        .A3(MULT_mult_6_n1645), .ZN(MULT_mult_6_CARRYB_3__10_) );
  NAND2_X2 MULT_mult_6_U4205 ( .A1(MULT_mult_6_SUMB_2__11_), .A2(
        MULT_mult_6_n1203), .ZN(MULT_mult_6_n1647) );
  NAND2_X2 MULT_mult_6_U4204 ( .A1(MULT_mult_6_SUMB_2__11_), .A2(
        MULT_mult_6_ab_3__10_), .ZN(MULT_mult_6_n1646) );
  NAND3_X4 MULT_mult_6_U4203 ( .A1(MULT_mult_6_n1638), .A2(MULT_mult_6_n1637), 
        .A3(MULT_mult_6_n1636), .ZN(MULT_mult_6_CARRYB_12__5_) );
  NAND2_X2 MULT_mult_6_U4202 ( .A1(MULT_mult_6_n1275), .A2(
        MULT_mult_6_CARRYB_11__5_), .ZN(MULT_mult_6_n1638) );
  INV_X1 MULT_mult_6_U4201 ( .A(MULT_mult_6_ab_14__4_), .ZN(MULT_mult_6_n1632)
         );
  NAND2_X2 MULT_mult_6_U4200 ( .A1(MULT_mult_6_ab_6__15_), .A2(
        MULT_mult_6_n847), .ZN(MULT_mult_6_n2032) );
  NAND2_X2 MULT_mult_6_U4199 ( .A1(MULT_mult_6_n1187), .A2(MULT_mult_6_n1881), 
        .ZN(MULT_mult_6_n1848) );
  NAND2_X4 MULT_mult_6_U4198 ( .A1(MULT_mult_6_n1630), .A2(MULT_mult_6_n1629), 
        .ZN(MULT_mult_6_SUMB_13__12_) );
  XOR2_X2 MULT_mult_6_U4197 ( .A(MULT_mult_6_net82532), .B(
        MULT_mult_6_SUMB_16__2_), .Z(MULT_mult_6_SUMB_17__1_) );
  NAND2_X1 MULT_mult_6_U4196 ( .A1(MULT_mult_6_ab_18__12_), .A2(
        MULT_mult_6_SUMB_17__13_), .ZN(MULT_mult_6_n2255) );
  XNOR2_X2 MULT_mult_6_U4195 ( .A(MULT_mult_6_SUMB_6__23_), .B(
        MULT_mult_6_n1626), .ZN(MULT_mult_6_SUMB_7__22_) );
  XNOR2_X2 MULT_mult_6_U4194 ( .A(MULT_mult_6_CARRYB_4__23_), .B(
        MULT_mult_6_ab_5__23_), .ZN(MULT_mult_6_n1625) );
  XNOR2_X2 MULT_mult_6_U4193 ( .A(MULT_mult_6_SUMB_4__24_), .B(
        MULT_mult_6_n1625), .ZN(MULT_mult_6_SUMB_5__23_) );
  NAND3_X2 MULT_mult_6_U4192 ( .A1(MULT_mult_6_net80838), .A2(
        MULT_mult_6_net80839), .A3(MULT_mult_6_net80840), .ZN(
        MULT_mult_6_CARRYB_5__15_) );
  NAND2_X2 MULT_mult_6_U4191 ( .A1(MULT_mult_6_ab_16__14_), .A2(
        MULT_mult_6_CARRYB_15__14_), .ZN(MULT_mult_6_n1952) );
  NAND3_X4 MULT_mult_6_U4190 ( .A1(MULT_mult_6_net84308), .A2(
        MULT_mult_6_net84309), .A3(MULT_mult_6_n1623), .ZN(
        MULT_mult_6_CARRYB_15__14_) );
  NAND2_X1 MULT_mult_6_U4189 ( .A1(MULT_mult_6_ab_15__14_), .A2(
        MULT_mult_6_CARRYB_14__14_), .ZN(MULT_mult_6_n1623) );
  NAND2_X4 MULT_mult_6_U4188 ( .A1(MULT_mult_6_net84305), .A2(
        MULT_mult_6_n1622), .ZN(MULT_mult_6_SUMB_25__5_) );
  NAND3_X4 MULT_mult_6_U4187 ( .A1(MULT_mult_6_net84302), .A2(
        MULT_mult_6_net84301), .A3(MULT_mult_6_net84300), .ZN(
        MULT_mult_6_CARRYB_3__23_) );
  XNOR2_X2 MULT_mult_6_U4186 ( .A(MULT_mult_6_n1207), .B(MULT_mult_6_ab_3__12_), .ZN(MULT_mult_6_n1928) );
  XNOR2_X2 MULT_mult_6_U4185 ( .A(MULT_mult_6_CARRYB_7__9_), .B(
        MULT_mult_6_ab_8__9_), .ZN(MULT_mult_6_n1836) );
  NAND3_X4 MULT_mult_6_U4184 ( .A1(MULT_mult_6_net80350), .A2(
        MULT_mult_6_net80348), .A3(MULT_mult_6_net80349), .ZN(
        MULT_mult_6_CARRYB_9__13_) );
  NOR2_X1 MULT_mult_6_U4183 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__9_) );
  NAND2_X4 MULT_mult_6_U4182 ( .A1(MULT_mult_6_n1756), .A2(MULT_mult_6_n1757), 
        .ZN(MULT_mult_6_SUMB_13__8_) );
  NAND3_X4 MULT_mult_6_U4181 ( .A1(MULT_mult_6_net81066), .A2(
        MULT_mult_6_net81065), .A3(MULT_mult_6_n2118), .ZN(
        MULT_mult_6_CARRYB_18__7_) );
  INV_X1 MULT_mult_6_U4180 ( .A(MULT_mult_6_ab_19__7_), .ZN(MULT_mult_6_n1614)
         );
  NAND3_X4 MULT_mult_6_U4179 ( .A1(MULT_mult_6_n2158), .A2(
        MULT_mult_6_net80836), .A3(MULT_mult_6_net80835), .ZN(
        MULT_mult_6_CARRYB_4__16_) );
  NAND2_X2 MULT_mult_6_U4178 ( .A1(MULT_mult_6_CARRYB_18__7_), .A2(
        MULT_mult_6_SUMB_18__8_), .ZN(MULT_mult_6_n2012) );
  NAND2_X2 MULT_mult_6_U4177 ( .A1(MULT_mult_6_CARRYB_13__3_), .A2(
        MULT_mult_6_SUMB_13__4_), .ZN(MULT_mult_6_n1969) );
  NAND2_X2 MULT_mult_6_U4176 ( .A1(MULT_mult_6_n1424), .A2(
        MULT_mult_6_SUMB_1__21_), .ZN(MULT_mult_6_n1684) );
  INV_X1 MULT_mult_6_U4175 ( .A(MULT_mult_6_ab_7__16_), .ZN(MULT_mult_6_n1900)
         );
  INV_X4 MULT_mult_6_U4174 ( .A(MULT_mult_6_CARRYB_6__16_), .ZN(
        MULT_mult_6_n1611) );
  INV_X4 MULT_mult_6_U4173 ( .A(MULT_mult_6_n1900), .ZN(MULT_mult_6_n1610) );
  NAND2_X4 MULT_mult_6_U4172 ( .A1(MULT_mult_6_n1611), .A2(MULT_mult_6_n1610), 
        .ZN(MULT_mult_6_n1613) );
  NAND2_X2 MULT_mult_6_U4171 ( .A1(MULT_mult_6_n1900), .A2(
        MULT_mult_6_CARRYB_6__16_), .ZN(MULT_mult_6_n1612) );
  XNOR2_X2 MULT_mult_6_U4170 ( .A(MULT_mult_6_ab_3__21_), .B(
        MULT_mult_6_CARRYB_2__21_), .ZN(MULT_mult_6_n1609) );
  XNOR2_X2 MULT_mult_6_U4169 ( .A(MULT_mult_6_n557), .B(MULT_mult_6_n866), 
        .ZN(MULT_mult_6_SUMB_3__21_) );
  XNOR2_X2 MULT_mult_6_U4168 ( .A(MULT_mult_6_ab_8__16_), .B(
        MULT_mult_6_CARRYB_7__16_), .ZN(MULT_mult_6_n1608) );
  XNOR2_X2 MULT_mult_6_U4167 ( .A(MULT_mult_6_CARRYB_13__6_), .B(
        MULT_mult_6_n1607), .ZN(MULT_mult_6_n1973) );
  NAND2_X1 MULT_mult_6_U4166 ( .A1(MULT_mult_6_ab_5__16_), .A2(
        MULT_mult_6_CARRYB_4__16_), .ZN(MULT_mult_6_n1896) );
  INV_X8 MULT_mult_6_U4165 ( .A(MULT_mult_6_n2342), .ZN(
        MULT_mult_6_SUMB_1__20_) );
  XNOR2_X2 MULT_mult_6_U4164 ( .A(MULT_mult_6_SUMB_12__15_), .B(
        MULT_mult_6_net84481), .ZN(MULT_mult_6_SUMB_13__14_) );
  NAND2_X4 MULT_mult_6_U4163 ( .A1(MULT_mult_6_n1612), .A2(MULT_mult_6_n1613), 
        .ZN(MULT_mult_6_n2248) );
  XNOR2_X2 MULT_mult_6_U4162 ( .A(MULT_mult_6_ab_19__11_), .B(
        MULT_mult_6_CARRYB_18__11_), .ZN(MULT_mult_6_n1606) );
  INV_X4 MULT_mult_6_U4161 ( .A(MULT_mult_6_n1766), .ZN(MULT_mult_6_n1603) );
  NAND2_X4 MULT_mult_6_U4160 ( .A1(MULT_mult_6_n1597), .A2(MULT_mult_6_n1598), 
        .ZN(MULT_mult_6_SUMB_25__4_) );
  NAND2_X4 MULT_mult_6_U4159 ( .A1(MULT_mult_6_n340), .A2(MULT_mult_6_n1596), 
        .ZN(MULT_mult_6_n1598) );
  NAND2_X2 MULT_mult_6_U4158 ( .A1(MULT_mult_6_n1301), .A2(MULT_mult_6_n145), 
        .ZN(MULT_mult_6_n1597) );
  NAND2_X2 MULT_mult_6_U4157 ( .A1(MULT_mult_6_CARRYB_8__20_), .A2(
        MULT_mult_6_n1278), .ZN(MULT_mult_6_n2218) );
  NAND3_X4 MULT_mult_6_U4156 ( .A1(MULT_mult_6_n2218), .A2(MULT_mult_6_n2217), 
        .A3(MULT_mult_6_n2216), .ZN(MULT_mult_6_CARRYB_9__20_) );
  NAND2_X4 MULT_mult_6_U4155 ( .A1(MULT_mult_6_n1594), .A2(MULT_mult_6_n1595), 
        .ZN(MULT_mult_6_SUMB_7__16_) );
  NAND2_X2 MULT_mult_6_U4154 ( .A1(MULT_mult_6_ab_0__13_), .A2(
        MULT_mult_6_n237), .ZN(MULT_mult_6_n2336) );
  INV_X1 MULT_mult_6_U4153 ( .A(MULT_mult_6_ab_6__10_), .ZN(MULT_mult_6_n1589)
         );
  XNOR2_X2 MULT_mult_6_U4152 ( .A(MULT_mult_6_n1587), .B(
        MULT_mult_6_SUMB_8__15_), .ZN(MULT_mult_6_SUMB_9__14_) );
  NAND2_X2 MULT_mult_6_U4151 ( .A1(MULT_mult_6_ab_2__21_), .A2(
        MULT_mult_6_n1692), .ZN(MULT_mult_6_n2190) );
  NAND2_X2 MULT_mult_6_U4150 ( .A1(MULT_mult_6_SUMB_18__1_), .A2(
        MULT_mult_6_CARRYB_18__0_), .ZN(MULT_mult_6_n1815) );
  XOR2_X1 MULT_mult_6_U4149 ( .A(MULT_mult_6_n1812), .B(
        MULT_mult_6_CARRYB_18__0_), .Z(multOut[12]) );
  NAND2_X2 MULT_mult_6_U4148 ( .A1(MULT_mult_6_ab_2__22_), .A2(
        MULT_mult_6_SUMB_1__23_), .ZN(MULT_mult_6_n1931) );
  NAND2_X2 MULT_mult_6_U4147 ( .A1(MULT_mult_6_CARRYB_1__22_), .A2(
        MULT_mult_6_SUMB_1__23_), .ZN(MULT_mult_6_n1932) );
  XNOR2_X2 MULT_mult_6_U4146 ( .A(MULT_mult_6_CARRYB_11__5_), .B(
        MULT_mult_6_ab_12__5_), .ZN(MULT_mult_6_n1586) );
  XNOR2_X2 MULT_mult_6_U4145 ( .A(MULT_mult_6_n1586), .B(MULT_mult_6_n1275), 
        .ZN(MULT_mult_6_SUMB_12__5_) );
  XNOR2_X2 MULT_mult_6_U4144 ( .A(MULT_mult_6_n1585), .B(MULT_mult_6_n1236), 
        .ZN(MULT_mult_6_SUMB_16__5_) );
  XNOR2_X2 MULT_mult_6_U4143 ( .A(MULT_mult_6_CARRYB_19__6_), .B(
        MULT_mult_6_ab_20__6_), .ZN(MULT_mult_6_net84348) );
  XNOR2_X2 MULT_mult_6_U4142 ( .A(MULT_mult_6_n1584), .B(MULT_mult_6_n1202), 
        .ZN(MULT_mult_6_SUMB_14__5_) );
  INV_X4 MULT_mult_6_U4141 ( .A(MULT_mult_6_net80694), .ZN(
        MULT_mult_6_net84711) );
  NAND2_X4 MULT_mult_6_U4140 ( .A1(MULT_mult_6_net84712), .A2(
        MULT_mult_6_n1583), .ZN(MULT_mult_6_n2243) );
  NAND2_X4 MULT_mult_6_U4139 ( .A1(MULT_mult_6_net84710), .A2(
        MULT_mult_6_net84711), .ZN(MULT_mult_6_n1583) );
  INV_X1 MULT_mult_6_U4138 ( .A(MULT_mult_6_ab_19__5_), .ZN(
        MULT_mult_6_net84706) );
  NAND2_X2 MULT_mult_6_U4137 ( .A1(MULT_mult_6_SUMB_8__15_), .A2(
        MULT_mult_6_ab_9__14_), .ZN(MULT_mult_6_n2293) );
  XNOR2_X2 MULT_mult_6_U4136 ( .A(MULT_mult_6_n1581), .B(MULT_mult_6_n1225), 
        .ZN(MULT_mult_6_SUMB_15__4_) );
  NOR2_X1 MULT_mult_6_U4135 ( .A1(MULT_mult_6_net91660), .A2(
        MULT_mult_6_net70461), .ZN(MULT_mult_6_ab_17__10_) );
  NAND2_X4 MULT_mult_6_U4134 ( .A1(MULT_mult_6_n1577), .A2(MULT_mult_6_n1578), 
        .ZN(MULT_mult_6_SUMB_5__18_) );
  NAND2_X1 MULT_mult_6_U4133 ( .A1(MULT_mult_6_ab_13__13_), .A2(
        MULT_mult_6_CARRYB_12__13_), .ZN(MULT_mult_6_n1573) );
  NAND2_X2 MULT_mult_6_U4132 ( .A1(MULT_mult_6_ab_18__7_), .A2(
        MULT_mult_6_net87619), .ZN(MULT_mult_6_n2118) );
  NAND3_X4 MULT_mult_6_U4131 ( .A1(MULT_mult_6_net82408), .A2(
        MULT_mult_6_net82407), .A3(MULT_mult_6_n1882), .ZN(
        MULT_mult_6_CARRYB_21__4_) );
  NAND2_X4 MULT_mult_6_U4130 ( .A1(MULT_mult_6_n1771), .A2(MULT_mult_6_n1772), 
        .ZN(MULT_mult_6_net81169) );
  XOR2_X1 MULT_mult_6_U4129 ( .A(MULT_mult_6_n2099), .B(
        MULT_mult_6_SUMB_19__1_), .Z(multOut[11]) );
  XNOR2_X2 MULT_mult_6_U4128 ( .A(MULT_mult_6_ab_3__27_), .B(
        MULT_mult_6_CARRYB_2__27_), .ZN(MULT_mult_6_n1572) );
  XNOR2_X2 MULT_mult_6_U4127 ( .A(MULT_mult_6_n1572), .B(
        MULT_mult_6_SUMB_2__28_), .ZN(MULT_mult_6_SUMB_3__27_) );
  NAND2_X4 MULT_mult_6_U4126 ( .A1(MULT_mult_6_net83796), .A2(
        MULT_mult_6_net83797), .ZN(MULT_mult_6_n1696) );
  NAND2_X2 MULT_mult_6_U4125 ( .A1(MULT_mult_6_n1769), .A2(
        MULT_mult_6_CARRYB_14__11_), .ZN(MULT_mult_6_n1772) );
  NOR2_X4 MULT_mult_6_U4124 ( .A1(MULT_mult_6_net70478), .A2(
        MULT_mult_6_net82149), .ZN(MULT_mult_6_ab_0__22_) );
  XNOR2_X2 MULT_mult_6_U4123 ( .A(MULT_mult_6_CARRYB_12__5_), .B(
        MULT_mult_6_ab_13__5_), .ZN(MULT_mult_6_n1837) );
  NAND2_X2 MULT_mult_6_U4122 ( .A1(MULT_mult_6_ab_22__0_), .A2(
        MULT_mult_6_CARRYB_21__0_), .ZN(MULT_mult_6_n1796) );
  NAND2_X2 MULT_mult_6_U4121 ( .A1(MULT_mult_6_ab_0__22_), .A2(
        MULT_mult_6_ab_1__21_), .ZN(MULT_mult_6_n2343) );
  NOR2_X2 MULT_mult_6_U4120 ( .A1(MULT_mult_6_net70492), .A2(
        MULT_mult_6_net83263), .ZN(MULT_mult_6_ab_1__29_) );
  NOR2_X2 MULT_mult_6_U4119 ( .A1(MULT_mult_6_net77858), .A2(
        MULT_mult_6_net70447), .ZN(MULT_mult_6_ab_24__0_) );
  NOR2_X1 MULT_mult_6_U4118 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net77938), .ZN(MULT_mult_6_ab_6__3_) );
  NAND2_X2 MULT_mult_6_U4117 ( .A1(MULT_mult_6_CARRYB_23__0_), .A2(
        MULT_mult_6_n23), .ZN(MULT_mult_6_n1568) );
  NAND2_X2 MULT_mult_6_U4116 ( .A1(MULT_mult_6_ab_6__3_), .A2(
        MULT_mult_6_SUMB_5__4_), .ZN(MULT_mult_6_n1565) );
  NAND3_X4 MULT_mult_6_U4115 ( .A1(MULT_mult_6_net81069), .A2(
        MULT_mult_6_net81068), .A3(MULT_mult_6_net81067), .ZN(
        MULT_mult_6_CARRYB_19__6_) );
  XNOR2_X2 MULT_mult_6_U4114 ( .A(MULT_mult_6_n1649), .B(
        MULT_mult_6_SUMB_3__8_), .ZN(MULT_mult_6_SUMB_4__7_) );
  NAND2_X4 MULT_mult_6_U4113 ( .A1(MULT_mult_6_net84212), .A2(
        MULT_mult_6_net84211), .ZN(MULT_mult_6_n1937) );
  NOR2_X1 MULT_mult_6_U4112 ( .A1(MULT_mult_6_net77948), .A2(
        MULT_mult_6_net70486), .ZN(MULT_mult_6_ab_5__26_) );
  NOR2_X1 MULT_mult_6_U4111 ( .A1(MULT_mult_6_net77940), .A2(
        MULT_mult_6_net82239), .ZN(MULT_mult_6_ab_6__25_) );
  XOR2_X2 MULT_mult_6_U4110 ( .A(MULT_mult_6_SUMB_4__27_), .B(
        MULT_mult_6_n1561), .Z(MULT_mult_6_SUMB_5__26_) );
  XOR2_X2 MULT_mult_6_U4109 ( .A(MULT_mult_6_CARRYB_4__26_), .B(
        MULT_mult_6_ab_5__26_), .Z(MULT_mult_6_n1561) );
  XOR2_X2 MULT_mult_6_U4108 ( .A(MULT_mult_6_SUMB_5__26_), .B(
        MULT_mult_6_n1560), .Z(MULT_mult_6_SUMB_6__25_) );
  XOR2_X2 MULT_mult_6_U4107 ( .A(MULT_mult_6_CARRYB_5__25_), .B(
        MULT_mult_6_ab_6__25_), .Z(MULT_mult_6_n1560) );
  NAND2_X2 MULT_mult_6_U4106 ( .A1(MULT_mult_6_CARRYB_7__8_), .A2(
        MULT_mult_6_ab_8__8_), .ZN(MULT_mult_6_n2004) );
  NAND2_X2 MULT_mult_6_U4105 ( .A1(MULT_mult_6_CARRYB_13__6_), .A2(
        MULT_mult_6_ab_14__6_), .ZN(MULT_mult_6_n1974) );
  XNOR2_X2 MULT_mult_6_U4104 ( .A(MULT_mult_6_CARRYB_13__5_), .B(
        MULT_mult_6_ab_14__5_), .ZN(MULT_mult_6_n1584) );
  NAND2_X4 MULT_mult_6_U4103 ( .A1(MULT_mult_6_n1558), .A2(MULT_mult_6_n1559), 
        .ZN(MULT_mult_6_SUMB_3__14_) );
  NAND3_X4 MULT_mult_6_U4102 ( .A1(MULT_mult_6_n2024), .A2(MULT_mult_6_n2023), 
        .A3(MULT_mult_6_n2022), .ZN(MULT_mult_6_CARRYB_13__7_) );
  NOR2_X1 MULT_mult_6_U4101 ( .A1(MULT_mult_6_net77914), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__7_) );
  NAND3_X2 MULT_mult_6_U4100 ( .A1(MULT_mult_6_net85000), .A2(
        MULT_mult_6_net84999), .A3(MULT_mult_6_net84998), .ZN(
        MULT_mult_6_CARRYB_14__7_) );
  INV_X4 MULT_mult_6_U4099 ( .A(MULT_mult_6_n2343), .ZN(
        MULT_mult_6_CARRYB_1__21_) );
  NAND3_X4 MULT_mult_6_U4098 ( .A1(MULT_mult_6_net80813), .A2(
        MULT_mult_6_net80812), .A3(MULT_mult_6_net80814), .ZN(
        MULT_mult_6_CARRYB_17__9_) );
  INV_X1 MULT_mult_6_U4097 ( .A(MULT_mult_6_ab_18__9_), .ZN(
        MULT_mult_6_net85017) );
  NAND2_X4 MULT_mult_6_U4096 ( .A1(MULT_mult_6_net83850), .A2(
        MULT_mult_6_net85017), .ZN(MULT_mult_6_n1555) );
  NOR2_X1 MULT_mult_6_U4095 ( .A1(MULT_mult_6_net85716), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__11_) );
  NOR2_X1 MULT_mult_6_U4094 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net77956), .ZN(MULT_mult_6_ab_4__9_) );
  XNOR2_X2 MULT_mult_6_U4093 ( .A(MULT_mult_6_CARRYB_13__7_), .B(
        MULT_mult_6_ab_14__7_), .ZN(MULT_mult_6_n1553) );
  NAND2_X4 MULT_mult_6_U4092 ( .A1(MULT_mult_6_n1554), .A2(MULT_mult_6_n1555), 
        .ZN(MULT_mult_6_net81782) );
  NAND2_X4 MULT_mult_6_U4091 ( .A1(MULT_mult_6_n1818), .A2(MULT_mult_6_n1819), 
        .ZN(MULT_mult_6_n2135) );
  NAND3_X4 MULT_mult_6_U4090 ( .A1(MULT_mult_6_n2232), .A2(MULT_mult_6_n2233), 
        .A3(MULT_mult_6_n2231), .ZN(MULT_mult_6_CARRYB_18__5_) );
  NAND2_X2 MULT_mult_6_U4089 ( .A1(MULT_mult_6_ab_5__20_), .A2(
        MULT_mult_6_SUMB_4__21_), .ZN(MULT_mult_6_n1884) );
  NAND3_X2 MULT_mult_6_U4088 ( .A1(MULT_mult_6_n2276), .A2(MULT_mult_6_n2277), 
        .A3(MULT_mult_6_n2278), .ZN(MULT_mult_6_CARRYB_4__21_) );
  NAND3_X2 MULT_mult_6_U4087 ( .A1(MULT_mult_6_n2266), .A2(MULT_mult_6_n2267), 
        .A3(MULT_mult_6_n2268), .ZN(MULT_mult_6_CARRYB_7__23_) );
  NAND2_X2 MULT_mult_6_U4086 ( .A1(MULT_mult_6_n1501), .A2(
        MULT_mult_6_ab_14__5_), .ZN(MULT_mult_6_n1702) );
  NAND3_X4 MULT_mult_6_U4085 ( .A1(MULT_mult_6_n1643), .A2(MULT_mult_6_n1644), 
        .A3(MULT_mult_6_n1642), .ZN(MULT_mult_6_CARRYB_2__11_) );
  XOR2_X2 MULT_mult_6_U4084 ( .A(MULT_mult_6_SUMB_9__22_), .B(
        MULT_mult_6_n2321), .Z(MULT_mult_6_SUMB_10__21_) );
  NAND2_X2 MULT_mult_6_U4083 ( .A1(MULT_mult_6_SUMB_3__9_), .A2(
        MULT_mult_6_CARRYB_3__8_), .ZN(MULT_mult_6_n1946) );
  NAND2_X4 MULT_mult_6_U4082 ( .A1(MULT_mult_6_SUMB_1__12_), .A2(
        MULT_mult_6_n289), .ZN(MULT_mult_6_n1643) );
  NOR2_X4 MULT_mult_6_U4081 ( .A1(MULT_mult_6_net70456), .A2(
        MULT_mult_6_net77970), .ZN(MULT_mult_6_ab_2__11_) );
  NAND2_X2 MULT_mult_6_U4080 ( .A1(MULT_mult_6_SUMB_4__9_), .A2(
        MULT_mult_6_ab_5__8_), .ZN(MULT_mult_6_n1965) );
  NOR2_X4 MULT_mult_6_U4079 ( .A1(MULT_mult_6_net70454), .A2(
        MULT_mult_6_net77970), .ZN(MULT_mult_6_ab_2__10_) );
  NAND2_X4 MULT_mult_6_U4078 ( .A1(MULT_mult_6_n1616), .A2(MULT_mult_6_n2010), 
        .ZN(MULT_mult_6_n1943) );
  NAND2_X2 MULT_mult_6_U4077 ( .A1(MULT_mult_6_ab_16__8_), .A2(
        MULT_mult_6_CARRYB_15__8_), .ZN(MULT_mult_6_n2299) );
  XNOR2_X2 MULT_mult_6_U4076 ( .A(MULT_mult_6_ab_10__20_), .B(
        MULT_mult_6_CARRYB_9__20_), .ZN(MULT_mult_6_n1550) );
  XNOR2_X2 MULT_mult_6_U4075 ( .A(MULT_mult_6_n1550), .B(
        MULT_mult_6_SUMB_9__21_), .ZN(MULT_mult_6_SUMB_10__20_) );
  NAND2_X2 MULT_mult_6_U4074 ( .A1(MULT_mult_6_CARRYB_2__24_), .A2(
        MULT_mult_6_SUMB_2__25_), .ZN(MULT_mult_6_n2170) );
  NAND2_X2 MULT_mult_6_U4073 ( .A1(MULT_mult_6_CARRYB_2__8_), .A2(
        MULT_mult_6_n1427), .ZN(MULT_mult_6_n1907) );
  NAND2_X2 MULT_mult_6_U4072 ( .A1(MULT_mult_6_ab_11__7_), .A2(
        MULT_mult_6_SUMB_10__8_), .ZN(MULT_mult_6_n1778) );
  NAND2_X2 MULT_mult_6_U4071 ( .A1(MULT_mult_6_n1501), .A2(
        MULT_mult_6_SUMB_13__6_), .ZN(MULT_mult_6_n1704) );
  NAND2_X2 MULT_mult_6_U4070 ( .A1(MULT_mult_6_n1301), .A2(
        MULT_mult_6_net90433), .ZN(MULT_mult_6_n2115) );
  INV_X4 MULT_mult_6_U4069 ( .A(MULT_mult_6_n1792), .ZN(MULT_mult_6_n1556) );
  NAND3_X2 MULT_mult_6_U4068 ( .A1(MULT_mult_6_net80796), .A2(
        MULT_mult_6_net80795), .A3(MULT_mult_6_net80794), .ZN(
        MULT_mult_6_CARRYB_5__22_) );
  NAND2_X2 MULT_mult_6_U4067 ( .A1(MULT_mult_6_ab_19__4_), .A2(
        MULT_mult_6_CARRYB_18__4_), .ZN(MULT_mult_6_n2234) );
  NAND3_X4 MULT_mult_6_U4066 ( .A1(MULT_mult_6_n1713), .A2(MULT_mult_6_n1712), 
        .A3(MULT_mult_6_n1711), .ZN(MULT_mult_6_CARRYB_2__18_) );
  NAND2_X2 MULT_mult_6_U4065 ( .A1(MULT_mult_6_n1546), .A2(MULT_mult_6_n1547), 
        .ZN(MULT_mult_6_n1549) );
  NAND2_X2 MULT_mult_6_U4064 ( .A1(MULT_mult_6_ab_3__18_), .A2(
        MULT_mult_6_CARRYB_2__18_), .ZN(MULT_mult_6_n1548) );
  INV_X1 MULT_mult_6_U4063 ( .A(MULT_mult_6_n1770), .ZN(MULT_mult_6_n1545) );
  INV_X2 MULT_mult_6_U4062 ( .A(MULT_mult_6_ab_5__13_), .ZN(MULT_mult_6_n1845)
         );
  NAND2_X2 MULT_mult_6_U4061 ( .A1(MULT_mult_6_CARRYB_6__12_), .A2(
        MULT_mult_6_ab_7__12_), .ZN(MULT_mult_6_n1544) );
  INV_X4 MULT_mult_6_U4060 ( .A(MULT_mult_6_n1845), .ZN(MULT_mult_6_n1540) );
  XNOR2_X2 MULT_mult_6_U4059 ( .A(MULT_mult_6_ab_4__25_), .B(
        MULT_mult_6_CARRYB_3__25_), .ZN(MULT_mult_6_n1539) );
  INV_X2 MULT_mult_6_U4058 ( .A(MULT_mult_6_n2345), .ZN(
        MULT_mult_6_CARRYB_1__22_) );
  NOR2_X4 MULT_mult_6_U4057 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70441), .ZN(MULT_mult_6_ab_27__3_) );
  INV_X4 MULT_mult_6_U4056 ( .A(MULT_mult_6_n1537), .ZN(MULT_mult_6_n1538) );
  NAND2_X4 MULT_mult_6_U4055 ( .A1(MULT_mult_6_n1538), .A2(
        MULT_mult_6_net81053), .ZN(MULT_mult_6_CARRYB_26__3_) );
  NAND2_X2 MULT_mult_6_U4054 ( .A1(MULT_mult_6_net81052), .A2(
        MULT_mult_6_n2116), .ZN(MULT_mult_6_n1537) );
  INV_X1 MULT_mult_6_U4053 ( .A(MULT_mult_6_ab_27__3_), .ZN(MULT_mult_6_n1534)
         );
  XOR2_X2 MULT_mult_6_U4052 ( .A(MULT_mult_6_SUMB_13__18_), .B(
        MULT_mult_6_n1532), .Z(MULT_mult_6_SUMB_14__17_) );
  XOR2_X2 MULT_mult_6_U4051 ( .A(MULT_mult_6_SUMB_8__23_), .B(
        MULT_mult_6_n1531), .Z(MULT_mult_6_SUMB_9__22_) );
  XOR2_X2 MULT_mult_6_U4050 ( .A(MULT_mult_6_CARRYB_8__22_), .B(
        MULT_mult_6_ab_9__22_), .Z(MULT_mult_6_n1531) );
  XNOR2_X2 MULT_mult_6_U4049 ( .A(MULT_mult_6_n1530), .B(
        MULT_mult_6_CARRYB_12__4_), .ZN(MULT_mult_6_n1635) );
  INV_X4 MULT_mult_6_U4048 ( .A(MULT_mult_6_n1528), .ZN(MULT_mult_6_n1529) );
  INV_X1 MULT_mult_6_U4047 ( .A(MULT_mult_6_ab_2__19_), .ZN(MULT_mult_6_n1525)
         );
  NAND2_X4 MULT_mult_6_U4046 ( .A1(MULT_mult_6_n1527), .A2(MULT_mult_6_n1526), 
        .ZN(MULT_mult_6_SUMB_2__19_) );
  NAND2_X4 MULT_mult_6_U4045 ( .A1(MULT_mult_6_n1524), .A2(MULT_mult_6_n1525), 
        .ZN(MULT_mult_6_n1527) );
  NAND3_X2 MULT_mult_6_U4044 ( .A1(MULT_mult_6_n2201), .A2(MULT_mult_6_n2202), 
        .A3(MULT_mult_6_n2203), .ZN(MULT_mult_6_CARRYB_5__17_) );
  NAND2_X1 MULT_mult_6_U4043 ( .A1(MULT_mult_6_ab_14__12_), .A2(
        MULT_mult_6_CARRYB_13__12_), .ZN(MULT_mult_6_n2122) );
  NAND2_X4 MULT_mult_6_U4042 ( .A1(MULT_mult_6_SUMB_12__12_), .A2(
        MULT_mult_6_net121285), .ZN(MULT_mult_6_net82159) );
  NAND2_X4 MULT_mult_6_U4041 ( .A1(MULT_mult_6_n1523), .A2(MULT_mult_6_n1522), 
        .ZN(MULT_mult_6_SUMB_11__10_) );
  NOR2_X1 MULT_mult_6_U4040 ( .A1(MULT_mult_6_net77898), .A2(
        MULT_mult_6_net77930), .ZN(MULT_mult_6_ab_7__5_) );
  NAND3_X2 MULT_mult_6_U4039 ( .A1(MULT_mult_6_n1519), .A2(MULT_mult_6_n1520), 
        .A3(MULT_mult_6_n1521), .ZN(MULT_mult_6_CARRYB_7__5_) );
  NAND2_X2 MULT_mult_6_U4038 ( .A1(MULT_mult_6_ab_7__5_), .A2(
        MULT_mult_6_CARRYB_6__5_), .ZN(MULT_mult_6_n1520) );
  INV_X4 MULT_mult_6_U4037 ( .A(MULT_mult_6_ab_1__9_), .ZN(MULT_mult_6_n1516)
         );
  NAND2_X2 MULT_mult_6_U4036 ( .A1(MULT_mult_6_n1518), .A2(MULT_mult_6_n1517), 
        .ZN(MULT_mult_6_n2331) );
  NOR2_X4 MULT_mult_6_U4035 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net86101), .ZN(MULT_mult_6_ab_1__9_) );
  NAND3_X4 MULT_mult_6_U4034 ( .A1(MULT_mult_6_n2076), .A2(MULT_mult_6_n2075), 
        .A3(MULT_mult_6_n2074), .ZN(MULT_mult_6_CARRYB_17__4_) );
  INV_X2 MULT_mult_6_U4033 ( .A(MULT_mult_6_ab_5__8_), .ZN(MULT_mult_6_n1513)
         );
  NAND2_X2 MULT_mult_6_U4032 ( .A1(MULT_mult_6_ab_2__20_), .A2(
        MULT_mult_6_CARRYB_1__20_), .ZN(MULT_mult_6_n2051) );
  XOR2_X2 MULT_mult_6_U4031 ( .A(MULT_mult_6_CARRYB_21__9_), .B(
        MULT_mult_6_n1929), .Z(MULT_mult_6_n1512) );
  XNOR2_X2 MULT_mult_6_U4030 ( .A(MULT_mult_6_SUMB_21__10_), .B(
        MULT_mult_6_n1512), .ZN(MULT_mult_6_SUMB_22__9_) );
  NAND2_X4 MULT_mult_6_U4029 ( .A1(MULT_mult_6_net84825), .A2(
        MULT_mult_6_net84826), .ZN(MULT_mult_6_net83866) );
  INV_X4 MULT_mult_6_U4028 ( .A(MULT_mult_6_n1943), .ZN(MULT_mult_6_n1509) );
  NAND2_X4 MULT_mult_6_U4027 ( .A1(MULT_mult_6_n1509), .A2(
        MULT_mult_6_net85469), .ZN(MULT_mult_6_n1511) );
  NAND2_X2 MULT_mult_6_U4026 ( .A1(MULT_mult_6_n1937), .A2(
        MULT_mult_6_net85465), .ZN(MULT_mult_6_n1507) );
  NAND2_X4 MULT_mult_6_U4025 ( .A1(MULT_mult_6_net85457), .A2(
        MULT_mult_6_n1505), .ZN(MULT_mult_6_SUMB_12__11_) );
  NAND3_X4 MULT_mult_6_U4024 ( .A1(MULT_mult_6_n2042), .A2(MULT_mult_6_n2041), 
        .A3(MULT_mult_6_n2040), .ZN(MULT_mult_6_CARRYB_18__4_) );
  XNOR2_X2 MULT_mult_6_U4023 ( .A(MULT_mult_6_CARRYB_14__4_), .B(
        MULT_mult_6_ab_15__4_), .ZN(MULT_mult_6_n1581) );
  NAND2_X2 MULT_mult_6_U4022 ( .A1(MULT_mult_6_ab_8__6_), .A2(
        MULT_mult_6_CARRYB_7__6_), .ZN(MULT_mult_6_n1825) );
  NAND2_X2 MULT_mult_6_U4021 ( .A1(MULT_mult_6_SUMB_12__5_), .A2(
        MULT_mult_6_ab_13__4_), .ZN(MULT_mult_6_n1640) );
  NAND2_X4 MULT_mult_6_U4020 ( .A1(MULT_mult_6_n1816), .A2(MULT_mult_6_n1817), 
        .ZN(MULT_mult_6_n1819) );
  XNOR2_X2 MULT_mult_6_U4019 ( .A(MULT_mult_6_ab_16__14_), .B(
        MULT_mult_6_CARRYB_15__14_), .ZN(MULT_mult_6_n1502) );
  XNOR2_X2 MULT_mult_6_U4018 ( .A(MULT_mult_6_n1502), .B(
        MULT_mult_6_SUMB_15__15_), .ZN(MULT_mult_6_SUMB_16__14_) );
  NAND3_X2 MULT_mult_6_U4017 ( .A1(MULT_mult_6_n1922), .A2(MULT_mult_6_n1921), 
        .A3(MULT_mult_6_n1920), .ZN(MULT_mult_6_n1501) );
  NAND2_X4 MULT_mult_6_U4016 ( .A1(MULT_mult_6_n287), .A2(MULT_mult_6_n1498), 
        .ZN(MULT_mult_6_net85603) );
  NAND2_X2 MULT_mult_6_U4015 ( .A1(MULT_mult_6_n397), .A2(
        MULT_mult_6_SUMB_1__19_), .ZN(MULT_mult_6_net85602) );
  NAND2_X4 MULT_mult_6_U4014 ( .A1(MULT_mult_6_n1496), .A2(MULT_mult_6_n1497), 
        .ZN(MULT_mult_6_SUMB_6__16_) );
  XNOR2_X2 MULT_mult_6_U4013 ( .A(MULT_mult_6_CARRYB_5__3_), .B(
        MULT_mult_6_ab_6__3_), .ZN(MULT_mult_6_n1495) );
  XNOR2_X2 MULT_mult_6_U4012 ( .A(MULT_mult_6_SUMB_5__4_), .B(
        MULT_mult_6_n1495), .ZN(MULT_mult_6_SUMB_6__3_) );
  NOR2_X4 MULT_mult_6_U4011 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net70451), .ZN(MULT_mult_6_ab_22__8_) );
  INV_X2 MULT_mult_6_U4010 ( .A(MULT_mult_6_CARRYB_3__18_), .ZN(
        MULT_mult_6_n1492) );
  INV_X4 MULT_mult_6_U4009 ( .A(MULT_mult_6_n1693), .ZN(MULT_mult_6_n1491) );
  NAND2_X4 MULT_mult_6_U4008 ( .A1(MULT_mult_6_n1493), .A2(MULT_mult_6_n1494), 
        .ZN(MULT_mult_6_SUMB_4__18_) );
  NAND2_X4 MULT_mult_6_U4007 ( .A1(MULT_mult_6_n1491), .A2(MULT_mult_6_n1492), 
        .ZN(MULT_mult_6_n1494) );
  NAND2_X2 MULT_mult_6_U4006 ( .A1(MULT_mult_6_CARRYB_3__18_), .A2(
        MULT_mult_6_n1693), .ZN(MULT_mult_6_n1493) );
  NAND3_X2 MULT_mult_6_U4005 ( .A1(MULT_mult_6_n2201), .A2(MULT_mult_6_n2202), 
        .A3(MULT_mult_6_n2203), .ZN(MULT_mult_6_n1490) );
  NAND2_X4 MULT_mult_6_U4004 ( .A1(MULT_mult_6_n2116), .A2(MULT_mult_6_n1696), 
        .ZN(MULT_mult_6_net81663) );
  NOR2_X2 MULT_mult_6_U4003 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__12_) );
  INV_X2 MULT_mult_6_U4002 ( .A(MULT_mult_6_ab_14__12_), .ZN(MULT_mult_6_n1487) );
  NAND2_X2 MULT_mult_6_U4001 ( .A1(MULT_mult_6_CARRYB_8__5_), .A2(
        MULT_mult_6_SUMB_8__6_), .ZN(MULT_mult_6_n1785) );
  XNOR2_X2 MULT_mult_6_U4000 ( .A(MULT_mult_6_n1485), .B(
        MULT_mult_6_SUMB_1__12_), .ZN(MULT_mult_6_SUMB_2__11_) );
  NAND3_X4 MULT_mult_6_U3999 ( .A1(MULT_mult_6_n1999), .A2(MULT_mult_6_n1998), 
        .A3(MULT_mult_6_n2000), .ZN(MULT_mult_6_CARRYB_13__6_) );
  XNOR2_X2 MULT_mult_6_U3998 ( .A(MULT_mult_6_net85734), .B(
        MULT_mult_6_net85036), .ZN(MULT_mult_6_SUMB_3__7_) );
  NOR2_X2 MULT_mult_6_U3997 ( .A1(MULT_mult_6_net77882), .A2(
        MULT_mult_6_net77970), .ZN(MULT_mult_6_ab_2__3_) );
  NAND3_X2 MULT_mult_6_U3996 ( .A1(MULT_mult_6_n1482), .A2(MULT_mult_6_n1483), 
        .A3(MULT_mult_6_n1484), .ZN(MULT_mult_6_CARRYB_5__1_) );
  NAND2_X1 MULT_mult_6_U3995 ( .A1(MULT_mult_6_SUMB_4__2_), .A2(
        MULT_mult_6_CARRYB_4__1_), .ZN(MULT_mult_6_n1484) );
  NAND2_X2 MULT_mult_6_U3994 ( .A1(MULT_mult_6_ab_5__1_), .A2(
        MULT_mult_6_CARRYB_4__1_), .ZN(MULT_mult_6_n1483) );
  NAND2_X1 MULT_mult_6_U3993 ( .A1(MULT_mult_6_ab_5__1_), .A2(
        MULT_mult_6_SUMB_4__2_), .ZN(MULT_mult_6_n1482) );
  XOR2_X2 MULT_mult_6_U3992 ( .A(MULT_mult_6_n1481), .B(
        MULT_mult_6_CARRYB_4__1_), .Z(MULT_mult_6_SUMB_5__1_) );
  NAND3_X2 MULT_mult_6_U3991 ( .A1(MULT_mult_6_n1478), .A2(MULT_mult_6_n1479), 
        .A3(MULT_mult_6_n1480), .ZN(MULT_mult_6_CARRYB_4__1_) );
  NAND2_X1 MULT_mult_6_U3990 ( .A1(MULT_mult_6_CARRYB_3__1_), .A2(
        MULT_mult_6_SUMB_3__2_), .ZN(MULT_mult_6_n1480) );
  NAND2_X2 MULT_mult_6_U3989 ( .A1(MULT_mult_6_ab_4__1_), .A2(
        MULT_mult_6_SUMB_3__2_), .ZN(MULT_mult_6_n1479) );
  NAND2_X1 MULT_mult_6_U3988 ( .A1(MULT_mult_6_ab_4__1_), .A2(
        MULT_mult_6_CARRYB_3__1_), .ZN(MULT_mult_6_n1478) );
  NAND3_X2 MULT_mult_6_U3987 ( .A1(MULT_mult_6_n1475), .A2(MULT_mult_6_n1476), 
        .A3(MULT_mult_6_n1477), .ZN(MULT_mult_6_CARRYB_2__3_) );
  NAND2_X1 MULT_mult_6_U3986 ( .A1(MULT_mult_6_ab_2__3_), .A2(
        MULT_mult_6_CARRYB_1__3_), .ZN(MULT_mult_6_n1477) );
  NAND2_X2 MULT_mult_6_U3985 ( .A1(MULT_mult_6_ab_2__3_), .A2(
        MULT_mult_6_SUMB_1__4_), .ZN(MULT_mult_6_n1476) );
  NAND2_X1 MULT_mult_6_U3984 ( .A1(MULT_mult_6_CARRYB_1__3_), .A2(
        MULT_mult_6_SUMB_1__4_), .ZN(MULT_mult_6_n1475) );
  XOR2_X2 MULT_mult_6_U3983 ( .A(MULT_mult_6_SUMB_1__4_), .B(MULT_mult_6_n1474), .Z(MULT_mult_6_SUMB_2__3_) );
  XOR2_X2 MULT_mult_6_U3982 ( .A(MULT_mult_6_CARRYB_1__3_), .B(
        MULT_mult_6_ab_2__3_), .Z(MULT_mult_6_n1474) );
  NAND2_X1 MULT_mult_6_U3981 ( .A1(MULT_mult_6_ab_5__23_), .A2(
        MULT_mult_6_SUMB_4__24_), .ZN(MULT_mult_6_n1959) );
  NOR2_X1 MULT_mult_6_U3980 ( .A1(MULT_mult_6_net70454), .A2(
        MULT_mult_6_net119855), .ZN(MULT_mult_6_ab_4__10_) );
  NAND3_X2 MULT_mult_6_U3979 ( .A1(MULT_mult_6_n2072), .A2(MULT_mult_6_n2073), 
        .A3(MULT_mult_6_n2071), .ZN(MULT_mult_6_CARRYB_16__5_) );
  NAND3_X2 MULT_mult_6_U3978 ( .A1(MULT_mult_6_n2289), .A2(MULT_mult_6_n2290), 
        .A3(MULT_mult_6_n2291), .ZN(MULT_mult_6_CARRYB_9__19_) );
  NAND2_X2 MULT_mult_6_U3977 ( .A1(MULT_mult_6_SUMB_9__2_), .A2(
        MULT_mult_6_CARRYB_9__1_), .ZN(MULT_mult_6_n1473) );
  NAND2_X2 MULT_mult_6_U3976 ( .A1(MULT_mult_6_SUMB_9__2_), .A2(
        MULT_mult_6_ab_10__1_), .ZN(MULT_mult_6_n1472) );
  NAND2_X2 MULT_mult_6_U3975 ( .A1(MULT_mult_6_ab_11__4_), .A2(
        MULT_mult_6_n2370), .ZN(MULT_mult_6_n1834) );
  XNOR2_X2 MULT_mult_6_U3974 ( .A(MULT_mult_6_ab_4__24_), .B(
        MULT_mult_6_CARRYB_3__24_), .ZN(MULT_mult_6_n1469) );
  XNOR2_X2 MULT_mult_6_U3973 ( .A(MULT_mult_6_n1469), .B(
        MULT_mult_6_SUMB_3__25_), .ZN(MULT_mult_6_SUMB_4__24_) );
  NAND2_X1 MULT_mult_6_U3972 ( .A1(MULT_mult_6_CARRYB_11__17_), .A2(
        MULT_mult_6_SUMB_11__18_), .ZN(MULT_mult_6_n1467) );
  NAND2_X1 MULT_mult_6_U3971 ( .A1(MULT_mult_6_CARRYB_11__17_), .A2(
        MULT_mult_6_ab_12__17_), .ZN(MULT_mult_6_n1466) );
  NAND3_X2 MULT_mult_6_U3970 ( .A1(MULT_mult_6_n1463), .A2(MULT_mult_6_n1464), 
        .A3(MULT_mult_6_n1465), .ZN(MULT_mult_6_CARRYB_11__18_) );
  NAND2_X1 MULT_mult_6_U3969 ( .A1(MULT_mult_6_CARRYB_10__18_), .A2(
        MULT_mult_6_SUMB_10__19_), .ZN(MULT_mult_6_n1465) );
  NAND2_X1 MULT_mult_6_U3968 ( .A1(MULT_mult_6_ab_11__18_), .A2(
        MULT_mult_6_SUMB_10__19_), .ZN(MULT_mult_6_n1464) );
  NAND2_X1 MULT_mult_6_U3967 ( .A1(MULT_mult_6_ab_11__18_), .A2(
        MULT_mult_6_CARRYB_10__18_), .ZN(MULT_mult_6_n1463) );
  XOR2_X2 MULT_mult_6_U3966 ( .A(MULT_mult_6_n1462), .B(
        MULT_mult_6_SUMB_10__19_), .Z(MULT_mult_6_SUMB_11__18_) );
  XOR2_X2 MULT_mult_6_U3965 ( .A(MULT_mult_6_ab_11__18_), .B(
        MULT_mult_6_CARRYB_10__18_), .Z(MULT_mult_6_n1462) );
  NAND2_X2 MULT_mult_6_U3964 ( .A1(MULT_mult_6_n173), .A2(
        MULT_mult_6_ab_11__7_), .ZN(MULT_mult_6_n1777) );
  XNOR2_X2 MULT_mult_6_U3963 ( .A(MULT_mult_6_ab_4__9_), .B(
        MULT_mult_6_CARRYB_3__9_), .ZN(MULT_mult_6_n1461) );
  XNOR2_X2 MULT_mult_6_U3962 ( .A(MULT_mult_6_n1461), .B(MULT_mult_6_n1259), 
        .ZN(MULT_mult_6_SUMB_4__9_) );
  NAND3_X4 MULT_mult_6_U3961 ( .A1(MULT_mult_6_n1777), .A2(MULT_mult_6_n1779), 
        .A3(MULT_mult_6_n1778), .ZN(MULT_mult_6_CARRYB_11__7_) );
  NAND2_X4 MULT_mult_6_U3960 ( .A1(MULT_mult_6_SUMB_1__12_), .A2(
        MULT_mult_6_CARRYB_1__11_), .ZN(MULT_mult_6_n1644) );
  INV_X4 MULT_mult_6_U3959 ( .A(MULT_mult_6_CARRYB_23__5_), .ZN(
        MULT_mult_6_n2155) );
  NAND2_X2 MULT_mult_6_U3958 ( .A1(MULT_mult_6_SUMB_23__6_), .A2(
        MULT_mult_6_n1251), .ZN(MULT_mult_6_net79968) );
  NOR2_X2 MULT_mult_6_U3957 ( .A1(MULT_mult_6_net70491), .A2(
        MULT_mult_6_net70478), .ZN(MULT_mult_6_ab_2__22_) );
  XNOR2_X2 MULT_mult_6_U3956 ( .A(MULT_mult_6_n1457), .B(
        MULT_mult_6_SUMB_1__23_), .ZN(MULT_mult_6_SUMB_2__22_) );
  NAND2_X2 MULT_mult_6_U3955 ( .A1(MULT_mult_6_CARRYB_17__9_), .A2(
        MULT_mult_6_ab_18__9_), .ZN(MULT_mult_6_n1554) );
  NAND3_X2 MULT_mult_6_U3954 ( .A1(MULT_mult_6_net81034), .A2(
        MULT_mult_6_net81035), .A3(MULT_mult_6_net81033), .ZN(
        MULT_mult_6_CARRYB_20__9_) );
  NAND2_X2 MULT_mult_6_U3953 ( .A1(MULT_mult_6_ab_4__9_), .A2(
        MULT_mult_6_SUMB_3__10_), .ZN(MULT_mult_6_n1962) );
  INV_X1 MULT_mult_6_U3952 ( .A(MULT_mult_6_ab_16__5_), .ZN(MULT_mult_6_n1453)
         );
  NAND2_X2 MULT_mult_6_U3951 ( .A1(MULT_mult_6_n1514), .A2(MULT_mult_6_n1513), 
        .ZN(MULT_mult_6_n1515) );
  XNOR2_X2 MULT_mult_6_U3950 ( .A(MULT_mult_6_n1452), .B(MULT_mult_6_n1427), 
        .ZN(MULT_mult_6_SUMB_3__8_) );
  NAND2_X4 MULT_mult_6_U3949 ( .A1(MULT_mult_6_n1450), .A2(MULT_mult_6_n1451), 
        .ZN(MULT_mult_6_SUMB_16__8_) );
  NAND2_X2 MULT_mult_6_U3948 ( .A1(MULT_mult_6_n1279), .A2(MULT_mult_6_n1449), 
        .ZN(MULT_mult_6_n1450) );
  NAND2_X2 MULT_mult_6_U3947 ( .A1(MULT_mult_6_n194), .A2(MULT_mult_6_n2060), 
        .ZN(MULT_mult_6_n1459) );
  XNOR2_X2 MULT_mult_6_U3946 ( .A(MULT_mult_6_n1448), .B(MULT_mult_6_n1206), 
        .ZN(MULT_mult_6_SUMB_9__5_) );
  XOR2_X2 MULT_mult_6_U3945 ( .A(MULT_mult_6_SUMB_4__2_), .B(
        MULT_mult_6_ab_5__1_), .Z(MULT_mult_6_n1481) );
  NAND2_X2 MULT_mult_6_U3944 ( .A1(MULT_mult_6_ab_18__0_), .A2(
        MULT_mult_6_CARRYB_17__0_), .ZN(MULT_mult_6_n1809) );
  NAND2_X2 MULT_mult_6_U3943 ( .A1(MULT_mult_6_CARRYB_17__0_), .A2(
        MULT_mult_6_SUMB_17__1_), .ZN(MULT_mult_6_n1811) );
  NAND2_X4 MULT_mult_6_U3942 ( .A1(MULT_mult_6_ab_21__0_), .A2(
        MULT_mult_6_n1237), .ZN(MULT_mult_6_n1807) );
  XNOR2_X2 MULT_mult_6_U3941 ( .A(MULT_mult_6_CARRYB_14__14_), .B(
        MULT_mult_6_ab_15__14_), .ZN(MULT_mult_6_net86054) );
  NAND2_X4 MULT_mult_6_U3940 ( .A1(MULT_mult_6_n1447), .A2(MULT_mult_6_n1446), 
        .ZN(MULT_mult_6_SUMB_13__7_) );
  NAND2_X4 MULT_mult_6_U3939 ( .A1(MULT_mult_6_n1444), .A2(MULT_mult_6_n1445), 
        .ZN(MULT_mult_6_n1447) );
  NAND2_X4 MULT_mult_6_U3938 ( .A1(MULT_mult_6_n1556), .A2(MULT_mult_6_n1557), 
        .ZN(MULT_mult_6_n1559) );
  INV_X1 MULT_mult_6_U3937 ( .A(MULT_mult_6_ab_7__7_), .ZN(MULT_mult_6_n1499)
         );
  NAND2_X4 MULT_mult_6_U3935 ( .A1(MULT_mult_6_n1763), .A2(MULT_mult_6_n1762), 
        .ZN(MULT_mult_6_n2001) );
  NOR2_X1 MULT_mult_6_U3934 ( .A1(MULT_mult_6_net77898), .A2(
        MULT_mult_6_net77938), .ZN(MULT_mult_6_ab_6__5_) );
  NAND3_X2 MULT_mult_6_U3933 ( .A1(MULT_mult_6_n1440), .A2(MULT_mult_6_n1441), 
        .A3(MULT_mult_6_n1442), .ZN(MULT_mult_6_CARRYB_6__5_) );
  NAND2_X1 MULT_mult_6_U3932 ( .A1(MULT_mult_6_ab_6__5_), .A2(
        MULT_mult_6_CARRYB_5__5_), .ZN(MULT_mult_6_n1442) );
  NAND2_X1 MULT_mult_6_U3931 ( .A1(MULT_mult_6_SUMB_5__6_), .A2(
        MULT_mult_6_ab_6__5_), .ZN(MULT_mult_6_n1441) );
  NAND2_X1 MULT_mult_6_U3930 ( .A1(MULT_mult_6_SUMB_5__6_), .A2(
        MULT_mult_6_CARRYB_5__5_), .ZN(MULT_mult_6_n1440) );
  NAND3_X2 MULT_mult_6_U3929 ( .A1(MULT_mult_6_n1839), .A2(MULT_mult_6_n1840), 
        .A3(MULT_mult_6_n1841), .ZN(MULT_mult_6_CARRYB_10__15_) );
  NAND2_X4 MULT_mult_6_U3928 ( .A1(MULT_mult_6_n1858), .A2(MULT_mult_6_n1857), 
        .ZN(MULT_mult_6_n1860) );
  NAND2_X2 MULT_mult_6_U3927 ( .A1(MULT_mult_6_ab_5__7_), .A2(
        MULT_mult_6_SUMB_4__8_), .ZN(MULT_mult_6_n1947) );
  NAND2_X2 MULT_mult_6_U3926 ( .A1(MULT_mult_6_CARRYB_4__7_), .A2(
        MULT_mult_6_SUMB_4__8_), .ZN(MULT_mult_6_n1948) );
  NAND2_X4 MULT_mult_6_U3925 ( .A1(MULT_mult_6_n1460), .A2(MULT_mult_6_n1459), 
        .ZN(MULT_mult_6_SUMB_11__5_) );
  NOR2_X4 MULT_mult_6_U3924 ( .A1(MULT_mult_6_net84698), .A2(
        MULT_mult_6_net70491), .ZN(MULT_mult_6_ab_2__14_) );
  NOR2_X2 MULT_mult_6_U3923 ( .A1(MULT_mult_6_net77908), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__6_) );
  NAND3_X4 MULT_mult_6_U3922 ( .A1(MULT_mult_6_n1974), .A2(MULT_mult_6_n1976), 
        .A3(MULT_mult_6_n1975), .ZN(MULT_mult_6_CARRYB_14__6_) );
  NAND3_X2 MULT_mult_6_U3921 ( .A1(MULT_mult_6_net86170), .A2(
        MULT_mult_6_net86171), .A3(MULT_mult_6_net86172), .ZN(
        MULT_mult_6_CARRYB_2__14_) );
  NAND3_X2 MULT_mult_6_U3920 ( .A1(MULT_mult_6_n1437), .A2(MULT_mult_6_n1436), 
        .A3(MULT_mult_6_n1438), .ZN(MULT_mult_6_CARRYB_15__6_) );
  NAND2_X2 MULT_mult_6_U3919 ( .A1(MULT_mult_6_CARRYB_14__6_), .A2(
        MULT_mult_6_SUMB_14__7_), .ZN(MULT_mult_6_n1436) );
  NAND3_X2 MULT_mult_6_U3918 ( .A1(MULT_mult_6_n1964), .A2(MULT_mult_6_n1966), 
        .A3(MULT_mult_6_n1965), .ZN(MULT_mult_6_CARRYB_5__8_) );
  XNOR2_X2 MULT_mult_6_U3917 ( .A(MULT_mult_6_SUMB_4__22_), .B(
        MULT_mult_6_n1435), .ZN(MULT_mult_6_SUMB_5__21_) );
  NAND3_X4 MULT_mult_6_U3916 ( .A1(MULT_mult_6_n2237), .A2(MULT_mult_6_n2239), 
        .A3(MULT_mult_6_n2238), .ZN(MULT_mult_6_CARRYB_4__20_) );
  NAND2_X4 MULT_mult_6_U3915 ( .A1(MULT_mult_6_ab_4__19_), .A2(
        MULT_mult_6_SUMB_3__20_), .ZN(MULT_mult_6_n2137) );
  INV_X4 MULT_mult_6_U3914 ( .A(MULT_mult_6_n1765), .ZN(MULT_mult_6_n1431) );
  NAND2_X4 MULT_mult_6_U3913 ( .A1(MULT_mult_6_n1433), .A2(MULT_mult_6_n1434), 
        .ZN(MULT_mult_6_SUMB_3__20_) );
  NAND3_X2 MULT_mult_6_U3912 ( .A1(MULT_mult_6_net86158), .A2(
        MULT_mult_6_net86159), .A3(MULT_mult_6_n1019), .ZN(
        MULT_mult_6_CARRYB_12__12_) );
  NAND3_X4 MULT_mult_6_U3911 ( .A1(MULT_mult_6_net81513), .A2(
        MULT_mult_6_net81514), .A3(MULT_mult_6_net81515), .ZN(
        MULT_mult_6_CARRYB_3__13_) );
  XNOR2_X2 MULT_mult_6_U3910 ( .A(MULT_mult_6_n1246), .B(MULT_mult_6_ab_3__9_), 
        .ZN(MULT_mult_6_n1428) );
  XNOR2_X2 MULT_mult_6_U3909 ( .A(MULT_mult_6_n1428), .B(
        MULT_mult_6_SUMB_2__10_), .ZN(MULT_mult_6_SUMB_3__9_) );
  INV_X2 MULT_mult_6_U3908 ( .A(MULT_mult_6_SUMB_2__9_), .ZN(MULT_mult_6_n1426) );
  NAND2_X2 MULT_mult_6_U3907 ( .A1(MULT_mult_6_CARRYB_15__5_), .A2(
        MULT_mult_6_SUMB_15__6_), .ZN(MULT_mult_6_n2073) );
  NAND3_X2 MULT_mult_6_U3906 ( .A1(MULT_mult_6_n2150), .A2(MULT_mult_6_n2151), 
        .A3(MULT_mult_6_n2152), .ZN(MULT_mult_6_CARRYB_14__4_) );
  XOR2_X1 MULT_mult_6_U3905 ( .A(MULT_mult_6_CARRYB_17__0_), .B(
        MULT_mult_6_ab_18__0_), .Z(MULT_mult_6_n1808) );
  NOR2_X4 MULT_mult_6_U3904 ( .A1(MULT_mult_6_net123000), .A2(
        MULT_mult_6_net70491), .ZN(MULT_mult_6_ab_2__17_) );
  NAND2_X2 MULT_mult_6_U3903 ( .A1(MULT_mult_6_ab_8__9_), .A2(
        MULT_mult_6_CARRYB_7__9_), .ZN(MULT_mult_6_n2083) );
  NOR2_X2 MULT_mult_6_U3902 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net77970), .ZN(MULT_mult_6_ab_2__9_) );
  XNOR2_X2 MULT_mult_6_U3901 ( .A(MULT_mult_6_ab_17__13_), .B(
        MULT_mult_6_CARRYB_16__13_), .ZN(MULT_mult_6_n1423) );
  XNOR2_X2 MULT_mult_6_U3900 ( .A(MULT_mult_6_SUMB_16__14_), .B(
        MULT_mult_6_n1423), .ZN(MULT_mult_6_SUMB_17__13_) );
  NOR2_X4 MULT_mult_6_U3899 ( .A1(MULT_mult_6_net70472), .A2(
        MULT_mult_6_net82149), .ZN(MULT_mult_6_net81354) );
  INV_X8 MULT_mult_6_U3898 ( .A(MULT_mult_6_net81080), .ZN(
        MULT_mult_6_net80727) );
  NOR2_X4 MULT_mult_6_U3897 ( .A1(MULT_mult_6_net86565), .A2(
        MULT_mult_6_net77948), .ZN(MULT_mult_6_ab_5__19_) );
  NOR2_X4 MULT_mult_6_U3896 ( .A1(MULT_mult_6_net70472), .A2(
        MULT_mult_6_net80409), .ZN(MULT_mult_6_ab_1__19_) );
  NAND3_X4 MULT_mult_6_U3895 ( .A1(MULT_mult_6_n2085), .A2(MULT_mult_6_n2084), 
        .A3(MULT_mult_6_n2083), .ZN(MULT_mult_6_CARRYB_8__9_) );
  INV_X4 MULT_mult_6_U3894 ( .A(MULT_mult_6_SUMB_4__19_), .ZN(
        MULT_mult_6_n1576) );
  NAND2_X2 MULT_mult_6_U3893 ( .A1(MULT_mult_6_n708), .A2(
        MULT_mult_6_SUMB_4__19_), .ZN(MULT_mult_6_n1577) );
  INV_X4 MULT_mult_6_U3892 ( .A(MULT_mult_6_n2135), .ZN(MULT_mult_6_n1419) );
  NAND2_X4 MULT_mult_6_U3891 ( .A1(MULT_mult_6_n1421), .A2(MULT_mult_6_n1422), 
        .ZN(MULT_mult_6_SUMB_4__19_) );
  NAND2_X2 MULT_mult_6_U3890 ( .A1(MULT_mult_6_n2135), .A2(MULT_mult_6_n1420), 
        .ZN(MULT_mult_6_n1421) );
  NAND3_X2 MULT_mult_6_U3889 ( .A1(MULT_mult_6_net86412), .A2(
        MULT_mult_6_net86413), .A3(MULT_mult_6_net86414), .ZN(
        MULT_mult_6_CARRYB_23__7_) );
  NAND2_X4 MULT_mult_6_U3888 ( .A1(MULT_mult_6_CARRYB_24__4_), .A2(
        MULT_mult_6_ab_25__4_), .ZN(MULT_mult_6_n1854) );
  XNOR2_X2 MULT_mult_6_U3887 ( .A(MULT_mult_6_net86427), .B(
        MULT_mult_6_net88656), .ZN(MULT_mult_6_SUMB_26__1_) );
  INV_X8 MULT_mult_6_U3886 ( .A(MULT_mult_6_CARRYB_24__4_), .ZN(
        MULT_mult_6_net82551) );
  NAND2_X4 MULT_mult_6_U3885 ( .A1(MULT_mult_6_n1190), .A2(
        MULT_mult_6_ab_20__6_), .ZN(MULT_mult_6_n2212) );
  INV_X4 MULT_mult_6_U3884 ( .A(MULT_mult_6_n1732), .ZN(MULT_mult_6_n1444) );
  NOR2_X2 MULT_mult_6_U3883 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net77940), .ZN(MULT_mult_6_ab_6__12_) );
  INV_X1 MULT_mult_6_U3882 ( .A(MULT_mult_6_ab_6__12_), .ZN(
        MULT_mult_6_net86440) );
  NAND2_X2 MULT_mult_6_U3881 ( .A1(MULT_mult_6_ab_6__12_), .A2(
        MULT_mult_6_CARRYB_5__12_), .ZN(MULT_mult_6_n1983) );
  NAND3_X4 MULT_mult_6_U3880 ( .A1(MULT_mult_6_n2106), .A2(MULT_mult_6_n2108), 
        .A3(MULT_mult_6_n2107), .ZN(MULT_mult_6_CARRYB_17__3_) );
  NOR2_X2 MULT_mult_6_U3879 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70459), .ZN(MULT_mult_6_ab_18__3_) );
  NAND3_X4 MULT_mult_6_U3878 ( .A1(MULT_mult_6_net80247), .A2(
        MULT_mult_6_net80248), .A3(MULT_mult_6_net80246), .ZN(
        MULT_mult_6_CARRYB_10__13_) );
  NAND3_X4 MULT_mult_6_U3877 ( .A1(MULT_mult_6_n2293), .A2(MULT_mult_6_n2292), 
        .A3(MULT_mult_6_n2294), .ZN(MULT_mult_6_CARRYB_9__14_) );
  NAND2_X1 MULT_mult_6_U3876 ( .A1(MULT_mult_6_CARRYB_8__21_), .A2(
        MULT_mult_6_SUMB_8__22_), .ZN(MULT_mult_6_n1688) );
  NAND2_X4 MULT_mult_6_U3875 ( .A1(MULT_mult_6_ab_0__5_), .A2(
        MULT_mult_6_ab_1__4_), .ZN(MULT_mult_6_n2327) );
  XNOR2_X2 MULT_mult_6_U3874 ( .A(MULT_mult_6_n1413), .B(MULT_mult_6_n2142), 
        .ZN(MULT_mult_6_SUMB_20__11_) );
  NAND2_X4 MULT_mult_6_U3873 ( .A1(MULT_mult_6_n1488), .A2(MULT_mult_6_n1489), 
        .ZN(MULT_mult_6_net83535) );
  NAND2_X1 MULT_mult_6_U3872 ( .A1(MULT_mult_6_ab_3__19_), .A2(
        MULT_mult_6_CARRYB_2__19_), .ZN(MULT_mult_6_n2054) );
  NOR2_X2 MULT_mult_6_U3871 ( .A1(MULT_mult_6_net70436), .A2(
        MULT_mult_6_net83263), .ZN(MULT_mult_6_ab_1__0_) );
  NOR2_X2 MULT_mult_6_U3870 ( .A1(MULT_mult_6_net77900), .A2(MULT_mult_6_n242), 
        .ZN(MULT_mult_6_ab_1__5_) );
  NAND2_X4 MULT_mult_6_U3869 ( .A1(MULT_mult_6_net86630), .A2(
        MULT_mult_6_n1412), .ZN(MULT_mult_6_SUMB_14__13_) );
  NAND3_X2 MULT_mult_6_U3868 ( .A1(MULT_mult_6_n2209), .A2(MULT_mult_6_n2210), 
        .A3(MULT_mult_6_n2208), .ZN(MULT_mult_6_CARRYB_7__15_) );
  NAND3_X4 MULT_mult_6_U3867 ( .A1(MULT_mult_6_n2160), .A2(
        MULT_mult_6_net80852), .A3(MULT_mult_6_net80850), .ZN(
        MULT_mult_6_CARRYB_20__1_) );
  NAND2_X2 MULT_mult_6_U3866 ( .A1(MULT_mult_6_ab_20__6_), .A2(
        MULT_mult_6_CARRYB_19__6_), .ZN(MULT_mult_6_n2213) );
  NAND3_X4 MULT_mult_6_U3865 ( .A1(MULT_mult_6_n2211), .A2(MULT_mult_6_n2212), 
        .A3(MULT_mult_6_n2213), .ZN(MULT_mult_6_CARRYB_20__6_) );
  NOR2_X2 MULT_mult_6_U3864 ( .A1(MULT_mult_6_net77860), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__0_) );
  NOR2_X1 MULT_mult_6_U3863 ( .A1(MULT_mult_6_net77866), .A2(
        MULT_mult_6_net77938), .ZN(MULT_mult_6_ab_6__1_) );
  NAND2_X2 MULT_mult_6_U3862 ( .A1(MULT_mult_6_CARRYB_14__0_), .A2(
        MULT_mult_6_ab_15__0_), .ZN(MULT_mult_6_n1410) );
  XOR2_X2 MULT_mult_6_U3861 ( .A(MULT_mult_6_n846), .B(MULT_mult_6_n1408), .Z(
        multOut[16]) );
  XOR2_X1 MULT_mult_6_U3860 ( .A(MULT_mult_6_SUMB_14__1_), .B(
        MULT_mult_6_ab_15__0_), .Z(MULT_mult_6_n1408) );
  NAND3_X2 MULT_mult_6_U3859 ( .A1(MULT_mult_6_net86654), .A2(
        MULT_mult_6_n1407), .A3(MULT_mult_6_net86656), .ZN(
        MULT_mult_6_CARRYB_17__0_) );
  NAND2_X2 MULT_mult_6_U3858 ( .A1(MULT_mult_6_ab_17__0_), .A2(
        MULT_mult_6_CARRYB_16__0_), .ZN(MULT_mult_6_n1407) );
  XOR2_X1 MULT_mult_6_U3857 ( .A(MULT_mult_6_net86653), .B(
        MULT_mult_6_CARRYB_16__0_), .Z(multOut[14]) );
  NAND2_X2 MULT_mult_6_U3856 ( .A1(MULT_mult_6_ab_16__0_), .A2(
        MULT_mult_6_CARRYB_15__0_), .ZN(MULT_mult_6_n1406) );
  XOR2_X1 MULT_mult_6_U3855 ( .A(MULT_mult_6_CARRYB_15__0_), .B(
        MULT_mult_6_ab_16__0_), .Z(MULT_mult_6_net86649) );
  NAND3_X2 MULT_mult_6_U3854 ( .A1(MULT_mult_6_n1403), .A2(MULT_mult_6_n1404), 
        .A3(MULT_mult_6_n1405), .ZN(MULT_mult_6_CARRYB_6__1_) );
  NAND2_X2 MULT_mult_6_U3853 ( .A1(MULT_mult_6_ab_6__1_), .A2(
        MULT_mult_6_CARRYB_5__1_), .ZN(MULT_mult_6_n1405) );
  NAND2_X2 MULT_mult_6_U3852 ( .A1(MULT_mult_6_ab_6__1_), .A2(
        MULT_mult_6_SUMB_5__2_), .ZN(MULT_mult_6_n1404) );
  NAND2_X2 MULT_mult_6_U3851 ( .A1(MULT_mult_6_CARRYB_5__1_), .A2(
        MULT_mult_6_SUMB_5__2_), .ZN(MULT_mult_6_n1403) );
  XOR2_X2 MULT_mult_6_U3850 ( .A(MULT_mult_6_SUMB_5__2_), .B(MULT_mult_6_n1402), .Z(MULT_mult_6_SUMB_6__1_) );
  XOR2_X2 MULT_mult_6_U3849 ( .A(MULT_mult_6_CARRYB_5__1_), .B(
        MULT_mult_6_ab_6__1_), .Z(MULT_mult_6_n1402) );
  NAND2_X2 MULT_mult_6_U3848 ( .A1(MULT_mult_6_ab_12__6_), .A2(
        MULT_mult_6_SUMB_11__7_), .ZN(MULT_mult_6_n1918) );
  NAND2_X4 MULT_mult_6_U3847 ( .A1(MULT_mult_6_net86704), .A2(
        MULT_mult_6_n1401), .ZN(MULT_mult_6_SUMB_21__7_) );
  INV_X4 MULT_mult_6_U3846 ( .A(MULT_mult_6_CARRYB_24__5_), .ZN(
        MULT_mult_6_net86698) );
  NAND2_X4 MULT_mult_6_U3845 ( .A1(MULT_mult_6_net86699), .A2(
        MULT_mult_6_n1400), .ZN(MULT_mult_6_net81815) );
  NAND2_X4 MULT_mult_6_U3844 ( .A1(MULT_mult_6_net86697), .A2(
        MULT_mult_6_net86698), .ZN(MULT_mult_6_n1400) );
  NAND2_X2 MULT_mult_6_U3843 ( .A1(MULT_mult_6_n6), .A2(
        MULT_mult_6_SUMB_16__8_), .ZN(MULT_mult_6_net81267) );
  NAND2_X2 MULT_mult_6_U3842 ( .A1(MULT_mult_6_ab_3__21_), .A2(
        MULT_mult_6_SUMB_2__22_), .ZN(MULT_mult_6_n1934) );
  XNOR2_X2 MULT_mult_6_U3841 ( .A(MULT_mult_6_n128), .B(MULT_mult_6_n1399), 
        .ZN(MULT_mult_6_SUMB_3__10_) );
  NAND3_X2 MULT_mult_6_U3840 ( .A1(MULT_mult_6_n2077), .A2(MULT_mult_6_n2078), 
        .A3(MULT_mult_6_n2079), .ZN(MULT_mult_6_n1425) );
  NAND2_X2 MULT_mult_6_U3839 ( .A1(MULT_mult_6_n572), .A2(MULT_mult_6_ab_5__9_), .ZN(MULT_mult_6_n1397) );
  NAND3_X4 MULT_mult_6_U3838 ( .A1(MULT_mult_6_n1395), .A2(MULT_mult_6_n1394), 
        .A3(MULT_mult_6_n1393), .ZN(MULT_mult_6_CARRYB_4__10_) );
  NAND2_X1 MULT_mult_6_U3837 ( .A1(MULT_mult_6_ab_19__8_), .A2(
        MULT_mult_6_CARRYB_18__8_), .ZN(MULT_mult_6_n1392) );
  NAND3_X4 MULT_mult_6_U3836 ( .A1(MULT_mult_6_n1982), .A2(MULT_mult_6_n1981), 
        .A3(MULT_mult_6_n1980), .ZN(MULT_mult_6_CARRYB_5__13_) );
  NAND3_X4 MULT_mult_6_U3835 ( .A1(MULT_mult_6_n2127), .A2(MULT_mult_6_n2126), 
        .A3(MULT_mult_6_n2128), .ZN(MULT_mult_6_CARRYB_8__11_) );
  NAND3_X4 MULT_mult_6_U3834 ( .A1(MULT_mult_6_n2027), .A2(
        MULT_mult_6_net81535), .A3(MULT_mult_6_net81533), .ZN(
        MULT_mult_6_CARRYB_26__0_) );
  NAND2_X4 MULT_mult_6_U3833 ( .A1(MULT_mult_6_CARRYB_26__0_), .A2(
        MULT_mult_6_ab_27__0_), .ZN(MULT_mult_6_net80767) );
  NAND3_X4 MULT_mult_6_U3832 ( .A1(MULT_mult_6_net80805), .A2(
        MULT_mult_6_net80806), .A3(MULT_mult_6_n2164), .ZN(
        MULT_mult_6_CARRYB_10__16_) );
  XNOR2_X2 MULT_mult_6_U3831 ( .A(MULT_mult_6_CARRYB_2__8_), .B(
        MULT_mult_6_ab_3__8_), .ZN(MULT_mult_6_n1452) );
  NAND2_X2 MULT_mult_6_U3830 ( .A1(MULT_mult_6_ab_3__8_), .A2(
        MULT_mult_6_CARRYB_2__8_), .ZN(MULT_mult_6_n1905) );
  NAND2_X4 MULT_mult_6_U3829 ( .A1(MULT_mult_6_n1859), .A2(MULT_mult_6_n1860), 
        .ZN(MULT_mult_6_n2109) );
  NOR2_X4 MULT_mult_6_U3828 ( .A1(MULT_mult_6_net124723), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__16_) );
  NOR2_X4 MULT_mult_6_U3827 ( .A1(MULT_mult_6_net124723), .A2(
        MULT_mult_6_net77926), .ZN(MULT_mult_6_ab_8__16_) );
  NOR2_X1 MULT_mult_6_U3826 ( .A1(MULT_mult_6_net124723), .A2(
        MULT_mult_6_net77932), .ZN(MULT_mult_6_ab_7__16_) );
  NAND2_X2 MULT_mult_6_U3825 ( .A1(MULT_mult_6_n1453), .A2(MULT_mult_6_n1454), 
        .ZN(MULT_mult_6_n1455) );
  NAND2_X4 MULT_mult_6_U3824 ( .A1(MULT_mult_6_n1515), .A2(MULT_mult_6_n1964), 
        .ZN(MULT_mult_6_n1880) );
  NAND2_X4 MULT_mult_6_U3823 ( .A1(MULT_mult_6_net83121), .A2(
        MULT_mult_6_n1759), .ZN(MULT_mult_6_net80264) );
  NAND2_X4 MULT_mult_6_U3822 ( .A1(MULT_mult_6_n2046), .A2(MULT_mult_6_n2047), 
        .ZN(MULT_mult_6_n2112) );
  NOR2_X2 MULT_mult_6_U3821 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net70463), .ZN(MULT_mult_6_ab_16__12_) );
  INV_X4 MULT_mult_6_U3820 ( .A(MULT_mult_6_n1608), .ZN(MULT_mult_6_n1386) );
  NAND2_X2 MULT_mult_6_U3819 ( .A1(MULT_mult_6_ab_17__11_), .A2(
        MULT_mult_6_SUMB_16__12_), .ZN(MULT_mult_6_net87012) );
  NAND2_X1 MULT_mult_6_U3818 ( .A1(MULT_mult_6_CARRYB_16__11_), .A2(
        MULT_mult_6_ab_17__11_), .ZN(MULT_mult_6_net87010) );
  NAND2_X2 MULT_mult_6_U3817 ( .A1(MULT_mult_6_net87003), .A2(
        MULT_mult_6_net87004), .ZN(MULT_mult_6_n1385) );
  NAND3_X2 MULT_mult_6_U3816 ( .A1(MULT_mult_6_net84926), .A2(
        MULT_mult_6_net84925), .A3(MULT_mult_6_net84924), .ZN(
        MULT_mult_6_CARRYB_3__6_) );
  XNOR2_X2 MULT_mult_6_U3815 ( .A(MULT_mult_6_CARRYB_17__4_), .B(
        MULT_mult_6_ab_18__4_), .ZN(MULT_mult_6_n1384) );
  XNOR2_X2 MULT_mult_6_U3814 ( .A(MULT_mult_6_n1384), .B(MULT_mult_6_n1189), 
        .ZN(MULT_mult_6_SUMB_18__4_) );
  NAND2_X2 MULT_mult_6_U3813 ( .A1(MULT_mult_6_ab_1__10_), .A2(
        MULT_mult_6_ab_0__11_), .ZN(MULT_mult_6_n2332) );
  NAND2_X2 MULT_mult_6_U3812 ( .A1(MULT_mult_6_CARRYB_18__3_), .A2(
        MULT_mult_6_n1209), .ZN(MULT_mult_6_n2273) );
  XNOR2_X2 MULT_mult_6_U3811 ( .A(MULT_mult_6_CARRYB_5__6_), .B(
        MULT_mult_6_ab_6__6_), .ZN(MULT_mult_6_n1552) );
  NAND2_X4 MULT_mult_6_U3810 ( .A1(MULT_mult_6_SUMB_20__2_), .A2(
        MULT_mult_6_CARRYB_20__1_), .ZN(MULT_mult_6_n2163) );
  INV_X4 MULT_mult_6_U3809 ( .A(MULT_mult_6_ab_17__5_), .ZN(MULT_mult_6_n1381)
         );
  NAND2_X4 MULT_mult_6_U3808 ( .A1(MULT_mult_6_n1380), .A2(MULT_mult_6_n1381), 
        .ZN(MULT_mult_6_n1383) );
  NAND2_X2 MULT_mult_6_U3807 ( .A1(MULT_mult_6_SUMB_7__16_), .A2(
        MULT_mult_6_n858), .ZN(MULT_mult_6_n2254) );
  NAND2_X2 MULT_mult_6_U3806 ( .A1(MULT_mult_6_ab_14__7_), .A2(
        MULT_mult_6_CARRYB_13__7_), .ZN(MULT_mult_6_net85000) );
  XNOR2_X2 MULT_mult_6_U3805 ( .A(MULT_mult_6_n1936), .B(MULT_mult_6_n863), 
        .ZN(MULT_mult_6_SUMB_17__4_) );
  NOR2_X2 MULT_mult_6_U3804 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__12_) );
  INV_X4 MULT_mult_6_U3803 ( .A(MULT_mult_6_n2204), .ZN(MULT_mult_6_n1376) );
  INV_X2 MULT_mult_6_U3802 ( .A(MULT_mult_6_ab_13__12_), .ZN(MULT_mult_6_n1372) );
  NAND2_X4 MULT_mult_6_U3801 ( .A1(MULT_mult_6_n935), .A2(MULT_mult_6_net87136), .ZN(MULT_mult_6_net85979) );
  XNOR2_X2 MULT_mult_6_U3800 ( .A(MULT_mult_6_ab_20__4_), .B(
        MULT_mult_6_CARRYB_19__4_), .ZN(MULT_mult_6_n1371) );
  XNOR2_X2 MULT_mult_6_U3799 ( .A(MULT_mult_6_CARRYB_14__6_), .B(
        MULT_mult_6_ab_15__6_), .ZN(MULT_mult_6_n1370) );
  XNOR2_X2 MULT_mult_6_U3798 ( .A(MULT_mult_6_n1370), .B(MULT_mult_6_n1123), 
        .ZN(MULT_mult_6_SUMB_15__6_) );
  NAND2_X4 MULT_mult_6_U3797 ( .A1(MULT_mult_6_net87309), .A2(
        MULT_mult_6_net87308), .ZN(MULT_mult_6_n1367) );
  NAND2_X1 MULT_mult_6_U3796 ( .A1(MULT_mult_6_ab_5__17_), .A2(
        MULT_mult_6_CARRYB_4__17_), .ZN(MULT_mult_6_n2203) );
  NAND2_X1 MULT_mult_6_U3795 ( .A1(MULT_mult_6_ab_27__3_), .A2(
        MULT_mult_6_n1272), .ZN(MULT_mult_6_net80818) );
  NAND3_X4 MULT_mult_6_U3794 ( .A1(MULT_mult_6_n2302), .A2(
        MULT_mult_6_net79993), .A3(MULT_mult_6_net79992), .ZN(
        MULT_mult_6_CARRYB_22__4_) );
  NAND3_X2 MULT_mult_6_U3793 ( .A1(MULT_mult_6_n2037), .A2(MULT_mult_6_n2038), 
        .A3(MULT_mult_6_n2039), .ZN(MULT_mult_6_CARRYB_17__5_) );
  NAND3_X4 MULT_mult_6_U3792 ( .A1(MULT_mult_6_n1702), .A2(MULT_mult_6_n1704), 
        .A3(MULT_mult_6_n1703), .ZN(MULT_mult_6_CARRYB_14__5_) );
  NAND3_X4 MULT_mult_6_U3791 ( .A1(MULT_mult_6_n1707), .A2(MULT_mult_6_n1706), 
        .A3(MULT_mult_6_n1705), .ZN(MULT_mult_6_n1500) );
  NAND2_X2 MULT_mult_6_U3790 ( .A1(MULT_mult_6_ab_12__2_), .A2(
        MULT_mult_6_CARRYB_11__2_), .ZN(MULT_mult_6_n1997) );
  NAND3_X4 MULT_mult_6_U3789 ( .A1(MULT_mult_6_n1801), .A2(MULT_mult_6_n1800), 
        .A3(MULT_mult_6_n1799), .ZN(MULT_mult_6_CARRYB_23__0_) );
  INV_X4 MULT_mult_6_U3788 ( .A(MULT_mult_6_n2244), .ZN(MULT_mult_6_n1363) );
  NAND2_X4 MULT_mult_6_U3787 ( .A1(MULT_mult_6_n1364), .A2(MULT_mult_6_n1365), 
        .ZN(MULT_mult_6_SUMB_21__3_) );
  NOR2_X2 MULT_mult_6_U3786 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net77948), .ZN(MULT_mult_6_ab_5__12_) );
  INV_X1 MULT_mult_6_U3785 ( .A(MULT_mult_6_ab_5__12_), .ZN(
        MULT_mult_6_net87464) );
  NAND2_X4 MULT_mult_6_U3784 ( .A1(MULT_mult_6_net87064), .A2(
        MULT_mult_6_n1506), .ZN(MULT_mult_6_n1508) );
  NAND2_X4 MULT_mult_6_U3783 ( .A1(MULT_mult_6_net84706), .A2(
        MULT_mult_6_net84707), .ZN(MULT_mult_6_n1582) );
  NAND3_X2 MULT_mult_6_U3782 ( .A1(MULT_mult_6_net81205), .A2(
        MULT_mult_6_net81204), .A3(MULT_mult_6_net81206), .ZN(
        MULT_mult_6_n1439) );
  INV_X4 MULT_mult_6_U3781 ( .A(MULT_mult_6_n1439), .ZN(MULT_mult_6_n1362) );
  NAND3_X2 MULT_mult_6_U3780 ( .A1(MULT_mult_6_n2056), .A2(MULT_mult_6_n2055), 
        .A3(MULT_mult_6_n2054), .ZN(MULT_mult_6_CARRYB_3__19_) );
  NAND2_X1 MULT_mult_6_U3779 ( .A1(MULT_mult_6_CARRYB_11__16_), .A2(
        MULT_mult_6_SUMB_11__17_), .ZN(MULT_mult_6_n2309) );
  NAND2_X1 MULT_mult_6_U3778 ( .A1(MULT_mult_6_ab_12__16_), .A2(
        MULT_mult_6_SUMB_11__17_), .ZN(MULT_mult_6_n2308) );
  NAND3_X2 MULT_mult_6_U3777 ( .A1(MULT_mult_6_net80478), .A2(
        MULT_mult_6_net80479), .A3(MULT_mult_6_net80480), .ZN(
        MULT_mult_6_CARRYB_14__14_) );
  NAND2_X1 MULT_mult_6_U3776 ( .A1(MULT_mult_6_CARRYB_13__16_), .A2(
        MULT_mult_6_n1250), .ZN(MULT_mult_6_n2227) );
  XNOR2_X2 MULT_mult_6_U3775 ( .A(MULT_mult_6_ab_7__23_), .B(
        MULT_mult_6_CARRYB_6__23_), .ZN(MULT_mult_6_n1360) );
  XNOR2_X2 MULT_mult_6_U3774 ( .A(MULT_mult_6_n1360), .B(
        MULT_mult_6_SUMB_6__24_), .ZN(MULT_mult_6_SUMB_7__23_) );
  NOR2_X2 MULT_mult_6_U3773 ( .A1(MULT_mult_6_net77868), .A2(MULT_mult_6_n242), 
        .ZN(MULT_mult_6_ab_1__1_) );
  XNOR2_X2 MULT_mult_6_U3772 ( .A(MULT_mult_6_ab_6__23_), .B(
        MULT_mult_6_CARRYB_5__23_), .ZN(MULT_mult_6_n1359) );
  XNOR2_X2 MULT_mult_6_U3771 ( .A(MULT_mult_6_SUMB_5__24_), .B(
        MULT_mult_6_n1359), .ZN(MULT_mult_6_SUMB_6__23_) );
  INV_X2 MULT_mult_6_U3770 ( .A(MULT_mult_6_net83151), .ZN(
        MULT_mult_6_net87573) );
  NAND2_X4 MULT_mult_6_U3769 ( .A1(MULT_mult_6_SUMB_7__12_), .A2(
        MULT_mult_6_CARRYB_7__11_), .ZN(MULT_mult_6_n2126) );
  INV_X4 MULT_mult_6_U3768 ( .A(MULT_mult_6_n362), .ZN(MULT_mult_6_n1355) );
  NAND2_X4 MULT_mult_6_U3767 ( .A1(MULT_mult_6_n1357), .A2(MULT_mult_6_n1358), 
        .ZN(MULT_mult_6_SUMB_5__13_) );
  NAND2_X2 MULT_mult_6_U3766 ( .A1(MULT_mult_6_n362), .A2(MULT_mult_6_n1356), 
        .ZN(MULT_mult_6_n1357) );
  NAND2_X4 MULT_mult_6_U3765 ( .A1(MULT_mult_6_n1353), .A2(MULT_mult_6_n1354), 
        .ZN(MULT_mult_6_SUMB_2__15_) );
  NAND2_X4 MULT_mult_6_U3764 ( .A1(MULT_mult_6_n1351), .A2(MULT_mult_6_n1352), 
        .ZN(MULT_mult_6_n1354) );
  NAND3_X2 MULT_mult_6_U3763 ( .A1(MULT_mult_6_net84297), .A2(
        MULT_mult_6_net84298), .A3(MULT_mult_6_net84299), .ZN(
        MULT_mult_6_CARRYB_2__24_) );
  XNOR2_X2 MULT_mult_6_U3762 ( .A(MULT_mult_6_n1258), .B(MULT_mult_6_n1350), 
        .ZN(MULT_mult_6_SUMB_5__9_) );
  INV_X4 MULT_mult_6_U3761 ( .A(MULT_mult_6_net93878), .ZN(
        MULT_mult_6_net85540) );
  NAND2_X4 MULT_mult_6_U3760 ( .A1(MULT_mult_6_n1455), .A2(MULT_mult_6_n2071), 
        .ZN(MULT_mult_6_n1585) );
  INV_X4 MULT_mult_6_U3759 ( .A(MULT_mult_6_n2109), .ZN(MULT_mult_6_n1346) );
  INV_X2 MULT_mult_6_U3758 ( .A(MULT_mult_6_ab_2__17_), .ZN(
        MULT_mult_6_net87682) );
  XNOR2_X2 MULT_mult_6_U3757 ( .A(MULT_mult_6_ab_3__24_), .B(
        MULT_mult_6_CARRYB_2__24_), .ZN(MULT_mult_6_n1342) );
  XNOR2_X2 MULT_mult_6_U3756 ( .A(MULT_mult_6_n1342), .B(
        MULT_mult_6_SUMB_2__25_), .ZN(MULT_mult_6_SUMB_3__24_) );
  NAND2_X2 MULT_mult_6_U3755 ( .A1(MULT_mult_6_net87683), .A2(
        MULT_mult_6_ab_2__17_), .ZN(MULT_mult_6_n1941) );
  NAND2_X1 MULT_mult_6_U3754 ( .A1(MULT_mult_6_ab_13__12_), .A2(
        MULT_mult_6_CARRYB_12__12_), .ZN(MULT_mult_6_n2125) );
  NAND2_X2 MULT_mult_6_U3753 ( .A1(MULT_mult_6_net88704), .A2(
        MULT_mult_6_CARRYB_8__16_), .ZN(MULT_mult_6_n2304) );
  INV_X2 MULT_mult_6_U3752 ( .A(MULT_mult_6_CARRYB_6__9_), .ZN(
        MULT_mult_6_n1699) );
  XNOR2_X2 MULT_mult_6_U3751 ( .A(MULT_mult_6_n165), .B(MULT_mult_6_n1831), 
        .ZN(MULT_mult_6_n1340) );
  XNOR2_X2 MULT_mult_6_U3750 ( .A(MULT_mult_6_n1340), .B(MULT_mult_6_n1864), 
        .ZN(MULT_mult_6_SUMB_8__7_) );
  XNOR2_X2 MULT_mult_6_U3749 ( .A(MULT_mult_6_CARRYB_8__14_), .B(
        MULT_mult_6_ab_9__14_), .ZN(MULT_mult_6_n1587) );
  XNOR2_X2 MULT_mult_6_U3748 ( .A(MULT_mult_6_CARRYB_5__15_), .B(
        MULT_mult_6_ab_6__15_), .ZN(MULT_mult_6_n1695) );
  NAND2_X2 MULT_mult_6_U3747 ( .A1(MULT_mult_6_n2197), .A2(MULT_mult_6_n848), 
        .ZN(MULT_mult_6_n1790) );
  NAND2_X4 MULT_mult_6_U3746 ( .A1(MULT_mult_6_ab_2__20_), .A2(
        MULT_mult_6_SUMB_1__21_), .ZN(MULT_mult_6_n2052) );
  NAND3_X2 MULT_mult_6_U3745 ( .A1(MULT_mult_6_n1746), .A2(MULT_mult_6_n1745), 
        .A3(MULT_mult_6_n1744), .ZN(MULT_mult_6_CARRYB_5__10_) );
  XNOR2_X2 MULT_mult_6_U3744 ( .A(MULT_mult_6_n1339), .B(MULT_mult_6_n1229), 
        .ZN(MULT_mult_6_SUMB_4__10_) );
  OR2_X1 MULT_mult_6_U3743 ( .A1(MULT_mult_6_net70461), .A2(
        MULT_mult_6_net84698), .ZN(MULT_mult_6_n1338) );
  XNOR2_X2 MULT_mult_6_U3742 ( .A(MULT_mult_6_CARRYB_16__14_), .B(
        MULT_mult_6_n1338), .ZN(MULT_mult_6_n1369) );
  NAND2_X4 MULT_mult_6_U3741 ( .A1(MULT_mult_6_n1790), .A2(MULT_mult_6_n1791), 
        .ZN(MULT_mult_6_SUMB_5__19_) );
  NAND2_X4 MULT_mult_6_U3740 ( .A1(MULT_mult_6_n2044), .A2(MULT_mult_6_n2045), 
        .ZN(MULT_mult_6_n2047) );
  NAND2_X4 MULT_mult_6_U3739 ( .A1(MULT_mult_6_n1336), .A2(MULT_mult_6_n1337), 
        .ZN(MULT_mult_6_SUMB_21__4_) );
  NAND3_X4 MULT_mult_6_U3737 ( .A1(MULT_mult_6_net80565), .A2(
        MULT_mult_6_net83296), .A3(MULT_mult_6_net80566), .ZN(
        MULT_mult_6_CARRYB_16__7_) );
  NAND2_X4 MULT_mult_6_U3736 ( .A1(MULT_mult_6_ab_21__1_), .A2(
        MULT_mult_6_CARRYB_20__1_), .ZN(MULT_mult_6_n2162) );
  INV_X4 MULT_mult_6_U3735 ( .A(MULT_mult_6_n621), .ZN(MULT_mult_6_n1761) );
  NOR2_X1 MULT_mult_6_U3734 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net77948), .ZN(MULT_mult_6_ab_5__13_) );
  NAND2_X2 MULT_mult_6_U3733 ( .A1(MULT_mult_6_ab_9__16_), .A2(
        MULT_mult_6_net88704), .ZN(MULT_mult_6_n2305) );
  NAND3_X4 MULT_mult_6_U3732 ( .A1(MULT_mult_6_n1335), .A2(MULT_mult_6_n1334), 
        .A3(MULT_mult_6_n1333), .ZN(MULT_mult_6_CARRYB_7__6_) );
  NAND2_X2 MULT_mult_6_U3731 ( .A1(MULT_mult_6_n29), .A2(
        MULT_mult_6_SUMB_5__8_), .ZN(MULT_mult_6_n1332) );
  NAND2_X1 MULT_mult_6_U3729 ( .A1(MULT_mult_6_CARRYB_5__7_), .A2(
        MULT_mult_6_ab_6__7_), .ZN(MULT_mult_6_n1330) );
  XOR2_X2 MULT_mult_6_U3728 ( .A(MULT_mult_6_n1329), .B(MULT_mult_6_n853), .Z(
        MULT_mult_6_SUMB_6__7_) );
  INV_X4 MULT_mult_6_U3727 ( .A(MULT_mult_6_CARRYB_3__8_), .ZN(
        MULT_mult_6_n1327) );
  INV_X4 MULT_mult_6_U3726 ( .A(MULT_mult_6_ab_4__8_), .ZN(MULT_mult_6_n1326)
         );
  NAND2_X2 MULT_mult_6_U3725 ( .A1(MULT_mult_6_n1326), .A2(MULT_mult_6_n1327), 
        .ZN(MULT_mult_6_n1328) );
  NAND3_X4 MULT_mult_6_U3724 ( .A1(MULT_mult_6_n2028), .A2(MULT_mult_6_n2029), 
        .A3(MULT_mult_6_n2030), .ZN(MULT_mult_6_CARRYB_3__11_) );
  NAND2_X4 MULT_mult_6_U3723 ( .A1(MULT_mult_6_n1662), .A2(MULT_mult_6_n1661), 
        .ZN(MULT_mult_6_net80993) );
  NAND2_X2 MULT_mult_6_U3722 ( .A1(MULT_mult_6_SUMB_8__15_), .A2(
        MULT_mult_6_n1235), .ZN(MULT_mult_6_n2292) );
  NOR2_X1 MULT_mult_6_U3721 ( .A1(MULT_mult_6_net124723), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__16_) );
  NAND2_X4 MULT_mult_6_U3720 ( .A1(MULT_mult_6_net84948), .A2(
        MULT_mult_6_net84947), .ZN(MULT_mult_6_n1901) );
  XNOR2_X2 MULT_mult_6_U3719 ( .A(MULT_mult_6_CARRYB_4__9_), .B(
        MULT_mult_6_ab_5__9_), .ZN(MULT_mult_6_n1350) );
  XNOR2_X2 MULT_mult_6_U3718 ( .A(MULT_mult_6_ab_13__13_), .B(
        MULT_mult_6_CARRYB_12__13_), .ZN(MULT_mult_6_n1323) );
  NAND2_X4 MULT_mult_6_U3717 ( .A1(MULT_mult_6_net83120), .A2(
        MULT_mult_6_ab_22__7_), .ZN(MULT_mult_6_n1759) );
  NAND2_X2 MULT_mult_6_U3716 ( .A1(MULT_mult_6_ab_6__17_), .A2(
        MULT_mult_6_SUMB_5__18_), .ZN(MULT_mult_6_n2246) );
  NAND3_X2 MULT_mult_6_U3715 ( .A1(MULT_mult_6_n1715), .A2(MULT_mult_6_n1714), 
        .A3(MULT_mult_6_n1716), .ZN(MULT_mult_6_CARRYB_3__17_) );
  INV_X8 MULT_mult_6_U3714 ( .A(MULT_mult_6_CARRYB_17__9_), .ZN(
        MULT_mult_6_net83850) );
  NAND2_X4 MULT_mult_6_U3713 ( .A1(MULT_mult_6_SUMB_1__20_), .A2(
        MULT_mult_6_ab_2__19_), .ZN(MULT_mult_6_n2144) );
  NAND2_X4 MULT_mult_6_U3712 ( .A1(MULT_mult_6_n1541), .A2(MULT_mult_6_n1540), 
        .ZN(MULT_mult_6_n1543) );
  XNOR2_X2 MULT_mult_6_U3711 ( .A(MULT_mult_6_ab_3__25_), .B(
        MULT_mult_6_CARRYB_2__25_), .ZN(MULT_mult_6_n1322) );
  XNOR2_X2 MULT_mult_6_U3710 ( .A(MULT_mult_6_n1219), .B(MULT_mult_6_n1322), 
        .ZN(MULT_mult_6_SUMB_3__25_) );
  NAND3_X2 MULT_mult_6_U3709 ( .A1(MULT_mult_6_net82099), .A2(
        MULT_mult_6_n1923), .A3(MULT_mult_6_net82101), .ZN(
        MULT_mult_6_CARRYB_9__4_) );
  NOR2_X4 MULT_mult_6_U3708 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net77932), .ZN(MULT_mult_6_ab_7__13_) );
  INV_X1 MULT_mult_6_U3707 ( .A(MULT_mult_6_ab_7__13_), .ZN(
        MULT_mult_6_net88156) );
  NAND2_X2 MULT_mult_6_U3706 ( .A1(MULT_mult_6_n1246), .A2(
        MULT_mult_6_ab_3__9_), .ZN(MULT_mult_6_n1655) );
  XNOR2_X2 MULT_mult_6_U3705 ( .A(MULT_mult_6_net88165), .B(
        MULT_mult_6_SUMB_17__13_), .ZN(MULT_mult_6_SUMB_18__12_) );
  NAND2_X4 MULT_mult_6_U3704 ( .A1(MULT_mult_6_n1318), .A2(MULT_mult_6_n1319), 
        .ZN(MULT_mult_6_SUMB_7__12_) );
  NAND2_X2 MULT_mult_6_U3703 ( .A1(MULT_mult_6_n2095), .A2(MULT_mult_6_n1733), 
        .ZN(MULT_mult_6_n1727) );
  NAND3_X2 MULT_mult_6_U3702 ( .A1(MULT_mult_6_net82557), .A2(
        MULT_mult_6_net82558), .A3(MULT_mult_6_net82556), .ZN(
        MULT_mult_6_CARRYB_14__11_) );
  NAND2_X1 MULT_mult_6_U3701 ( .A1(MULT_mult_6_ab_20__8_), .A2(
        MULT_mult_6_CARRYB_19__8_), .ZN(MULT_mult_6_net81955) );
  NAND3_X4 MULT_mult_6_U3700 ( .A1(MULT_mult_6_net88209), .A2(
        MULT_mult_6_net88210), .A3(MULT_mult_6_net88211), .ZN(
        MULT_mult_6_CARRYB_5__5_) );
  NAND3_X2 MULT_mult_6_U3699 ( .A1(MULT_mult_6_net88206), .A2(
        MULT_mult_6_net88207), .A3(MULT_mult_6_net88208), .ZN(
        MULT_mult_6_CARRYB_4__6_) );
  XOR2_X2 MULT_mult_6_U3698 ( .A(MULT_mult_6_n1316), .B(MULT_mult_6_SUMB_6__4_), .Z(MULT_mult_6_SUMB_7__3_) );
  XOR2_X2 MULT_mult_6_U3697 ( .A(MULT_mult_6_ab_7__3_), .B(
        MULT_mult_6_CARRYB_6__3_), .Z(MULT_mult_6_n1316) );
  NAND3_X2 MULT_mult_6_U3696 ( .A1(MULT_mult_6_n2091), .A2(MULT_mult_6_n2090), 
        .A3(MULT_mult_6_n2089), .ZN(MULT_mult_6_CARRYB_4__13_) );
  NAND2_X4 MULT_mult_6_U3695 ( .A1(MULT_mult_6_n952), .A2(MULT_mult_6_n1282), 
        .ZN(MULT_mult_6_n1451) );
  INV_X4 MULT_mult_6_U3694 ( .A(MULT_mult_6_CARRYB_14__11_), .ZN(
        MULT_mult_6_n1770) );
  NAND2_X2 MULT_mult_6_U3693 ( .A1(MULT_mult_6_CARRYB_8__16_), .A2(
        MULT_mult_6_n1600), .ZN(MULT_mult_6_n1601) );
  INV_X4 MULT_mult_6_U3692 ( .A(MULT_mult_6_CARRYB_26__3_), .ZN(
        MULT_mult_6_n1533) );
  NAND2_X1 MULT_mult_6_U3691 ( .A1(MULT_mult_6_ab_9__21_), .A2(
        MULT_mult_6_SUMB_8__22_), .ZN(MULT_mult_6_n1687) );
  NAND2_X4 MULT_mult_6_U3690 ( .A1(MULT_mult_6_ab_3__8_), .A2(
        MULT_mult_6_n1427), .ZN(MULT_mult_6_n1906) );
  XNOR2_X2 MULT_mult_6_U3689 ( .A(MULT_mult_6_ab_9__21_), .B(
        MULT_mult_6_CARRYB_8__21_), .ZN(MULT_mult_6_n1314) );
  XNOR2_X2 MULT_mult_6_U3688 ( .A(MULT_mult_6_n1314), .B(
        MULT_mult_6_SUMB_8__22_), .ZN(MULT_mult_6_SUMB_9__21_) );
  NOR2_X1 MULT_mult_6_U3687 ( .A1(MULT_mult_6_net124723), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__16_) );
  NOR2_X2 MULT_mult_6_U3686 ( .A1(MULT_mult_6_net88344), .A2(
        MULT_mult_6_net77940), .ZN(MULT_mult_6_ab_6__16_) );
  INV_X4 MULT_mult_6_U3685 ( .A(MULT_mult_6_net85465), .ZN(
        MULT_mult_6_net87064) );
  INV_X2 MULT_mult_6_U3684 ( .A(MULT_mult_6_net70474), .ZN(
        MULT_mult_6_net81080) );
  XNOR2_X2 MULT_mult_6_U3683 ( .A(MULT_mult_6_n1312), .B(MULT_mult_6_n1369), 
        .ZN(MULT_mult_6_SUMB_17__14_) );
  XNOR2_X2 MULT_mult_6_U3682 ( .A(MULT_mult_6_CARRYB_3__11_), .B(
        MULT_mult_6_ab_4__11_), .ZN(MULT_mult_6_n1311) );
  XNOR2_X2 MULT_mult_6_U3681 ( .A(MULT_mult_6_net121785), .B(MULT_mult_6_n1311), .ZN(MULT_mult_6_SUMB_4__11_) );
  NAND2_X4 MULT_mult_6_U3680 ( .A1(MULT_mult_6_SUMB_3__21_), .A2(
        MULT_mult_6_n1009), .ZN(MULT_mult_6_n2239) );
  INV_X4 MULT_mult_6_U3679 ( .A(MULT_mult_6_ab_3__18_), .ZN(MULT_mult_6_n1546)
         );
  NOR2_X1 MULT_mult_6_U3677 ( .A1(MULT_mult_6_net70454), .A2(
        MULT_mult_6_net77946), .ZN(MULT_mult_6_ab_5__10_) );
  NOR2_X1 MULT_mult_6_U3676 ( .A1(MULT_mult_6_net91660), .A2(
        MULT_mult_6_net70455), .ZN(MULT_mult_6_ab_20__10_) );
  NAND3_X2 MULT_mult_6_U3675 ( .A1(MULT_mult_6_n2011), .A2(MULT_mult_6_n2012), 
        .A3(MULT_mult_6_n2376), .ZN(MULT_mult_6_CARRYB_19__7_) );
  NAND3_X2 MULT_mult_6_U3674 ( .A1(MULT_mult_6_net80676), .A2(
        MULT_mult_6_net80675), .A3(MULT_mult_6_net80674), .ZN(
        MULT_mult_6_CARRYB_21__6_) );
  XNOR2_X2 MULT_mult_6_U3673 ( .A(MULT_mult_6_SUMB_25__5_), .B(
        MULT_mult_6_n1310), .ZN(MULT_mult_6_SUMB_26__4_) );
  XNOR2_X2 MULT_mult_6_U3671 ( .A(MULT_mult_6_n1973), .B(MULT_mult_6_n1308), 
        .ZN(MULT_mult_6_SUMB_14__6_) );
  NAND3_X4 MULT_mult_6_U3670 ( .A1(MULT_mult_6_n1832), .A2(MULT_mult_6_n1833), 
        .A3(MULT_mult_6_n1834), .ZN(MULT_mult_6_CARRYB_11__4_) );
  NAND2_X4 MULT_mult_6_U3669 ( .A1(MULT_mult_6_n1780), .A2(MULT_mult_6_n896), 
        .ZN(MULT_mult_6_n2149) );
  NAND3_X4 MULT_mult_6_U3668 ( .A1(MULT_mult_6_n1307), .A2(MULT_mult_6_n1306), 
        .A3(MULT_mult_6_n1305), .ZN(MULT_mult_6_CARRYB_11__13_) );
  NAND2_X2 MULT_mult_6_U3667 ( .A1(MULT_mult_6_SUMB_10__14_), .A2(
        MULT_mult_6_ab_11__13_), .ZN(MULT_mult_6_n1307) );
  NAND2_X2 MULT_mult_6_U3666 ( .A1(MULT_mult_6_SUMB_10__14_), .A2(
        MULT_mult_6_CARRYB_10__13_), .ZN(MULT_mult_6_n1306) );
  NAND2_X1 MULT_mult_6_U3665 ( .A1(MULT_mult_6_CARRYB_10__13_), .A2(
        MULT_mult_6_ab_11__13_), .ZN(MULT_mult_6_n1305) );
  NAND2_X2 MULT_mult_6_U3664 ( .A1(MULT_mult_6_SUMB_9__15_), .A2(
        MULT_mult_6_CARRYB_9__14_), .ZN(MULT_mult_6_n1304) );
  NAND2_X2 MULT_mult_6_U3663 ( .A1(MULT_mult_6_SUMB_9__15_), .A2(
        MULT_mult_6_ab_10__14_), .ZN(MULT_mult_6_n1303) );
  INV_X8 MULT_mult_6_U3662 ( .A(MULT_mult_6_CARRYB_6__13_), .ZN(
        MULT_mult_6_net88157) );
  INV_X1 MULT_mult_6_U3661 ( .A(MULT_mult_6_net88157), .ZN(
        MULT_mult_6_net88444) );
  NAND3_X2 MULT_mult_6_U3660 ( .A1(MULT_mult_6_n2061), .A2(MULT_mult_6_n2062), 
        .A3(MULT_mult_6_n2063), .ZN(MULT_mult_6_CARRYB_11__5_) );
  NAND2_X2 MULT_mult_6_U3659 ( .A1(MULT_mult_6_ab_13__4_), .A2(
        MULT_mult_6_CARRYB_12__4_), .ZN(MULT_mult_6_n1639) );
  NAND2_X2 MULT_mult_6_U3658 ( .A1(MULT_mult_6_CARRYB_12__4_), .A2(
        MULT_mult_6_SUMB_12__5_), .ZN(MULT_mult_6_n1641) );
  NAND2_X2 MULT_mult_6_U3657 ( .A1(MULT_mult_6_SUMB_6__8_), .A2(
        MULT_mult_6_ab_7__7_), .ZN(MULT_mult_6_n1823) );
  NAND2_X2 MULT_mult_6_U3656 ( .A1(MULT_mult_6_CARRYB_6__7_), .A2(
        MULT_mult_6_SUMB_6__8_), .ZN(MULT_mult_6_n1824) );
  NAND3_X4 MULT_mult_6_U3655 ( .A1(MULT_mult_6_n1826), .A2(MULT_mult_6_n1827), 
        .A3(MULT_mult_6_n1825), .ZN(MULT_mult_6_CARRYB_8__6_) );
  INV_X1 MULT_mult_6_U3654 ( .A(MULT_mult_6_SUMB_12__5_), .ZN(
        MULT_mult_6_n1298) );
  INV_X4 MULT_mult_6_U3653 ( .A(MULT_mult_6_n1635), .ZN(MULT_mult_6_n1297) );
  NAND2_X4 MULT_mult_6_U3652 ( .A1(MULT_mult_6_n1299), .A2(MULT_mult_6_n1300), 
        .ZN(MULT_mult_6_SUMB_13__4_) );
  NAND2_X2 MULT_mult_6_U3651 ( .A1(MULT_mult_6_n1297), .A2(MULT_mult_6_n1194), 
        .ZN(MULT_mult_6_n1300) );
  NAND2_X2 MULT_mult_6_U3650 ( .A1(MULT_mult_6_n1635), .A2(MULT_mult_6_n1298), 
        .ZN(MULT_mult_6_n1299) );
  NAND2_X2 MULT_mult_6_U3649 ( .A1(MULT_mult_6_ab_9__6_), .A2(
        MULT_mult_6_SUMB_8__7_), .ZN(MULT_mult_6_n1293) );
  NAND2_X2 MULT_mult_6_U3648 ( .A1(MULT_mult_6_n1375), .A2(MULT_mult_6_n2204), 
        .ZN(MULT_mult_6_n1378) );
  NAND2_X4 MULT_mult_6_U3647 ( .A1(MULT_mult_6_n1377), .A2(MULT_mult_6_n1378), 
        .ZN(MULT_mult_6_SUMB_7__15_) );
  NAND2_X4 MULT_mult_6_U3646 ( .A1(MULT_mult_6_n1755), .A2(
        MULT_mult_6_net87573), .ZN(MULT_mult_6_n1756) );
  NAND2_X4 MULT_mult_6_U3645 ( .A1(MULT_mult_6_CARRYB_26__0_), .A2(
        MULT_mult_6_n1281), .ZN(MULT_mult_6_net80769) );
  NAND2_X4 MULT_mult_6_U3644 ( .A1(MULT_mult_6_SUMB_26__1_), .A2(
        MULT_mult_6_ab_27__0_), .ZN(MULT_mult_6_net80768) );
  NAND2_X4 MULT_mult_6_U3643 ( .A1(MULT_mult_6_n1430), .A2(
        MULT_mult_6_ab_7__8_), .ZN(MULT_mult_6_n2058) );
  INV_X1 MULT_mult_6_U3642 ( .A(MULT_mult_6_ab_10__8_), .ZN(MULT_mult_6_n1503)
         );
  NOR2_X2 MULT_mult_6_U3641 ( .A1(MULT_mult_6_net77914), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__7_) );
  INV_X8 MULT_mult_6_U3640 ( .A(MULT_mult_6_n1503), .ZN(MULT_mult_6_n1288) );
  NAND2_X4 MULT_mult_6_U3639 ( .A1(MULT_mult_6_n1288), .A2(MULT_mult_6_n1289), 
        .ZN(MULT_mult_6_n1291) );
  NAND2_X2 MULT_mult_6_U3638 ( .A1(MULT_mult_6_CARRYB_9__8_), .A2(
        MULT_mult_6_n1503), .ZN(MULT_mult_6_n1290) );
  INV_X2 MULT_mult_6_U3637 ( .A(MULT_mult_6_ab_12__7_), .ZN(MULT_mult_6_n1285)
         );
  NAND2_X4 MULT_mult_6_U3636 ( .A1(MULT_mult_6_n1287), .A2(MULT_mult_6_n2019), 
        .ZN(MULT_mult_6_n1902) );
  NAND2_X4 MULT_mult_6_U3635 ( .A1(MULT_mult_6_n1286), .A2(MULT_mult_6_n1285), 
        .ZN(MULT_mult_6_n1287) );
  NAND2_X2 MULT_mult_6_U3634 ( .A1(MULT_mult_6_CARRYB_4__19_), .A2(
        MULT_mult_6_SUMB_4__20_), .ZN(MULT_mult_6_n2242) );
  NAND3_X2 MULT_mult_6_U3633 ( .A1(MULT_mult_6_net80957), .A2(
        MULT_mult_6_net80956), .A3(MULT_mult_6_net80958), .ZN(
        MULT_mult_6_net88525) );
  NAND2_X2 MULT_mult_6_U3632 ( .A1(MULT_mult_6_ab_3__10_), .A2(
        MULT_mult_6_n1203), .ZN(MULT_mult_6_n1645) );
  NAND2_X2 MULT_mult_6_U3631 ( .A1(MULT_mult_6_SUMB_13__10_), .A2(
        MULT_mult_6_net85043), .ZN(MULT_mult_6_n1940) );
  OR2_X1 MULT_mult_6_U3630 ( .A1(MULT_mult_6_net70455), .A2(
        MULT_mult_6_net85716), .ZN(MULT_mult_6_n1283) );
  XNOR2_X2 MULT_mult_6_U3629 ( .A(MULT_mult_6_CARRYB_19__11_), .B(
        MULT_mult_6_n1283), .ZN(MULT_mult_6_n2142) );
  INV_X4 MULT_mult_6_U3628 ( .A(MULT_mult_6_n1449), .ZN(MULT_mult_6_n1282) );
  INV_X2 MULT_mult_6_U3627 ( .A(MULT_mult_6_net88655), .ZN(
        MULT_mult_6_net88656) );
  XNOR2_X2 MULT_mult_6_U3626 ( .A(MULT_mult_6_net86427), .B(
        MULT_mult_6_net88656), .ZN(MULT_mult_6_n1281) );
  INV_X2 MULT_mult_6_U3624 ( .A(MULT_mult_6_SUMB_8__21_), .ZN(
        MULT_mult_6_n1277) );
  XNOR2_X2 MULT_mult_6_U3623 ( .A(MULT_mult_6_CARRYB_10__4_), .B(
        MULT_mult_6_ab_11__4_), .ZN(MULT_mult_6_n1276) );
  NAND2_X1 MULT_mult_6_U3622 ( .A1(MULT_mult_6_CARRYB_12__17_), .A2(
        MULT_mult_6_n1240), .ZN(MULT_mult_6_n2224) );
  NAND2_X1 MULT_mult_6_U3621 ( .A1(MULT_mult_6_ab_13__17_), .A2(
        MULT_mult_6_n1240), .ZN(MULT_mult_6_n2223) );
  XNOR2_X2 MULT_mult_6_U3620 ( .A(MULT_mult_6_CARRYB_25__4_), .B(
        MULT_mult_6_ab_26__4_), .ZN(MULT_mult_6_n1310) );
  XNOR2_X2 MULT_mult_6_U3619 ( .A(MULT_mult_6_CARRYB_22__8_), .B(
        MULT_mult_6_ab_23__8_), .ZN(MULT_mult_6_n1273) );
  NAND3_X2 MULT_mult_6_U3618 ( .A1(MULT_mult_6_n1575), .A2(MULT_mult_6_n1574), 
        .A3(MULT_mult_6_n1573), .ZN(MULT_mult_6_CARRYB_13__13_) );
  INV_X4 MULT_mult_6_U3617 ( .A(MULT_mult_6_CARRYB_10__5_), .ZN(
        MULT_mult_6_n1781) );
  INV_X4 MULT_mult_6_U3616 ( .A(MULT_mult_6_n1781), .ZN(MULT_mult_6_n1271) );
  FA_X1 MULT_mult_6_U3615 ( .A(MULT_mult_6_ab_15__15_), .B(
        MULT_mult_6_CARRYB_14__15_), .CI(MULT_mult_6_SUMB_14__16_), .S(
        MULT_mult_6_n1269) );
  INV_X2 MULT_mult_6_U3614 ( .A(MULT_mult_6_net88859), .ZN(
        MULT_mult_6_net88860) );
  INV_X2 MULT_mult_6_U3613 ( .A(MULT_mult_6_net88867), .ZN(
        MULT_mult_6_net88868) );
  XNOR2_X2 MULT_mult_6_U3612 ( .A(MULT_mult_6_n1268), .B(MULT_mult_6_n1241), 
        .ZN(MULT_mult_6_SUMB_18__3_) );
  XNOR2_X2 MULT_mult_6_U3611 ( .A(MULT_mult_6_ab_13__2_), .B(
        MULT_mult_6_CARRYB_12__2_), .ZN(MULT_mult_6_n1267) );
  XNOR2_X2 MULT_mult_6_U3610 ( .A(MULT_mult_6_n1267), .B(
        MULT_mult_6_SUMB_12__3_), .ZN(MULT_mult_6_SUMB_13__2_) );
  XNOR2_X2 MULT_mult_6_U3609 ( .A(MULT_mult_6_ab_10__4_), .B(
        MULT_mult_6_SUMB_9__5_), .ZN(MULT_mult_6_n1903) );
  XNOR2_X2 MULT_mult_6_U3608 ( .A(MULT_mult_6_n1903), .B(
        MULT_mult_6_CARRYB_9__4_), .ZN(MULT_mult_6_SUMB_10__4_) );
  INV_X4 MULT_mult_6_U3607 ( .A(MULT_mult_6_n1263), .ZN(MULT_mult_6_n1264) );
  INV_X4 MULT_mult_6_U3606 ( .A(MULT_mult_6_net124563), .ZN(
        MULT_mult_6_net85456) );
  INV_X4 MULT_mult_6_U3605 ( .A(MULT_mult_6_n1730), .ZN(MULT_mult_6_n1627) );
  NAND2_X4 MULT_mult_6_U3604 ( .A1(MULT_mult_6_CARRYB_18__7_), .A2(
        MULT_mult_6_ab_19__7_), .ZN(MULT_mult_6_n2010) );
  XNOR2_X2 MULT_mult_6_U3601 ( .A(MULT_mult_6_ab_9__19_), .B(
        MULT_mult_6_CARRYB_8__19_), .ZN(MULT_mult_6_n1257) );
  XNOR2_X2 MULT_mult_6_U3600 ( .A(MULT_mult_6_SUMB_8__20_), .B(
        MULT_mult_6_n1257), .ZN(MULT_mult_6_SUMB_9__19_) );
  NAND2_X1 MULT_mult_6_U3599 ( .A1(MULT_mult_6_ab_7__23_), .A2(
        MULT_mult_6_n1213), .ZN(MULT_mult_6_n2267) );
  NAND2_X1 MULT_mult_6_U3598 ( .A1(MULT_mult_6_CARRYB_6__23_), .A2(
        MULT_mult_6_n1213), .ZN(MULT_mult_6_n2268) );
  NAND3_X2 MULT_mult_6_U3597 ( .A1(MULT_mult_6_net79906), .A2(
        MULT_mult_6_net79905), .A3(MULT_mult_6_net79904), .ZN(
        MULT_mult_6_CARRYB_23__5_) );
  NOR2_X2 MULT_mult_6_U3596 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net77956), .ZN(MULT_mult_6_ab_4__12_) );
  NAND3_X2 MULT_mult_6_U3595 ( .A1(MULT_mult_6_n2091), .A2(MULT_mult_6_n2090), 
        .A3(MULT_mult_6_n2089), .ZN(MULT_mult_6_n1255) );
  NAND2_X4 MULT_mult_6_U3594 ( .A1(MULT_mult_6_SUMB_9__12_), .A2(
        MULT_mult_6_net82678), .ZN(MULT_mult_6_net80956) );
  XNOR2_X2 MULT_mult_6_U3593 ( .A(MULT_mult_6_n1254), .B(MULT_mult_6_n24), 
        .ZN(MULT_mult_6_SUMB_19__2_) );
  NAND2_X4 MULT_mult_6_U3592 ( .A1(MULT_mult_6_net86662), .A2(
        MULT_mult_6_ab_18__5_), .ZN(MULT_mult_6_n2232) );
  NAND3_X2 MULT_mult_6_U3591 ( .A1(MULT_mult_6_n1673), .A2(MULT_mult_6_n1674), 
        .A3(MULT_mult_6_n1675), .ZN(MULT_mult_6_CARRYB_12__3_) );
  NAND2_X2 MULT_mult_6_U3590 ( .A1(MULT_mult_6_ab_13__3_), .A2(
        MULT_mult_6_CARRYB_12__3_), .ZN(MULT_mult_6_n1678) );
  NAND3_X2 MULT_mult_6_U3589 ( .A1(MULT_mult_6_net79906), .A2(
        MULT_mult_6_net79905), .A3(MULT_mult_6_net79904), .ZN(
        MULT_mult_6_n1251) );
  INV_X2 MULT_mult_6_U3588 ( .A(MULT_mult_6_n615), .ZN(MULT_mult_6_n1250) );
  NOR2_X2 MULT_mult_6_U3587 ( .A1(MULT_mult_6_net81424), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__15_) );
  NAND2_X2 MULT_mult_6_U3586 ( .A1(MULT_mult_6_CARRYB_14__12_), .A2(
        MULT_mult_6_ab_15__12_), .ZN(MULT_mult_6_n1852) );
  XNOR2_X2 MULT_mult_6_U3584 ( .A(MULT_mult_6_CARRYB_5__20_), .B(
        MULT_mult_6_ab_6__20_), .ZN(MULT_mult_6_n1247) );
  XNOR2_X2 MULT_mult_6_U3583 ( .A(MULT_mult_6_SUMB_5__21_), .B(
        MULT_mult_6_n1247), .ZN(MULT_mult_6_SUMB_6__20_) );
  NAND3_X2 MULT_mult_6_U3582 ( .A1(MULT_mult_6_n2241), .A2(MULT_mult_6_n2240), 
        .A3(MULT_mult_6_n2242), .ZN(MULT_mult_6_CARRYB_5__19_) );
  INV_X4 MULT_mult_6_U3581 ( .A(MULT_mult_6_n1245), .ZN(MULT_mult_6_n1246) );
  XNOR2_X2 MULT_mult_6_U3580 ( .A(MULT_mult_6_ab_2__25_), .B(MULT_mult_6_n349), 
        .ZN(MULT_mult_6_n1244) );
  XNOR2_X2 MULT_mult_6_U3579 ( .A(MULT_mult_6_n1244), .B(
        MULT_mult_6_SUMB_1__26_), .ZN(MULT_mult_6_SUMB_2__25_) );
  XNOR2_X2 MULT_mult_6_U3578 ( .A(MULT_mult_6_SUMB_11__5_), .B(
        MULT_mult_6_n1243), .ZN(MULT_mult_6_SUMB_12__4_) );
  XNOR2_X2 MULT_mult_6_U3577 ( .A(MULT_mult_6_CARRYB_16__11_), .B(
        MULT_mult_6_ab_17__11_), .ZN(MULT_mult_6_n1239) );
  XNOR2_X2 MULT_mult_6_U3576 ( .A(MULT_mult_6_SUMB_16__12_), .B(
        MULT_mult_6_n1239), .ZN(MULT_mult_6_SUMB_17__11_) );
  XNOR2_X2 MULT_mult_6_U3575 ( .A(MULT_mult_6_n1371), .B(MULT_mult_6_net88800), 
        .ZN(MULT_mult_6_net89876) );
  XNOR2_X2 MULT_mult_6_U3574 ( .A(MULT_mult_6_ab_4__1_), .B(
        MULT_mult_6_CARRYB_3__1_), .ZN(MULT_mult_6_n1238) );
  XNOR2_X2 MULT_mult_6_U3573 ( .A(MULT_mult_6_n1238), .B(
        MULT_mult_6_SUMB_3__2_), .ZN(MULT_mult_6_SUMB_4__1_) );
  XOR2_X2 MULT_mult_6_U3572 ( .A(MULT_mult_6_SUMB_9__20_), .B(
        MULT_mult_6_n2215), .Z(MULT_mult_6_SUMB_10__19_) );
  NAND2_X2 MULT_mult_6_U3571 ( .A1(MULT_mult_6_n1121), .A2(MULT_mult_6_n2149), 
        .ZN(MULT_mult_6_n1301) );
  NAND3_X2 MULT_mult_6_U3570 ( .A1(MULT_mult_6_n2102), .A2(MULT_mult_6_n2101), 
        .A3(MULT_mult_6_n2100), .ZN(MULT_mult_6_n1237) );
  XNOR2_X2 MULT_mult_6_U3569 ( .A(MULT_mult_6_CARRYB_22__6_), .B(
        MULT_mult_6_n1234), .ZN(MULT_mult_6_n2282) );
  NAND2_X2 MULT_mult_6_U3568 ( .A1(MULT_mult_6_n1627), .A2(MULT_mult_6_n1628), 
        .ZN(MULT_mult_6_n1630) );
  NAND2_X2 MULT_mult_6_U3567 ( .A1(MULT_mult_6_ab_7__6_), .A2(
        MULT_mult_6_SUMB_6__7_), .ZN(MULT_mult_6_n1334) );
  XNOR2_X2 MULT_mult_6_U3566 ( .A(MULT_mult_6_CARRYB_20__2_), .B(
        MULT_mult_6_ab_21__2_), .ZN(MULT_mult_6_n2171) );
  XNOR2_X2 MULT_mult_6_U3565 ( .A(MULT_mult_6_n1232), .B(MULT_mult_6_n20), 
        .ZN(MULT_mult_6_SUMB_20__2_) );
  FA_X1 MULT_mult_6_U3564 ( .A(MULT_mult_6_ab_5__24_), .B(
        MULT_mult_6_CARRYB_4__24_), .CI(MULT_mult_6_n844), .S(
        MULT_mult_6_n1231) );
  NAND2_X2 MULT_mult_6_U3563 ( .A1(MULT_mult_6_net91088), .A2(
        MULT_mult_6_CARRYB_11__9_), .ZN(MULT_mult_6_net88295) );
  XNOR2_X2 MULT_mult_6_U3562 ( .A(MULT_mult_6_n1227), .B(MULT_mult_6_n367), 
        .ZN(MULT_mult_6_SUMB_10__14_) );
  XNOR2_X2 MULT_mult_6_U3561 ( .A(MULT_mult_6_ab_11__14_), .B(
        MULT_mult_6_CARRYB_10__14_), .ZN(MULT_mult_6_n1226) );
  XNOR2_X2 MULT_mult_6_U3560 ( .A(MULT_mult_6_CARRYB_11__17_), .B(
        MULT_mult_6_ab_12__17_), .ZN(MULT_mult_6_n1223) );
  XNOR2_X2 MULT_mult_6_U3559 ( .A(MULT_mult_6_n1223), .B(
        MULT_mult_6_SUMB_11__18_), .ZN(MULT_mult_6_SUMB_12__17_) );
  XNOR2_X2 MULT_mult_6_U3558 ( .A(MULT_mult_6_n1993), .B(MULT_mult_6_n1253), 
        .ZN(MULT_mult_6_n1222) );
  NAND3_X2 MULT_mult_6_U3557 ( .A1(MULT_mult_6_n1437), .A2(MULT_mult_6_n1436), 
        .A3(MULT_mult_6_n1438), .ZN(MULT_mult_6_net90347) );
  XNOR2_X2 MULT_mult_6_U3556 ( .A(MULT_mult_6_n1221), .B(
        MULT_mult_6_SUMB_10__14_), .ZN(MULT_mult_6_SUMB_11__13_) );
  INV_X2 MULT_mult_6_U3555 ( .A(MULT_mult_6_SUMB_2__26_), .ZN(
        MULT_mult_6_n1218) );
  NAND2_X2 MULT_mult_6_U3554 ( .A1(MULT_mult_6_n1943), .A2(
        MULT_mult_6_SUMB_18__8_), .ZN(MULT_mult_6_n1510) );
  XNOR2_X2 MULT_mult_6_U3553 ( .A(MULT_mult_6_CARRYB_9__15_), .B(
        MULT_mult_6_n1624), .ZN(MULT_mult_6_n1216) );
  XNOR2_X2 MULT_mult_6_U3552 ( .A(MULT_mult_6_n1216), .B(MULT_mult_6_n1220), 
        .ZN(MULT_mult_6_SUMB_10__15_) );
  XNOR2_X2 MULT_mult_6_U3551 ( .A(MULT_mult_6_ab_12__16_), .B(
        MULT_mult_6_CARRYB_11__16_), .ZN(MULT_mult_6_n1215) );
  XNOR2_X2 MULT_mult_6_U3550 ( .A(MULT_mult_6_n1215), .B(
        MULT_mult_6_SUMB_11__17_), .ZN(MULT_mult_6_SUMB_12__16_) );
  INV_X4 MULT_mult_6_U3547 ( .A(MULT_mult_6_CARRYB_4__13_), .ZN(
        MULT_mult_6_n1541) );
  CLKBUF_X2 MULT_mult_6_U3546 ( .A(MULT_mult_6_SUMB_6__24_), .Z(
        MULT_mult_6_n1213) );
  XNOR2_X2 MULT_mult_6_U3545 ( .A(MULT_mult_6_CARRYB_5__18_), .B(
        MULT_mult_6_ab_6__18_), .ZN(MULT_mult_6_n1212) );
  XNOR2_X2 MULT_mult_6_U3544 ( .A(MULT_mult_6_SUMB_5__19_), .B(
        MULT_mult_6_n1212), .ZN(MULT_mult_6_net90702) );
  NAND2_X2 MULT_mult_6_U3543 ( .A1(MULT_mult_6_n943), .A2(MULT_mult_6_ab_5__9_), .ZN(MULT_mult_6_n1396) );
  CLKBUF_X3 MULT_mult_6_U3542 ( .A(MULT_mult_6_SUMB_13__5_), .Z(
        MULT_mult_6_n1253) );
  NAND3_X2 MULT_mult_6_U3541 ( .A1(MULT_mult_6_n2150), .A2(MULT_mult_6_n2151), 
        .A3(MULT_mult_6_n2152), .ZN(MULT_mult_6_n1211) );
  CLKBUF_X3 MULT_mult_6_U3540 ( .A(MULT_mult_6_SUMB_15__6_), .Z(
        MULT_mult_6_n1236) );
  XNOR2_X2 MULT_mult_6_U3539 ( .A(MULT_mult_6_n1210), .B(
        MULT_mult_6_SUMB_4__21_), .ZN(MULT_mult_6_SUMB_5__20_) );
  NAND3_X2 MULT_mult_6_U3538 ( .A1(MULT_mult_6_n1409), .A2(MULT_mult_6_n1410), 
        .A3(MULT_mult_6_n1411), .ZN(MULT_mult_6_CARRYB_15__0_) );
  NOR2_X2 MULT_mult_6_U3535 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__13_) );
  INV_X2 MULT_mult_6_U3534 ( .A(MULT_mult_6_n1767), .ZN(MULT_mult_6_n1768) );
  NAND3_X2 MULT_mult_6_U3533 ( .A1(MULT_mult_6_net81365), .A2(
        MULT_mult_6_net81367), .A3(MULT_mult_6_n2035), .ZN(
        MULT_mult_6_CARRYB_7__14_) );
  NAND3_X2 MULT_mult_6_U3532 ( .A1(MULT_mult_6_n1958), .A2(MULT_mult_6_n1959), 
        .A3(MULT_mult_6_n1960), .ZN(MULT_mult_6_CARRYB_5__23_) );
  XNOR2_X2 MULT_mult_6_U3531 ( .A(MULT_mult_6_n1204), .B(
        MULT_mult_6_SUMB_19__11_), .ZN(MULT_mult_6_SUMB_20__10_) );
  NAND3_X2 MULT_mult_6_U3530 ( .A1(MULT_mult_6_n1652), .A2(MULT_mult_6_n1653), 
        .A3(MULT_mult_6_n1654), .ZN(MULT_mult_6_n1203) );
  NAND2_X4 MULT_mult_6_U3529 ( .A1(MULT_mult_6_n1617), .A2(
        MULT_mult_6_net91243), .ZN(MULT_mult_6_n1522) );
  NAND3_X2 MULT_mult_6_U3528 ( .A1(MULT_mult_6_n2071), .A2(MULT_mult_6_n2072), 
        .A3(MULT_mult_6_n2073), .ZN(MULT_mult_6_n1201) );
  XNOR2_X2 MULT_mult_6_U3527 ( .A(MULT_mult_6_n1200), .B(MULT_mult_6_n842), 
        .ZN(MULT_mult_6_SUMB_11__3_) );
  NAND2_X4 MULT_mult_6_U3526 ( .A1(MULT_mult_6_net85373), .A2(
        MULT_mult_6_net85732), .ZN(MULT_mult_6_n1523) );
  NAND2_X4 MULT_mult_6_U3525 ( .A1(MULT_mult_6_CARRYB_18__5_), .A2(
        MULT_mult_6_ab_19__5_), .ZN(MULT_mult_6_net84708) );
  XNOR2_X2 MULT_mult_6_U3524 ( .A(MULT_mult_6_n1198), .B(
        MULT_mult_6_SUMB_8__7_), .ZN(MULT_mult_6_SUMB_9__6_) );
  INV_X4 MULT_mult_6_U3523 ( .A(MULT_mult_6_SUMB_2__27_), .ZN(
        MULT_mult_6_n1196) );
  NAND3_X2 MULT_mult_6_U3522 ( .A1(MULT_mult_6_n2198), .A2(MULT_mult_6_n2199), 
        .A3(MULT_mult_6_n2200), .ZN(MULT_mult_6_CARRYB_15__12_) );
  NAND2_X1 MULT_mult_6_U3521 ( .A1(MULT_mult_6_CARRYB_14__12_), .A2(
        MULT_mult_6_SUMB_14__13_), .ZN(MULT_mult_6_n2198) );
  NAND2_X4 MULT_mult_6_U3519 ( .A1(MULT_mult_6_net87310), .A2(
        MULT_mult_6_n1367), .ZN(MULT_mult_6_net85212) );
  XNOR2_X2 MULT_mult_6_U3518 ( .A(MULT_mult_6_n1585), .B(MULT_mult_6_n1236), 
        .ZN(MULT_mult_6_n1195) );
  INV_X2 MULT_mult_6_U3517 ( .A(MULT_mult_6_n1298), .ZN(MULT_mult_6_n1194) );
  INV_X4 MULT_mult_6_U3516 ( .A(MULT_mult_6_n1192), .ZN(MULT_mult_6_n1193) );
  XNOR2_X2 MULT_mult_6_U3515 ( .A(MULT_mult_6_CARRYB_10__13_), .B(
        MULT_mult_6_ab_11__13_), .ZN(MULT_mult_6_n1221) );
  NAND3_X2 MULT_mult_6_U3514 ( .A1(MULT_mult_6_n2279), .A2(MULT_mult_6_n2280), 
        .A3(MULT_mult_6_n2281), .ZN(MULT_mult_6_CARRYB_6__19_) );
  CLKBUF_X3 MULT_mult_6_U3513 ( .A(MULT_mult_6_SUMB_16__6_), .Z(
        MULT_mult_6_n1270) );
  INV_X4 MULT_mult_6_U3512 ( .A(MULT_mult_6_n1188), .ZN(MULT_mult_6_SUMB_7__7_) );
  XNOR2_X2 MULT_mult_6_U3511 ( .A(MULT_mult_6_n1821), .B(
        MULT_mult_6_SUMB_6__8_), .ZN(MULT_mult_6_n1188) );
  XNOR2_X2 MULT_mult_6_U3510 ( .A(MULT_mult_6_n2065), .B(
        MULT_mult_6_SUMB_14__13_), .ZN(MULT_mult_6_n1187) );
  NAND2_X4 MULT_mult_6_U3509 ( .A1(MULT_mult_6_ab_3__20_), .A2(
        MULT_mult_6_CARRYB_2__20_), .ZN(MULT_mult_6_n2192) );
  NAND2_X4 MULT_mult_6_U3508 ( .A1(MULT_mult_6_ab_15__4_), .A2(
        MULT_mult_6_n1211), .ZN(MULT_mult_6_n1705) );
  XNOR2_X2 MULT_mult_6_U3507 ( .A(MULT_mult_6_n1184), .B(MULT_mult_6_net92341), 
        .ZN(MULT_mult_6_n1183) );
  XNOR2_X2 MULT_mult_6_U3506 ( .A(MULT_mult_6_n1182), .B(MULT_mult_6_n1183), 
        .ZN(MULT_mult_6_net92322) );
  NAND2_X4 MULT_mult_6_U3505 ( .A1(MULT_mult_6_n176), .A2(
        MULT_mult_6_ab_17__4_), .ZN(MULT_mult_6_n2074) );
  NAND3_X4 MULT_mult_6_U3504 ( .A1(MULT_mult_6_n1302), .A2(MULT_mult_6_n1303), 
        .A3(MULT_mult_6_n1304), .ZN(MULT_mult_6_CARRYB_10__14_) );
  NAND3_X2 MULT_mult_6_U3503 ( .A1(MULT_mult_6_n1796), .A2(MULT_mult_6_n1797), 
        .A3(MULT_mult_6_n1798), .ZN(MULT_mult_6_CARRYB_22__0_) );
  NAND3_X1 MULT_mult_6_U3502 ( .A1(MULT_mult_6_n2011), .A2(MULT_mult_6_n2376), 
        .A3(MULT_mult_6_n2012), .ZN(MULT_mult_6_net91001) );
  NAND3_X4 MULT_mult_6_U3501 ( .A1(MULT_mult_6_net84116), .A2(
        MULT_mult_6_n1648), .A3(MULT_mult_6_net84118), .ZN(
        MULT_mult_6_CARRYB_3__7_) );
  XNOR2_X2 MULT_mult_6_U3500 ( .A(MULT_mult_6_net92378), .B(MULT_mult_6_n284), 
        .ZN(multOut[3]) );
  NAND2_X4 MULT_mult_6_U3499 ( .A1(MULT_mult_6_n1544), .A2(
        MULT_mult_6_net85254), .ZN(MULT_mult_6_n1679) );
  NAND3_X4 MULT_mult_6_U3498 ( .A1(MULT_mult_6_net80920), .A2(
        MULT_mult_6_net80922), .A3(MULT_mult_6_net80921), .ZN(
        MULT_mult_6_CARRYB_24__1_) );
  NOR2_X1 MULT_mult_6_U3497 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net77966), .ZN(MULT_mult_6_ab_3__9_) );
  NAND2_X2 MULT_mult_6_U3496 ( .A1(MULT_mult_6_SUMB_22__1_), .A2(
        MULT_mult_6_ab_23__0_), .ZN(MULT_mult_6_n1799) );
  CLKBUF_X3 MULT_mult_6_U3495 ( .A(MULT_mult_6_SUMB_4__9_), .Z(
        MULT_mult_6_n1217) );
  NAND2_X2 MULT_mult_6_U3494 ( .A1(MULT_mult_6_SUMB_4__9_), .A2(
        MULT_mult_6_CARRYB_4__8_), .ZN(MULT_mult_6_n1966) );
  NAND3_X2 MULT_mult_6_U3493 ( .A1(MULT_mult_6_n1670), .A2(MULT_mult_6_n1671), 
        .A3(MULT_mult_6_n1672), .ZN(MULT_mult_6_CARRYB_11__3_) );
  NAND2_X4 MULT_mult_6_U3492 ( .A1(MULT_mult_6_ab_24__2_), .A2(
        MULT_mult_6_CARRYB_23__2_), .ZN(MULT_mult_6_net80258) );
  NAND2_X2 MULT_mult_6_U3491 ( .A1(MULT_mult_6_CARRYB_6__6_), .A2(
        MULT_mult_6_ab_7__6_), .ZN(MULT_mult_6_n1333) );
  NAND2_X4 MULT_mult_6_U3490 ( .A1(MULT_mult_6_n1201), .A2(
        MULT_mult_6_ab_17__5_), .ZN(MULT_mult_6_n1382) );
  NAND2_X2 MULT_mult_6_U3489 ( .A1(MULT_mult_6_ab_12__3_), .A2(
        MULT_mult_6_CARRYB_11__3_), .ZN(MULT_mult_6_n1674) );
  INV_X4 MULT_mult_6_U3488 ( .A(MULT_mult_6_SUMB_15__9_), .ZN(
        MULT_mult_6_n1449) );
  NAND2_X4 MULT_mult_6_U3487 ( .A1(MULT_mult_6_n1275), .A2(
        MULT_mult_6_ab_12__5_), .ZN(MULT_mult_6_n1637) );
  NAND2_X4 MULT_mult_6_U3486 ( .A1(MULT_mult_6_SUMB_16__5_), .A2(
        MULT_mult_6_ab_17__4_), .ZN(MULT_mult_6_n2075) );
  NAND2_X4 MULT_mult_6_U3485 ( .A1(MULT_mult_6_n1195), .A2(MULT_mult_6_n176), 
        .ZN(MULT_mult_6_n2076) );
  NAND3_X1 MULT_mult_6_U3484 ( .A1(MULT_mult_6_net80355), .A2(
        MULT_mult_6_net80356), .A3(MULT_mult_6_n2272), .ZN(MULT_mult_6_n1235)
         );
  NAND2_X4 MULT_mult_6_U3483 ( .A1(MULT_mult_6_n1373), .A2(MULT_mult_6_n1374), 
        .ZN(MULT_mult_6_n1730) );
  INV_X4 MULT_mult_6_U3482 ( .A(MULT_mult_6_net88702), .ZN(
        MULT_mult_6_net85469) );
  NAND2_X2 MULT_mult_6_U3481 ( .A1(MULT_mult_6_CARRYB_6__13_), .A2(
        MULT_mult_6_ab_7__13_), .ZN(MULT_mult_6_n1320) );
  INV_X1 MULT_mult_6_U3480 ( .A(MULT_mult_6_ab_9__8_), .ZN(MULT_mult_6_n1178)
         );
  NAND2_X2 MULT_mult_6_U3479 ( .A1(MULT_mult_6_CARRYB_8__8_), .A2(
        MULT_mult_6_ab_9__8_), .ZN(MULT_mult_6_n1179) );
  INV_X4 MULT_mult_6_U3478 ( .A(MULT_mult_6_n2243), .ZN(MULT_mult_6_n1755) );
  XNOR2_X2 MULT_mult_6_U3477 ( .A(MULT_mult_6_n1176), .B(MULT_mult_6_n946), 
        .ZN(MULT_mult_6_SUMB_9__7_) );
  NAND2_X4 MULT_mult_6_U3476 ( .A1(MULT_mult_6_SUMB_7__12_), .A2(
        MULT_mult_6_ab_8__11_), .ZN(MULT_mult_6_n2127) );
  NAND2_X4 MULT_mult_6_U3475 ( .A1(MULT_mult_6_n1345), .A2(
        MULT_mult_6_ab_14__12_), .ZN(MULT_mult_6_n1488) );
  INV_X2 MULT_mult_6_U3474 ( .A(MULT_mult_6_ab_9__9_), .ZN(MULT_mult_6_n1563)
         );
  INV_X4 MULT_mult_6_U3473 ( .A(MULT_mult_6_n1563), .ZN(MULT_mult_6_n1173) );
  NAND2_X4 MULT_mult_6_U3472 ( .A1(MULT_mult_6_n1172), .A2(MULT_mult_6_n1173), 
        .ZN(MULT_mult_6_n1175) );
  NAND2_X2 MULT_mult_6_U3471 ( .A1(MULT_mult_6_n1563), .A2(
        MULT_mult_6_CARRYB_8__9_), .ZN(MULT_mult_6_n1174) );
  NAND3_X4 MULT_mult_6_U3470 ( .A1(MULT_mult_6_n2080), .A2(MULT_mult_6_n2081), 
        .A3(MULT_mult_6_n2082), .ZN(MULT_mult_6_n1207) );
  INV_X1 MULT_mult_6_U3469 ( .A(MULT_mult_6_CARRYB_5__10_), .ZN(
        MULT_mult_6_n1169) );
  INV_X4 MULT_mult_6_U3468 ( .A(MULT_mult_6_n1694), .ZN(MULT_mult_6_n1168) );
  NAND2_X4 MULT_mult_6_U3467 ( .A1(MULT_mult_6_n1170), .A2(MULT_mult_6_n1171), 
        .ZN(MULT_mult_6_SUMB_6__10_) );
  INV_X4 MULT_mult_6_U3466 ( .A(MULT_mult_6_n1260), .ZN(MULT_mult_6_n1165) );
  INV_X4 MULT_mult_6_U3465 ( .A(MULT_mult_6_n1837), .ZN(MULT_mult_6_n1164) );
  NAND2_X4 MULT_mult_6_U3464 ( .A1(MULT_mult_6_n1166), .A2(MULT_mult_6_n1167), 
        .ZN(MULT_mult_6_SUMB_13__5_) );
  NAND2_X4 MULT_mult_6_U3463 ( .A1(MULT_mult_6_n1164), .A2(MULT_mult_6_n1165), 
        .ZN(MULT_mult_6_n1167) );
  NAND2_X2 MULT_mult_6_U3462 ( .A1(MULT_mult_6_n1837), .A2(MULT_mult_6_n1260), 
        .ZN(MULT_mult_6_n1166) );
  NOR2_X1 MULT_mult_6_U3461 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net70457), .ZN(MULT_mult_6_ab_19__9_) );
  NOR2_X1 MULT_mult_6_U3460 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net70453), .ZN(MULT_mult_6_ab_21__9_) );
  OR2_X1 MULT_mult_6_U3459 ( .A1(MULT_mult_6_net70451), .A2(
        MULT_mult_6_net70452), .ZN(MULT_mult_6_n1929) );
  NAND2_X4 MULT_mult_6_U3458 ( .A1(MULT_mult_6_net85455), .A2(
        MULT_mult_6_net85456), .ZN(MULT_mult_6_n1505) );
  INV_X4 MULT_mult_6_U3457 ( .A(MULT_mult_6_n1361), .ZN(MULT_mult_6_n1351) );
  NAND2_X2 MULT_mult_6_U3456 ( .A1(MULT_mult_6_n1361), .A2(
        MULT_mult_6_SUMB_1__16_), .ZN(MULT_mult_6_n1353) );
  NOR2_X4 MULT_mult_6_U3455 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net77940), .ZN(MULT_mult_6_ab_6__13_) );
  NAND3_X4 MULT_mult_6_U3454 ( .A1(MULT_mult_6_n1988), .A2(MULT_mult_6_n1987), 
        .A3(MULT_mult_6_n1989), .ZN(MULT_mult_6_CARRYB_3__14_) );
  NOR2_X2 MULT_mult_6_U3453 ( .A1(MULT_mult_6_net84698), .A2(
        MULT_mult_6_net119855), .ZN(MULT_mult_6_ab_4__14_) );
  INV_X2 MULT_mult_6_U3452 ( .A(MULT_mult_6_ab_2__15_), .ZN(
        MULT_mult_6_net92724) );
  NAND2_X4 MULT_mult_6_U3451 ( .A1(MULT_mult_6_n1984), .A2(MULT_mult_6_n1163), 
        .ZN(MULT_mult_6_n1361) );
  INV_X1 MULT_mult_6_U3450 ( .A(MULT_mult_6_ab_6__13_), .ZN(MULT_mult_6_n1159)
         );
  INV_X4 MULT_mult_6_U3449 ( .A(MULT_mult_6_CARRYB_3__14_), .ZN(
        MULT_mult_6_net92717) );
  NAND2_X4 MULT_mult_6_U3448 ( .A1(MULT_mult_6_n1158), .A2(
        MULT_mult_6_net92718), .ZN(MULT_mult_6_n1720) );
  NAND2_X4 MULT_mult_6_U3447 ( .A1(MULT_mult_6_net92716), .A2(
        MULT_mult_6_net92717), .ZN(MULT_mult_6_n1158) );
  INV_X8 MULT_mult_6_U3446 ( .A(MULT_mult_6_n2335), .ZN(
        MULT_mult_6_SUMB_1__11_) );
  INV_X4 MULT_mult_6_U3445 ( .A(MULT_mult_6_ab_2__10_), .ZN(MULT_mult_6_n1154)
         );
  NAND2_X2 MULT_mult_6_U3444 ( .A1(MULT_mult_6_ab_2__10_), .A2(
        MULT_mult_6_n2332), .ZN(MULT_mult_6_n1155) );
  NAND2_X2 MULT_mult_6_U3443 ( .A1(MULT_mult_6_CARRYB_6__6_), .A2(
        MULT_mult_6_SUMB_6__7_), .ZN(MULT_mult_6_n1335) );
  XNOR2_X1 MULT_mult_6_U3442 ( .A(MULT_mult_6_CARRYB_2__11_), .B(
        MULT_mult_6_ab_3__11_), .ZN(MULT_mult_6_n1869) );
  XNOR2_X2 MULT_mult_6_U3441 ( .A(MULT_mult_6_ab_20__10_), .B(
        MULT_mult_6_CARRYB_19__10_), .ZN(MULT_mult_6_n1204) );
  NAND2_X2 MULT_mult_6_U3440 ( .A1(MULT_mult_6_ab_9__6_), .A2(
        MULT_mult_6_CARRYB_8__6_), .ZN(MULT_mult_6_n1294) );
  INV_X4 MULT_mult_6_U3439 ( .A(MULT_mult_6_n1721), .ZN(MULT_mult_6_n1150) );
  NAND2_X4 MULT_mult_6_U3438 ( .A1(MULT_mult_6_n1153), .A2(MULT_mult_6_n1152), 
        .ZN(MULT_mult_6_SUMB_15__5_) );
  NAND2_X4 MULT_mult_6_U3437 ( .A1(MULT_mult_6_n1150), .A2(MULT_mult_6_n1151), 
        .ZN(MULT_mult_6_n1153) );
  NAND3_X4 MULT_mult_6_U3436 ( .A1(MULT_mult_6_n2229), .A2(MULT_mult_6_n2230), 
        .A3(MULT_mult_6_n2228), .ZN(MULT_mult_6_CARRYB_20__4_) );
  NAND2_X2 MULT_mult_6_U3435 ( .A1(MULT_mult_6_CARRYB_9__1_), .A2(
        MULT_mult_6_ab_10__1_), .ZN(MULT_mult_6_n1471) );
  NAND2_X2 MULT_mult_6_U3434 ( .A1(MULT_mult_6_n1783), .A2(MULT_mult_6_n1784), 
        .ZN(MULT_mult_6_n2060) );
  NAND2_X1 MULT_mult_6_U3433 ( .A1(MULT_mult_6_ab_5__20_), .A2(
        MULT_mult_6_CARRYB_4__20_), .ZN(MULT_mult_6_n1885) );
  NAND3_X4 MULT_mult_6_U3432 ( .A1(MULT_mult_6_n1620), .A2(MULT_mult_6_n1619), 
        .A3(MULT_mult_6_n1621), .ZN(MULT_mult_6_CARRYB_9__9_) );
  NAND2_X2 MULT_mult_6_U3431 ( .A1(MULT_mult_6_n2244), .A2(
        MULT_mult_6_net148233), .ZN(MULT_mult_6_n1364) );
  NOR2_X1 MULT_mult_6_U3430 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net77966), .ZN(MULT_mult_6_ab_3__4_) );
  NOR2_X2 MULT_mult_6_U3429 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net77970), .ZN(MULT_mult_6_ab_2__4_) );
  NAND3_X2 MULT_mult_6_U3428 ( .A1(MULT_mult_6_n1147), .A2(MULT_mult_6_n1148), 
        .A3(MULT_mult_6_n1149), .ZN(MULT_mult_6_CARRYB_3__4_) );
  NAND2_X1 MULT_mult_6_U3427 ( .A1(MULT_mult_6_ab_3__4_), .A2(
        MULT_mult_6_CARRYB_2__4_), .ZN(MULT_mult_6_n1149) );
  NAND2_X2 MULT_mult_6_U3426 ( .A1(MULT_mult_6_ab_3__4_), .A2(
        MULT_mult_6_SUMB_2__5_), .ZN(MULT_mult_6_n1148) );
  NAND3_X2 MULT_mult_6_U3425 ( .A1(MULT_mult_6_n1144), .A2(MULT_mult_6_n1145), 
        .A3(MULT_mult_6_n1146), .ZN(MULT_mult_6_CARRYB_12__0_) );
  NAND2_X2 MULT_mult_6_U3424 ( .A1(MULT_mult_6_ab_12__0_), .A2(
        MULT_mult_6_CARRYB_11__0_), .ZN(MULT_mult_6_n1145) );
  XOR2_X2 MULT_mult_6_U3423 ( .A(MULT_mult_6_n1143), .B(
        MULT_mult_6_CARRYB_11__0_), .Z(multOut[19]) );
  XOR2_X1 MULT_mult_6_U3422 ( .A(MULT_mult_6_ab_12__0_), .B(
        MULT_mult_6_SUMB_11__1_), .Z(MULT_mult_6_n1143) );
  NAND3_X2 MULT_mult_6_U3421 ( .A1(MULT_mult_6_n1140), .A2(MULT_mult_6_n1141), 
        .A3(MULT_mult_6_n1142), .ZN(MULT_mult_6_CARRYB_11__0_) );
  NAND3_X2 MULT_mult_6_U3420 ( .A1(MULT_mult_6_n1136), .A2(MULT_mult_6_n1137), 
        .A3(MULT_mult_6_n1138), .ZN(MULT_mult_6_CARRYB_2__4_) );
  NAND2_X1 MULT_mult_6_U3419 ( .A1(MULT_mult_6_ab_2__4_), .A2(
        MULT_mult_6_CARRYB_1__4_), .ZN(MULT_mult_6_n1138) );
  NAND2_X2 MULT_mult_6_U3418 ( .A1(MULT_mult_6_ab_2__4_), .A2(
        MULT_mult_6_SUMB_1__5_), .ZN(MULT_mult_6_n1137) );
  NAND2_X1 MULT_mult_6_U3417 ( .A1(MULT_mult_6_CARRYB_1__4_), .A2(
        MULT_mult_6_SUMB_1__5_), .ZN(MULT_mult_6_n1136) );
  XOR2_X2 MULT_mult_6_U3416 ( .A(MULT_mult_6_SUMB_1__5_), .B(MULT_mult_6_n1135), .Z(MULT_mult_6_SUMB_2__4_) );
  NOR2_X1 MULT_mult_6_U3415 ( .A1(MULT_mult_6_net70482), .A2(
        MULT_mult_6_net77966), .ZN(MULT_mult_6_ab_3__24_) );
  NAND2_X4 MULT_mult_6_U3414 ( .A1(MULT_mult_6_CARRYB_19__6_), .A2(
        MULT_mult_6_n1190), .ZN(MULT_mult_6_n2211) );
  NAND2_X4 MULT_mult_6_U3413 ( .A1(MULT_mult_6_net88166), .A2(
        MULT_mult_6_n1317), .ZN(MULT_mult_6_n1319) );
  NAND2_X2 MULT_mult_6_U3412 ( .A1(MULT_mult_6_CARRYB_10__3_), .A2(
        MULT_mult_6_SUMB_10__4_), .ZN(MULT_mult_6_n1672) );
  NAND2_X2 MULT_mult_6_U3411 ( .A1(MULT_mult_6_CARRYB_8__6_), .A2(
        MULT_mult_6_SUMB_8__7_), .ZN(MULT_mult_6_n1292) );
  NAND2_X4 MULT_mult_6_U3410 ( .A1(MULT_mult_6_n1523), .A2(MULT_mult_6_n1522), 
        .ZN(MULT_mult_6_net91088) );
  INV_X8 MULT_mult_6_U3409 ( .A(n10909), .ZN(MULT_mult_6_n2355) );
  NOR2_X1 MULT_mult_6_U3408 ( .A1(MULT_mult_6_net70486), .A2(
        MULT_mult_6_net77956), .ZN(MULT_mult_6_ab_4__26_) );
  XNOR2_X2 MULT_mult_6_U3407 ( .A(MULT_mult_6_n558), .B(MULT_mult_6_n1869), 
        .ZN(MULT_mult_6_n1229) );
  XNOR2_X2 MULT_mult_6_U3406 ( .A(MULT_mult_6_CARRYB_18__3_), .B(
        MULT_mult_6_ab_19__3_), .ZN(MULT_mult_6_n2110) );
  XNOR2_X2 MULT_mult_6_U3405 ( .A(MULT_mult_6_CARRYB_15__15_), .B(
        MULT_mult_6_ab_16__15_), .ZN(MULT_mult_6_n1133) );
  XNOR2_X2 MULT_mult_6_U3404 ( .A(MULT_mult_6_n2066), .B(
        MULT_mult_6_SUMB_14__17_), .ZN(MULT_mult_6_n1132) );
  XNOR2_X2 MULT_mult_6_U3403 ( .A(MULT_mult_6_n1132), .B(MULT_mult_6_n1133), 
        .ZN(MULT_mult_6_n1312) );
  NAND3_X4 MULT_mult_6_U3402 ( .A1(MULT_mult_6_n1990), .A2(MULT_mult_6_n1991), 
        .A3(MULT_mult_6_n1992), .ZN(MULT_mult_6_CARRYB_15__3_) );
  NAND2_X2 MULT_mult_6_U3401 ( .A1(MULT_mult_6_ab_16__3_), .A2(
        MULT_mult_6_SUMB_15__4_), .ZN(MULT_mult_6_n1130) );
  NAND2_X2 MULT_mult_6_U3400 ( .A1(MULT_mult_6_n1732), .A2(MULT_mult_6_n1588), 
        .ZN(MULT_mult_6_n1446) );
  NAND2_X2 MULT_mult_6_U3399 ( .A1(MULT_mult_6_CARRYB_1__18_), .A2(
        MULT_mult_6_ab_2__18_), .ZN(MULT_mult_6_n1711) );
  NAND2_X2 MULT_mult_6_U3398 ( .A1(MULT_mult_6_SUMB_9__4_), .A2(
        MULT_mult_6_CARRYB_9__3_), .ZN(MULT_mult_6_n1804) );
  NAND3_X4 MULT_mult_6_U3397 ( .A1(MULT_mult_6_n1813), .A2(MULT_mult_6_n1814), 
        .A3(MULT_mult_6_n1815), .ZN(MULT_mult_6_CARRYB_19__0_) );
  NAND2_X4 MULT_mult_6_U3394 ( .A1(MULT_mult_6_n1500), .A2(
        MULT_mult_6_SUMB_15__5_), .ZN(MULT_mult_6_n2103) );
  NAND2_X2 MULT_mult_6_U3393 ( .A1(MULT_mult_6_n1193), .A2(
        MULT_mult_6_SUMB_11__7_), .ZN(MULT_mult_6_n1919) );
  NAND2_X4 MULT_mult_6_U3392 ( .A1(MULT_mult_6_n288), .A2(MULT_mult_6_n1157), 
        .ZN(MULT_mult_6_n2057) );
  XNOR2_X2 MULT_mult_6_U3391 ( .A(MULT_mult_6_n1539), .B(
        MULT_mult_6_SUMB_3__26_), .ZN(MULT_mult_6_n1185) );
  NAND3_X2 MULT_mult_6_U3390 ( .A1(MULT_mult_6_n2307), .A2(MULT_mult_6_n2308), 
        .A3(MULT_mult_6_n2309), .ZN(MULT_mult_6_CARRYB_12__16_) );
  NAND2_X4 MULT_mult_6_U3389 ( .A1(MULT_mult_6_SUMB_15__5_), .A2(
        MULT_mult_6_ab_16__4_), .ZN(MULT_mult_6_n2104) );
  INV_X4 MULT_mult_6_U3388 ( .A(MULT_mult_6_net82548), .ZN(
        MULT_mult_6_net93308) );
  NAND2_X4 MULT_mult_6_U3387 ( .A1(MULT_mult_6_n1125), .A2(MULT_mult_6_n1124), 
        .ZN(MULT_mult_6_SUMB_12__8_) );
  NAND2_X4 MULT_mult_6_U3385 ( .A1(MULT_mult_6_net86662), .A2(
        MULT_mult_6_n1719), .ZN(MULT_mult_6_n2233) );
  NAND2_X4 MULT_mult_6_U3384 ( .A1(MULT_mult_6_ab_3__7_), .A2(
        MULT_mult_6_net85036), .ZN(MULT_mult_6_n1648) );
  INV_X8 MULT_mult_6_U3383 ( .A(MULT_mult_6_net86661), .ZN(
        MULT_mult_6_net86662) );
  NAND3_X2 MULT_mult_6_U3382 ( .A1(MULT_mult_6_net80817), .A2(
        MULT_mult_6_net80818), .A3(MULT_mult_6_net80816), .ZN(
        MULT_mult_6_n1184) );
  NAND2_X2 MULT_mult_6_U3380 ( .A1(MULT_mult_6_n596), .A2(
        MULT_mult_6_SUMB_20__3_), .ZN(MULT_mult_6_n2185) );
  NAND2_X1 MULT_mult_6_U3378 ( .A1(MULT_mult_6_ab_18__9_), .A2(
        MULT_mult_6_CARRYB_17__9_), .ZN(MULT_mult_6_n2154) );
  NAND2_X2 MULT_mult_6_U3377 ( .A1(MULT_mult_6_SUMB_7__10_), .A2(
        MULT_mult_6_ab_8__9_), .ZN(MULT_mult_6_n2084) );
  NOR2_X2 MULT_mult_6_U3376 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net77924), .ZN(MULT_mult_6_ab_8__9_) );
  NOR2_X2 MULT_mult_6_U3375 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net77946), .ZN(MULT_mult_6_ab_5__9_) );
  XNOR2_X2 MULT_mult_6_U3374 ( .A(MULT_mult_6_n1122), .B(MULT_mult_6_n1389), 
        .ZN(MULT_mult_6_SUMB_5__7_) );
  XNOR2_X2 MULT_mult_6_U3373 ( .A(MULT_mult_6_CARRYB_15__8_), .B(
        MULT_mult_6_n2153), .ZN(MULT_mult_6_n1279) );
  XNOR2_X2 MULT_mult_6_U3372 ( .A(MULT_mult_6_net93713), .B(
        MULT_mult_6_net83358), .ZN(MULT_mult_6_SUMB_23__1_) );
  INV_X1 MULT_mult_6_U3371 ( .A(MULT_mult_6_net83850), .ZN(
        MULT_mult_6_net93747) );
  NAND2_X2 MULT_mult_6_U3370 ( .A1(MULT_mult_6_SUMB_6__16_), .A2(
        MULT_mult_6_n676), .ZN(MULT_mult_6_n2210) );
  XNOR2_X2 MULT_mult_6_U3369 ( .A(MULT_mult_6_net124618), .B(
        MULT_mult_6_SUMB_1__14_), .ZN(MULT_mult_6_n1120) );
  INV_X8 MULT_mult_6_U3368 ( .A(n10915), .ZN(MULT_mult_6_net70474) );
  XNOR2_X2 MULT_mult_6_U3367 ( .A(MULT_mult_6_net93880), .B(
        MULT_mult_6_SUMB_24__2_), .ZN(MULT_mult_6_SUMB_25__1_) );
  NAND2_X1 MULT_mult_6_U3366 ( .A1(MULT_mult_6_SUMB_4__22_), .A2(
        MULT_mult_6_CARRYB_4__21_), .ZN(MULT_mult_6_n1115) );
  NAND3_X2 MULT_mult_6_U3365 ( .A1(MULT_mult_6_n1115), .A2(MULT_mult_6_n1116), 
        .A3(MULT_mult_6_n1117), .ZN(MULT_mult_6_CARRYB_5__21_) );
  NOR2_X1 MULT_mult_6_U3364 ( .A1(MULT_mult_6_net80643), .A2(
        MULT_mult_6_net77940), .ZN(MULT_mult_6_ab_6__21_) );
  INV_X16 MULT_mult_6_U3363 ( .A(n10910), .ZN(MULT_mult_6_net70486) );
  XNOR2_X2 MULT_mult_6_U3362 ( .A(MULT_mult_6_ab_0__26_), .B(
        MULT_mult_6_ab_1__25_), .ZN(MULT_mult_6__UDW__112644_net78437) );
  NAND2_X2 MULT_mult_6_U3361 ( .A1(MULT_mult_6_SUMB_1__25_), .A2(
        MULT_mult_6_n39), .ZN(MULT_mult_6_net84297) );
  XNOR2_X2 MULT_mult_6_U3360 ( .A(MULT_mult_6_SUMB_1__25_), .B(MULT_mult_6_n39), .ZN(MULT_mult_6_net84883) );
  NOR2_X1 MULT_mult_6_U3359 ( .A1(MULT_mult_6_net91660), .A2(
        MULT_mult_6_net70457), .ZN(MULT_mult_6_ab_19__10_) );
  NAND2_X1 MULT_mult_6_U3358 ( .A1(MULT_mult_6_CARRYB_17__10_), .A2(
        MULT_mult_6_ab_18__10_), .ZN(MULT_mult_6_n1112) );
  NAND2_X2 MULT_mult_6_U3357 ( .A1(MULT_mult_6_CARRYB_17__10_), .A2(
        MULT_mult_6_SUMB_17__11_), .ZN(MULT_mult_6_n1113) );
  NAND2_X2 MULT_mult_6_U3356 ( .A1(MULT_mult_6_ab_18__10_), .A2(
        MULT_mult_6_SUMB_17__11_), .ZN(MULT_mult_6_n1114) );
  NAND2_X1 MULT_mult_6_U3355 ( .A1(MULT_mult_6_CARRYB_18__10_), .A2(
        MULT_mult_6_ab_19__10_), .ZN(MULT_mult_6_net82667) );
  NAND3_X4 MULT_mult_6_U3354 ( .A1(MULT_mult_6_n1114), .A2(MULT_mult_6_n1113), 
        .A3(MULT_mult_6_n1112), .ZN(MULT_mult_6_CARRYB_18__10_) );
  NOR2_X2 MULT_mult_6_U3353 ( .A1(MULT_mult_6_n1111), .A2(MULT_mult_6_net80409), .ZN(MULT_mult_6_ab_1__25_) );
  INV_X8 MULT_mult_6_U3352 ( .A(n10911), .ZN(MULT_mult_6_n1111) );
  NAND2_X2 MULT_mult_6_U3351 ( .A1(MULT_mult_6_ab_7__18_), .A2(
        MULT_mult_6_CARRYB_6__18_), .ZN(MULT_mult_6_net80302) );
  NOR2_X1 MULT_mult_6_U3350 ( .A1(MULT_mult_6_n182), .A2(MULT_mult_6_net70477), 
        .ZN(MULT_mult_6_ab_9__18_) );
  NAND2_X2 MULT_mult_6_U3349 ( .A1(MULT_mult_6_SUMB_7__19_), .A2(
        MULT_mult_6_ab_8__18_), .ZN(MULT_mult_6_n1106) );
  NAND2_X1 MULT_mult_6_U3348 ( .A1(MULT_mult_6_SUMB_6__19_), .A2(
        MULT_mult_6_CARRYB_6__18_), .ZN(MULT_mult_6_n1110) );
  NAND3_X2 MULT_mult_6_U3347 ( .A1(MULT_mult_6_n1110), .A2(
        MULT_mult_6_net80303), .A3(MULT_mult_6_net80302), .ZN(
        MULT_mult_6_CARRYB_7__18_) );
  XNOR2_X2 MULT_mult_6_U3346 ( .A(MULT_mult_6_ab_8__18_), .B(MULT_mult_6_n1108), .ZN(MULT_mult_6_net79939) );
  INV_X4 MULT_mult_6_U3345 ( .A(MULT_mult_6_CARRYB_7__18_), .ZN(
        MULT_mult_6_n1108) );
  INV_X4 MULT_mult_6_U3344 ( .A(MULT_mult_6_n1108), .ZN(MULT_mult_6_n1109) );
  NAND2_X2 MULT_mult_6_U3343 ( .A1(MULT_mult_6_SUMB_7__19_), .A2(
        MULT_mult_6_n1109), .ZN(MULT_mult_6_n1107) );
  CLKBUF_X2 MULT_mult_6_U3342 ( .A(MULT_mult_6_CARRYB_12__15_), .Z(
        MULT_mult_6_net93674) );
  NAND2_X1 MULT_mult_6_U3341 ( .A1(MULT_mult_6_ab_13__15_), .A2(
        MULT_mult_6_net93674), .ZN(MULT_mult_6_net79891) );
  NAND2_X1 MULT_mult_6_U3340 ( .A1(MULT_mult_6_net93674), .A2(
        MULT_mult_6_SUMB_12__16_), .ZN(MULT_mult_6_net79893) );
  NAND2_X1 MULT_mult_6_U3339 ( .A1(MULT_mult_6_ab_13__15_), .A2(
        MULT_mult_6_SUMB_12__16_), .ZN(MULT_mult_6_net79892) );
  NOR2_X1 MULT_mult_6_U3338 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net70463), .ZN(MULT_mult_6_ab_16__13_) );
  NAND3_X4 MULT_mult_6_U3337 ( .A1(MULT_mult_6_net87011), .A2(
        MULT_mult_6_net87010), .A3(MULT_mult_6_net87012), .ZN(
        MULT_mult_6_CARRYB_17__11_) );
  NAND2_X1 MULT_mult_6_U3336 ( .A1(MULT_mult_6_ab_18__11_), .A2(
        MULT_mult_6_CARRYB_17__11_), .ZN(MULT_mult_6_net82664) );
  NOR2_X1 MULT_mult_6_U3335 ( .A1(MULT_mult_6_net85716), .A2(
        MULT_mult_6_net70459), .ZN(MULT_mult_6_ab_18__11_) );
  XNOR2_X2 MULT_mult_6_U3334 ( .A(MULT_mult_6_ab_18__11_), .B(
        MULT_mult_6_CARRYB_17__11_), .ZN(MULT_mult_6_net89353) );
  NAND2_X1 MULT_mult_6_U3333 ( .A1(MULT_mult_6_SUMB_18__11_), .A2(
        MULT_mult_6_CARRYB_18__10_), .ZN(MULT_mult_6_net82668) );
  NAND2_X1 MULT_mult_6_U3332 ( .A1(MULT_mult_6_ab_19__10_), .A2(
        MULT_mult_6_SUMB_18__11_), .ZN(MULT_mult_6_net82669) );
  XNOR2_X2 MULT_mult_6_U3331 ( .A(MULT_mult_6_n1104), .B(
        MULT_mult_6_SUMB_6__20_), .ZN(MULT_mult_6_SUMB_7__19_) );
  XNOR2_X2 MULT_mult_6_U3330 ( .A(MULT_mult_6_CARRYB_6__19_), .B(
        MULT_mult_6_ab_7__19_), .ZN(MULT_mult_6_n1104) );
  NAND2_X1 MULT_mult_6_U3329 ( .A1(MULT_mult_6_ab_7__20_), .A2(
        MULT_mult_6_CARRYB_6__20_), .ZN(MULT_mult_6_net79961) );
  NAND2_X1 MULT_mult_6_U3328 ( .A1(MULT_mult_6_CARRYB_6__20_), .A2(
        MULT_mult_6_n840), .ZN(MULT_mult_6_net79959) );
  NAND2_X2 MULT_mult_6_U3327 ( .A1(MULT_mult_6_ab_7__20_), .A2(
        MULT_mult_6_n840), .ZN(MULT_mult_6_net79960) );
  INV_X8 MULT_mult_6_U3326 ( .A(n5943), .ZN(MULT_mult_6_net86565) );
  NOR2_X1 MULT_mult_6_U3325 ( .A1(MULT_mult_6_net86565), .A2(
        MULT_mult_6_net77926), .ZN(MULT_mult_6_ab_8__19_) );
  NAND2_X2 MULT_mult_6_U3324 ( .A1(MULT_mult_6_ab_7__19_), .A2(
        MULT_mult_6_SUMB_6__20_), .ZN(MULT_mult_6_n1102) );
  NAND2_X1 MULT_mult_6_U3323 ( .A1(MULT_mult_6_ab_7__19_), .A2(
        MULT_mult_6_CARRYB_6__19_), .ZN(MULT_mult_6_n1101) );
  NAND2_X2 MULT_mult_6_U3322 ( .A1(MULT_mult_6_ab_8__19_), .A2(
        MULT_mult_6_CARRYB_7__19_), .ZN(MULT_mult_6_net79957) );
  NAND3_X4 MULT_mult_6_U3321 ( .A1(MULT_mult_6_n1103), .A2(MULT_mult_6_n1102), 
        .A3(MULT_mult_6_n1101), .ZN(MULT_mult_6_CARRYB_7__19_) );
  NAND2_X1 MULT_mult_6_U3320 ( .A1(MULT_mult_6_CARRYB_7__19_), .A2(
        MULT_mult_6_SUMB_7__20_), .ZN(MULT_mult_6_net79955) );
  XNOR2_X2 MULT_mult_6_U3319 ( .A(MULT_mult_6_CARRYB_7__19_), .B(
        MULT_mult_6_ab_8__19_), .ZN(MULT_mult_6_net86231) );
  XNOR2_X2 MULT_mult_6_U3318 ( .A(MULT_mult_6_SUMB_7__20_), .B(
        MULT_mult_6_net86231), .ZN(MULT_mult_6_SUMB_8__19_) );
  NAND2_X1 MULT_mult_6_U3317 ( .A1(MULT_mult_6_ab_9__18_), .A2(
        MULT_mult_6_CARRYB_8__18_), .ZN(MULT_mult_6_net79953) );
  NAND2_X1 MULT_mult_6_U3316 ( .A1(MULT_mult_6_CARRYB_8__18_), .A2(
        MULT_mult_6_n32), .ZN(MULT_mult_6_net79951) );
  NAND2_X1 MULT_mult_6_U3315 ( .A1(MULT_mult_6_ab_9__18_), .A2(
        MULT_mult_6_SUMB_8__19_), .ZN(MULT_mult_6_net79952) );
  XOR2_X2 MULT_mult_6_U3314 ( .A(MULT_mult_6_n32), .B(MULT_mult_6_net79950), 
        .Z(MULT_mult_6_SUMB_9__18_) );
  NAND2_X2 MULT_mult_6_U3313 ( .A1(MULT_mult_6_net89467), .A2(
        MULT_mult_6_net89289), .ZN(MULT_mult_6_n1100) );
  NAND3_X4 MULT_mult_6_U3312 ( .A1(MULT_mult_6_n1100), .A2(
        MULT_mult_6_net81956), .A3(MULT_mult_6_net81955), .ZN(
        MULT_mult_6_CARRYB_20__8_) );
  NOR2_X4 MULT_mult_6_U3311 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net70453), .ZN(MULT_mult_6_ab_21__8_) );
  NAND2_X1 MULT_mult_6_U3310 ( .A1(MULT_mult_6_ab_22__8_), .A2(
        MULT_mult_6_CARRYB_21__8_), .ZN(MULT_mult_6_net81180) );
  NAND2_X1 MULT_mult_6_U3309 ( .A1(MULT_mult_6_n856), .A2(
        MULT_mult_6_CARRYB_21__8_), .ZN(MULT_mult_6_net81178) );
  NAND2_X2 MULT_mult_6_U3308 ( .A1(MULT_mult_6_CARRYB_21__8_), .A2(
        MULT_mult_6_ab_22__8_), .ZN(MULT_mult_6_n1098) );
  INV_X4 MULT_mult_6_U3307 ( .A(MULT_mult_6_CARRYB_21__8_), .ZN(
        MULT_mult_6_n1096) );
  INV_X1 MULT_mult_6_U3306 ( .A(MULT_mult_6_ab_22__8_), .ZN(MULT_mult_6_n1097)
         );
  NAND2_X4 MULT_mult_6_U3305 ( .A1(MULT_mult_6_n1096), .A2(MULT_mult_6_n1097), 
        .ZN(MULT_mult_6_n1099) );
  NAND2_X4 MULT_mult_6_U3304 ( .A1(MULT_mult_6_n1098), .A2(MULT_mult_6_n1099), 
        .ZN(MULT_mult_6_n1095) );
  XNOR2_X2 MULT_mult_6_U3303 ( .A(MULT_mult_6_n1095), .B(
        MULT_mult_6_SUMB_21__9_), .ZN(MULT_mult_6_SUMB_22__8_) );
  NOR2_X1 MULT_mult_6_U3302 ( .A1(MULT_mult_6_net84698), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__14_) );
  INV_X1 MULT_mult_6_U3301 ( .A(MULT_mult_6_ab_22__7_), .ZN(
        MULT_mult_6_net81491) );
  NAND2_X1 MULT_mult_6_U3300 ( .A1(MULT_mult_6_ab_23__7_), .A2(
        MULT_mult_6_CARRYB_22__7_), .ZN(MULT_mult_6_net86414) );
  NOR2_X1 MULT_mult_6_U3299 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__13_) );
  XNOR2_X2 MULT_mult_6_U3298 ( .A(MULT_mult_6_CARRYB_10__15_), .B(
        MULT_mult_6_ab_11__15_), .ZN(MULT_mult_6_n1094) );
  NOR2_X2 MULT_mult_6_U3297 ( .A1(MULT_mult_6_net81424), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__15_) );
  NAND2_X2 MULT_mult_6_U3296 ( .A1(MULT_mult_6_ab_11__15_), .A2(
        MULT_mult_6_SUMB_10__16_), .ZN(MULT_mult_6_n1092) );
  NAND2_X1 MULT_mult_6_U3295 ( .A1(MULT_mult_6_ab_11__15_), .A2(
        MULT_mult_6_CARRYB_10__15_), .ZN(MULT_mult_6_n1093) );
  NAND3_X2 MULT_mult_6_U3294 ( .A1(MULT_mult_6_n1091), .A2(MULT_mult_6_n1092), 
        .A3(MULT_mult_6_n1093), .ZN(MULT_mult_6_CARRYB_11__15_) );
  NAND2_X1 MULT_mult_6_U3293 ( .A1(MULT_mult_6_SUMB_22__8_), .A2(
        MULT_mult_6_CARRYB_22__7_), .ZN(MULT_mult_6_net86412) );
  XNOR2_X2 MULT_mult_6_U3292 ( .A(MULT_mult_6_SUMB_22__8_), .B(
        MULT_mult_6_net88961), .ZN(MULT_mult_6_SUMB_23__7_) );
  NAND2_X2 MULT_mult_6_U3291 ( .A1(MULT_mult_6_ab_24__6_), .A2(
        MULT_mult_6_CARRYB_23__6_), .ZN(MULT_mult_6_net79863) );
  XNOR2_X2 MULT_mult_6_U3290 ( .A(MULT_mult_6_n949), .B(MULT_mult_6_n867), 
        .ZN(MULT_mult_6_net89094) );
  INV_X2 MULT_mult_6_U3289 ( .A(MULT_mult_6_ab_24__6_), .ZN(
        MULT_mult_6_net83115) );
  INV_X4 MULT_mult_6_U3288 ( .A(MULT_mult_6_CARRYB_23__6_), .ZN(
        MULT_mult_6_net83116) );
  NAND2_X4 MULT_mult_6_U3287 ( .A1(MULT_mult_6_net83116), .A2(
        MULT_mult_6_net83115), .ZN(MULT_mult_6_n1090) );
  NAND2_X2 MULT_mult_6_U3286 ( .A1(MULT_mult_6_CARRYB_3__23_), .A2(
        MULT_mult_6_ab_4__23_), .ZN(MULT_mult_6_net80791) );
  NAND2_X2 MULT_mult_6_U3285 ( .A1(MULT_mult_6_CARRYB_3__23_), .A2(
        MULT_mult_6_SUMB_3__24_), .ZN(MULT_mult_6_net80792) );
  NAND2_X2 MULT_mult_6_U3284 ( .A1(MULT_mult_6_ab_4__23_), .A2(
        MULT_mult_6_SUMB_3__24_), .ZN(MULT_mult_6_net80793) );
  XNOR2_X2 MULT_mult_6_U3283 ( .A(MULT_mult_6_CARRYB_3__23_), .B(
        MULT_mult_6_ab_4__23_), .ZN(MULT_mult_6_n1088) );
  INV_X16 MULT_mult_6_U3282 ( .A(net36479), .ZN(MULT_mult_6_net70482) );
  NOR2_X1 MULT_mult_6_U3281 ( .A1(MULT_mult_6_net84698), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__14_) );
  NAND2_X1 MULT_mult_6_U3280 ( .A1(MULT_mult_6_ab_16__13_), .A2(
        MULT_mult_6_CARRYB_15__13_), .ZN(MULT_mult_6_net80275) );
  NAND2_X1 MULT_mult_6_U3279 ( .A1(MULT_mult_6_CARRYB_15__13_), .A2(
        MULT_mult_6_net90525), .ZN(MULT_mult_6_net80273) );
  NAND2_X1 MULT_mult_6_U3278 ( .A1(MULT_mult_6_CARRYB_14__14_), .A2(
        MULT_mult_6_SUMB_14__15_), .ZN(MULT_mult_6_net84308) );
  NAND2_X1 MULT_mult_6_U3277 ( .A1(MULT_mult_6_ab_15__14_), .A2(
        MULT_mult_6_SUMB_14__15_), .ZN(MULT_mult_6_net84309) );
  INV_X1 MULT_mult_6_U3276 ( .A(MULT_mult_6_ab_16__12_), .ZN(
        MULT_mult_6_net87003) );
  XNOR2_X2 MULT_mult_6_U3275 ( .A(MULT_mult_6_net82641), .B(
        MULT_mult_6_SUMB_15__13_), .ZN(MULT_mult_6_SUMB_16__12_) );
  NAND2_X2 MULT_mult_6_U3274 ( .A1(MULT_mult_6_ab_16__12_), .A2(
        MULT_mult_6_CARRYB_15__12_), .ZN(MULT_mult_6_net87005) );
  XNOR2_X2 MULT_mult_6_U3273 ( .A(MULT_mult_6_CARRYB_15__13_), .B(
        MULT_mult_6_ab_16__13_), .ZN(MULT_mult_6_net81290) );
  NAND2_X1 MULT_mult_6_U3272 ( .A1(MULT_mult_6_ab_16__13_), .A2(
        MULT_mult_6_SUMB_15__14_), .ZN(MULT_mult_6_net80274) );
  XNOR2_X2 MULT_mult_6_U3271 ( .A(MULT_mult_6_SUMB_14__15_), .B(
        MULT_mult_6_net86054), .ZN(MULT_mult_6_SUMB_15__14_) );
  NAND2_X1 MULT_mult_6_U3270 ( .A1(MULT_mult_6_ab_16__12_), .A2(
        MULT_mult_6_CARRYB_15__12_), .ZN(MULT_mult_6_n1085) );
  XNOR2_X2 MULT_mult_6_U3269 ( .A(MULT_mult_6_SUMB_15__14_), .B(
        MULT_mult_6_net81290), .ZN(MULT_mult_6_SUMB_16__13_) );
  XNOR2_X2 MULT_mult_6_U3268 ( .A(MULT_mult_6_SUMB_17__12_), .B(
        MULT_mult_6_net89353), .ZN(MULT_mult_6_SUMB_18__11_) );
  NAND2_X1 MULT_mult_6_U3267 ( .A1(MULT_mult_6_ab_18__12_), .A2(
        MULT_mult_6_CARRYB_17__12_), .ZN(MULT_mult_6_net80449) );
  NAND2_X1 MULT_mult_6_U3266 ( .A1(MULT_mult_6_CARRYB_17__12_), .A2(
        MULT_mult_6_SUMB_17__13_), .ZN(MULT_mult_6_net80451) );
  XNOR2_X2 MULT_mult_6_U3265 ( .A(MULT_mult_6_ab_18__12_), .B(
        MULT_mult_6_CARRYB_17__12_), .ZN(MULT_mult_6_net88165) );
  NOR2_X2 MULT_mult_6_U3264 ( .A1(MULT_mult_6_net70480), .A2(
        MULT_mult_6_net86101), .ZN(MULT_mult_6_ab_1__23_) );
  INV_X8 MULT_mult_6_U3263 ( .A(n10912), .ZN(MULT_mult_6_net70480) );
  INV_X2 MULT_mult_6_U3262 ( .A(MULT_mult_6_net70480), .ZN(
        MULT_mult_6_net84357) );
  NOR2_X2 MULT_mult_6_U3261 ( .A1(MULT_mult_6_net84358), .A2(
        MULT_mult_6_net77964), .ZN(MULT_mult_6_ab_3__23_) );
  NOR2_X1 MULT_mult_6_U3260 ( .A1(MULT_mult_6_net70447), .A2(
        MULT_mult_6_net77912), .ZN(MULT_mult_6_ab_24__7_) );
  XOR2_X2 MULT_mult_6_U3259 ( .A(MULT_mult_6_CARRYB_23__7_), .B(
        MULT_mult_6_ab_24__7_), .Z(MULT_mult_6_n1084) );
  NAND3_X2 MULT_mult_6_U3258 ( .A1(MULT_mult_6_net79865), .A2(
        MULT_mult_6_net79864), .A3(MULT_mult_6_net79863), .ZN(
        MULT_mult_6_CARRYB_24__6_) );
  OR2_X2 MULT_mult_6_U3257 ( .A1(MULT_mult_6_net70445), .A2(
        MULT_mult_6_net77906), .ZN(MULT_mult_6_net81946) );
  XNOR2_X2 MULT_mult_6_U3256 ( .A(MULT_mult_6_CARRYB_24__6_), .B(
        MULT_mult_6_net81946), .ZN(MULT_mult_6_n1083) );
  NOR2_X1 MULT_mult_6_U3255 ( .A1(MULT_mult_6_net70443), .A2(
        MULT_mult_6_net77898), .ZN(MULT_mult_6_ab_26__5_) );
  NAND2_X1 MULT_mult_6_U3254 ( .A1(MULT_mult_6_n1082), .A2(
        MULT_mult_6_SUMB_25__5_), .ZN(MULT_mult_6_n1079) );
  BUF_X8 MULT_mult_6_U3253 ( .A(MULT_mult_6_CARRYB_25__4_), .Z(
        MULT_mult_6_n1082) );
  NAND2_X1 MULT_mult_6_U3252 ( .A1(MULT_mult_6_ab_26__4_), .A2(
        MULT_mult_6_n1082), .ZN(MULT_mult_6_n1081) );
  NAND3_X2 MULT_mult_6_U3251 ( .A1(MULT_mult_6_n1079), .A2(MULT_mult_6_n1080), 
        .A3(MULT_mult_6_n1081), .ZN(MULT_mult_6_CARRYB_26__4_) );
  NOR2_X1 MULT_mult_6_U3250 ( .A1(MULT_mult_6_net70441), .A2(
        MULT_mult_6_net77892), .ZN(MULT_mult_6_ab_27__4_) );
  XOR2_X2 MULT_mult_6_U3249 ( .A(MULT_mult_6_CARRYB_26__4_), .B(
        MULT_mult_6_ab_27__4_), .Z(MULT_mult_6_net82807) );
  XNOR2_X2 MULT_mult_6_U3248 ( .A(MULT_mult_6_SUMB_26__5_), .B(
        MULT_mult_6_net82807), .ZN(MULT_mult_6_net86937) );
  INV_X4 MULT_mult_6_U3247 ( .A(net70534), .ZN(MULT_mult_6_n1078) );
  XNOR2_X2 MULT_mult_6_U3246 ( .A(MULT_mult_6_ab_31__0_), .B(
        MULT_mult_6_net92320), .ZN(MULT_mult_6_net92319) );
  XNOR2_X2 MULT_mult_6_U3245 ( .A(MULT_mult_6_net86937), .B(
        MULT_mult_6_net92319), .ZN(MULT_mult_6_net92323) );
  XNOR2_X2 MULT_mult_6_U3244 ( .A(MULT_mult_6_net88004), .B(MULT_mult_6_n2357), 
        .ZN(MULT_mult_6_SUMB_2__23_) );
  XOR2_X2 MULT_mult_6_U3243 ( .A(MULT_mult_6_ab_1__24_), .B(
        MULT_mult_6_ab_0__25_), .Z(MULT_mult_6_net83044) );
  INV_X4 MULT_mult_6_U3242 ( .A(MULT_mult_6_ab_1__23_), .ZN(
        MULT_mult_6_net82043) );
  NAND2_X2 MULT_mult_6_U3241 ( .A1(MULT_mult_6_net82043), .A2(
        MULT_mult_6_net82044), .ZN(MULT_mult_6_net82046) );
  NAND2_X1 MULT_mult_6_U3240 ( .A1(MULT_mult_6_ab_2__23_), .A2(
        MULT_mult_6_net82124), .ZN(MULT_mult_6_n1077) );
  XNOR2_X2 MULT_mult_6_U3239 ( .A(MULT_mult_6_ab_2__23_), .B(
        MULT_mult_6_net82124), .ZN(MULT_mult_6_net88004) );
  NAND3_X2 MULT_mult_6_U3238 ( .A1(MULT_mult_6_net83575), .A2(
        MULT_mult_6_n1077), .A3(MULT_mult_6_net83576), .ZN(
        MULT_mult_6_CARRYB_2__23_) );
  XNOR2_X2 MULT_mult_6_U3237 ( .A(MULT_mult_6_ab_21__8_), .B(
        MULT_mult_6_CARRYB_20__8_), .ZN(MULT_mult_6_net90801) );
  NAND2_X1 MULT_mult_6_U3236 ( .A1(MULT_mult_6_ab_21__8_), .A2(
        MULT_mult_6_CARRYB_20__8_), .ZN(MULT_mult_6_net81036) );
  XNOR2_X2 MULT_mult_6_U3235 ( .A(MULT_mult_6_CARRYB_20__7_), .B(
        MULT_mult_6_ab_21__7_), .ZN(MULT_mult_6_net83134) );
  XNOR2_X2 MULT_mult_6_U3234 ( .A(MULT_mult_6_ab_21__8_), .B(
        MULT_mult_6_CARRYB_20__8_), .ZN(MULT_mult_6_net81113) );
  NAND2_X2 MULT_mult_6_U3231 ( .A1(MULT_mult_6_CARRYB_20__7_), .A2(
        MULT_mult_6_SUMB_20__8_), .ZN(MULT_mult_6_n1074) );
  NAND2_X2 MULT_mult_6_U3230 ( .A1(MULT_mult_6_SUMB_20__8_), .A2(
        MULT_mult_6_ab_21__7_), .ZN(MULT_mult_6_n1073) );
  NAND2_X1 MULT_mult_6_U3229 ( .A1(MULT_mult_6_ab_21__7_), .A2(
        MULT_mult_6_CARRYB_20__7_), .ZN(MULT_mult_6_n1072) );
  NAND2_X1 MULT_mult_6_U3228 ( .A1(MULT_mult_6_CARRYB_21__7_), .A2(
        MULT_mult_6_ab_22__7_), .ZN(MULT_mult_6_n1071) );
  NAND3_X4 MULT_mult_6_U3227 ( .A1(MULT_mult_6_n1074), .A2(MULT_mult_6_n1073), 
        .A3(MULT_mult_6_n1072), .ZN(MULT_mult_6_CARRYB_21__7_) );
  NAND2_X2 MULT_mult_6_U3226 ( .A1(MULT_mult_6_CARRYB_2__23_), .A2(
        MULT_mult_6_SUMB_2__24_), .ZN(MULT_mult_6_net84302) );
  NAND2_X1 MULT_mult_6_U3225 ( .A1(MULT_mult_6_n262), .A2(
        MULT_mult_6_SUMB_23__7_), .ZN(MULT_mult_6_net79865) );
  NAND2_X2 MULT_mult_6_U3224 ( .A1(MULT_mult_6_ab_25__5_), .A2(
        MULT_mult_6_CARRYB_24__5_), .ZN(MULT_mult_6_net86699) );
  INV_X1 MULT_mult_6_U3223 ( .A(MULT_mult_6_ab_25__5_), .ZN(
        MULT_mult_6_net86697) );
  NOR2_X4 MULT_mult_6_U3222 ( .A1(MULT_mult_6_net77898), .A2(
        MULT_mult_6_net70445), .ZN(MULT_mult_6_ab_25__5_) );
  NAND2_X2 MULT_mult_6_U3221 ( .A1(MULT_mult_6_SUMB_2__24_), .A2(
        MULT_mult_6_ab_3__23_), .ZN(MULT_mult_6_net84301) );
  NAND2_X1 MULT_mult_6_U3220 ( .A1(MULT_mult_6_ab_3__23_), .A2(
        MULT_mult_6_CARRYB_2__23_), .ZN(MULT_mult_6_net84300) );
  NAND2_X2 MULT_mult_6_U3219 ( .A1(MULT_mult_6_SUMB_1__25_), .A2(
        MULT_mult_6_n838), .ZN(MULT_mult_6_net84298) );
  NAND2_X1 MULT_mult_6_U3218 ( .A1(MULT_mult_6_n39), .A2(MULT_mult_6_ab_2__24_), .ZN(MULT_mult_6_net84299) );
  XNOR2_X2 MULT_mult_6_U3217 ( .A(MULT_mult_6_net84883), .B(
        MULT_mult_6_ab_2__24_), .ZN(MULT_mult_6_SUMB_2__24_) );
  XNOR2_X2 MULT_mult_6_U3216 ( .A(MULT_mult_6_ab_3__23_), .B(
        MULT_mult_6_CARRYB_2__23_), .ZN(MULT_mult_6_net87855) );
  XNOR2_X2 MULT_mult_6_U3215 ( .A(MULT_mult_6_net87855), .B(
        MULT_mult_6_net90671), .ZN(MULT_mult_6_SUMB_3__23_) );
  NAND2_X2 MULT_mult_6_U3214 ( .A1(MULT_mult_6_ab_3__22_), .A2(
        MULT_mult_6_SUMB_2__23_), .ZN(MULT_mult_6_n1069) );
  NOR2_X1 MULT_mult_6_U3213 ( .A1(MULT_mult_6_net70478), .A2(
        MULT_mult_6_net77956), .ZN(MULT_mult_6_ab_4__22_) );
  XNOR2_X2 MULT_mult_6_U3212 ( .A(MULT_mult_6_net80825), .B(
        MULT_mult_6_SUMB_4__23_), .ZN(MULT_mult_6_SUMB_5__22_) );
  XNOR2_X2 MULT_mult_6_U3211 ( .A(MULT_mult_6_ab_12__14_), .B(
        MULT_mult_6_CARRYB_11__14_), .ZN(MULT_mult_6_n1067) );
  FA_X1 MULT_mult_6_U3210 ( .A(MULT_mult_6_n111), .B(MULT_mult_6_ab_12__15_), 
        .CI(MULT_mult_6_SUMB_11__16_), .S(MULT_mult_6_net88756) );
  NAND2_X2 MULT_mult_6_U3209 ( .A1(MULT_mult_6_ab_12__14_), .A2(
        MULT_mult_6_SUMB_11__15_), .ZN(MULT_mult_6_n1065) );
  NAND2_X1 MULT_mult_6_U3208 ( .A1(MULT_mult_6_ab_12__14_), .A2(
        MULT_mult_6_CARRYB_11__14_), .ZN(MULT_mult_6_n1064) );
  NAND2_X1 MULT_mult_6_U3207 ( .A1(MULT_mult_6_ab_13__14_), .A2(
        MULT_mult_6_CARRYB_12__14_), .ZN(MULT_mult_6_n1063) );
  XNOR2_X2 MULT_mult_6_U3206 ( .A(MULT_mult_6_ab_13__14_), .B(
        MULT_mult_6_CARRYB_12__14_), .ZN(MULT_mult_6_net84481) );
  NAND3_X4 MULT_mult_6_U3205 ( .A1(MULT_mult_6_n1066), .A2(MULT_mult_6_n1065), 
        .A3(MULT_mult_6_n1064), .ZN(MULT_mult_6_CARRYB_12__14_) );
  NAND3_X2 MULT_mult_6_U3204 ( .A1(MULT_mult_6_net82658), .A2(
        MULT_mult_6_net82657), .A3(MULT_mult_6_n1063), .ZN(
        MULT_mult_6_CARRYB_13__14_) );
  NAND3_X2 MULT_mult_6_U3203 ( .A1(MULT_mult_6_net79969), .A2(
        MULT_mult_6_net79968), .A3(MULT_mult_6_net79970), .ZN(
        MULT_mult_6_CARRYB_24__5_) );
  NAND2_X1 MULT_mult_6_U3202 ( .A1(MULT_mult_6_ab_24__6_), .A2(
        MULT_mult_6_net89094), .ZN(MULT_mult_6_net79864) );
  XNOR2_X2 MULT_mult_6_U3201 ( .A(MULT_mult_6_net80110), .B(
        MULT_mult_6_SUMB_23__7_), .ZN(MULT_mult_6_SUMB_24__6_) );
  NAND2_X1 MULT_mult_6_U3200 ( .A1(MULT_mult_6_ab_25__5_), .A2(
        MULT_mult_6_net86696), .ZN(MULT_mult_6_n1062) );
  NAND3_X1 MULT_mult_6_U3199 ( .A1(MULT_mult_6_net79969), .A2(
        MULT_mult_6_net79970), .A3(MULT_mult_6_net79968), .ZN(
        MULT_mult_6_net86696) );
  NAND2_X2 MULT_mult_6_U3198 ( .A1(MULT_mult_6_net81815), .A2(
        MULT_mult_6_net88916), .ZN(MULT_mult_6_net84305) );
  XNOR2_X2 MULT_mult_6_U3197 ( .A(MULT_mult_6_net89094), .B(
        MULT_mult_6_net80110), .ZN(MULT_mult_6_net88916) );
  NAND2_X1 MULT_mult_6_U3196 ( .A1(MULT_mult_6_ab_14__14_), .A2(
        MULT_mult_6_CARRYB_13__14_), .ZN(MULT_mult_6_net80480) );
  NAND2_X1 MULT_mult_6_U3195 ( .A1(MULT_mult_6_CARRYB_13__14_), .A2(
        MULT_mult_6_SUMB_13__15_), .ZN(MULT_mult_6_net80478) );
  NAND2_X2 MULT_mult_6_U3194 ( .A1(MULT_mult_6_SUMB_13__14_), .A2(
        MULT_mult_6_n695), .ZN(MULT_mult_6_n1061) );
  NAND2_X1 MULT_mult_6_U3193 ( .A1(MULT_mult_6_ab_14__13_), .A2(
        MULT_mult_6_CARRYB_13__13_), .ZN(MULT_mult_6_n1059) );
  NAND2_X1 MULT_mult_6_U3192 ( .A1(MULT_mult_6_ab_15__13_), .A2(
        MULT_mult_6_CARRYB_14__13_), .ZN(MULT_mult_6_n1058) );
  XNOR2_X2 MULT_mult_6_U3191 ( .A(MULT_mult_6_CARRYB_14__13_), .B(
        MULT_mult_6_ab_15__13_), .ZN(MULT_mult_6_net93107) );
  XNOR2_X2 MULT_mult_6_U3190 ( .A(MULT_mult_6_CARRYB_13__14_), .B(
        MULT_mult_6_ab_14__14_), .ZN(MULT_mult_6_net85119) );
  XOR2_X2 MULT_mult_6_U3189 ( .A(MULT_mult_6_SUMB_3__23_), .B(
        MULT_mult_6_net84311), .Z(MULT_mult_6_SUMB_4__22_) );
  XOR2_X2 MULT_mult_6_U3188 ( .A(MULT_mult_6_CARRYB_3__22_), .B(
        MULT_mult_6_ab_4__22_), .Z(MULT_mult_6_net84311) );
  NAND2_X2 MULT_mult_6_U3187 ( .A1(MULT_mult_6_CARRYB_3__22_), .A2(
        MULT_mult_6_SUMB_3__23_), .ZN(MULT_mult_6_net84312) );
  NAND2_X1 MULT_mult_6_U3186 ( .A1(MULT_mult_6_ab_4__22_), .A2(
        MULT_mult_6_CARRYB_3__22_), .ZN(MULT_mult_6_n1057) );
  NAND2_X1 MULT_mult_6_U3185 ( .A1(MULT_mult_6_CARRYB_4__22_), .A2(
        MULT_mult_6_SUMB_4__23_), .ZN(MULT_mult_6_net80796) );
  INV_X16 MULT_mult_6_U3184 ( .A(n10913), .ZN(MULT_mult_6_net70478) );
  NOR2_X1 MULT_mult_6_U3183 ( .A1(MULT_mult_6_net70478), .A2(
        MULT_mult_6_net77948), .ZN(MULT_mult_6_ab_5__22_) );
  INV_X4 MULT_mult_6_U3182 ( .A(MULT_mult_6_CARRYB_4__22_), .ZN(
        MULT_mult_6_net81285) );
  INV_X1 MULT_mult_6_U3181 ( .A(MULT_mult_6_ab_5__22_), .ZN(
        MULT_mult_6_net81284) );
  NAND2_X2 MULT_mult_6_U3180 ( .A1(MULT_mult_6_net80794), .A2(
        MULT_mult_6_n1056), .ZN(MULT_mult_6_net80825) );
  NAND2_X2 MULT_mult_6_U3179 ( .A1(MULT_mult_6_net81285), .A2(
        MULT_mult_6_net81284), .ZN(MULT_mult_6_n1056) );
  NAND2_X1 MULT_mult_6_U3178 ( .A1(MULT_mult_6_ab_11__16_), .A2(
        MULT_mult_6_CARRYB_10__16_), .ZN(MULT_mult_6_net80521) );
  NAND2_X1 MULT_mult_6_U3177 ( .A1(MULT_mult_6_ab_10__17_), .A2(
        MULT_mult_6_CARRYB_9__17_), .ZN(MULT_mult_6_net80518) );
  NAND2_X1 MULT_mult_6_U3176 ( .A1(MULT_mult_6_CARRYB_9__17_), .A2(
        MULT_mult_6_n573), .ZN(MULT_mult_6_net80520) );
  NAND2_X1 MULT_mult_6_U3175 ( .A1(MULT_mult_6_ab_10__17_), .A2(
        MULT_mult_6_n573), .ZN(MULT_mult_6_net80519) );
  INV_X4 MULT_mult_6_U3174 ( .A(MULT_mult_6_ab_11__16_), .ZN(
        MULT_mult_6_net81394) );
  XNOR2_X2 MULT_mult_6_U3173 ( .A(MULT_mult_6_CARRYB_10__16_), .B(
        MULT_mult_6_net81394), .ZN(MULT_mult_6_net80517) );
  NAND2_X2 MULT_mult_6_U3172 ( .A1(MULT_mult_6_net80517), .A2(
        MULT_mult_6_net88225), .ZN(MULT_mult_6_net86409) );
  XNOR2_X2 MULT_mult_6_U3171 ( .A(MULT_mult_6_net88226), .B(
        MULT_mult_6_SUMB_9__18_), .ZN(MULT_mult_6_net88225) );
  NAND2_X1 MULT_mult_6_U3170 ( .A1(MULT_mult_6_ab_11__16_), .A2(
        MULT_mult_6_SUMB_10__17_), .ZN(MULT_mult_6_net80522) );
  NAND2_X1 MULT_mult_6_U3169 ( .A1(MULT_mult_6_CARRYB_10__16_), .A2(
        MULT_mult_6_SUMB_10__17_), .ZN(MULT_mult_6_net80523) );
  INV_X4 MULT_mult_6_U3168 ( .A(MULT_mult_6_net88225), .ZN(
        MULT_mult_6_SUMB_10__17_) );
  NAND2_X4 MULT_mult_6_U3167 ( .A1(MULT_mult_6_net86409), .A2(
        MULT_mult_6_n1055), .ZN(MULT_mult_6_SUMB_11__16_) );
  NAND2_X4 MULT_mult_6_U3166 ( .A1(MULT_mult_6_net86407), .A2(
        MULT_mult_6_SUMB_10__17_), .ZN(MULT_mult_6_n1055) );
  NAND3_X2 MULT_mult_6_U3165 ( .A1(MULT_mult_6_net80257), .A2(MULT_mult_6_n500), .A3(MULT_mult_6_net80258), .ZN(MULT_mult_6_net93840) );
  XNOR2_X2 MULT_mult_6_U3164 ( .A(MULT_mult_6_CARRYB_14__7_), .B(
        MULT_mult_6_ab_15__7_), .ZN(MULT_mult_6_net83755) );
  XNOR2_X2 MULT_mult_6_U3163 ( .A(MULT_mult_6_CARRYB_25__2_), .B(
        MULT_mult_6_net93792), .ZN(MULT_mult_6_net93791) );
  NAND2_X4 MULT_mult_6_U3162 ( .A1(MULT_mult_6_SUMB_26__2_), .A2(
        MULT_mult_6_CARRYB_26__1_), .ZN(MULT_mult_6_net80992) );
  XNOR2_X2 MULT_mult_6_U3161 ( .A(MULT_mult_6_net121859), .B(
        MULT_mult_6_net149611), .ZN(MULT_mult_6_net119817) );
  NOR2_X4 MULT_mult_6_U3160 ( .A1(MULT_mult_6_n1111), .A2(MULT_mult_6_net81673), .ZN(MULT_mult_6_ab_0__25_) );
  INV_X4 MULT_mult_6_U3159 ( .A(MULT_mult_6_CARRYB_11__9_), .ZN(
        MULT_mult_6_net119979) );
  NAND2_X4 MULT_mult_6_U3158 ( .A1(MULT_mult_6_net119979), .A2(
        MULT_mult_6_n1054), .ZN(MULT_mult_6_net119982) );
  NAND2_X2 MULT_mult_6_U3157 ( .A1(MULT_mult_6_ab_4__21_), .A2(
        MULT_mult_6_SUMB_3__22_), .ZN(MULT_mult_6_n2277) );
  NAND2_X4 MULT_mult_6_U3156 ( .A1(MULT_mult_6_n1603), .A2(
        MULT_mult_6_net86601), .ZN(MULT_mult_6_n1605) );
  NAND2_X4 MULT_mult_6_U3155 ( .A1(MULT_mult_6_n1738), .A2(MULT_mult_6_n1739), 
        .ZN(MULT_mult_6_n1740) );
  NAND2_X4 MULT_mult_6_U3154 ( .A1(MULT_mult_6_n2192), .A2(MULT_mult_6_n1740), 
        .ZN(MULT_mult_6_n1765) );
  INV_X8 MULT_mult_6_U3153 ( .A(MULT_mult_6_n2338), .ZN(
        MULT_mult_6_SUMB_1__16_) );
  NAND2_X4 MULT_mult_6_U3152 ( .A1(MULT_mult_6_n1355), .A2(MULT_mult_6_n1262), 
        .ZN(MULT_mult_6_n1358) );
  NAND2_X4 MULT_mult_6_U3151 ( .A1(MULT_mult_6_CARRYB_1__10_), .A2(
        MULT_mult_6_SUMB_1__11_), .ZN(MULT_mult_6_n1654) );
  NAND2_X2 MULT_mult_6_U3150 ( .A1(MULT_mult_6_ab_5__13_), .A2(
        MULT_mult_6_CARRYB_4__13_), .ZN(MULT_mult_6_n1980) );
  NAND2_X2 MULT_mult_6_U3149 ( .A1(MULT_mult_6_ab_0__23_), .A2(
        MULT_mult_6_n2196), .ZN(MULT_mult_6_n2345) );
  INV_X1 MULT_mult_6_U3148 ( .A(MULT_mult_6_ab_9__18_), .ZN(MULT_mult_6_n1051)
         );
  NAND2_X2 MULT_mult_6_U3147 ( .A1(MULT_mult_6_n1052), .A2(MULT_mult_6_n1053), 
        .ZN(MULT_mult_6_net79950) );
  NAND2_X1 MULT_mult_6_U3146 ( .A1(MULT_mult_6_n1050), .A2(
        MULT_mult_6_ab_9__18_), .ZN(MULT_mult_6_n1053) );
  NAND2_X1 MULT_mult_6_U3145 ( .A1(MULT_mult_6_CARRYB_8__18_), .A2(
        MULT_mult_6_n1051), .ZN(MULT_mult_6_n1052) );
  INV_X2 MULT_mult_6_U3144 ( .A(MULT_mult_6_ab_2__22_), .ZN(MULT_mult_6_n1047)
         );
  NAND2_X2 MULT_mult_6_U3143 ( .A1(MULT_mult_6_n1048), .A2(MULT_mult_6_n1049), 
        .ZN(MULT_mult_6_n1457) );
  NAND2_X2 MULT_mult_6_U3142 ( .A1(MULT_mult_6_n1047), .A2(MULT_mult_6_n2345), 
        .ZN(MULT_mult_6_n1049) );
  NAND2_X2 MULT_mult_6_U3141 ( .A1(MULT_mult_6_ab_2__22_), .A2(
        MULT_mult_6_CARRYB_1__22_), .ZN(MULT_mult_6_n1048) );
  XNOR2_X2 MULT_mult_6_U3140 ( .A(MULT_mult_6_CARRYB_17__3_), .B(
        MULT_mult_6_ab_18__3_), .ZN(MULT_mult_6_n1268) );
  NAND2_X4 MULT_mult_6_U3139 ( .A1(MULT_mult_6_n2243), .A2(
        MULT_mult_6_net83151), .ZN(MULT_mult_6_n1757) );
  NAND3_X2 MULT_mult_6_U3138 ( .A1(MULT_mult_6_n1568), .A2(MULT_mult_6_n1569), 
        .A3(MULT_mult_6_n1570), .ZN(MULT_mult_6_CARRYB_24__0_) );
  NAND2_X2 MULT_mult_6_U3137 ( .A1(MULT_mult_6_CARRYB_11__14_), .A2(
        MULT_mult_6_SUMB_11__15_), .ZN(MULT_mult_6_n1066) );
  INV_X2 MULT_mult_6_U3136 ( .A(MULT_mult_6_n848), .ZN(MULT_mult_6_n1789) );
  NAND2_X4 MULT_mult_6_U3135 ( .A1(MULT_mult_6_n1788), .A2(MULT_mult_6_n1789), 
        .ZN(MULT_mult_6_n1791) );
  NAND2_X1 MULT_mult_6_U3134 ( .A1(MULT_mult_6_ab_22__8_), .A2(
        MULT_mult_6_SUMB_21__9_), .ZN(MULT_mult_6_net81179) );
  NAND2_X4 MULT_mult_6_U3133 ( .A1(MULT_mult_6_n1500), .A2(
        MULT_mult_6_ab_16__4_), .ZN(MULT_mult_6_n2105) );
  NAND3_X4 MULT_mult_6_U3132 ( .A1(MULT_mult_6_net79935), .A2(
        MULT_mult_6_net79936), .A3(MULT_mult_6_net79937), .ZN(
        MULT_mult_6_CARRYB_6__20_) );
  NAND2_X2 MULT_mult_6_U3131 ( .A1(MULT_mult_6_ab_2__12_), .A2(
        MULT_mult_6_CARRYB_1__12_), .ZN(MULT_mult_6_n1045) );
  XOR2_X1 MULT_mult_6_U3130 ( .A(MULT_mult_6_ab_11__1_), .B(
        MULT_mult_6_CARRYB_10__1_), .Z(MULT_mult_6_n1315) );
  NOR2_X2 MULT_mult_6_U3129 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__13_) );
  INV_X1 MULT_mult_6_U3128 ( .A(MULT_mult_6_ab_12__13_), .ZN(MULT_mult_6_n1042) );
  NAND2_X4 MULT_mult_6_U3127 ( .A1(MULT_mult_6_n1795), .A2(MULT_mult_6_n1043), 
        .ZN(MULT_mult_6_n1753) );
  NAND2_X4 MULT_mult_6_U3126 ( .A1(MULT_mult_6_n1041), .A2(MULT_mult_6_n1042), 
        .ZN(MULT_mult_6_n1043) );
  NAND2_X4 MULT_mult_6_U3125 ( .A1(MULT_mult_6_n1037), .A2(MULT_mult_6_n1038), 
        .ZN(MULT_mult_6_n1040) );
  NAND2_X4 MULT_mult_6_U3124 ( .A1(MULT_mult_6_CARRYB_8__11_), .A2(
        MULT_mult_6_ab_9__11_), .ZN(MULT_mult_6_net86895) );
  NAND2_X4 MULT_mult_6_U3123 ( .A1(MULT_mult_6_CARRYB_14__5_), .A2(
        MULT_mult_6_n864), .ZN(MULT_mult_6_n1979) );
  BUF_X8 MULT_mult_6_U3122 ( .A(MULT_mult_6_CARRYB_26__3_), .Z(
        MULT_mult_6_n1272) );
  XNOR2_X2 MULT_mult_6_U3121 ( .A(MULT_mult_6_CARRYB_10__3_), .B(
        MULT_mult_6_ab_11__3_), .ZN(MULT_mult_6_n1200) );
  NAND2_X2 MULT_mult_6_U3120 ( .A1(MULT_mult_6_n170), .A2(MULT_mult_6_n393), 
        .ZN(MULT_mult_6_n1036) );
  NAND2_X2 MULT_mult_6_U3119 ( .A1(MULT_mult_6_net84978), .A2(
        MULT_mult_6_net84979), .ZN(MULT_mult_6_n1035) );
  NAND2_X2 MULT_mult_6_U3118 ( .A1(MULT_mult_6_SUMB_2__15_), .A2(
        MULT_mult_6_n1792), .ZN(MULT_mult_6_n1558) );
  NAND2_X2 MULT_mult_6_U3117 ( .A1(MULT_mult_6_net120359), .A2(
        MULT_mult_6_net93792), .ZN(MULT_mult_6_n1034) );
  NAND2_X1 MULT_mult_6_U3116 ( .A1(MULT_mult_6_ab_7__15_), .A2(
        MULT_mult_6_CARRYB_6__15_), .ZN(MULT_mult_6_n2208) );
  INV_X1 MULT_mult_6_U3115 ( .A(MULT_mult_6_ab_5__10_), .ZN(MULT_mult_6_n1030)
         );
  NAND2_X2 MULT_mult_6_U3113 ( .A1(MULT_mult_6_n1694), .A2(
        MULT_mult_6_CARRYB_5__10_), .ZN(MULT_mult_6_n1170) );
  NAND3_X4 MULT_mult_6_U3112 ( .A1(MULT_mult_6_net82028), .A2(
        MULT_mult_6_net82027), .A3(MULT_mult_6_n1941), .ZN(
        MULT_mult_6_CARRYB_2__17_) );
  NAND2_X4 MULT_mult_6_U3111 ( .A1(MULT_mult_6_n645), .A2(MULT_mult_6_n1372), 
        .ZN(MULT_mult_6_n1374) );
  INV_X2 MULT_mult_6_U3110 ( .A(MULT_mult_6_n2327), .ZN(
        MULT_mult_6_CARRYB_1__4_) );
  XNOR2_X2 MULT_mult_6_U3109 ( .A(MULT_mult_6_n2327), .B(MULT_mult_6_ab_2__4_), 
        .ZN(MULT_mult_6_n1135) );
  NAND2_X2 MULT_mult_6_U3108 ( .A1(MULT_mult_6_SUMB_9__5_), .A2(
        MULT_mult_6_CARRYB_9__4_), .ZN(MULT_mult_6_n1926) );
  XNOR2_X2 MULT_mult_6_U3107 ( .A(MULT_mult_6_net84883), .B(MULT_mult_6_n838), 
        .ZN(MULT_mult_6_net90671) );
  NOR2_X4 MULT_mult_6_U3106 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__8_) );
  INV_X4 MULT_mult_6_U3105 ( .A(MULT_mult_6_net88928), .ZN(
        MULT_mult_6_net120467) );
  NAND2_X4 MULT_mult_6_U3104 ( .A1(MULT_mult_6_n1027), .A2(MULT_mult_6_n1028), 
        .ZN(MULT_mult_6_SUMB_11__8_) );
  NAND2_X4 MULT_mult_6_U3103 ( .A1(MULT_mult_6_net120467), .A2(
        MULT_mult_6_net120468), .ZN(MULT_mult_6_n1028) );
  NAND2_X2 MULT_mult_6_U3102 ( .A1(MULT_mult_6_net88928), .A2(
        MULT_mult_6_net86844), .ZN(MULT_mult_6_n1027) );
  INV_X4 MULT_mult_6_U3101 ( .A(MULT_mult_6_CARRYB_10__8_), .ZN(
        MULT_mult_6_net120463) );
  NAND2_X4 MULT_mult_6_U3100 ( .A1(MULT_mult_6_net120463), .A2(
        MULT_mult_6_net120464), .ZN(MULT_mult_6_net120466) );
  INV_X4 MULT_mult_6_U3099 ( .A(MULT_mult_6_CARRYB_16__5_), .ZN(
        MULT_mult_6_n1380) );
  NAND2_X4 MULT_mult_6_U3098 ( .A1(MULT_mult_6_n1321), .A2(MULT_mult_6_n1320), 
        .ZN(MULT_mult_6_net81756) );
  INV_X4 MULT_mult_6_U3097 ( .A(MULT_mult_6_SUMB_15__12_), .ZN(
        MULT_mult_6_n1847) );
  NAND2_X4 MULT_mult_6_U3096 ( .A1(MULT_mult_6_n1846), .A2(MULT_mult_6_n1847), 
        .ZN(MULT_mult_6_n1849) );
  NAND2_X2 MULT_mult_6_U3095 ( .A1(MULT_mult_6_SUMB_10__15_), .A2(
        MULT_mult_6_ab_11__14_), .ZN(MULT_mult_6_n1843) );
  INV_X8 MULT_mult_6_U3094 ( .A(MULT_mult_6_n1780), .ZN(
        MULT_mult_6_SUMB_23__6_) );
  NOR2_X4 MULT_mult_6_U3093 ( .A1(MULT_mult_6_net70456), .A2(
        MULT_mult_6_net80409), .ZN(MULT_mult_6_ab_1__11_) );
  NAND2_X4 MULT_mult_6_U3092 ( .A1(MULT_mult_6_net86893), .A2(
        MULT_mult_6_net86894), .ZN(MULT_mult_6_net86896) );
  BUF_X4 MULT_mult_6_U3091 ( .A(MULT_mult_6_SUMB_10__9_), .Z(
        MULT_mult_6_net88928) );
  NAND2_X4 MULT_mult_6_U3090 ( .A1(MULT_mult_6_net120519), .A2(
        MULT_mult_6_n1022), .ZN(MULT_mult_6_SUMB_15__7_) );
  NAND2_X4 MULT_mult_6_U3089 ( .A1(MULT_mult_6_net120517), .A2(
        MULT_mult_6_net120518), .ZN(MULT_mult_6_n1022) );
  NAND2_X4 MULT_mult_6_U3088 ( .A1(MULT_mult_6_n1021), .A2(
        MULT_mult_6_net120515), .ZN(MULT_mult_6_SUMB_10__9_) );
  NAND2_X4 MULT_mult_6_U3087 ( .A1(MULT_mult_6_net120513), .A2(
        MULT_mult_6_net120514), .ZN(MULT_mult_6_n1021) );
  NAND2_X1 MULT_mult_6_U3086 ( .A1(MULT_mult_6_ab_4__7_), .A2(
        MULT_mult_6_CARRYB_3__7_), .ZN(MULT_mult_6_n1908) );
  INV_X4 MULT_mult_6_U3085 ( .A(MULT_mult_6_ab_8__7_), .ZN(MULT_mult_6_n1831)
         );
  NAND2_X2 MULT_mult_6_U3084 ( .A1(MULT_mult_6_SUMB_8__8_), .A2(
        MULT_mult_6_ab_9__7_), .ZN(MULT_mult_6_n2017) );
  INV_X4 MULT_mult_6_U3083 ( .A(MULT_mult_6_ab_6__7_), .ZN(MULT_mult_6_n1313)
         );
  NAND2_X2 MULT_mult_6_U3082 ( .A1(MULT_mult_6_ab_17__7_), .A2(
        MULT_mult_6_CARRYB_16__7_), .ZN(MULT_mult_6_net81265) );
  NAND2_X2 MULT_mult_6_U3081 ( .A1(MULT_mult_6_SUMB_13__8_), .A2(
        MULT_mult_6_ab_14__7_), .ZN(MULT_mult_6_net84999) );
  NOR2_X2 MULT_mult_6_U3080 ( .A1(MULT_mult_6_net77912), .A2(
        MULT_mult_6_net77956), .ZN(MULT_mult_6_ab_4__7_) );
  NOR2_X2 MULT_mult_6_U3079 ( .A1(MULT_mult_6_net77912), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__7_) );
  NOR2_X2 MULT_mult_6_U3078 ( .A1(MULT_mult_6_net77912), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__7_) );
  NOR2_X2 MULT_mult_6_U3077 ( .A1(MULT_mult_6_net77914), .A2(
        MULT_mult_6_net70453), .ZN(MULT_mult_6_ab_21__7_) );
  NOR2_X2 MULT_mult_6_U3076 ( .A1(MULT_mult_6_net77914), .A2(
        MULT_mult_6_net70461), .ZN(MULT_mult_6_ab_17__7_) );
  NOR2_X2 MULT_mult_6_U3075 ( .A1(MULT_mult_6_net77914), .A2(
        MULT_mult_6_net70459), .ZN(MULT_mult_6_ab_18__7_) );
  NOR2_X2 MULT_mult_6_U3074 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__12_) );
  INV_X1 MULT_mult_6_U3073 ( .A(MULT_mult_6_ab_12__12_), .ZN(
        MULT_mult_6_net120586) );
  NAND2_X2 MULT_mult_6_U3072 ( .A1(MULT_mult_6_n1019), .A2(MULT_mult_6_n1020), 
        .ZN(MULT_mult_6_net89026) );
  INV_X2 MULT_mult_6_U3071 ( .A(MULT_mult_6_CARRYB_9__17_), .ZN(
        MULT_mult_6_n1016) );
  INV_X1 MULT_mult_6_U3070 ( .A(MULT_mult_6_ab_10__17_), .ZN(MULT_mult_6_n1015) );
  NAND2_X2 MULT_mult_6_U3069 ( .A1(MULT_mult_6_n1017), .A2(MULT_mult_6_n1018), 
        .ZN(MULT_mult_6_net88226) );
  NAND2_X1 MULT_mult_6_U3068 ( .A1(MULT_mult_6_n1015), .A2(
        MULT_mult_6_CARRYB_9__17_), .ZN(MULT_mult_6_n1018) );
  NAND2_X1 MULT_mult_6_U3067 ( .A1(MULT_mult_6_ab_10__17_), .A2(
        MULT_mult_6_n1016), .ZN(MULT_mult_6_n1017) );
  NAND2_X2 MULT_mult_6_U3066 ( .A1(MULT_mult_6_n1927), .A2(
        MULT_mult_6_ab_2__19_), .ZN(MULT_mult_6_n1526) );
  INV_X2 MULT_mult_6_U3065 ( .A(MULT_mult_6_CARRYB_1__19_), .ZN(
        MULT_mult_6_n1013) );
  NAND2_X4 MULT_mult_6_U3064 ( .A1(MULT_mult_6_n1014), .A2(MULT_mult_6_n2143), 
        .ZN(MULT_mult_6_n1927) );
  NAND2_X4 MULT_mult_6_U3063 ( .A1(MULT_mult_6_n1012), .A2(MULT_mult_6_n1013), 
        .ZN(MULT_mult_6_n1014) );
  NOR2_X2 MULT_mult_6_U3062 ( .A1(MULT_mult_6_net70470), .A2(
        MULT_mult_6_net77964), .ZN(MULT_mult_6_ab_3__18_) );
  NAND2_X2 MULT_mult_6_U3061 ( .A1(MULT_mult_6_CARRYB_1__5_), .A2(
        MULT_mult_6_SUMB_1__6_), .ZN(MULT_mult_6_n1866) );
  INV_X2 MULT_mult_6_U3060 ( .A(MULT_mult_6_net80983), .ZN(
        MULT_mult_6_net120651) );
  NAND2_X2 MULT_mult_6_U3059 ( .A1(MULT_mult_6_net120651), .A2(
        MULT_mult_6_net120652), .ZN(MULT_mult_6_n1011) );
  NAND3_X4 MULT_mult_6_U3058 ( .A1(MULT_mult_6_n1060), .A2(MULT_mult_6_n1061), 
        .A3(MULT_mult_6_n1059), .ZN(MULT_mult_6_CARRYB_14__13_) );
  NAND2_X2 MULT_mult_6_U3057 ( .A1(MULT_mult_6_ab_10__3_), .A2(
        MULT_mult_6_CARRYB_9__3_), .ZN(MULT_mult_6_n1803) );
  XNOR2_X2 MULT_mult_6_U3055 ( .A(MULT_mult_6_n1010), .B(
        MULT_mult_6_CARRYB_14__3_), .ZN(MULT_mult_6_SUMB_15__3_) );
  INV_X4 MULT_mult_6_U3054 ( .A(MULT_mult_6_n1426), .ZN(MULT_mult_6_n1427) );
  NAND2_X2 MULT_mult_6_U3053 ( .A1(MULT_mult_6_ab_20__4_), .A2(
        MULT_mult_6_CARRYB_19__4_), .ZN(MULT_mult_6_n2228) );
  NAND2_X2 MULT_mult_6_U3052 ( .A1(MULT_mult_6_ab_1__19_), .A2(
        MULT_mult_6_ab_0__20_), .ZN(MULT_mult_6_n2339) );
  INV_X4 MULT_mult_6_U3051 ( .A(MULT_mult_6_n2339), .ZN(
        MULT_mult_6_CARRYB_1__19_) );
  INV_X1 MULT_mult_6_U3050 ( .A(MULT_mult_6_ab_18__5_), .ZN(MULT_mult_6_n1006)
         );
  NAND2_X2 MULT_mult_6_U3049 ( .A1(MULT_mult_6_n1007), .A2(MULT_mult_6_n1008), 
        .ZN(MULT_mult_6_n1718) );
  NAND2_X2 MULT_mult_6_U3048 ( .A1(MULT_mult_6_n1005), .A2(MULT_mult_6_n1006), 
        .ZN(MULT_mult_6_n1008) );
  NAND2_X1 MULT_mult_6_U3047 ( .A1(MULT_mult_6_CARRYB_17__5_), .A2(
        MULT_mult_6_ab_18__5_), .ZN(MULT_mult_6_n1007) );
  NAND2_X1 MULT_mult_6_U3046 ( .A1(MULT_mult_6_ab_5__21_), .A2(
        MULT_mult_6_CARRYB_4__21_), .ZN(MULT_mult_6_n1117) );
  NAND2_X1 MULT_mult_6_U3045 ( .A1(MULT_mult_6_CARRYB_9__18_), .A2(
        MULT_mult_6_SUMB_9__19_), .ZN(MULT_mult_6_n1876) );
  XNOR2_X2 MULT_mult_6_U3044 ( .A(MULT_mult_6_ab_2__20_), .B(MULT_mult_6_n2341), .ZN(MULT_mult_6_n1004) );
  NAND3_X4 MULT_mult_6_U3043 ( .A1(MULT_mult_6_net119921), .A2(
        MULT_mult_6_net119920), .A3(MULT_mult_6_n209), .ZN(
        MULT_mult_6_net82031) );
  XNOR2_X2 MULT_mult_6_U3042 ( .A(MULT_mult_6_ab_2__20_), .B(
        MULT_mult_6_CARRYB_1__20_), .ZN(MULT_mult_6_n1424) );
  NOR2_X1 MULT_mult_6_U3041 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__9_) );
  NOR2_X1 MULT_mult_6_U3040 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__9_) );
  INV_X4 MULT_mult_6_U3039 ( .A(MULT_mult_6_n1005), .ZN(MULT_mult_6_n1719) );
  NAND2_X4 MULT_mult_6_U3038 ( .A1(MULT_mult_6_net120628), .A2(
        MULT_mult_6_net120627), .ZN(MULT_mult_6_net83202) );
  NAND3_X4 MULT_mult_6_U3037 ( .A1(MULT_mult_6_n1676), .A2(MULT_mult_6_n1677), 
        .A3(MULT_mult_6_n1678), .ZN(MULT_mult_6_CARRYB_13__3_) );
  NAND3_X2 MULT_mult_6_U3036 ( .A1(MULT_mult_6_n1398), .A2(MULT_mult_6_n1397), 
        .A3(MULT_mult_6_n1396), .ZN(MULT_mult_6_CARRYB_5__9_) );
  CLKBUF_X3 MULT_mult_6_U3035 ( .A(MULT_mult_6_n854), .Z(MULT_mult_6_n1379) );
  INV_X2 MULT_mult_6_U3034 ( .A(MULT_mult_6_CARRYB_8__18_), .ZN(
        MULT_mult_6_n1050) );
  NAND3_X4 MULT_mult_6_U3033 ( .A1(MULT_mult_6_n1793), .A2(MULT_mult_6_n1794), 
        .A3(MULT_mult_6_n1795), .ZN(MULT_mult_6_CARRYB_12__13_) );
  NAND2_X2 MULT_mult_6_U3032 ( .A1(MULT_mult_6_n849), .A2(MULT_mult_6_n215), 
        .ZN(MULT_mult_6_n1387) );
  INV_X4 MULT_mult_6_U3031 ( .A(MULT_mult_6_SUMB_24__6_), .ZN(
        MULT_mult_6_net84304) );
  INV_X8 MULT_mult_6_U3030 ( .A(MULT_mult_6_net84357), .ZN(
        MULT_mult_6_net84358) );
  NOR2_X1 MULT_mult_6_U3029 ( .A1(MULT_mult_6_net77906), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__6_) );
  NAND3_X4 MULT_mult_6_U3028 ( .A1(MULT_mult_6_n1292), .A2(MULT_mult_6_n1293), 
        .A3(MULT_mult_6_n1294), .ZN(MULT_mult_6_CARRYB_9__6_) );
  INV_X4 MULT_mult_6_U3027 ( .A(MULT_mult_6_n1214), .ZN(MULT_mult_6_n1000) );
  NAND2_X4 MULT_mult_6_U3026 ( .A1(MULT_mult_6_n1002), .A2(MULT_mult_6_n1003), 
        .ZN(MULT_mult_6_SUMB_6__8_) );
  NAND2_X4 MULT_mult_6_U3025 ( .A1(MULT_mult_6_n1000), .A2(MULT_mult_6_n1001), 
        .ZN(MULT_mult_6_n1003) );
  NAND2_X2 MULT_mult_6_U3024 ( .A1(MULT_mult_6_n1214), .A2(MULT_mult_6_n1994), 
        .ZN(MULT_mult_6_n1002) );
  NAND3_X2 MULT_mult_6_U3023 ( .A1(MULT_mult_6_n997), .A2(MULT_mult_6_n998), 
        .A3(MULT_mult_6_n999), .ZN(MULT_mult_6_CARRYB_10__6_) );
  NAND2_X1 MULT_mult_6_U3022 ( .A1(MULT_mult_6_ab_10__6_), .A2(
        MULT_mult_6_CARRYB_9__6_), .ZN(MULT_mult_6_n999) );
  NAND2_X2 MULT_mult_6_U3021 ( .A1(MULT_mult_6_ab_10__6_), .A2(
        MULT_mult_6_SUMB_9__7_), .ZN(MULT_mult_6_n998) );
  NAND2_X1 MULT_mult_6_U3020 ( .A1(MULT_mult_6_CARRYB_9__6_), .A2(
        MULT_mult_6_SUMB_9__7_), .ZN(MULT_mult_6_n997) );
  XOR2_X2 MULT_mult_6_U3019 ( .A(MULT_mult_6_CARRYB_9__6_), .B(
        MULT_mult_6_ab_10__6_), .Z(MULT_mult_6_n996) );
  XNOR2_X2 MULT_mult_6_U3018 ( .A(MULT_mult_6_SUMB_22__9_), .B(
        MULT_mult_6_n1273), .ZN(MULT_mult_6_SUMB_23__8_) );
  XNOR2_X1 MULT_mult_6_U3017 ( .A(MULT_mult_6_ab_13__17_), .B(
        MULT_mult_6_CARRYB_12__17_), .ZN(MULT_mult_6_n1571) );
  NAND2_X4 MULT_mult_6_U3016 ( .A1(MULT_mult_6_n994), .A2(MULT_mult_6_n995), 
        .ZN(MULT_mult_6_SUMB_13__17_) );
  NAND2_X4 MULT_mult_6_U3015 ( .A1(MULT_mult_6_n993), .A2(MULT_mult_6_n860), 
        .ZN(MULT_mult_6_n995) );
  NAND2_X2 MULT_mult_6_U3014 ( .A1(MULT_mult_6_SUMB_12__18_), .A2(
        MULT_mult_6_n1571), .ZN(MULT_mult_6_n994) );
  INV_X4 MULT_mult_6_U3013 ( .A(MULT_mult_6_n1089), .ZN(MULT_mult_6_n990) );
  INV_X4 MULT_mult_6_U3012 ( .A(MULT_mult_6_n1088), .ZN(MULT_mult_6_n989) );
  NAND2_X4 MULT_mult_6_U3011 ( .A1(MULT_mult_6_n991), .A2(MULT_mult_6_n992), 
        .ZN(MULT_mult_6_SUMB_4__23_) );
  NAND2_X4 MULT_mult_6_U3010 ( .A1(MULT_mult_6_n989), .A2(MULT_mult_6_n990), 
        .ZN(MULT_mult_6_n992) );
  NAND2_X2 MULT_mult_6_U3009 ( .A1(MULT_mult_6_n1088), .A2(MULT_mult_6_n1089), 
        .ZN(MULT_mult_6_n991) );
  NAND3_X2 MULT_mult_6_U3008 ( .A1(MULT_mult_6_n986), .A2(MULT_mult_6_n987), 
        .A3(MULT_mult_6_n988), .ZN(MULT_mult_6_CARRYB_7__21_) );
  NAND2_X1 MULT_mult_6_U3007 ( .A1(MULT_mult_6_ab_7__21_), .A2(
        MULT_mult_6_CARRYB_6__21_), .ZN(MULT_mult_6_n988) );
  NAND2_X1 MULT_mult_6_U3006 ( .A1(MULT_mult_6_CARRYB_6__21_), .A2(
        MULT_mult_6_SUMB_6__22_), .ZN(MULT_mult_6_n986) );
  NAND2_X2 MULT_mult_6_U3005 ( .A1(MULT_mult_6_CARRYB_11__2_), .A2(
        MULT_mult_6_SUMB_11__3_), .ZN(MULT_mult_6_n1995) );
  XNOR2_X2 MULT_mult_6_U3004 ( .A(MULT_mult_6_n985), .B(
        MULT_mult_6_CARRYB_11__3_), .ZN(MULT_mult_6_SUMB_12__3_) );
  INV_X2 MULT_mult_6_U3003 ( .A(MULT_mult_6_SUMB_2__21_), .ZN(
        MULT_mult_6_n1432) );
  INV_X4 MULT_mult_6_U3002 ( .A(MULT_mult_6_n1692), .ZN(MULT_mult_6_n982) );
  INV_X4 MULT_mult_6_U3001 ( .A(MULT_mult_6_n1828), .ZN(MULT_mult_6_n981) );
  NAND2_X4 MULT_mult_6_U3000 ( .A1(MULT_mult_6_n983), .A2(MULT_mult_6_n984), 
        .ZN(MULT_mult_6_SUMB_2__21_) );
  NAND2_X4 MULT_mult_6_U2999 ( .A1(MULT_mult_6_n981), .A2(MULT_mult_6_n982), 
        .ZN(MULT_mult_6_n984) );
  NAND2_X2 MULT_mult_6_U2998 ( .A1(MULT_mult_6_n57), .A2(MULT_mult_6_n1692), 
        .ZN(MULT_mult_6_n983) );
  NAND3_X2 MULT_mult_6_U2997 ( .A1(MULT_mult_6_n1883), .A2(MULT_mult_6_n1884), 
        .A3(MULT_mult_6_n1885), .ZN(MULT_mult_6_CARRYB_5__20_) );
  NAND2_X2 MULT_mult_6_U2996 ( .A1(MULT_mult_6_n1186), .A2(
        MULT_mult_6_ab_3__14_), .ZN(MULT_mult_6_n1987) );
  NAND2_X1 MULT_mult_6_U2995 ( .A1(MULT_mult_6_SUMB_2__22_), .A2(
        MULT_mult_6_CARRYB_2__21_), .ZN(MULT_mult_6_n1935) );
  NAND2_X2 MULT_mult_6_U2994 ( .A1(MULT_mult_6_SUMB_15__9_), .A2(
        MULT_mult_6_ab_16__8_), .ZN(MULT_mult_6_n2300) );
  NOR2_X2 MULT_mult_6_U2993 ( .A1(MULT_mult_6_net86565), .A2(
        MULT_mult_6_net70491), .ZN(MULT_mult_6_ab_2__19_) );
  NAND3_X2 MULT_mult_6_U2992 ( .A1(MULT_mult_6_n2019), .A2(MULT_mult_6_n2020), 
        .A3(MULT_mult_6_n2021), .ZN(MULT_mult_6_CARRYB_12__7_) );
  NAND2_X4 MULT_mult_6_U2991 ( .A1(MULT_mult_6_n1168), .A2(MULT_mult_6_n1169), 
        .ZN(MULT_mult_6_n1171) );
  NAND2_X2 MULT_mult_6_U2990 ( .A1(MULT_mult_6_CARRYB_9__14_), .A2(
        MULT_mult_6_ab_10__14_), .ZN(MULT_mult_6_n1039) );
  NAND2_X4 MULT_mult_6_U2989 ( .A1(MULT_mult_6_net85540), .A2(
        MULT_mult_6_net88934), .ZN(MULT_mult_6_net85543) );
  INV_X2 MULT_mult_6_U2988 ( .A(MULT_mult_6_net123291), .ZN(
        MULT_mult_6_net121150) );
  NOR2_X4 MULT_mult_6_U2987 ( .A1(MULT_mult_6_net86565), .A2(
        MULT_mult_6_net77940), .ZN(MULT_mult_6_ab_6__19_) );
  INV_X1 MULT_mult_6_U2986 ( .A(MULT_mult_6_ab_6__19_), .ZN(MULT_mult_6_n978)
         );
  INV_X4 MULT_mult_6_U2985 ( .A(MULT_mult_6_CARRYB_5__19_), .ZN(
        MULT_mult_6_n977) );
  NAND2_X2 MULT_mult_6_U2984 ( .A1(MULT_mult_6_n977), .A2(MULT_mult_6_n978), 
        .ZN(MULT_mult_6_n980) );
  NAND3_X4 MULT_mult_6_U2983 ( .A1(MULT_mult_6_n2253), .A2(MULT_mult_6_n2254), 
        .A3(MULT_mult_6_n2252), .ZN(MULT_mult_6_CARRYB_8__15_) );
  NAND2_X4 MULT_mult_6_U2982 ( .A1(MULT_mult_6_net93308), .A2(
        MULT_mult_6_net93309), .ZN(MULT_mult_6_n1125) );
  NAND2_X1 MULT_mult_6_U2981 ( .A1(MULT_mult_6_ab_10__3_), .A2(
        MULT_mult_6_SUMB_9__4_), .ZN(MULT_mult_6_n1802) );
  INV_X8 MULT_mult_6_U2980 ( .A(MULT_mult_6_CARRYB_5__13_), .ZN(
        MULT_mult_6_n1160) );
  INV_X4 MULT_mult_6_U2979 ( .A(MULT_mult_6_SUMB_3__15_), .ZN(MULT_mult_6_n974) );
  INV_X4 MULT_mult_6_U2978 ( .A(MULT_mult_6_n1720), .ZN(MULT_mult_6_n973) );
  NAND2_X4 MULT_mult_6_U2977 ( .A1(MULT_mult_6_n976), .A2(MULT_mult_6_n975), 
        .ZN(MULT_mult_6_SUMB_4__14_) );
  NAND2_X4 MULT_mult_6_U2976 ( .A1(MULT_mult_6_n973), .A2(MULT_mult_6_n974), 
        .ZN(MULT_mult_6_n976) );
  NAND2_X2 MULT_mult_6_U2975 ( .A1(MULT_mult_6_n1720), .A2(
        MULT_mult_6_SUMB_3__15_), .ZN(MULT_mult_6_n975) );
  NAND2_X4 MULT_mult_6_U2974 ( .A1(MULT_mult_6_net84304), .A2(
        MULT_mult_6_net84303), .ZN(MULT_mult_6_n1622) );
  NAND2_X2 MULT_mult_6_U2973 ( .A1(MULT_mult_6_SUMB_11__4_), .A2(
        MULT_mult_6_ab_12__3_), .ZN(MULT_mult_6_n1673) );
  NAND2_X4 MULT_mult_6_U2972 ( .A1(MULT_mult_6_SUMB_12__8_), .A2(
        MULT_mult_6_ab_13__7_), .ZN(MULT_mult_6_n2022) );
  CLKBUF_X3 MULT_mult_6_U2971 ( .A(MULT_mult_6_SUMB_5__16_), .Z(
        MULT_mult_6_n1119) );
  INV_X2 MULT_mult_6_U2970 ( .A(MULT_mult_6_SUMB_6__10_), .ZN(
        MULT_mult_6_n1263) );
  NAND2_X2 MULT_mult_6_U2969 ( .A1(MULT_mult_6_n67), .A2(
        MULT_mult_6_SUMB_6__10_), .ZN(MULT_mult_6_n2003) );
  INV_X4 MULT_mult_6_U2968 ( .A(MULT_mult_6_ab_2__12_), .ZN(
        MULT_mult_6_net120174) );
  NAND2_X4 MULT_mult_6_U2967 ( .A1(MULT_mult_6_n1177), .A2(MULT_mult_6_n1178), 
        .ZN(MULT_mult_6_n1180) );
  NAND2_X4 MULT_mult_6_U2966 ( .A1(MULT_mult_6_n1180), .A2(MULT_mult_6_n1179), 
        .ZN(MULT_mult_6_n2015) );
  NAND2_X4 MULT_mult_6_U2965 ( .A1(MULT_mult_6_net88156), .A2(
        MULT_mult_6_net88157), .ZN(MULT_mult_6_n1321) );
  NAND2_X2 MULT_mult_6_U2964 ( .A1(MULT_mult_6_n1261), .A2(
        MULT_mult_6_CARRYB_8__7_), .ZN(MULT_mult_6_n2016) );
  NAND2_X4 MULT_mult_6_U2963 ( .A1(MULT_mult_6_net120174), .A2(
        MULT_mult_6_n1044), .ZN(MULT_mult_6_n1046) );
  NAND2_X4 MULT_mult_6_U2962 ( .A1(MULT_mult_6_n1045), .A2(MULT_mult_6_n1046), 
        .ZN(MULT_mult_6_n1504) );
  NOR2_X1 MULT_mult_6_U2961 ( .A1(MULT_mult_6_net77866), .A2(
        MULT_mult_6_net77924), .ZN(MULT_mult_6_ab_8__1_) );
  NOR2_X1 MULT_mult_6_U2960 ( .A1(MULT_mult_6_net77866), .A2(
        MULT_mult_6_net77930), .ZN(MULT_mult_6_ab_7__1_) );
  NAND3_X2 MULT_mult_6_U2959 ( .A1(MULT_mult_6_n969), .A2(MULT_mult_6_n970), 
        .A3(MULT_mult_6_n971), .ZN(MULT_mult_6_CARRYB_8__1_) );
  NAND2_X1 MULT_mult_6_U2958 ( .A1(MULT_mult_6_ab_8__1_), .A2(
        MULT_mult_6_CARRYB_7__1_), .ZN(MULT_mult_6_n971) );
  NAND2_X2 MULT_mult_6_U2957 ( .A1(MULT_mult_6_ab_8__1_), .A2(
        MULT_mult_6_SUMB_7__2_), .ZN(MULT_mult_6_n970) );
  NAND2_X1 MULT_mult_6_U2956 ( .A1(MULT_mult_6_CARRYB_7__1_), .A2(
        MULT_mult_6_SUMB_7__2_), .ZN(MULT_mult_6_n969) );
  XOR2_X2 MULT_mult_6_U2955 ( .A(MULT_mult_6_SUMB_7__2_), .B(MULT_mult_6_n968), 
        .Z(MULT_mult_6_SUMB_8__1_) );
  XOR2_X2 MULT_mult_6_U2954 ( .A(MULT_mult_6_CARRYB_7__1_), .B(
        MULT_mult_6_ab_8__1_), .Z(MULT_mult_6_n968) );
  NAND3_X2 MULT_mult_6_U2953 ( .A1(MULT_mult_6_n965), .A2(MULT_mult_6_n966), 
        .A3(MULT_mult_6_n967), .ZN(MULT_mult_6_CARRYB_7__1_) );
  NAND2_X1 MULT_mult_6_U2952 ( .A1(MULT_mult_6_ab_7__1_), .A2(
        MULT_mult_6_CARRYB_6__1_), .ZN(MULT_mult_6_n967) );
  NAND2_X2 MULT_mult_6_U2951 ( .A1(MULT_mult_6_ab_7__1_), .A2(
        MULT_mult_6_SUMB_6__2_), .ZN(MULT_mult_6_n966) );
  NAND2_X2 MULT_mult_6_U2950 ( .A1(MULT_mult_6_CARRYB_6__1_), .A2(
        MULT_mult_6_SUMB_6__2_), .ZN(MULT_mult_6_n965) );
  XOR2_X1 MULT_mult_6_U2949 ( .A(MULT_mult_6_SUMB_6__2_), .B(MULT_mult_6_n964), 
        .Z(MULT_mult_6_SUMB_7__1_) );
  XOR2_X2 MULT_mult_6_U2948 ( .A(MULT_mult_6_CARRYB_6__1_), .B(
        MULT_mult_6_ab_7__1_), .Z(MULT_mult_6_n964) );
  NAND3_X4 MULT_mult_6_U2947 ( .A1(MULT_mult_6_net80255), .A2(
        MULT_mult_6_net80254), .A3(MULT_mult_6_n2295), .ZN(
        MULT_mult_6_CARRYB_23__2_) );
  NAND2_X1 MULT_mult_6_U2946 ( .A1(MULT_mult_6_ab_18__11_), .A2(
        MULT_mult_6_net88647), .ZN(MULT_mult_6_net82665) );
  NOR2_X2 MULT_mult_6_U2945 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net70461), .ZN(MULT_mult_6_ab_17__12_) );
  XNOR2_X1 MULT_mult_6_U2944 ( .A(MULT_mult_6_net90525), .B(
        MULT_mult_6_net81290), .ZN(MULT_mult_6_net90103) );
  NAND2_X2 MULT_mult_6_U2943 ( .A1(MULT_mult_6_ab_14__14_), .A2(
        MULT_mult_6_SUMB_13__15_), .ZN(MULT_mult_6_net80479) );
  NOR2_X2 MULT_mult_6_U2942 ( .A1(MULT_mult_6_net80643), .A2(
        MULT_mult_6_net77948), .ZN(MULT_mult_6_ab_5__21_) );
  XOR2_X2 MULT_mult_6_U2941 ( .A(MULT_mult_6_net90103), .B(MULT_mult_6_n961), 
        .Z(MULT_mult_6_net88647) );
  XOR2_X2 MULT_mult_6_U2940 ( .A(MULT_mult_6_CARRYB_16__12_), .B(
        MULT_mult_6_ab_17__12_), .Z(MULT_mult_6_n961) );
  INV_X2 MULT_mult_6_U2939 ( .A(MULT_mult_6_ab_5__21_), .ZN(MULT_mult_6_n958)
         );
  INV_X4 MULT_mult_6_U2938 ( .A(MULT_mult_6_CARRYB_4__21_), .ZN(
        MULT_mult_6_n957) );
  NAND2_X2 MULT_mult_6_U2937 ( .A1(MULT_mult_6_n959), .A2(MULT_mult_6_n960), 
        .ZN(MULT_mult_6_n1435) );
  NAND2_X1 MULT_mult_6_U2936 ( .A1(MULT_mult_6_CARRYB_4__21_), .A2(
        MULT_mult_6_ab_5__21_), .ZN(MULT_mult_6_n959) );
  NAND2_X4 MULT_mult_6_U2935 ( .A1(MULT_mult_6_net121455), .A2(
        MULT_mult_6_n956), .ZN(MULT_mult_6_net90731) );
  NAND2_X4 MULT_mult_6_U2934 ( .A1(MULT_mult_6_net121453), .A2(
        MULT_mult_6_net121454), .ZN(MULT_mult_6_n956) );
  INV_X8 MULT_mult_6_U2933 ( .A(n10914), .ZN(MULT_mult_6_net70476) );
  INV_X2 MULT_mult_6_U2932 ( .A(MULT_mult_6_net70476), .ZN(MULT_mult_6_n1118)
         );
  NAND2_X2 MULT_mult_6_U2931 ( .A1(MULT_mult_6_SUMB_23__1_), .A2(
        MULT_mult_6_ab_24__0_), .ZN(MULT_mult_6_n1570) );
  NAND2_X4 MULT_mult_6_U2930 ( .A1(MULT_mult_6_ab_18__5_), .A2(
        MULT_mult_6_n1719), .ZN(MULT_mult_6_n2231) );
  NAND2_X2 MULT_mult_6_U2929 ( .A1(MULT_mult_6_ab_18__0_), .A2(
        MULT_mult_6_SUMB_17__1_), .ZN(MULT_mult_6_n1810) );
  NAND2_X2 MULT_mult_6_U2928 ( .A1(MULT_mult_6_CARRYB_12__7_), .A2(
        MULT_mult_6_ab_13__7_), .ZN(MULT_mult_6_n2023) );
  BUF_X8 MULT_mult_6_U2927 ( .A(MULT_mult_6_CARRYB_12__7_), .Z(
        MULT_mult_6_n1588) );
  NAND2_X2 MULT_mult_6_U2926 ( .A1(MULT_mult_6_CARRYB_3__9_), .A2(
        MULT_mult_6_ab_4__9_), .ZN(MULT_mult_6_n1961) );
  NAND2_X4 MULT_mult_6_U2925 ( .A1(MULT_mult_6_SUMB_1__20_), .A2(
        MULT_mult_6_CARRYB_1__19_), .ZN(MULT_mult_6_n2143) );
  INV_X8 MULT_mult_6_U2924 ( .A(MULT_mult_6_CARRYB_14__12_), .ZN(
        MULT_mult_6_n1850) );
  XNOR2_X2 MULT_mult_6_U2923 ( .A(MULT_mult_6_n1742), .B(MULT_mult_6_n852), 
        .ZN(MULT_mult_6_n1242) );
  INV_X4 MULT_mult_6_U2922 ( .A(MULT_mult_6_net125375), .ZN(
        MULT_mult_6_net121607) );
  NAND2_X4 MULT_mult_6_U2921 ( .A1(MULT_mult_6_n953), .A2(MULT_mult_6_n954), 
        .ZN(MULT_mult_6_SUMB_9__10_) );
  NAND2_X4 MULT_mult_6_U2920 ( .A1(MULT_mult_6_net121606), .A2(
        MULT_mult_6_net121607), .ZN(MULT_mult_6_n954) );
  NAND2_X2 MULT_mult_6_U2919 ( .A1(MULT_mult_6_net83736), .A2(
        MULT_mult_6_net125375), .ZN(MULT_mult_6_n953) );
  NAND2_X2 MULT_mult_6_U2918 ( .A1(MULT_mult_6_ab_6__13_), .A2(
        MULT_mult_6_CARRYB_5__13_), .ZN(MULT_mult_6_n1161) );
  NAND2_X1 MULT_mult_6_U2917 ( .A1(MULT_mult_6_CARRYB_3__18_), .A2(
        MULT_mult_6_SUMB_3__19_), .ZN(MULT_mult_6_n1722) );
  NAND2_X1 MULT_mult_6_U2916 ( .A1(MULT_mult_6_n1187), .A2(
        MULT_mult_6_CARRYB_15__11_), .ZN(MULT_mult_6_n2098) );
  INV_X4 MULT_mult_6_U2915 ( .A(MULT_mult_6_ab_16__8_), .ZN(MULT_mult_6_n2153)
         );
  XNOR2_X2 MULT_mult_6_U2914 ( .A(MULT_mult_6_ab_16__8_), .B(
        MULT_mult_6_CARRYB_15__8_), .ZN(MULT_mult_6_n952) );
  NOR2_X2 MULT_mult_6_U2913 ( .A1(MULT_mult_6_net82890), .A2(
        MULT_mult_6_net77956), .ZN(MULT_mult_6_ab_4__17_) );
  XOR2_X2 MULT_mult_6_U2912 ( .A(MULT_mult_6_CARRYB_17__13_), .B(
        MULT_mult_6_ab_18__13_), .Z(MULT_mult_6_n951) );
  NAND2_X2 MULT_mult_6_U2911 ( .A1(MULT_mult_6_ab_16__5_), .A2(
        MULT_mult_6_SUMB_15__6_), .ZN(MULT_mult_6_n2072) );
  XNOR2_X2 MULT_mult_6_U2910 ( .A(MULT_mult_6_n2362), .B(MULT_mult_6_n1325), 
        .ZN(MULT_mult_6_n950) );
  XNOR2_X2 MULT_mult_6_U2909 ( .A(MULT_mult_6_n856), .B(MULT_mult_6_n1095), 
        .ZN(MULT_mult_6_n949) );
  INV_X2 MULT_mult_6_U2908 ( .A(MULT_mult_6_SUMB_3__9_), .ZN(MULT_mult_6_n947)
         );
  NAND3_X4 MULT_mult_6_U2907 ( .A1(MULT_mult_6_n2117), .A2(
        MULT_mult_6_net81060), .A3(MULT_mult_6_net81059), .ZN(
        MULT_mult_6_net85043) );
  INV_X4 MULT_mult_6_U2906 ( .A(MULT_mult_6_n66), .ZN(MULT_mult_6_n1341) );
  XNOR2_X2 MULT_mult_6_U2905 ( .A(MULT_mult_6_CARRYB_20__4_), .B(
        MULT_mult_6_n945), .ZN(MULT_mult_6_n944) );
  INV_X4 MULT_mult_6_U2904 ( .A(MULT_mult_6_ab_4__14_), .ZN(
        MULT_mult_6_net92716) );
  NOR2_X2 MULT_mult_6_U2903 ( .A1(MULT_mult_6_net84698), .A2(
        MULT_mult_6_net77964), .ZN(MULT_mult_6_ab_3__14_) );
  NAND3_X2 MULT_mult_6_U2902 ( .A1(MULT_mult_6_n1962), .A2(MULT_mult_6_n1961), 
        .A3(MULT_mult_6_n1963), .ZN(MULT_mult_6_n943) );
  XNOR2_X2 MULT_mult_6_U2901 ( .A(MULT_mult_6_n942), .B(
        MULT_mult_6_SUMB_13__4_), .ZN(MULT_mult_6_SUMB_14__3_) );
  CLKBUF_X2 MULT_mult_6_U2900 ( .A(MULT_mult_6_SUMB_8__5_), .Z(
        MULT_mult_6_net121926) );
  NAND2_X1 MULT_mult_6_U2899 ( .A1(MULT_mult_6_ab_15__0_), .A2(
        MULT_mult_6_SUMB_14__1_), .ZN(MULT_mult_6_n1411) );
  NAND2_X2 MULT_mult_6_U2898 ( .A1(MULT_mult_6_n682), .A2(MULT_mult_6_n390), 
        .ZN(MULT_mult_6_n1579) );
  INV_X4 MULT_mult_6_U2897 ( .A(MULT_mult_6_CARRYB_17__5_), .ZN(
        MULT_mult_6_n1005) );
  XNOR2_X2 MULT_mult_6_U2896 ( .A(MULT_mult_6_net124874), .B(
        MULT_mult_6_SUMB_24__2_), .ZN(MULT_mult_6_n940) );
  NAND3_X2 MULT_mult_6_U2895 ( .A1(MULT_mult_6_n1822), .A2(MULT_mult_6_n1823), 
        .A3(MULT_mult_6_n1824), .ZN(MULT_mult_6_CARRYB_7__7_) );
  XNOR2_X2 MULT_mult_6_U2894 ( .A(MULT_mult_6_n1820), .B(MULT_mult_6_n1264), 
        .ZN(MULT_mult_6_n939) );
  XNOR2_X2 MULT_mult_6_U2893 ( .A(MULT_mult_6_n1820), .B(MULT_mult_6_n1264), 
        .ZN(MULT_mult_6_n938) );
  NAND2_X4 MULT_mult_6_U2892 ( .A1(MULT_mult_6_SUMB_23__6_), .A2(
        MULT_mult_6_n2148), .ZN(MULT_mult_6_n1121) );
  NOR2_X1 MULT_mult_6_U2891 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net70455), .ZN(MULT_mult_6_ab_20__9_) );
  NAND2_X4 MULT_mult_6_U2890 ( .A1(MULT_mult_6_net87133), .A2(
        MULT_mult_6_net87134), .ZN(MULT_mult_6_net87136) );
  INV_X4 MULT_mult_6_U2889 ( .A(MULT_mult_6_CARRYB_18__9_), .ZN(
        MULT_mult_6_net87134) );
  INV_X1 MULT_mult_6_U2888 ( .A(MULT_mult_6_net87134), .ZN(
        MULT_mult_6_net90802) );
  NAND2_X2 MULT_mult_6_U2887 ( .A1(MULT_mult_6_net90802), .A2(MULT_mult_6_n936), .ZN(MULT_mult_6_net81954) );
  XNOR2_X2 MULT_mult_6_U2886 ( .A(MULT_mult_6_net85979), .B(MULT_mult_6_n936), 
        .ZN(MULT_mult_6_net89289) );
  XNOR2_X2 MULT_mult_6_U2885 ( .A(MULT_mult_6_net85979), .B(MULT_mult_6_n936), 
        .ZN(MULT_mult_6_SUMB_19__9_) );
  NAND2_X2 MULT_mult_6_U2884 ( .A1(MULT_mult_6_n936), .A2(
        MULT_mult_6_ab_19__9_), .ZN(MULT_mult_6_net81953) );
  BUF_X8 MULT_mult_6_U2883 ( .A(MULT_mult_6_CARRYB_19__9_), .Z(
        MULT_mult_6_net82255) );
  XNOR2_X2 MULT_mult_6_U2882 ( .A(MULT_mult_6_CARRYB_18__10_), .B(
        MULT_mult_6_ab_19__10_), .ZN(MULT_mult_6_n934) );
  NAND2_X1 MULT_mult_6_U2881 ( .A1(MULT_mult_6_ab_20__9_), .A2(
        MULT_mult_6_SUMB_19__10_), .ZN(MULT_mult_6_net81034) );
  XNOR2_X2 MULT_mult_6_U2880 ( .A(MULT_mult_6_SUMB_18__11_), .B(
        MULT_mult_6_n934), .ZN(MULT_mult_6_SUMB_19__10_) );
  INV_X1 MULT_mult_6_U2879 ( .A(MULT_mult_6_ab_20__9_), .ZN(
        MULT_mult_6_net86403) );
  INV_X4 MULT_mult_6_U2878 ( .A(MULT_mult_6_CARRYB_19__9_), .ZN(
        MULT_mult_6_net86404) );
  NAND2_X2 MULT_mult_6_U2877 ( .A1(MULT_mult_6_net86403), .A2(
        MULT_mult_6_net86404), .ZN(MULT_mult_6_n937) );
  XNOR2_X2 MULT_mult_6_U2876 ( .A(MULT_mult_6_net82396), .B(
        MULT_mult_6_SUMB_19__10_), .ZN(MULT_mult_6_SUMB_20__9_) );
  XNOR2_X2 MULT_mult_6_U2875 ( .A(MULT_mult_6_net86557), .B(
        MULT_mult_6_SUMB_5__20_), .ZN(MULT_mult_6_SUMB_6__19_) );
  INV_X1 MULT_mult_6_U2874 ( .A(MULT_mult_6_ab_7__18_), .ZN(
        MULT_mult_6_net80657) );
  INV_X4 MULT_mult_6_U2873 ( .A(MULT_mult_6_CARRYB_6__18_), .ZN(
        MULT_mult_6_net80658) );
  NAND2_X2 MULT_mult_6_U2872 ( .A1(MULT_mult_6_ab_7__17_), .A2(
        MULT_mult_6_net90702), .ZN(MULT_mult_6_n931) );
  NAND2_X1 MULT_mult_6_U2871 ( .A1(MULT_mult_6_ab_7__17_), .A2(
        MULT_mult_6_CARRYB_6__17_), .ZN(MULT_mult_6_n930) );
  NAND3_X2 MULT_mult_6_U2870 ( .A1(MULT_mult_6_n931), .A2(MULT_mult_6_n932), 
        .A3(MULT_mult_6_n930), .ZN(MULT_mult_6_CARRYB_7__17_) );
  XNOR2_X2 MULT_mult_6_U2869 ( .A(MULT_mult_6_n921), .B(MULT_mult_6_net81945), 
        .ZN(MULT_mult_6_SUMB_10__16_) );
  CLKBUF_X3 MULT_mult_6_U2868 ( .A(MULT_mult_6_n922), .Z(MULT_mult_6_n929) );
  INV_X2 MULT_mult_6_U2867 ( .A(MULT_mult_6_net123072), .ZN(
        MULT_mult_6_net82890) );
  XNOR2_X2 MULT_mult_6_U2866 ( .A(MULT_mult_6_n922), .B(MULT_mult_6_net123019), 
        .ZN(MULT_mult_6_n926) );
  INV_X4 MULT_mult_6_U2865 ( .A(MULT_mult_6_n924), .ZN(MULT_mult_6_n921) );
  INV_X4 MULT_mult_6_U2864 ( .A(MULT_mult_6_n923), .ZN(MULT_mult_6_n920) );
  INV_X4 MULT_mult_6_U2863 ( .A(MULT_mult_6_net123055), .ZN(
        MULT_mult_6_net123028) );
  OAI21_X4 MULT_mult_6_U2862 ( .B1(MULT_mult_6_n929), .B2(
        MULT_mult_6_net123062), .A(MULT_mult_6_CARRYB_7__17_), .ZN(
        MULT_mult_6_n919) );
  INV_X4 MULT_mult_6_U2861 ( .A(MULT_mult_6_net123019), .ZN(
        MULT_mult_6_net123062) );
  XNOR2_X2 MULT_mult_6_U2860 ( .A(MULT_mult_6_n923), .B(MULT_mult_6_n925), 
        .ZN(MULT_mult_6_n924) );
  XNOR2_X2 MULT_mult_6_U2859 ( .A(MULT_mult_6_SUMB_7__19_), .B(
        MULT_mult_6_net79939), .ZN(MULT_mult_6_n923) );
  XNOR2_X2 MULT_mult_6_U2858 ( .A(MULT_mult_6_net80366), .B(
        MULT_mult_6_SUMB_6__19_), .ZN(MULT_mult_6_n922) );
  NAND2_X2 MULT_mult_6_U2857 ( .A1(MULT_mult_6_n921), .A2(
        MULT_mult_6_CARRYB_9__16_), .ZN(MULT_mult_6_net80806) );
  NAND2_X2 MULT_mult_6_U2856 ( .A1(MULT_mult_6_n921), .A2(
        MULT_mult_6_ab_10__16_), .ZN(MULT_mult_6_net80805) );
  NAND2_X2 MULT_mult_6_U2855 ( .A1(MULT_mult_6_n920), .A2(
        MULT_mult_6_net123028), .ZN(MULT_mult_6_net80802) );
  NAND2_X2 MULT_mult_6_U2854 ( .A1(MULT_mult_6_n917), .A2(MULT_mult_6_n920), 
        .ZN(MULT_mult_6_net80803) );
  NAND2_X2 MULT_mult_6_U2853 ( .A1(MULT_mult_6_n917), .A2(
        MULT_mult_6_net123028), .ZN(MULT_mult_6_net80801) );
  OAI21_X4 MULT_mult_6_U2852 ( .B1(MULT_mult_6_n918), .B2(
        MULT_mult_6_net123019), .A(MULT_mult_6_n919), .ZN(MULT_mult_6_n917) );
  INV_X4 MULT_mult_6_U2851 ( .A(MULT_mult_6_CARRYB_2__18_), .ZN(
        MULT_mult_6_n1547) );
  NAND2_X4 MULT_mult_6_U2850 ( .A1(MULT_mult_6_CARRYB_4__12_), .A2(
        MULT_mult_6_ab_5__12_), .ZN(MULT_mult_6_net81204) );
  XNOR2_X2 MULT_mult_6_U2849 ( .A(MULT_mult_6_CARRYB_22__2_), .B(
        MULT_mult_6_ab_23__2_), .ZN(MULT_mult_6_net121523) );
  INV_X8 MULT_mult_6_U2848 ( .A(MULT_mult_6_net81815), .ZN(
        MULT_mult_6_net84303) );
  NAND2_X4 MULT_mult_6_U2847 ( .A1(MULT_mult_6_n1162), .A2(MULT_mult_6_n1161), 
        .ZN(MULT_mult_6_n1942) );
  NAND2_X2 MULT_mult_6_U2846 ( .A1(MULT_mult_6_ab_1__20_), .A2(
        MULT_mult_6_ab_0__21_), .ZN(MULT_mult_6_n2341) );
  NAND2_X4 MULT_mult_6_U2845 ( .A1(MULT_mult_6_n2374), .A2(
        MULT_mult_6_ab_6__10_), .ZN(MULT_mult_6_n1590) );
  INV_X2 MULT_mult_6_U2844 ( .A(MULT_mult_6_ab_3__11_), .ZN(MULT_mult_6_n914)
         );
  NAND2_X4 MULT_mult_6_U2843 ( .A1(MULT_mult_6_n913), .A2(MULT_mult_6_n914), 
        .ZN(MULT_mult_6_n916) );
  NAND2_X2 MULT_mult_6_U2842 ( .A1(MULT_mult_6_CARRYB_2__11_), .A2(
        MULT_mult_6_ab_3__11_), .ZN(MULT_mult_6_n915) );
  NAND2_X4 MULT_mult_6_U2841 ( .A1(MULT_mult_6_ab_0__12_), .A2(
        MULT_mult_6_ab_1__11_), .ZN(MULT_mult_6_n2334) );
  NAND2_X4 MULT_mult_6_U2840 ( .A1(MULT_mult_6_n1417), .A2(MULT_mult_6_n1418), 
        .ZN(MULT_mult_6_net82089) );
  NAND2_X4 MULT_mult_6_U2839 ( .A1(MULT_mult_6_n911), .A2(MULT_mult_6_n912), 
        .ZN(MULT_mult_6_SUMB_4__13_) );
  INV_X8 MULT_mult_6_U2838 ( .A(MULT_mult_6_n907), .ZN(MULT_mult_6_n908) );
  INV_X2 MULT_mult_6_U2837 ( .A(MULT_mult_6_SUMB_4__26_), .ZN(MULT_mult_6_n907) );
  NAND3_X4 MULT_mult_6_U2836 ( .A1(MULT_mult_6_n904), .A2(MULT_mult_6_n905), 
        .A3(MULT_mult_6_n906), .ZN(MULT_mult_6_CARRYB_6__24_) );
  NAND2_X1 MULT_mult_6_U2835 ( .A1(MULT_mult_6_CARRYB_5__24_), .A2(
        MULT_mult_6_SUMB_5__25_), .ZN(MULT_mult_6_n906) );
  NAND2_X1 MULT_mult_6_U2834 ( .A1(MULT_mult_6_ab_6__24_), .A2(
        MULT_mult_6_CARRYB_5__24_), .ZN(MULT_mult_6_n904) );
  NAND3_X4 MULT_mult_6_U2833 ( .A1(MULT_mult_6_n901), .A2(MULT_mult_6_n902), 
        .A3(MULT_mult_6_n903), .ZN(MULT_mult_6_CARRYB_5__25_) );
  NAND2_X2 MULT_mult_6_U2832 ( .A1(MULT_mult_6_CARRYB_4__25_), .A2(
        MULT_mult_6_n908), .ZN(MULT_mult_6_n903) );
  NAND2_X2 MULT_mult_6_U2831 ( .A1(MULT_mult_6_ab_5__25_), .A2(
        MULT_mult_6_n908), .ZN(MULT_mult_6_n902) );
  NAND2_X1 MULT_mult_6_U2830 ( .A1(MULT_mult_6_ab_5__25_), .A2(
        MULT_mult_6_CARRYB_4__25_), .ZN(MULT_mult_6_n901) );
  XOR2_X2 MULT_mult_6_U2829 ( .A(MULT_mult_6_n900), .B(MULT_mult_6_SUMB_5__25_), .Z(MULT_mult_6_SUMB_6__24_) );
  XOR2_X2 MULT_mult_6_U2828 ( .A(MULT_mult_6_ab_6__24_), .B(
        MULT_mult_6_CARRYB_5__24_), .Z(MULT_mult_6_n900) );
  XOR2_X2 MULT_mult_6_U2827 ( .A(MULT_mult_6_n899), .B(MULT_mult_6_n908), .Z(
        MULT_mult_6_SUMB_5__25_) );
  XOR2_X2 MULT_mult_6_U2826 ( .A(MULT_mult_6_ab_5__25_), .B(
        MULT_mult_6_CARRYB_4__25_), .Z(MULT_mult_6_n899) );
  INV_X8 MULT_mult_6_U2825 ( .A(MULT_mult_6_CARRYB_1__12_), .ZN(
        MULT_mult_6_n1044) );
  XNOR2_X2 MULT_mult_6_U2824 ( .A(MULT_mult_6_ab_13__15_), .B(
        MULT_mult_6_CARRYB_12__15_), .ZN(MULT_mult_6_n898) );
  XNOR2_X2 MULT_mult_6_U2823 ( .A(MULT_mult_6_n898), .B(
        MULT_mult_6_SUMB_12__16_), .ZN(MULT_mult_6_SUMB_13__15_) );
  XNOR2_X2 MULT_mult_6_U2822 ( .A(MULT_mult_6_CARRYB_17__10_), .B(
        MULT_mult_6_n897), .ZN(MULT_mult_6_net87009) );
  NAND2_X4 MULT_mult_6_U2821 ( .A1(MULT_mult_6_n2155), .A2(
        MULT_mult_6_ab_24__5_), .ZN(MULT_mult_6_n2157) );
  NAND2_X4 MULT_mult_6_U2820 ( .A1(MULT_mult_6_n1290), .A2(MULT_mult_6_n1291), 
        .ZN(MULT_mult_6_n1773) );
  NAND2_X4 MULT_mult_6_U2819 ( .A1(MULT_mult_6_n1346), .A2(MULT_mult_6_n1347), 
        .ZN(MULT_mult_6_n1349) );
  INV_X2 MULT_mult_6_U2818 ( .A(MULT_mult_6_SUMB_4__14_), .ZN(
        MULT_mult_6_n1356) );
  XNOR2_X2 MULT_mult_6_U2817 ( .A(MULT_mult_6_ab_21__1_), .B(
        MULT_mult_6_SUMB_20__2_), .ZN(MULT_mult_6_n1266) );
  NAND2_X4 MULT_mult_6_U2816 ( .A1(MULT_mult_6_SUMB_1__13_), .A2(
        MULT_mult_6_n588), .ZN(MULT_mult_6_n2081) );
  INV_X4 MULT_mult_6_U2815 ( .A(MULT_mult_6_net88449), .ZN(
        MULT_mult_6_net123428) );
  CLKBUF_X3 MULT_mult_6_U2814 ( .A(MULT_mult_6_CARRYB_3__20_), .Z(
        MULT_mult_6_n1009) );
  INV_X2 MULT_mult_6_U2813 ( .A(MULT_mult_6_ab_1__11_), .ZN(MULT_mult_6_n1023)
         );
  NAND3_X4 MULT_mult_6_U2812 ( .A1(MULT_mult_6_n1085), .A2(MULT_mult_6_n1086), 
        .A3(MULT_mult_6_n1087), .ZN(MULT_mult_6_CARRYB_16__12_) );
  NAND2_X1 MULT_mult_6_U2810 ( .A1(MULT_mult_6_ab_17__12_), .A2(
        MULT_mult_6_CARRYB_16__12_), .ZN(MULT_mult_6_n894) );
  XOR2_X2 MULT_mult_6_U2809 ( .A(MULT_mult_6_SUMB_16__13_), .B(
        MULT_mult_6_n891), .Z(MULT_mult_6_SUMB_17__12_) );
  XOR2_X2 MULT_mult_6_U2808 ( .A(MULT_mult_6_CARRYB_16__12_), .B(
        MULT_mult_6_ab_17__12_), .Z(MULT_mult_6_n891) );
  INV_X2 MULT_mult_6_U2807 ( .A(MULT_mult_6_SUMB_12__18_), .ZN(
        MULT_mult_6_n993) );
  NAND3_X2 MULT_mult_6_U2806 ( .A1(MULT_mult_6_n1466), .A2(MULT_mult_6_n1467), 
        .A3(MULT_mult_6_n1468), .ZN(MULT_mult_6_CARRYB_12__17_) );
  NAND2_X2 MULT_mult_6_U2805 ( .A1(MULT_mult_6_ab_6__20_), .A2(
        MULT_mult_6_SUMB_5__21_), .ZN(MULT_mult_6_net79936) );
  NAND2_X2 MULT_mult_6_U2804 ( .A1(MULT_mult_6_ab_4__17_), .A2(
        MULT_mult_6_n861), .ZN(MULT_mult_6_n1893) );
  NAND2_X1 MULT_mult_6_U2803 ( .A1(MULT_mult_6_ab_6__24_), .A2(
        MULT_mult_6_SUMB_5__25_), .ZN(MULT_mult_6_n905) );
  NAND2_X1 MULT_mult_6_U2802 ( .A1(MULT_mult_6_ab_1__23_), .A2(
        MULT_mult_6_ab_0__24_), .ZN(MULT_mult_6_net82045) );
  NOR2_X1 MULT_mult_6_U2801 ( .A1(MULT_mult_6_net77930), .A2(
        MULT_mult_6_net70482), .ZN(MULT_mult_6_ab_7__24_) );
  NOR2_X1 MULT_mult_6_U2800 ( .A1(MULT_mult_6_net70482), .A2(
        MULT_mult_6_net77940), .ZN(MULT_mult_6_ab_6__24_) );
  NOR2_X1 MULT_mult_6_U2799 ( .A1(MULT_mult_6_net70482), .A2(
        MULT_mult_6_net77948), .ZN(MULT_mult_6_ab_5__24_) );
  NOR2_X1 MULT_mult_6_U2798 ( .A1(MULT_mult_6_net70482), .A2(
        MULT_mult_6_net77956), .ZN(MULT_mult_6_ab_4__24_) );
  INV_X1 MULT_mult_6_U2797 ( .A(MULT_mult_6_ab_4__10_), .ZN(MULT_mult_6_n889)
         );
  NAND2_X4 MULT_mult_6_U2796 ( .A1(MULT_mult_6_n887), .A2(MULT_mult_6_n886), 
        .ZN(MULT_mult_6_SUMB_2__12_) );
  NAND2_X2 MULT_mult_6_U2795 ( .A1(MULT_mult_6_CARRYB_1__12_), .A2(
        MULT_mult_6_ab_2__12_), .ZN(MULT_mult_6_n2082) );
  NAND3_X2 MULT_mult_6_U2794 ( .A1(MULT_mult_6_net81954), .A2(
        MULT_mult_6_net81953), .A3(MULT_mult_6_n935), .ZN(
        MULT_mult_6_CARRYB_19__9_) );
  NAND2_X4 MULT_mult_6_U2793 ( .A1(MULT_mult_6_net80801), .A2(MULT_mult_6_n928), .ZN(MULT_mult_6_n925) );
  NAND3_X2 MULT_mult_6_U2792 ( .A1(MULT_mult_6_net80803), .A2(
        MULT_mult_6_net80802), .A3(MULT_mult_6_net80801), .ZN(
        MULT_mult_6_CARRYB_9__17_) );
  INV_X4 MULT_mult_6_U2791 ( .A(MULT_mult_6_net80517), .ZN(
        MULT_mult_6_net86407) );
  NAND3_X2 MULT_mult_6_U2790 ( .A1(MULT_mult_6_net82664), .A2(
        MULT_mult_6_net82665), .A3(MULT_mult_6_net82666), .ZN(
        MULT_mult_6_CARRYB_18__11_) );
  NOR2_X4 MULT_mult_6_U2789 ( .A1(MULT_mult_6_net124610), .A2(
        MULT_mult_6_net70486), .ZN(MULT_mult_6_ab_0__26_) );
  NAND2_X2 MULT_mult_6_U2788 ( .A1(MULT_mult_6_CARRYB_2__4_), .A2(
        MULT_mult_6_SUMB_2__5_), .ZN(MULT_mult_6_n1147) );
  NAND2_X2 MULT_mult_6_U2787 ( .A1(MULT_mult_6_ab_15__6_), .A2(
        MULT_mult_6_SUMB_14__7_), .ZN(MULT_mult_6_n1437) );
  XNOR2_X2 MULT_mult_6_U2786 ( .A(MULT_mult_6_CARRYB_6__6_), .B(
        MULT_mult_6_ab_7__6_), .ZN(MULT_mult_6_n1309) );
  INV_X4 MULT_mult_6_U2785 ( .A(MULT_mult_6_net88703), .ZN(
        MULT_mult_6_net88704) );
  XNOR2_X2 MULT_mult_6_U2784 ( .A(MULT_mult_6_n2303), .B(MULT_mult_6_net88703), 
        .ZN(MULT_mult_6_SUMB_9__16_) );
  INV_X4 MULT_mult_6_U2783 ( .A(MULT_mult_6_net86864), .ZN(
        MULT_mult_6_net123592) );
  INV_X4 MULT_mult_6_U2782 ( .A(MULT_mult_6_net93243), .ZN(
        MULT_mult_6_net123591) );
  NAND2_X4 MULT_mult_6_U2781 ( .A1(MULT_mult_6_n883), .A2(MULT_mult_6_n884), 
        .ZN(MULT_mult_6_SUMB_2__14_) );
  NAND2_X4 MULT_mult_6_U2780 ( .A1(MULT_mult_6_net123592), .A2(
        MULT_mult_6_net123591), .ZN(MULT_mult_6_n884) );
  NAND2_X2 MULT_mult_6_U2779 ( .A1(MULT_mult_6_net86864), .A2(
        MULT_mult_6_net93243), .ZN(MULT_mult_6_n883) );
  INV_X1 MULT_mult_6_U2778 ( .A(MULT_mult_6_SUMB_18__12_), .ZN(
        MULT_mult_6_n880) );
  INV_X4 MULT_mult_6_U2777 ( .A(MULT_mult_6_n1606), .ZN(MULT_mult_6_n879) );
  NAND2_X4 MULT_mult_6_U2776 ( .A1(MULT_mult_6_n881), .A2(MULT_mult_6_n882), 
        .ZN(MULT_mult_6_SUMB_19__11_) );
  NAND2_X2 MULT_mult_6_U2775 ( .A1(MULT_mult_6_n879), .A2(MULT_mult_6_n880), 
        .ZN(MULT_mult_6_n882) );
  NAND2_X1 MULT_mult_6_U2774 ( .A1(MULT_mult_6_n1606), .A2(
        MULT_mult_6_SUMB_18__12_), .ZN(MULT_mult_6_n881) );
  INV_X1 MULT_mult_6_U2773 ( .A(MULT_mult_6_ab_7__22_), .ZN(MULT_mult_6_n875)
         );
  NAND2_X2 MULT_mult_6_U2771 ( .A1(MULT_mult_6_n875), .A2(MULT_mult_6_n876), 
        .ZN(MULT_mult_6_n878) );
  NAND2_X2 MULT_mult_6_U2770 ( .A1(MULT_mult_6_ab_3__11_), .A2(
        MULT_mult_6_CARRYB_2__11_), .ZN(MULT_mult_6_n2030) );
  NAND2_X4 MULT_mult_6_U2769 ( .A1(MULT_mult_6_ab_3__11_), .A2(
        MULT_mult_6_SUMB_2__12_), .ZN(MULT_mult_6_n2029) );
  NAND2_X2 MULT_mult_6_U2768 ( .A1(MULT_mult_6_SUMB_13__8_), .A2(
        MULT_mult_6_CARRYB_13__7_), .ZN(MULT_mult_6_net84998) );
  INV_X4 MULT_mult_6_U2767 ( .A(MULT_mult_6_n1679), .ZN(MULT_mult_6_n1317) );
  NAND2_X2 MULT_mult_6_U2766 ( .A1(MULT_mult_6_n1504), .A2(
        MULT_mult_6_SUMB_1__13_), .ZN(MULT_mult_6_n886) );
  NAND2_X2 MULT_mult_6_U2765 ( .A1(MULT_mult_6_net124104), .A2(
        MULT_mult_6_n1679), .ZN(MULT_mult_6_n1318) );
  NAND2_X4 MULT_mult_6_U2764 ( .A1(MULT_mult_6_SUMB_8__10_), .A2(
        MULT_mult_6_CARRYB_8__9_), .ZN(MULT_mult_6_n1619) );
  NAND2_X4 MULT_mult_6_U2763 ( .A1(MULT_mult_6_SUMB_8__10_), .A2(
        MULT_mult_6_ab_9__9_), .ZN(MULT_mult_6_n1620) );
  INV_X2 MULT_mult_6_U2762 ( .A(MULT_mult_6_net120922), .ZN(
        MULT_mult_6_net123843) );
  NAND2_X4 MULT_mult_6_U2761 ( .A1(MULT_mult_6_n874), .A2(MULT_mult_6_n873), 
        .ZN(MULT_mult_6_SUMB_8__10_) );
  NAND2_X4 MULT_mult_6_U2760 ( .A1(MULT_mult_6_net123842), .A2(
        MULT_mult_6_net123843), .ZN(MULT_mult_6_n874) );
  NOR2_X1 MULT_mult_6_U2759 ( .A1(MULT_mult_6_n2354), .A2(MULT_mult_6_n242), 
        .ZN(MULT_mult_6_ab_1__28_) );
  NAND2_X1 MULT_mult_6_U2758 ( .A1(MULT_mult_6_ab_8__16_), .A2(
        MULT_mult_6_CARRYB_7__16_), .ZN(MULT_mult_6_n2297) );
  NAND2_X4 MULT_mult_6_U2757 ( .A1(MULT_mult_6_n1386), .A2(MULT_mult_6_n428), 
        .ZN(MULT_mult_6_n1388) );
  NAND2_X1 MULT_mult_6_U2756 ( .A1(MULT_mult_6_CARRYB_12__13_), .A2(
        MULT_mult_6_SUMB_12__14_), .ZN(MULT_mult_6_n1575) );
  INV_X2 MULT_mult_6_U2755 ( .A(MULT_mult_6_net82757), .ZN(
        MULT_mult_6_net123897) );
  NAND2_X4 MULT_mult_6_U2754 ( .A1(MULT_mult_6_net123899), .A2(
        MULT_mult_6_n872), .ZN(MULT_mult_6_n1456) );
  NAND3_X2 MULT_mult_6_U2753 ( .A1(MULT_mult_6_n1969), .A2(MULT_mult_6_n1968), 
        .A3(MULT_mult_6_n1967), .ZN(MULT_mult_6_CARRYB_14__3_) );
  XNOR2_X2 MULT_mult_6_U2752 ( .A(MULT_mult_6_n1942), .B(MULT_mult_6_n1256), 
        .ZN(MULT_mult_6_net124104) );
  NAND2_X2 MULT_mult_6_U2751 ( .A1(MULT_mult_6_CARRYB_11__12_), .A2(
        MULT_mult_6_ab_12__12_), .ZN(MULT_mult_6_n1019) );
  NAND2_X1 MULT_mult_6_U2750 ( .A1(MULT_mult_6_n1781), .A2(MULT_mult_6_n1782), 
        .ZN(MULT_mult_6_n1784) );
  NAND3_X2 MULT_mult_6_U2749 ( .A1(MULT_mult_6_n1910), .A2(MULT_mult_6_n1909), 
        .A3(MULT_mult_6_n1908), .ZN(MULT_mult_6_CARRYB_4__7_) );
  INV_X2 MULT_mult_6_U2748 ( .A(MULT_mult_6_n2060), .ZN(MULT_mult_6_n1458) );
  XOR2_X1 MULT_mult_6_U2747 ( .A(MULT_mult_6_n1139), .B(
        MULT_mult_6_SUMB_10__1_), .Z(multOut[20]) );
  NAND2_X1 MULT_mult_6_U2746 ( .A1(MULT_mult_6_ab_11__0_), .A2(
        MULT_mult_6_SUMB_10__1_), .ZN(MULT_mult_6_n1141) );
  NAND3_X2 MULT_mult_6_U2745 ( .A1(MULT_mult_6_net79867), .A2(
        MULT_mult_6_net79868), .A3(MULT_mult_6_n1062), .ZN(
        MULT_mult_6_CARRYB_25__5_) );
  XNOR2_X2 MULT_mult_6_U2744 ( .A(MULT_mult_6_n368), .B(
        MULT_mult_6_SUMB_19__9_), .ZN(MULT_mult_6_n869) );
  NAND2_X1 MULT_mult_6_U2743 ( .A1(MULT_mult_6_ab_8__19_), .A2(
        MULT_mult_6_SUMB_7__20_), .ZN(MULT_mult_6_net79956) );
  INV_X2 MULT_mult_6_U2742 ( .A(MULT_mult_6_ab_19__9_), .ZN(
        MULT_mult_6_net87133) );
  INV_X4 MULT_mult_6_U2741 ( .A(MULT_mult_6_n865), .ZN(MULT_mult_6_n866) );
  INV_X2 MULT_mult_6_U2740 ( .A(MULT_mult_6_SUMB_2__22_), .ZN(MULT_mult_6_n865) );
  INV_X4 MULT_mult_6_U2739 ( .A(MULT_mult_6_CARRYB_11__12_), .ZN(
        MULT_mult_6_net120585) );
  XNOR2_X2 MULT_mult_6_U2738 ( .A(MULT_mult_6_n862), .B(MULT_mult_6_n871), 
        .ZN(MULT_mult_6_SUMB_16__3_) );
  XNOR2_X2 MULT_mult_6_U2737 ( .A(MULT_mult_6_SUMB_8__6_), .B(
        MULT_mult_6_ab_9__5_), .ZN(MULT_mult_6_n1448) );
  INV_X4 MULT_mult_6_U2736 ( .A(MULT_mult_6_CARRYB_3__10_), .ZN(
        MULT_mult_6_n888) );
  NAND3_X2 MULT_mult_6_U2735 ( .A1(MULT_mult_6_n1933), .A2(MULT_mult_6_n1934), 
        .A3(MULT_mult_6_n1935), .ZN(MULT_mult_6_CARRYB_3__21_) );
  NAND2_X2 MULT_mult_6_U2733 ( .A1(MULT_mult_6_SUMB_6__17_), .A2(
        MULT_mult_6_n1368), .ZN(MULT_mult_6_n2251) );
  NAND2_X2 MULT_mult_6_U2732 ( .A1(MULT_mult_6_n299), .A2(
        MULT_mult_6_net123142), .ZN(MULT_mult_6_n909) );
  NOR2_X4 MULT_mult_6_U2731 ( .A1(MULT_mult_6_net82890), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__17_) );
  XOR2_X2 MULT_mult_6_U2730 ( .A(MULT_mult_6_ab_13__17_), .B(
        MULT_mult_6_CARRYB_12__17_), .Z(MULT_mult_6_n860) );
  NAND2_X4 MULT_mult_6_U2729 ( .A1(MULT_mult_6_net81033), .A2(MULT_mult_6_n937), .ZN(MULT_mult_6_net82396) );
  XNOR2_X2 MULT_mult_6_U2728 ( .A(MULT_mult_6_net82396), .B(
        MULT_mult_6_SUMB_19__10_), .ZN(MULT_mult_6_n859) );
  NAND3_X2 MULT_mult_6_U2727 ( .A1(MULT_mult_6_n2305), .A2(MULT_mult_6_n2304), 
        .A3(MULT_mult_6_n2306), .ZN(MULT_mult_6_CARRYB_9__16_) );
  NOR2_X1 MULT_mult_6_U2726 ( .A1(MULT_mult_6_net80727), .A2(
        MULT_mult_6_net77948), .ZN(MULT_mult_6_ab_5__20_) );
  XNOR2_X2 MULT_mult_6_U2725 ( .A(MULT_mult_6_CARRYB_4__20_), .B(
        MULT_mult_6_ab_5__20_), .ZN(MULT_mult_6_n1210) );
  NAND2_X4 MULT_mult_6_U2724 ( .A1(MULT_mult_6_CARRYB_3__14_), .A2(
        MULT_mult_6_ab_4__14_), .ZN(MULT_mult_6_net92718) );
  NAND3_X2 MULT_mult_6_U2723 ( .A1(MULT_mult_6_n2219), .A2(MULT_mult_6_n2220), 
        .A3(MULT_mult_6_n2221), .ZN(MULT_mult_6_CARRYB_10__19_) );
  BUF_X8 MULT_mult_6_U2722 ( .A(MULT_mult_6_SUMB_9__2_), .Z(
        MULT_mult_6_net124757) );
  XNOR2_X2 MULT_mult_6_U2721 ( .A(MULT_mult_6_n1663), .B(
        MULT_mult_6_SUMB_20__10_), .ZN(MULT_mult_6_n856) );
  XNOR2_X2 MULT_mult_6_U2720 ( .A(MULT_mult_6_CARRYB_6__21_), .B(
        MULT_mult_6_ab_7__21_), .ZN(MULT_mult_6_n855) );
  XNOR2_X1 MULT_mult_6_U2719 ( .A(MULT_mult_6_SUMB_6__22_), .B(
        MULT_mult_6_n855), .ZN(MULT_mult_6_SUMB_7__21_) );
  NAND3_X2 MULT_mult_6_U2718 ( .A1(MULT_mult_6_n1919), .A2(MULT_mult_6_n1918), 
        .A3(MULT_mult_6_n1917), .ZN(MULT_mult_6_n854) );
  NAND2_X2 MULT_mult_6_U2717 ( .A1(MULT_mult_6_net81491), .A2(
        MULT_mult_6_CARRYB_21__7_), .ZN(MULT_mult_6_net83121) );
  INV_X4 MULT_mult_6_U2716 ( .A(MULT_mult_6_CARRYB_21__7_), .ZN(
        MULT_mult_6_net83120) );
  XNOR2_X2 MULT_mult_6_U2715 ( .A(MULT_mult_6_n1880), .B(MULT_mult_6_n1217), 
        .ZN(MULT_mult_6_n853) );
  NAND2_X4 MULT_mult_6_U2714 ( .A1(MULT_mult_6_CARRYB_11__9_), .A2(
        MULT_mult_6_ab_12__9_), .ZN(MULT_mult_6_net88297) );
  INV_X2 MULT_mult_6_U2713 ( .A(MULT_mult_6_net91301), .ZN(
        MULT_mult_6_net83151) );
  NAND2_X2 MULT_mult_6_U2712 ( .A1(MULT_mult_6_CARRYB_26__3_), .A2(
        MULT_mult_6_ab_27__3_), .ZN(MULT_mult_6_n1535) );
  NAND2_X4 MULT_mult_6_U2711 ( .A1(MULT_mult_6_n1548), .A2(MULT_mult_6_n1549), 
        .ZN(MULT_mult_6_n2111) );
  INV_X8 MULT_mult_6_U2710 ( .A(MULT_mult_6_n850), .ZN(MULT_mult_6_n851) );
  INV_X4 MULT_mult_6_U2709 ( .A(MULT_mult_6_SUMB_7__21_), .ZN(MULT_mult_6_n850) );
  NAND2_X2 MULT_mult_6_U2708 ( .A1(MULT_mult_6_ab_19__9_), .A2(
        MULT_mult_6_CARRYB_18__9_), .ZN(MULT_mult_6_n935) );
  XNOR2_X2 MULT_mult_6_U2707 ( .A(MULT_mult_6_n2367), .B(MULT_mult_6_n1233), 
        .ZN(MULT_mult_6_n848) );
  CLKBUF_X3 MULT_mult_6_U2706 ( .A(MULT_mult_6_SUMB_14__12_), .Z(
        MULT_mult_6_net125062) );
  INV_X4 MULT_mult_6_U2705 ( .A(MULT_mult_6_net83134), .ZN(
        MULT_mult_6_net86702) );
  NAND3_X2 MULT_mult_6_U2704 ( .A1(MULT_mult_6_net80838), .A2(
        MULT_mult_6_net80839), .A3(MULT_mult_6_net80840), .ZN(MULT_mult_6_n847) );
  INV_X2 MULT_mult_6_U2703 ( .A(MULT_mult_6_n845), .ZN(MULT_mult_6_n846) );
  INV_X1 MULT_mult_6_U2702 ( .A(MULT_mult_6_CARRYB_14__0_), .ZN(
        MULT_mult_6_n845) );
  NOR2_X1 MULT_mult_6_U2701 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net77938), .ZN(MULT_mult_6_ab_6__9_) );
  NAND2_X4 MULT_mult_6_U2700 ( .A1(MULT_mult_6_n885), .A2(
        MULT_mult_6_net123509), .ZN(MULT_mult_6_n887) );
  XNOR2_X2 MULT_mult_6_U2699 ( .A(MULT_mult_6_net87855), .B(
        MULT_mult_6_net90671), .ZN(MULT_mult_6_n843) );
  INV_X4 MULT_mult_6_U2698 ( .A(MULT_mult_6_CARRYB_7__11_), .ZN(
        MULT_mult_6_n1659) );
  CLKBUF_X2 MULT_mult_6_U2697 ( .A(MULT_mult_6_SUMB_10__4_), .Z(
        MULT_mult_6_n842) );
  NAND2_X2 MULT_mult_6_U2696 ( .A1(MULT_mult_6_ab_7__22_), .A2(
        MULT_mult_6_CARRYB_6__22_), .ZN(MULT_mult_6_n877) );
  XNOR2_X2 MULT_mult_6_U2695 ( .A(MULT_mult_6_ab_3__22_), .B(
        MULT_mult_6_CARRYB_2__22_), .ZN(MULT_mult_6_n841) );
  XNOR2_X2 MULT_mult_6_U2694 ( .A(MULT_mult_6_n841), .B(MULT_mult_6_n34), .ZN(
        MULT_mult_6_SUMB_3__22_) );
  INV_X4 MULT_mult_6_U2693 ( .A(MULT_mult_6_n839), .ZN(MULT_mult_6_n840) );
  INV_X2 MULT_mult_6_U2692 ( .A(MULT_mult_6_SUMB_6__21_), .ZN(MULT_mult_6_n839) );
  NOR2_X1 MULT_mult_6_U2691 ( .A1(MULT_mult_6_net70482), .A2(MULT_mult_6_n331), 
        .ZN(MULT_mult_6_ab_2__24_) );
  NOR2_X1 MULT_mult_6_U2690 ( .A1(MULT_mult_6_net70482), .A2(MULT_mult_6_n331), 
        .ZN(MULT_mult_6_n838) );
  NAND2_X1 MULT_mult_6_U2689 ( .A1(MULT_mult_6_CARRYB_13__11_), .A2(
        MULT_mult_6_ab_14__11_), .ZN(MULT_mult_6_net82556) );
  XNOR2_X2 MULT_mult_6_U2688 ( .A(MULT_mult_6_CARRYB_13__11_), .B(
        MULT_mult_6_ab_14__11_), .ZN(MULT_mult_6_net90817) );
  INV_X4 MULT_mult_6_U2687 ( .A(MULT_mult_6_net93672), .ZN(
        MULT_mult_6_net87654) );
  INV_X2 MULT_mult_6_U2686 ( .A(MULT_mult_6_net81548), .ZN(
        MULT_mult_6_net87655) );
  NAND2_X4 MULT_mult_6_U2685 ( .A1(MULT_mult_6_net87654), .A2(
        MULT_mult_6_net87655), .ZN(MULT_mult_6_n837) );
  NAND2_X4 MULT_mult_6_U2684 ( .A1(MULT_mult_6_n837), .A2(MULT_mult_6_n836), 
        .ZN(MULT_mult_6_net81157) );
  INV_X4 MULT_mult_6_U2683 ( .A(MULT_mult_6_net81157), .ZN(
        MULT_mult_6_net92325) );
  NAND2_X4 MULT_mult_6_U2682 ( .A1(MULT_mult_6_n834), .A2(MULT_mult_6_n835), 
        .ZN(MULT_mult_6_net92317) );
  NAND2_X1 MULT_mult_6_U2681 ( .A1(MULT_mult_6_SUMB_25__4_), .A2(
        MULT_mult_6_net84891), .ZN(MULT_mult_6_net81053) );
  XNOR2_X2 MULT_mult_6_U2680 ( .A(MULT_mult_6_net81663), .B(MULT_mult_6_n91), 
        .ZN(MULT_mult_6_SUMB_26__3_) );
  NAND2_X2 MULT_mult_6_U2679 ( .A1(MULT_mult_6_ab_8__14_), .A2(
        MULT_mult_6_CARRYB_7__14_), .ZN(MULT_mult_6_net80356) );
  NAND2_X2 MULT_mult_6_U2678 ( .A1(MULT_mult_6_CARRYB_7__14_), .A2(
        MULT_mult_6_SUMB_7__15_), .ZN(MULT_mult_6_net80355) );
  XNOR2_X2 MULT_mult_6_U2677 ( .A(MULT_mult_6_net81995), .B(MULT_mult_6_n833), 
        .ZN(MULT_mult_6_SUMB_8__14_) );
  NAND2_X2 MULT_mult_6_U2676 ( .A1(MULT_mult_6_ab_9__13_), .A2(
        MULT_mult_6_CARRYB_8__13_), .ZN(MULT_mult_6_net80348) );
  NOR2_X2 MULT_mult_6_U2675 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__13_) );
  NAND2_X2 MULT_mult_6_U2674 ( .A1(MULT_mult_6_ab_10__13_), .A2(
        MULT_mult_6_CARRYB_9__13_), .ZN(MULT_mult_6_net80246) );
  NAND2_X2 MULT_mult_6_U2673 ( .A1(MULT_mult_6_ab_10__13_), .A2(
        MULT_mult_6_SUMB_9__14_), .ZN(MULT_mult_6_net80247) );
  XNOR2_X2 MULT_mult_6_U2672 ( .A(MULT_mult_6_CARRYB_9__13_), .B(
        MULT_mult_6_ab_10__13_), .ZN(MULT_mult_6_n832) );
  XNOR2_X2 MULT_mult_6_U2671 ( .A(MULT_mult_6_n832), .B(
        MULT_mult_6_SUMB_9__14_), .ZN(MULT_mult_6_SUMB_10__13_) );
  XNOR2_X2 MULT_mult_6_U2670 ( .A(MULT_mult_6_net84163), .B(
        MULT_mult_6_net87942), .ZN(MULT_mult_6_net89255) );
  NAND2_X2 MULT_mult_6_U2669 ( .A1(MULT_mult_6_net89255), .A2(
        MULT_mult_6_CARRYB_14__9_), .ZN(MULT_mult_6_n829) );
  INV_X4 MULT_mult_6_U2668 ( .A(MULT_mult_6_net120648), .ZN(
        MULT_mult_6_net82263) );
  XNOR2_X2 MULT_mult_6_U2667 ( .A(MULT_mult_6_net84163), .B(
        MULT_mult_6_net93756), .ZN(MULT_mult_6_SUMB_14__10_) );
  NAND3_X4 MULT_mult_6_U2666 ( .A1(MULT_mult_6_n829), .A2(MULT_mult_6_n828), 
        .A3(MULT_mult_6_n827), .ZN(MULT_mult_6_CARRYB_15__9_) );
  NAND2_X1 MULT_mult_6_U2665 ( .A1(MULT_mult_6_ab_18__9_), .A2(
        MULT_mult_6_SUMB_17__10_), .ZN(MULT_mult_6_net80880) );
  XNOR2_X2 MULT_mult_6_U2664 ( .A(MULT_mult_6_n150), .B(MULT_mult_6_n826), 
        .ZN(MULT_mult_6_net88692) );
  NOR2_X1 MULT_mult_6_U2663 ( .A1(MULT_mult_6_net91660), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__10_) );
  NAND3_X2 MULT_mult_6_U2662 ( .A1(MULT_mult_6_net81058), .A2(
        MULT_mult_6_net81057), .A3(MULT_mult_6_net81056), .ZN(
        MULT_mult_6_net124392) );
  INV_X4 MULT_mult_6_U2661 ( .A(MULT_mult_6_SUMB_12__11_), .ZN(
        MULT_mult_6_net85465) );
  NAND2_X2 MULT_mult_6_U2660 ( .A1(MULT_mult_6_net84007), .A2(
        MULT_mult_6_net124392), .ZN(MULT_mult_6_net84211) );
  INV_X4 MULT_mult_6_U2659 ( .A(MULT_mult_6_ab_13__10_), .ZN(
        MULT_mult_6_net84007) );
  INV_X2 MULT_mult_6_U2658 ( .A(MULT_mult_6_ab_8__13_), .ZN(
        MULT_mult_6_net87065) );
  NAND2_X4 MULT_mult_6_U2657 ( .A1(MULT_mult_6_net87067), .A2(
        MULT_mult_6_net87068), .ZN(MULT_mult_6_net81958) );
  NAND2_X4 MULT_mult_6_U2656 ( .A1(MULT_mult_6_CARRYB_7__13_), .A2(
        MULT_mult_6_ab_8__13_), .ZN(MULT_mult_6_net87067) );
  XNOR2_X2 MULT_mult_6_U2655 ( .A(MULT_mult_6_CARRYB_18__8_), .B(
        MULT_mult_6_ab_19__8_), .ZN(MULT_mult_6_net88700) );
  NOR2_X4 MULT_mult_6_U2654 ( .A1(MULT_mult_6_net81424), .A2(
        MULT_mult_6_net77948), .ZN(MULT_mult_6_ab_5__15_) );
  NAND2_X1 MULT_mult_6_U2653 ( .A1(MULT_mult_6_ab_5__15_), .A2(MULT_mult_6_n93), .ZN(MULT_mult_6_net80838) );
  NAND2_X4 MULT_mult_6_U2652 ( .A1(MULT_mult_6_net124908), .A2(
        MULT_mult_6_net120511), .ZN(MULT_mult_6_net88079) );
  NOR2_X2 MULT_mult_6_U2651 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__12_) );
  NAND3_X2 MULT_mult_6_U2650 ( .A1(MULT_mult_6_net80251), .A2(
        MULT_mult_6_net80250), .A3(MULT_mult_6_net83630), .ZN(
        MULT_mult_6_CARRYB_11__12_) );
  INV_X1 MULT_mult_6_U2649 ( .A(MULT_mult_6_ab_11__12_), .ZN(
        MULT_mult_6_net83628) );
  NAND2_X1 MULT_mult_6_U2647 ( .A1(MULT_mult_6_ab_22__6_), .A2(
        MULT_mult_6_CARRYB_21__6_), .ZN(MULT_mult_6_net80940) );
  NAND2_X2 MULT_mult_6_U2646 ( .A1(MULT_mult_6_ab_22__6_), .A2(
        MULT_mult_6_SUMB_21__7_), .ZN(MULT_mult_6_net80941) );
  NAND2_X2 MULT_mult_6_U2645 ( .A1(MULT_mult_6_SUMB_21__7_), .A2(
        MULT_mult_6_net89008), .ZN(MULT_mult_6_net80942) );
  INV_X4 MULT_mult_6_U2644 ( .A(MULT_mult_6_CARRYB_21__6_), .ZN(
        MULT_mult_6_n818) );
  NAND2_X2 MULT_mult_6_U2643 ( .A1(MULT_mult_6_n824), .A2(
        MULT_mult_6_CARRYB_21__6_), .ZN(MULT_mult_6_n819) );
  XNOR2_X2 MULT_mult_6_U2642 ( .A(MULT_mult_6_SUMB_21__7_), .B(
        MULT_mult_6_n822), .ZN(MULT_mult_6_n823) );
  XNOR2_X2 MULT_mult_6_U2641 ( .A(MULT_mult_6_net81983), .B(MULT_mult_6_n821), 
        .ZN(MULT_mult_6_net93813) );
  NAND2_X4 MULT_mult_6_U2640 ( .A1(MULT_mult_6_n821), .A2(
        MULT_mult_6_ab_23__5_), .ZN(MULT_mult_6_net79905) );
  NAND2_X4 MULT_mult_6_U2639 ( .A1(MULT_mult_6_net88860), .A2(MULT_mult_6_n821), .ZN(MULT_mult_6_net79906) );
  INV_X8 MULT_mult_6_U2638 ( .A(MULT_mult_6_n823), .ZN(MULT_mult_6_n821) );
  XNOR2_X2 MULT_mult_6_U2637 ( .A(MULT_mult_6_net81983), .B(MULT_mult_6_n821), 
        .ZN(MULT_mult_6_SUMB_23__5_) );
  NAND3_X2 MULT_mult_6_U2636 ( .A1(MULT_mult_6_net82030), .A2(
        MULT_mult_6_net82029), .A3(MULT_mult_6_net82031), .ZN(
        MULT_mult_6_net123303) );
  NAND2_X4 MULT_mult_6_U2635 ( .A1(MULT_mult_6_net119921), .A2(
        MULT_mult_6_n817), .ZN(MULT_mult_6_net82030) );
  XNOR2_X2 MULT_mult_6_U2634 ( .A(MULT_mult_6_net86799), .B(
        MULT_mult_6_net88668), .ZN(MULT_mult_6_SUMB_15__10_) );
  NOR2_X1 MULT_mult_6_U2633 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net70463), .ZN(MULT_mult_6_ab_16__9_) );
  NOR2_X1 MULT_mult_6_U2632 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70449), .ZN(MULT_mult_6_ab_23__4_) );
  NAND2_X2 MULT_mult_6_U2631 ( .A1(MULT_mult_6_n816), .A2(MULT_mult_6_net81169), .ZN(MULT_mult_6_net87688) );
  INV_X4 MULT_mult_6_U2630 ( .A(MULT_mult_6_net81169), .ZN(MULT_mult_6_n814)
         );
  NAND2_X4 MULT_mult_6_U2629 ( .A1(MULT_mult_6_net87688), .A2(MULT_mult_6_n815), .ZN(MULT_mult_6_SUMB_15__11_) );
  NOR2_X1 MULT_mult_6_U2628 ( .A1(MULT_mult_6_net91660), .A2(
        MULT_mult_6_net70463), .ZN(MULT_mult_6_ab_16__10_) );
  XNOR2_X2 MULT_mult_6_U2627 ( .A(MULT_mult_6_net86801), .B(
        MULT_mult_6_net90817), .ZN(MULT_mult_6_net88668) );
  BUF_X4 MULT_mult_6_U2626 ( .A(MULT_mult_6_SUMB_13__12_), .Z(
        MULT_mult_6_net86801) );
  NAND2_X2 MULT_mult_6_U2625 ( .A1(MULT_mult_6_SUMB_14__11_), .A2(
        MULT_mult_6_ab_15__10_), .ZN(MULT_mult_6_net82560) );
  NAND3_X2 MULT_mult_6_U2624 ( .A1(MULT_mult_6_net82561), .A2(
        MULT_mult_6_net82560), .A3(MULT_mult_6_net82559), .ZN(
        MULT_mult_6_CARRYB_15__10_) );
  NAND2_X1 MULT_mult_6_U2623 ( .A1(MULT_mult_6_ab_17__10_), .A2(
        MULT_mult_6_n390), .ZN(MULT_mult_6_net84746) );
  XNOR2_X2 MULT_mult_6_U2622 ( .A(MULT_mult_6_n390), .B(MULT_mult_6_ab_17__10_), .ZN(MULT_mult_6_net85325) );
  NAND2_X2 MULT_mult_6_U2621 ( .A1(MULT_mult_6_net87944), .A2(
        MULT_mult_6_net85807), .ZN(MULT_mult_6_n813) );
  NAND2_X4 MULT_mult_6_U2620 ( .A1(MULT_mult_6_net85808), .A2(
        MULT_mult_6_net89819), .ZN(MULT_mult_6_net80812) );
  INV_X8 MULT_mult_6_U2619 ( .A(MULT_mult_6_net85807), .ZN(
        MULT_mult_6_net85808) );
  NAND2_X4 MULT_mult_6_U2618 ( .A1(MULT_mult_6_n813), .A2(MULT_mult_6_net87945), .ZN(MULT_mult_6_SUMB_17__9_) );
  NAND2_X1 MULT_mult_6_U2617 ( .A1(MULT_mult_6_ab_17__8_), .A2(
        MULT_mult_6_CARRYB_16__8_), .ZN(MULT_mult_6_n810) );
  NAND3_X4 MULT_mult_6_U2616 ( .A1(MULT_mult_6_n812), .A2(MULT_mult_6_n811), 
        .A3(MULT_mult_6_n810), .ZN(MULT_mult_6_CARRYB_17__8_) );
  INV_X16 MULT_mult_6_U2615 ( .A(WIRE_ALU_A_MUX2TO1_32BIT_13__MUX_N1), .ZN(
        MULT_mult_6_net70459) );
  NOR2_X4 MULT_mult_6_U2614 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net70459), .ZN(MULT_mult_6_ab_18__8_) );
  NAND2_X4 MULT_mult_6_U2613 ( .A1(MULT_mult_6_net83628), .A2(
        MULT_mult_6_net83629), .ZN(MULT_mult_6_net83631) );
  NAND2_X4 MULT_mult_6_U2612 ( .A1(MULT_mult_6_net83630), .A2(
        MULT_mult_6_net83631), .ZN(MULT_mult_6_net81087) );
  NAND2_X1 MULT_mult_6_U2611 ( .A1(MULT_mult_6_ab_11__11_), .A2(
        MULT_mult_6_net88525), .ZN(MULT_mult_6_net81168) );
  NAND2_X2 MULT_mult_6_U2610 ( .A1(MULT_mult_6_SUMB_10__12_), .A2(
        MULT_mult_6_net87490), .ZN(MULT_mult_6_net81166) );
  NAND3_X2 MULT_mult_6_U2609 ( .A1(MULT_mult_6_net79991), .A2(
        MULT_mult_6_net79990), .A3(MULT_mult_6_net79989), .ZN(
        MULT_mult_6_CARRYB_21__5_) );
  NAND3_X2 MULT_mult_6_U2608 ( .A1(MULT_mult_6_net80686), .A2(MULT_mult_6_n809), .A3(MULT_mult_6_net93918), .ZN(MULT_mult_6_CARRYB_27__2_) );
  NAND2_X2 MULT_mult_6_U2607 ( .A1(MULT_mult_6_net89453), .A2(
        MULT_mult_6_net87797), .ZN(MULT_mult_6_net80472) );
  NAND3_X4 MULT_mult_6_U2606 ( .A1(MULT_mult_6_net80262), .A2(
        MULT_mult_6_net80261), .A3(MULT_mult_6_net80263), .ZN(
        MULT_mult_6_CARRYB_25__2_) );
  INV_X4 MULT_mult_6_U2605 ( .A(WIRE_ALU_A_MUX2TO1_32BIT_5__MUX_N1), .ZN(
        MULT_mult_6_net70443) );
  NOR2_X4 MULT_mult_6_U2604 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70443), .ZN(MULT_mult_6_ab_26__2_) );
  NAND2_X2 MULT_mult_6_U2603 ( .A1(MULT_mult_6_ab_26__2_), .A2(
        MULT_mult_6_CARRYB_25__2_), .ZN(MULT_mult_6_net80987) );
  NAND2_X4 MULT_mult_6_U2602 ( .A1(MULT_mult_6_CARRYB_26__2_), .A2(
        MULT_mult_6_ab_27__2_), .ZN(MULT_mult_6_net93918) );
  NAND3_X4 MULT_mult_6_U2601 ( .A1(MULT_mult_6_net80989), .A2(
        MULT_mult_6_net80988), .A3(MULT_mult_6_net80987), .ZN(
        MULT_mult_6_CARRYB_26__2_) );
  NAND2_X2 MULT_mult_6_U2600 ( .A1(MULT_mult_6_net83866), .A2(
        MULT_mult_6_SUMB_11__12_), .ZN(MULT_mult_6_net85457) );
  NAND2_X2 MULT_mult_6_U2599 ( .A1(MULT_mult_6_ab_11__12_), .A2(
        MULT_mult_6_SUMB_10__13_), .ZN(MULT_mult_6_net80250) );
  NAND3_X2 MULT_mult_6_U2598 ( .A1(MULT_mult_6_net81166), .A2(
        MULT_mult_6_net81167), .A3(MULT_mult_6_net81168), .ZN(
        MULT_mult_6_net90604) );
  NOR2_X4 MULT_mult_6_U2597 ( .A1(MULT_mult_6_net85716), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__11_) );
  NAND2_X4 MULT_mult_6_U2596 ( .A1(MULT_mult_6_SUMB_11__12_), .A2(
        MULT_mult_6_ab_12__11_), .ZN(MULT_mult_6_net82022) );
  XNOR2_X2 MULT_mult_6_U2595 ( .A(MULT_mult_6_net90262), .B(
        MULT_mult_6_net81087), .ZN(MULT_mult_6_SUMB_11__12_) );
  XNOR2_X2 MULT_mult_6_U2594 ( .A(MULT_mult_6_net90262), .B(
        MULT_mult_6_net81087), .ZN(MULT_mult_6_net124563) );
  NAND3_X2 MULT_mult_6_U2593 ( .A1(MULT_mult_6_net81166), .A2(
        MULT_mult_6_net81167), .A3(MULT_mult_6_net81168), .ZN(
        MULT_mult_6_CARRYB_11__11_) );
  NAND2_X4 MULT_mult_6_U2592 ( .A1(MULT_mult_6_n807), .A2(MULT_mult_6_net84824), .ZN(MULT_mult_6_net84826) );
  INV_X4 MULT_mult_6_U2591 ( .A(MULT_mult_6_CARRYB_11__11_), .ZN(
        MULT_mult_6_n807) );
  INV_X1 MULT_mult_6_U2590 ( .A(MULT_mult_6_n807), .ZN(MULT_mult_6_n808) );
  NAND2_X4 MULT_mult_6_U2589 ( .A1(MULT_mult_6_net89670), .A2(MULT_mult_6_n808), .ZN(MULT_mult_6_net82021) );
  NAND3_X4 MULT_mult_6_U2588 ( .A1(MULT_mult_6_net82022), .A2(
        MULT_mult_6_net82021), .A3(MULT_mult_6_n806), .ZN(
        MULT_mult_6_CARRYB_12__11_) );
  NAND2_X2 MULT_mult_6_U2587 ( .A1(MULT_mult_6_n565), .A2(
        MULT_mult_6_CARRYB_8__13_), .ZN(MULT_mult_6_net80350) );
  NAND3_X2 MULT_mult_6_U2586 ( .A1(MULT_mult_6_net84678), .A2(
        MULT_mult_6_net84679), .A3(MULT_mult_6_net84680), .ZN(
        MULT_mult_6_CARRYB_24__3_) );
  NAND3_X4 MULT_mult_6_U2585 ( .A1(MULT_mult_6_net80992), .A2(
        MULT_mult_6_net80991), .A3(MULT_mult_6_net80990), .ZN(
        MULT_mult_6_CARRYB_27__1_) );
  NAND2_X2 MULT_mult_6_U2584 ( .A1(MULT_mult_6_n2356), .A2(
        MULT_mult_6_net86884), .ZN(MULT_mult_6_net80686) );
  INV_X1 MULT_mult_6_U2583 ( .A(MULT_mult_6_ab_10__12_), .ZN(
        MULT_mult_6_net84819) );
  NOR2_X2 MULT_mult_6_U2582 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__12_) );
  NAND2_X1 MULT_mult_6_U2581 ( .A1(MULT_mult_6_SUMB_9__13_), .A2(
        MULT_mult_6_net80983), .ZN(MULT_mult_6_net120653) );
  XNOR2_X2 MULT_mult_6_U2580 ( .A(MULT_mult_6_net85399), .B(
        MULT_mult_6_net80346), .ZN(MULT_mult_6_SUMB_9__13_) );
  XNOR2_X2 MULT_mult_6_U2578 ( .A(MULT_mult_6_net85399), .B(
        MULT_mult_6_net80346), .ZN(MULT_mult_6_net89065) );
  NAND2_X4 MULT_mult_6_U2577 ( .A1(MULT_mult_6_net80351), .A2(
        MULT_mult_6_net84822), .ZN(MULT_mult_6_net80983) );
  NAND2_X2 MULT_mult_6_U2576 ( .A1(MULT_mult_6_CARRYB_9__12_), .A2(
        MULT_mult_6_ab_10__12_), .ZN(MULT_mult_6_net80351) );
  NAND2_X4 MULT_mult_6_U2575 ( .A1(MULT_mult_6_SUMB_9__13_), .A2(
        MULT_mult_6_ab_10__12_), .ZN(MULT_mult_6_net80352) );
  NAND2_X4 MULT_mult_6_U2574 ( .A1(MULT_mult_6_net84819), .A2(
        MULT_mult_6_net84820), .ZN(MULT_mult_6_net84822) );
  INV_X4 MULT_mult_6_U2573 ( .A(MULT_mult_6_CARRYB_9__12_), .ZN(
        MULT_mult_6_net84820) );
  INV_X1 MULT_mult_6_U2572 ( .A(MULT_mult_6_net84820), .ZN(
        MULT_mult_6_net89982) );
  NAND2_X4 MULT_mult_6_U2571 ( .A1(MULT_mult_6_net89065), .A2(
        MULT_mult_6_net89982), .ZN(MULT_mult_6_net80353) );
  BUF_X4 MULT_mult_6_U2570 ( .A(MULT_mult_6_net80351), .Z(MULT_mult_6_net90996) );
  NAND2_X2 MULT_mult_6_U2569 ( .A1(MULT_mult_6_SUMB_10__13_), .A2(
        MULT_mult_6_CARRYB_10__12_), .ZN(MULT_mult_6_net80251) );
  NAND2_X2 MULT_mult_6_U2568 ( .A1(MULT_mult_6_CARRYB_10__12_), .A2(
        MULT_mult_6_ab_11__12_), .ZN(MULT_mult_6_net83630) );
  NAND3_X4 MULT_mult_6_U2567 ( .A1(MULT_mult_6_net80352), .A2(
        MULT_mult_6_net90996), .A3(MULT_mult_6_net80353), .ZN(
        MULT_mult_6_CARRYB_10__12_) );
  INV_X2 MULT_mult_6_U2566 ( .A(MULT_mult_6_net93813), .ZN(
        MULT_mult_6_net86022) );
  NAND2_X4 MULT_mult_6_U2565 ( .A1(MULT_mult_6_net86024), .A2(
        MULT_mult_6_net86023), .ZN(MULT_mult_6_SUMB_24__4_) );
  INV_X4 MULT_mult_6_U2564 ( .A(WIRE_ALU_A_MUX2TO1_32BIT_6__MUX_N1), .ZN(
        MULT_mult_6_net70445) );
  NOR2_X4 MULT_mult_6_U2563 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70445), .ZN(MULT_mult_6_ab_25__3_) );
  NAND3_X2 MULT_mult_6_U2562 ( .A1(MULT_mult_6_net81006), .A2(
        MULT_mult_6_net81007), .A3(MULT_mult_6_net87940), .ZN(
        MULT_mult_6_CARRYB_25__3_) );
  NAND3_X2 MULT_mult_6_U2561 ( .A1(MULT_mult_6_net81007), .A2(
        MULT_mult_6_net81006), .A3(MULT_mult_6_net87940), .ZN(
        MULT_mult_6_net123427) );
  NAND2_X4 MULT_mult_6_U2560 ( .A1(MULT_mult_6_n3), .A2(MULT_mult_6_ab_25__3_), 
        .ZN(MULT_mult_6_net87940) );
  INV_X1 MULT_mult_6_U2559 ( .A(MULT_mult_6_ab_25__3_), .ZN(
        MULT_mult_6_net87939) );
  NAND2_X4 MULT_mult_6_U2558 ( .A1(MULT_mult_6_net87941), .A2(
        MULT_mult_6_net87940), .ZN(MULT_mult_6_net82544) );
  NAND3_X4 MULT_mult_6_U2557 ( .A1(MULT_mult_6_net79909), .A2(
        MULT_mult_6_net79908), .A3(MULT_mult_6_net79907), .ZN(
        MULT_mult_6_CARRYB_24__4_) );
  NAND2_X2 MULT_mult_6_U2556 ( .A1(MULT_mult_6_ab_16__9_), .A2(
        MULT_mult_6_SUMB_15__10_), .ZN(MULT_mult_6_net79980) );
  CLKBUF_X3 MULT_mult_6_U2555 ( .A(MULT_mult_6_CARRYB_15__9_), .Z(
        MULT_mult_6_net121214) );
  NAND2_X2 MULT_mult_6_U2554 ( .A1(MULT_mult_6_SUMB_15__10_), .A2(
        MULT_mult_6_net121214), .ZN(MULT_mult_6_net79981) );
  NAND3_X2 MULT_mult_6_U2553 ( .A1(MULT_mult_6_net79980), .A2(
        MULT_mult_6_net79981), .A3(MULT_mult_6_n805), .ZN(
        MULT_mult_6_CARRYB_16__9_) );
  NAND2_X1 MULT_mult_6_U2552 ( .A1(MULT_mult_6_ab_17__9_), .A2(
        MULT_mult_6_CARRYB_16__9_), .ZN(MULT_mult_6_net80814) );
  NOR2_X1 MULT_mult_6_U2551 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net70461), .ZN(MULT_mult_6_ab_17__9_) );
  INV_X1 MULT_mult_6_U2550 ( .A(MULT_mult_6_ab_17__9_), .ZN(
        MULT_mult_6_net120656) );
  INV_X4 MULT_mult_6_U2549 ( .A(MULT_mult_6_net84208), .ZN(
        MULT_mult_6_net87944) );
  NAND2_X4 MULT_mult_6_U2548 ( .A1(MULT_mult_6_net120657), .A2(
        MULT_mult_6_n804), .ZN(MULT_mult_6_net84208) );
  NAND3_X2 MULT_mult_6_U2547 ( .A1(MULT_mult_6_net80667), .A2(
        MULT_mult_6_net80668), .A3(MULT_mult_6_net149917), .ZN(
        MULT_mult_6_net93672) );
  NAND3_X2 MULT_mult_6_U2546 ( .A1(MULT_mult_6_net80668), .A2(
        MULT_mult_6_net80667), .A3(MULT_mult_6_net149917), .ZN(
        MULT_mult_6_CARRYB_29__1_) );
  NAND2_X4 MULT_mult_6_U2545 ( .A1(MULT_mult_6_SUMB_3__17_), .A2(
        MULT_mult_6_ab_4__16_), .ZN(MULT_mult_6_net80836) );
  NOR2_X2 MULT_mult_6_U2544 ( .A1(MULT_mult_6_net88344), .A2(
        MULT_mult_6_net119855), .ZN(MULT_mult_6_ab_4__16_) );
  NAND2_X2 MULT_mult_6_U2543 ( .A1(MULT_mult_6_CARRYB_2__17_), .A2(
        MULT_mult_6_ab_3__17_), .ZN(MULT_mult_6_n800) );
  INV_X1 MULT_mult_6_U2542 ( .A(MULT_mult_6_ab_3__17_), .ZN(MULT_mult_6_n798)
         );
  NAND2_X4 MULT_mult_6_U2541 ( .A1(MULT_mult_6_n798), .A2(MULT_mult_6_n799), 
        .ZN(MULT_mult_6_n801) );
  XNOR2_X2 MULT_mult_6_U2540 ( .A(MULT_mult_6_n802), .B(
        MULT_mult_6_SUMB_2__18_), .ZN(MULT_mult_6_SUMB_3__17_) );
  XNOR2_X2 MULT_mult_6_U2539 ( .A(MULT_mult_6_n802), .B(
        MULT_mult_6_SUMB_2__18_), .ZN(MULT_mult_6_net124367) );
  NAND2_X4 MULT_mult_6_U2538 ( .A1(MULT_mult_6_n800), .A2(MULT_mult_6_n801), 
        .ZN(MULT_mult_6_n802) );
  INV_X4 MULT_mult_6_U2537 ( .A(MULT_mult_6_ab_5__15_), .ZN(
        MULT_mult_6_net119953) );
  XNOR2_X2 MULT_mult_6_U2536 ( .A(MULT_mult_6_net88079), .B(
        MULT_mult_6_net119953), .ZN(MULT_mult_6_net80834) );
  XNOR2_X2 MULT_mult_6_U2535 ( .A(MULT_mult_6_net88079), .B(
        MULT_mult_6_ab_5__15_), .ZN(MULT_mult_6_net119976) );
  NAND2_X1 MULT_mult_6_U2534 ( .A1(MULT_mult_6_net88881), .A2(
        MULT_mult_6_ab_7__14_), .ZN(MULT_mult_6_net81365) );
  INV_X4 MULT_mult_6_U2533 ( .A(MULT_mult_6_net88880), .ZN(
        MULT_mult_6_net88881) );
  XNOR2_X2 MULT_mult_6_U2532 ( .A(MULT_mult_6_n797), .B(MULT_mult_6_net93800), 
        .ZN(MULT_mult_6_net89356) );
  NAND2_X4 MULT_mult_6_U2531 ( .A1(MULT_mult_6_net87066), .A2(
        MULT_mult_6_net87065), .ZN(MULT_mult_6_net87068) );
  INV_X8 MULT_mult_6_U2530 ( .A(MULT_mult_6_CARRYB_7__13_), .ZN(
        MULT_mult_6_net87066) );
  INV_X2 MULT_mult_6_U2529 ( .A(MULT_mult_6_net87066), .ZN(
        MULT_mult_6_net88943) );
  NAND3_X2 MULT_mult_6_U2528 ( .A1(MULT_mult_6_net81372), .A2(
        MULT_mult_6_net81371), .A3(MULT_mult_6_n555), .ZN(MULT_mult_6_net84447) );
  NAND3_X2 MULT_mult_6_U2527 ( .A1(MULT_mult_6_net81372), .A2(
        MULT_mult_6_net81371), .A3(MULT_mult_6_n555), .ZN(
        MULT_mult_6_CARRYB_8__13_) );
  INV_X1 MULT_mult_6_U2525 ( .A(MULT_mult_6_ab_27__2_), .ZN(
        MULT_mult_6_net83055) );
  NAND2_X4 MULT_mult_6_U2524 ( .A1(MULT_mult_6_net83054), .A2(
        MULT_mult_6_net83055), .ZN(MULT_mult_6_net83057) );
  NAND2_X4 MULT_mult_6_U2523 ( .A1(MULT_mult_6_net83057), .A2(
        MULT_mult_6_net93918), .ZN(MULT_mult_6_net80927) );
  NAND3_X2 MULT_mult_6_U2522 ( .A1(MULT_mult_6_net80992), .A2(
        MULT_mult_6_net80991), .A3(MULT_mult_6_net80990), .ZN(
        MULT_mult_6_net123363) );
  NAND2_X4 MULT_mult_6_U2521 ( .A1(MULT_mult_6_n199), .A2(
        MULT_mult_6_net121451), .ZN(MULT_mult_6_SUMB_25__3_) );
  NAND3_X2 MULT_mult_6_U2520 ( .A1(MULT_mult_6_net81058), .A2(
        MULT_mult_6_net81057), .A3(MULT_mult_6_net81056), .ZN(
        MULT_mult_6_CARRYB_12__10_) );
  INV_X4 MULT_mult_6_U2519 ( .A(MULT_mult_6_CARRYB_12__10_), .ZN(
        MULT_mult_6_n795) );
  NAND2_X4 MULT_mult_6_U2518 ( .A1(MULT_mult_6_n796), .A2(
        MULT_mult_6_SUMB_12__11_), .ZN(MULT_mult_6_n794) );
  NAND2_X4 MULT_mult_6_U2517 ( .A1(MULT_mult_6_SUMB_12__11_), .A2(
        MULT_mult_6_ab_13__10_), .ZN(MULT_mult_6_n793) );
  NAND2_X2 MULT_mult_6_U2516 ( .A1(MULT_mult_6_ab_13__10_), .A2(
        MULT_mult_6_net124392), .ZN(MULT_mult_6_n792) );
  NAND3_X4 MULT_mult_6_U2515 ( .A1(MULT_mult_6_n794), .A2(MULT_mult_6_n793), 
        .A3(MULT_mult_6_n792), .ZN(MULT_mult_6_CARRYB_13__10_) );
  INV_X1 MULT_mult_6_U2514 ( .A(MULT_mult_6_ab_14__10_), .ZN(
        MULT_mult_6_net88407) );
  NOR2_X2 MULT_mult_6_U2513 ( .A1(MULT_mult_6_net91660), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__10_) );
  NAND2_X4 MULT_mult_6_U2512 ( .A1(MULT_mult_6_net82160), .A2(
        MULT_mult_6_net88410), .ZN(MULT_mult_6_net84163) );
  NAND2_X4 MULT_mult_6_U2511 ( .A1(MULT_mult_6_CARRYB_13__10_), .A2(
        MULT_mult_6_ab_14__10_), .ZN(MULT_mult_6_net82160) );
  NAND2_X2 MULT_mult_6_U2510 ( .A1(MULT_mult_6_net88668), .A2(
        MULT_mult_6_CARRYB_14__10_), .ZN(MULT_mult_6_net82561) );
  NAND2_X1 MULT_mult_6_U2509 ( .A1(MULT_mult_6_CARRYB_14__10_), .A2(
        MULT_mult_6_ab_15__10_), .ZN(MULT_mult_6_net82559) );
  XNOR2_X2 MULT_mult_6_U2508 ( .A(MULT_mult_6_CARRYB_14__10_), .B(
        MULT_mult_6_ab_15__10_), .ZN(MULT_mult_6_net86799) );
  NAND3_X4 MULT_mult_6_U2507 ( .A1(MULT_mult_6_net82162), .A2(
        MULT_mult_6_net82161), .A3(MULT_mult_6_net82160), .ZN(
        MULT_mult_6_CARRYB_14__10_) );
  XNOR2_X2 MULT_mult_6_U2506 ( .A(MULT_mult_6_net93277), .B(
        MULT_mult_6_net82263), .ZN(MULT_mult_6_net93756) );
  XNOR2_X2 MULT_mult_6_U2505 ( .A(MULT_mult_6_net93277), .B(
        MULT_mult_6_net82263), .ZN(MULT_mult_6_net87942) );
  NAND2_X2 MULT_mult_6_U2504 ( .A1(MULT_mult_6_net93277), .A2(
        MULT_mult_6_SUMB_12__12_), .ZN(MULT_mult_6_net120649) );
  XNOR2_X2 MULT_mult_6_U2503 ( .A(MULT_mult_6_net88906), .B(
        MULT_mult_6_SUMB_17__9_), .ZN(MULT_mult_6_net88702) );
  XNOR2_X2 MULT_mult_6_U2502 ( .A(MULT_mult_6_net84349), .B(
        MULT_mult_6_SUMB_17__9_), .ZN(MULT_mult_6_SUMB_18__8_) );
  XNOR2_X2 MULT_mult_6_U2501 ( .A(MULT_mult_6_CARRYB_17__8_), .B(
        MULT_mult_6_ab_18__8_), .ZN(MULT_mult_6_net84349) );
  XNOR2_X2 MULT_mult_6_U2500 ( .A(MULT_mult_6_ab_18__8_), .B(
        MULT_mult_6_CARRYB_17__8_), .ZN(MULT_mult_6_net88906) );
  NAND2_X2 MULT_mult_6_U2499 ( .A1(MULT_mult_6_SUMB_17__9_), .A2(
        MULT_mult_6_ab_18__8_), .ZN(MULT_mult_6_net81559) );
  NAND2_X2 MULT_mult_6_U2498 ( .A1(MULT_mult_6_SUMB_17__9_), .A2(
        MULT_mult_6_CARRYB_17__8_), .ZN(MULT_mult_6_net81560) );
  NAND2_X1 MULT_mult_6_U2497 ( .A1(MULT_mult_6_ab_18__8_), .A2(
        MULT_mult_6_CARRYB_17__8_), .ZN(MULT_mult_6_n791) );
  NAND3_X4 MULT_mult_6_U2496 ( .A1(MULT_mult_6_net81559), .A2(
        MULT_mult_6_net81560), .A3(MULT_mult_6_n791), .ZN(
        MULT_mult_6_CARRYB_18__8_) );
  NOR2_X4 MULT_mult_6_U2495 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net70457), .ZN(MULT_mult_6_ab_19__8_) );
  NAND2_X4 MULT_mult_6_U2494 ( .A1(MULT_mult_6_SUMB_12__12_), .A2(
        MULT_mult_6_ab_13__11_), .ZN(MULT_mult_6_net82158) );
  NAND3_X4 MULT_mult_6_U2493 ( .A1(MULT_mult_6_net82158), .A2(
        MULT_mult_6_net82159), .A3(MULT_mult_6_n97), .ZN(
        MULT_mult_6_CARRYB_13__11_) );
  NAND2_X4 MULT_mult_6_U2492 ( .A1(MULT_mult_6_CARRYB_12__11_), .A2(
        MULT_mult_6_ab_13__11_), .ZN(MULT_mult_6_net87936) );
  INV_X2 MULT_mult_6_U2491 ( .A(MULT_mult_6_ab_13__11_), .ZN(
        MULT_mult_6_net87934) );
  INV_X8 MULT_mult_6_U2490 ( .A(MULT_mult_6_CARRYB_12__11_), .ZN(
        MULT_mult_6_net87935) );
  NAND2_X4 MULT_mult_6_U2489 ( .A1(MULT_mult_6_net87936), .A2(
        MULT_mult_6_net87937), .ZN(MULT_mult_6_net93277) );
  NAND2_X4 MULT_mult_6_U2488 ( .A1(MULT_mult_6_net87935), .A2(
        MULT_mult_6_net87934), .ZN(MULT_mult_6_net87937) );
  NAND2_X2 MULT_mult_6_U2487 ( .A1(MULT_mult_6_n790), .A2(MULT_mult_6_net89026), .ZN(MULT_mult_6_n787) );
  INV_X2 MULT_mult_6_U2486 ( .A(MULT_mult_6_n785), .ZN(MULT_mult_6_n790) );
  INV_X2 MULT_mult_6_U2485 ( .A(MULT_mult_6_net89026), .ZN(MULT_mult_6_n786)
         );
  NAND2_X2 MULT_mult_6_U2484 ( .A1(MULT_mult_6_n786), .A2(MULT_mult_6_n785), 
        .ZN(MULT_mult_6_n788) );
  NAND2_X4 MULT_mult_6_U2483 ( .A1(MULT_mult_6_n787), .A2(MULT_mult_6_n788), 
        .ZN(MULT_mult_6_SUMB_12__12_) );
  NAND2_X2 MULT_mult_6_U2482 ( .A1(MULT_mult_6_net87937), .A2(
        MULT_mult_6_net87936), .ZN(MULT_mult_6_net84059) );
  INV_X4 MULT_mult_6_U2481 ( .A(MULT_mult_6_net84059), .ZN(
        MULT_mult_6_net120647) );
  NAND2_X4 MULT_mult_6_U2480 ( .A1(MULT_mult_6_net120649), .A2(
        MULT_mult_6_n789), .ZN(MULT_mult_6_SUMB_13__11_) );
  NAND2_X4 MULT_mult_6_U2479 ( .A1(MULT_mult_6_net120647), .A2(
        MULT_mult_6_net120648), .ZN(MULT_mult_6_n789) );
  NAND2_X4 MULT_mult_6_U2478 ( .A1(MULT_mult_6_net124635), .A2(
        MULT_mult_6_ab_23__4_), .ZN(MULT_mult_6_n782) );
  NAND2_X2 MULT_mult_6_U2477 ( .A1(MULT_mult_6_ab_23__4_), .A2(
        MULT_mult_6_CARRYB_22__4_), .ZN(MULT_mult_6_n783) );
  NAND3_X4 MULT_mult_6_U2476 ( .A1(MULT_mult_6_net80290), .A2(MULT_mult_6_n782), .A3(MULT_mult_6_n783), .ZN(MULT_mult_6_CARRYB_23__4_) );
  NOR2_X4 MULT_mult_6_U2475 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70445), .ZN(MULT_mult_6_ab_25__4_) );
  NAND2_X4 MULT_mult_6_U2474 ( .A1(MULT_mult_6_CARRYB_23__4_), .A2(
        MULT_mult_6_ab_24__4_), .ZN(MULT_mult_6_net79907) );
  NOR2_X4 MULT_mult_6_U2473 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70447), .ZN(MULT_mult_6_ab_24__4_) );
  INV_X8 MULT_mult_6_U2472 ( .A(MULT_mult_6_CARRYB_23__4_), .ZN(
        MULT_mult_6_net84000) );
  INV_X2 MULT_mult_6_U2471 ( .A(MULT_mult_6_ab_24__4_), .ZN(
        MULT_mult_6_net84001) );
  NAND2_X4 MULT_mult_6_U2470 ( .A1(MULT_mult_6_net79907), .A2(MULT_mult_6_n784), .ZN(MULT_mult_6_net80021) );
  NAND2_X4 MULT_mult_6_U2469 ( .A1(MULT_mult_6_net84000), .A2(
        MULT_mult_6_net84001), .ZN(MULT_mult_6_n784) );
  NAND2_X1 MULT_mult_6_U2468 ( .A1(MULT_mult_6_ab_21__6_), .A2(
        MULT_mult_6_CARRYB_20__6_), .ZN(MULT_mult_6_net80674) );
  NAND2_X1 MULT_mult_6_U2467 ( .A1(MULT_mult_6_ab_21__6_), .A2(
        MULT_mult_6_net149530), .ZN(MULT_mult_6_net80675) );
  NAND2_X1 MULT_mult_6_U2466 ( .A1(MULT_mult_6_net149530), .A2(MULT_mult_6_n69), .ZN(MULT_mult_6_net80676) );
  NAND2_X4 MULT_mult_6_U2465 ( .A1(MULT_mult_6_net81553), .A2(
        MULT_mult_6_net81552), .ZN(MULT_mult_6_net81555) );
  INV_X4 MULT_mult_6_U2464 ( .A(MULT_mult_6_net81042), .ZN(
        MULT_mult_6_net81552) );
  INV_X1 MULT_mult_6_U2463 ( .A(MULT_mult_6_ab_21__6_), .ZN(
        MULT_mult_6_net81042) );
  NAND2_X4 MULT_mult_6_U2462 ( .A1(MULT_mult_6_net81555), .A2(MULT_mult_6_n781), .ZN(MULT_mult_6_net87681) );
  NAND2_X2 MULT_mult_6_U2461 ( .A1(MULT_mult_6_net90818), .A2(
        MULT_mult_6_ab_20__7_), .ZN(MULT_mult_6_net80672) );
  NAND2_X1 MULT_mult_6_U2460 ( .A1(MULT_mult_6_ab_20__7_), .A2(
        MULT_mult_6_net91001), .ZN(MULT_mult_6_net80671) );
  INV_X4 MULT_mult_6_U2459 ( .A(MULT_mult_6_CARRYB_19__7_), .ZN(
        MULT_mult_6_n778) );
  NAND2_X2 MULT_mult_6_U2458 ( .A1(MULT_mult_6_ab_20__7_), .A2(
        MULT_mult_6_CARRYB_19__7_), .ZN(MULT_mult_6_n779) );
  INV_X4 MULT_mult_6_U2457 ( .A(MULT_mult_6_ab_20__7_), .ZN(
        MULT_mult_6_net93279) );
  NAND2_X4 MULT_mult_6_U2456 ( .A1(MULT_mult_6_n778), .A2(MULT_mult_6_net93279), .ZN(MULT_mult_6_n780) );
  NAND2_X4 MULT_mult_6_U2455 ( .A1(MULT_mult_6_n779), .A2(MULT_mult_6_n780), 
        .ZN(MULT_mult_6_net90022) );
  INV_X4 MULT_mult_6_U2454 ( .A(MULT_mult_6_CARRYB_18__8_), .ZN(
        MULT_mult_6_net123291) );
  INV_X1 MULT_mult_6_U2453 ( .A(MULT_mult_6_ab_19__8_), .ZN(MULT_mult_6_n775)
         );
  INV_X4 MULT_mult_6_U2451 ( .A(MULT_mult_6_net88699), .ZN(
        MULT_mult_6_net87391) );
  NAND2_X4 MULT_mult_6_U2450 ( .A1(MULT_mult_6_net89109), .A2(
        MULT_mult_6_net123363), .ZN(MULT_mult_6_net79882) );
  XNOR2_X2 MULT_mult_6_U2449 ( .A(MULT_mult_6_net80927), .B(
        MULT_mult_6_net89104), .ZN(MULT_mult_6_net89109) );
  NAND3_X4 MULT_mult_6_U2448 ( .A1(MULT_mult_6_net79882), .A2(
        MULT_mult_6_net79881), .A3(MULT_mult_6_net79880), .ZN(
        MULT_mult_6_CARRYB_28__1_) );
  NAND2_X1 MULT_mult_6_U2447 ( .A1(MULT_mult_6_ab_4__6_), .A2(
        MULT_mult_6_SUMB_3__7_), .ZN(MULT_mult_6_net88207) );
  XNOR2_X2 MULT_mult_6_U2446 ( .A(MULT_mult_6_n774), .B(MULT_mult_6_SUMB_3__7_), .ZN(MULT_mult_6_SUMB_4__6_) );
  CLKBUF_X3 MULT_mult_6_U2445 ( .A(MULT_mult_6_SUMB_4__6_), .Z(
        MULT_mult_6_net125691) );
  XNOR2_X2 MULT_mult_6_U2444 ( .A(MULT_mult_6_net92884), .B(
        MULT_mult_6_SUMB_5__5_), .ZN(MULT_mult_6_SUMB_6__4_) );
  NAND2_X1 MULT_mult_6_U2443 ( .A1(MULT_mult_6_ab_7__3_), .A2(
        MULT_mult_6_CARRYB_6__3_), .ZN(MULT_mult_6_n771) );
  NAND2_X2 MULT_mult_6_U2442 ( .A1(MULT_mult_6_ab_7__3_), .A2(
        MULT_mult_6_SUMB_6__4_), .ZN(MULT_mult_6_n772) );
  NAND2_X2 MULT_mult_6_U2441 ( .A1(MULT_mult_6_CARRYB_6__3_), .A2(
        MULT_mult_6_SUMB_6__4_), .ZN(MULT_mult_6_n773) );
  NAND3_X2 MULT_mult_6_U2440 ( .A1(MULT_mult_6_n771), .A2(MULT_mult_6_n772), 
        .A3(MULT_mult_6_n773), .ZN(MULT_mult_6_CARRYB_7__3_) );
  NAND2_X2 MULT_mult_6_U2439 ( .A1(MULT_mult_6_ab_6__4_), .A2(MULT_mult_6_n343), .ZN(MULT_mult_6_net88198) );
  NAND2_X2 MULT_mult_6_U2438 ( .A1(MULT_mult_6_ab_6__4_), .A2(
        MULT_mult_6_SUMB_5__5_), .ZN(MULT_mult_6_net88199) );
  NAND2_X2 MULT_mult_6_U2437 ( .A1(MULT_mult_6_ab_5__5_), .A2(
        MULT_mult_6_SUMB_4__6_), .ZN(MULT_mult_6_net88210) );
  NOR2_X4 MULT_mult_6_U2436 ( .A1(MULT_mult_6_net77898), .A2(
        MULT_mult_6_net77946), .ZN(MULT_mult_6_ab_5__5_) );
  XNOR2_X2 MULT_mult_6_U2435 ( .A(MULT_mult_6_net89958), .B(
        MULT_mult_6_net125691), .ZN(MULT_mult_6_SUMB_5__5_) );
  NAND2_X2 MULT_mult_6_U2434 ( .A1(MULT_mult_6_SUMB_22__3_), .A2(
        MULT_mult_6_ab_23__2_), .ZN(MULT_mult_6_net80254) );
  NAND2_X2 MULT_mult_6_U2433 ( .A1(MULT_mult_6_n394), .A2(
        MULT_mult_6_SUMB_22__3_), .ZN(MULT_mult_6_net80255) );
  XNOR2_X2 MULT_mult_6_U2432 ( .A(MULT_mult_6_net121523), .B(MULT_mult_6_n564), 
        .ZN(MULT_mult_6_SUMB_23__2_) );
  XNOR2_X2 MULT_mult_6_U2431 ( .A(MULT_mult_6_net121523), .B(MULT_mult_6_n564), 
        .ZN(MULT_mult_6_net122156) );
  NOR2_X1 MULT_mult_6_U2430 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__2_) );
  XNOR2_X2 MULT_mult_6_U2429 ( .A(MULT_mult_6_SUMB_9__4_), .B(
        MULT_mult_6_ab_10__3_), .ZN(MULT_mult_6_n770) );
  NAND2_X2 MULT_mult_6_U2428 ( .A1(MULT_mult_6_ab_11__2_), .A2(
        MULT_mult_6_SUMB_10__3_), .ZN(MULT_mult_6_net81616) );
  XNOR2_X2 MULT_mult_6_U2427 ( .A(MULT_mult_6_n770), .B(
        MULT_mult_6_CARRYB_9__3_), .ZN(MULT_mult_6_SUMB_10__3_) );
  NAND2_X2 MULT_mult_6_U2426 ( .A1(MULT_mult_6_n343), .A2(
        MULT_mult_6_SUMB_5__5_), .ZN(MULT_mult_6_net88200) );
  NAND3_X4 MULT_mult_6_U2425 ( .A1(MULT_mult_6_net88198), .A2(
        MULT_mult_6_net88199), .A3(MULT_mult_6_net88200), .ZN(
        MULT_mult_6_CARRYB_6__4_) );
  XNOR2_X2 MULT_mult_6_U2424 ( .A(MULT_mult_6_CARRYB_5__5_), .B(
        MULT_mult_6_ab_6__5_), .ZN(MULT_mult_6_n768) );
  XNOR2_X2 MULT_mult_6_U2423 ( .A(MULT_mult_6_SUMB_5__6_), .B(MULT_mult_6_n768), .ZN(MULT_mult_6_SUMB_6__5_) );
  INV_X32 MULT_mult_6_U2422 ( .A(n10929), .ZN(MULT_mult_6_net77892) );
  XNOR2_X2 MULT_mult_6_U2421 ( .A(MULT_mult_6_SUMB_6__6_), .B(
        MULT_mult_6_ab_7__5_), .ZN(MULT_mult_6_n769) );
  XNOR2_X2 MULT_mult_6_U2420 ( .A(MULT_mult_6_n769), .B(
        MULT_mult_6_CARRYB_6__5_), .ZN(MULT_mult_6_SUMB_7__5_) );
  XNOR2_X2 MULT_mult_6_U2419 ( .A(MULT_mult_6_CARRYB_8__4_), .B(
        MULT_mult_6_ab_9__4_), .ZN(MULT_mult_6_net82601) );
  NOR2_X4 MULT_mult_6_U2418 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__2_) );
  XNOR2_X2 MULT_mult_6_U2417 ( .A(MULT_mult_6_n51), .B(MULT_mult_6_ab_13__3_), 
        .ZN(MULT_mult_6_n767) );
  XNOR2_X2 MULT_mult_6_U2416 ( .A(MULT_mult_6_SUMB_12__4_), .B(
        MULT_mult_6_n767), .ZN(MULT_mult_6_SUMB_13__3_) );
  NAND2_X2 MULT_mult_6_U2415 ( .A1(MULT_mult_6_ab_13__2_), .A2(
        MULT_mult_6_SUMB_12__3_), .ZN(MULT_mult_6_n763) );
  NAND2_X2 MULT_mult_6_U2414 ( .A1(MULT_mult_6_n19), .A2(
        MULT_mult_6_SUMB_12__3_), .ZN(MULT_mult_6_n764) );
  NAND2_X4 MULT_mult_6_U2413 ( .A1(MULT_mult_6_ab_14__2_), .A2(
        MULT_mult_6_CARRYB_13__2_), .ZN(MULT_mult_6_net81780) );
  NAND3_X4 MULT_mult_6_U2412 ( .A1(MULT_mult_6_n764), .A2(MULT_mult_6_n763), 
        .A3(MULT_mult_6_n762), .ZN(MULT_mult_6_CARRYB_13__2_) );
  INV_X16 MULT_mult_6_U2411 ( .A(aluA[16]), .ZN(MULT_mult_6_net70465) );
  NAND2_X2 MULT_mult_6_U2410 ( .A1(MULT_mult_6_SUMB_13__2_), .A2(
        MULT_mult_6_ab_14__1_), .ZN(MULT_mult_6_n766) );
  XOR2_X1 MULT_mult_6_U2409 ( .A(MULT_mult_6_net86649), .B(
        MULT_mult_6_SUMB_15__1_), .Z(multOut[15]) );
  NAND2_X2 MULT_mult_6_U2408 ( .A1(MULT_mult_6_ab_16__0_), .A2(
        MULT_mult_6_SUMB_15__1_), .ZN(MULT_mult_6_net86651) );
  NAND2_X2 MULT_mult_6_U2407 ( .A1(MULT_mult_6_CARRYB_15__0_), .A2(
        MULT_mult_6_SUMB_15__1_), .ZN(MULT_mult_6_net86652) );
  NOR2_X2 MULT_mult_6_U2406 ( .A1(MULT_mult_6_net124610), .A2(
        MULT_mult_6_net70492), .ZN(MULT_mult_6_ab_0__29_) );
  XNOR2_X2 MULT_mult_6_U2405 ( .A(MULT_mult_6_ab_1__6_), .B(
        MULT_mult_6_ab_0__7_), .ZN(MULT_mult_6__UDW__112739_net78703) );
  NOR2_X2 MULT_mult_6_U2404 ( .A1(MULT_mult_6_net77906), .A2(
        MULT_mult_6_net77970), .ZN(MULT_mult_6_ab_2__6_) );
  XNOR2_X1 MULT_mult_6_U2403 ( .A(MULT_mult_6_ab_1__7_), .B(
        MULT_mult_6_ab_0__8_), .ZN(MULT_mult_6_n757) );
  XNOR2_X2 MULT_mult_6_U2402 ( .A(MULT_mult_6_SUMB_1__7_), .B(MULT_mult_6_n758), .ZN(MULT_mult_6_SUMB_2__6_) );
  INV_X4 MULT_mult_6_U2401 ( .A(MULT_mult_6_n757), .ZN(MULT_mult_6_SUMB_1__7_)
         );
  NAND2_X2 MULT_mult_6_U2400 ( .A1(MULT_mult_6_n350), .A2(
        MULT_mult_6_SUMB_1__7_), .ZN(MULT_mult_6_n759) );
  NAND2_X1 MULT_mult_6_U2399 ( .A1(MULT_mult_6_ab_2__6_), .A2(MULT_mult_6_n350), .ZN(MULT_mult_6_n761) );
  NAND2_X2 MULT_mult_6_U2398 ( .A1(MULT_mult_6_ab_3__6_), .A2(
        MULT_mult_6_CARRYB_2__6_), .ZN(MULT_mult_6_net84924) );
  NAND3_X2 MULT_mult_6_U2397 ( .A1(MULT_mult_6_n759), .A2(MULT_mult_6_n760), 
        .A3(MULT_mult_6_n761), .ZN(MULT_mult_6_CARRYB_2__6_) );
  NAND2_X2 MULT_mult_6_U2396 ( .A1(MULT_mult_6_ab_18__2_), .A2(
        MULT_mult_6_CARRYB_17__2_), .ZN(MULT_mult_6_net81110) );
  NAND2_X2 MULT_mult_6_U2395 ( .A1(MULT_mult_6_ab_18__2_), .A2(
        MULT_mult_6_SUMB_17__3_), .ZN(MULT_mult_6_net81111) );
  NAND2_X2 MULT_mult_6_U2394 ( .A1(MULT_mult_6_CARRYB_17__2_), .A2(
        MULT_mult_6_SUMB_17__3_), .ZN(MULT_mult_6_net81112) );
  NOR2_X4 MULT_mult_6_U2393 ( .A1(MULT_mult_6_net77868), .A2(
        MULT_mult_6_net70457), .ZN(MULT_mult_6_ab_19__1_) );
  BUF_X8 MULT_mult_6_U2392 ( .A(MULT_mult_6_SUMB_17__3_), .Z(MULT_mult_6_n755)
         );
  XNOR2_X2 MULT_mult_6_U2391 ( .A(MULT_mult_6_net93676), .B(MULT_mult_6_n359), 
        .ZN(MULT_mult_6_SUMB_19__1_) );
  XNOR2_X2 MULT_mult_6_U2390 ( .A(MULT_mult_6_n754), .B(MULT_mult_6_n755), 
        .ZN(MULT_mult_6_SUMB_18__2_) );
  NAND2_X2 MULT_mult_6_U2389 ( .A1(MULT_mult_6_ab_19__1_), .A2(
        MULT_mult_6_SUMB_18__2_), .ZN(MULT_mult_6_n756) );
  NAND2_X2 MULT_mult_6_U2388 ( .A1(MULT_mult_6_CARRYB_19__1_), .A2(
        MULT_mult_6_SUMB_19__2_), .ZN(MULT_mult_6_net80852) );
  NAND2_X2 MULT_mult_6_U2387 ( .A1(MULT_mult_6_ab_20__1_), .A2(
        MULT_mult_6_CARRYB_19__1_), .ZN(MULT_mult_6_net80850) );
  NAND3_X2 MULT_mult_6_U2386 ( .A1(MULT_mult_6_net81095), .A2(MULT_mult_6_n756), .A3(MULT_mult_6_net81097), .ZN(MULT_mult_6_CARRYB_19__1_) );
  NAND2_X2 MULT_mult_6_U2385 ( .A1(MULT_mult_6_SUMB_21__3_), .A2(
        MULT_mult_6_n372), .ZN(MULT_mult_6_net80924) );
  XNOR2_X2 MULT_mult_6_U2384 ( .A(MULT_mult_6_SUMB_21__2_), .B(
        MULT_mult_6_ab_22__1_), .ZN(MULT_mult_6_n753) );
  XNOR2_X2 MULT_mult_6_U2383 ( .A(MULT_mult_6_n753), .B(
        MULT_mult_6_CARRYB_21__1_), .ZN(MULT_mult_6_SUMB_22__1_) );
  XNOR2_X2 MULT_mult_6_U2382 ( .A(MULT_mult_6_CARRYB_21__2_), .B(
        MULT_mult_6_ab_22__2_), .ZN(MULT_mult_6_n749) );
  INV_X1 MULT_mult_6_U2381 ( .A(MULT_mult_6_SUMB_22__2_), .ZN(
        MULT_mult_6_net83357) );
  XNOR2_X2 MULT_mult_6_U2380 ( .A(MULT_mult_6_SUMB_21__3_), .B(
        MULT_mult_6_n749), .ZN(MULT_mult_6_SUMB_22__2_) );
  NAND3_X2 MULT_mult_6_U2378 ( .A1(MULT_mult_6_net82541), .A2(
        MULT_mult_6_net82542), .A3(MULT_mult_6_net82543), .ZN(MULT_mult_6_n748) );
  NAND2_X2 MULT_mult_6_U2377 ( .A1(MULT_mult_6_CARRYB_21__1_), .A2(
        MULT_mult_6_SUMB_21__2_), .ZN(MULT_mult_6_net82541) );
  XNOR2_X2 MULT_mult_6_U2376 ( .A(MULT_mult_6_n748), .B(MULT_mult_6_ab_23__1_), 
        .ZN(MULT_mult_6_net93713) );
  NOR2_X2 MULT_mult_6_U2375 ( .A1(MULT_mult_6_net77866), .A2(
        MULT_mult_6_net70449), .ZN(MULT_mult_6_ab_23__1_) );
  NAND2_X2 MULT_mult_6_U2374 ( .A1(MULT_mult_6_n748), .A2(
        MULT_mult_6_SUMB_22__2_), .ZN(MULT_mult_6_n750) );
  NAND3_X2 MULT_mult_6_U2373 ( .A1(MULT_mult_6_net82541), .A2(
        MULT_mult_6_net82542), .A3(MULT_mult_6_net82543), .ZN(
        MULT_mult_6_CARRYB_22__1_) );
  NAND2_X2 MULT_mult_6_U2372 ( .A1(MULT_mult_6_ab_23__1_), .A2(
        MULT_mult_6_CARRYB_22__1_), .ZN(MULT_mult_6_n752) );
  NAND3_X2 MULT_mult_6_U2371 ( .A1(MULT_mult_6_n750), .A2(MULT_mult_6_n751), 
        .A3(MULT_mult_6_n752), .ZN(MULT_mult_6_CARRYB_23__1_) );
  NOR2_X4 MULT_mult_6_U2370 ( .A1(MULT_mult_6_net77868), .A2(
        MULT_mult_6_net70463), .ZN(MULT_mult_6_ab_16__1_) );
  XOR2_X1 MULT_mult_6_U2369 ( .A(MULT_mult_6_ab_17__0_), .B(
        MULT_mult_6_SUMB_16__1_), .Z(MULT_mult_6_net86653) );
  NAND2_X2 MULT_mult_6_U2368 ( .A1(MULT_mult_6_SUMB_16__1_), .A2(
        MULT_mult_6_CARRYB_16__0_), .ZN(MULT_mult_6_net86656) );
  XNOR2_X2 MULT_mult_6_U2367 ( .A(MULT_mult_6_CARRYB_16__1_), .B(
        MULT_mult_6_net88712), .ZN(MULT_mult_6_net82532) );
  XNOR2_X2 MULT_mult_6_U2366 ( .A(MULT_mult_6_n742), .B(
        MULT_mult_6_CARRYB_16__2_), .ZN(MULT_mult_6_SUMB_17__2_) );
  NAND2_X2 MULT_mult_6_U2365 ( .A1(MULT_mult_6_CARRYB_17__1_), .A2(
        MULT_mult_6_SUMB_17__2_), .ZN(MULT_mult_6_n747) );
  XNOR2_X1 MULT_mult_6_U2364 ( .A(MULT_mult_6_CARRYB_18__1_), .B(
        MULT_mult_6_ab_19__1_), .ZN(MULT_mult_6_net93676) );
  NAND2_X2 MULT_mult_6_U2363 ( .A1(MULT_mult_6_ab_19__1_), .A2(
        MULT_mult_6_CARRYB_18__1_), .ZN(MULT_mult_6_net81095) );
  NOR2_X4 MULT_mult_6_U2362 ( .A1(MULT_mult_6_net77868), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__1_) );
  XNOR2_X2 MULT_mult_6_U2361 ( .A(MULT_mult_6_CARRYB_11__2_), .B(
        MULT_mult_6_ab_12__2_), .ZN(MULT_mult_6_n741) );
  XNOR2_X2 MULT_mult_6_U2360 ( .A(MULT_mult_6_n741), .B(
        MULT_mult_6_SUMB_11__3_), .ZN(MULT_mult_6_SUMB_12__2_) );
  NAND2_X2 MULT_mult_6_U2359 ( .A1(MULT_mult_6_CARRYB_10__1_), .A2(
        MULT_mult_6_ab_11__1_), .ZN(MULT_mult_6_n738) );
  NAND2_X2 MULT_mult_6_U2358 ( .A1(MULT_mult_6_ab_11__1_), .A2(
        MULT_mult_6_SUMB_10__2_), .ZN(MULT_mult_6_n739) );
  NAND2_X2 MULT_mult_6_U2357 ( .A1(MULT_mult_6_CARRYB_10__1_), .A2(
        MULT_mult_6_SUMB_10__2_), .ZN(MULT_mult_6_n740) );
  XNOR2_X2 MULT_mult_6_U2356 ( .A(MULT_mult_6_SUMB_10__3_), .B(
        MULT_mult_6_net122130), .ZN(MULT_mult_6_SUMB_11__2_) );
  NAND2_X2 MULT_mult_6_U2355 ( .A1(MULT_mult_6_CARRYB_12__1_), .A2(
        MULT_mult_6_ab_13__1_), .ZN(MULT_mult_6_net86129) );
  NAND2_X2 MULT_mult_6_U2354 ( .A1(MULT_mult_6_ab_13__1_), .A2(
        MULT_mult_6_SUMB_12__2_), .ZN(MULT_mult_6_n737) );
  NAND2_X2 MULT_mult_6_U2353 ( .A1(MULT_mult_6_CARRYB_12__1_), .A2(
        MULT_mult_6_SUMB_12__2_), .ZN(MULT_mult_6_net86131) );
  NAND2_X2 MULT_mult_6_U2352 ( .A1(MULT_mult_6_CARRYB_13__1_), .A2(
        MULT_mult_6_SUMB_13__2_), .ZN(MULT_mult_6_net86135) );
  NAND2_X2 MULT_mult_6_U2351 ( .A1(MULT_mult_6_ab_14__1_), .A2(
        MULT_mult_6_CARRYB_13__1_), .ZN(MULT_mult_6_net86134) );
  NAND3_X2 MULT_mult_6_U2350 ( .A1(MULT_mult_6_net86129), .A2(MULT_mult_6_n737), .A3(MULT_mult_6_net86131), .ZN(MULT_mult_6_CARRYB_13__1_) );
  INV_X16 MULT_mult_6_U2349 ( .A(MULT_mult_6_n26), .ZN(MULT_mult_6_net77970)
         );
  NOR2_X2 MULT_mult_6_U2348 ( .A1(MULT_mult_6_net77912), .A2(
        MULT_mult_6_net77970), .ZN(MULT_mult_6_ab_2__7_) );
  NAND2_X2 MULT_mult_6_U2347 ( .A1(MULT_mult_6_ab_0__8_), .A2(
        MULT_mult_6_ab_1__7_), .ZN(MULT_mult_6__UDW__112734_net78687) );
  INV_X4 MULT_mult_6_U2346 ( .A(MULT_mult_6__UDW__112734_net78687), .ZN(
        MULT_mult_6_CARRYB_1__7_) );
  XNOR2_X2 MULT_mult_6_U2345 ( .A(MULT_mult_6_ab_1__8_), .B(
        MULT_mult_6_ab_0__9_), .ZN(MULT_mult_6_n731) );
  INV_X4 MULT_mult_6_U2344 ( .A(MULT_mult_6_n731), .ZN(MULT_mult_6_SUMB_1__8_)
         );
  NAND2_X2 MULT_mult_6_U2343 ( .A1(MULT_mult_6_ab_3__7_), .A2(MULT_mult_6_n567), .ZN(MULT_mult_6_net84118) );
  NAND2_X2 MULT_mult_6_U2342 ( .A1(MULT_mult_6_net85036), .A2(MULT_mult_6_n567), .ZN(MULT_mult_6_net84116) );
  INV_X2 MULT_mult_6_U2341 ( .A(MULT_mult_6_SUMB_2__7_), .ZN(
        MULT_mult_6_net87961) );
  NAND2_X2 MULT_mult_6_U2340 ( .A1(MULT_mult_6_CARRYB_2__6_), .A2(
        MULT_mult_6_net87962), .ZN(MULT_mult_6_net84926) );
  NAND2_X2 MULT_mult_6_U2339 ( .A1(MULT_mult_6_ab_3__6_), .A2(
        MULT_mult_6_net87962), .ZN(MULT_mult_6_net84925) );
  NAND2_X2 MULT_mult_6_U2337 ( .A1(MULT_mult_6_ab_3__5_), .A2(
        MULT_mult_6_SUMB_2__6_), .ZN(MULT_mult_6_n733) );
  NAND2_X1 MULT_mult_6_U2336 ( .A1(MULT_mult_6_ab_3__5_), .A2(
        MULT_mult_6_CARRYB_2__5_), .ZN(MULT_mult_6_n734) );
  NAND2_X1 MULT_mult_6_U2334 ( .A1(MULT_mult_6_ab_4__5_), .A2(
        MULT_mult_6_CARRYB_3__5_), .ZN(MULT_mult_6_n735) );
  NAND2_X1 MULT_mult_6_U2333 ( .A1(MULT_mult_6_ab_4__5_), .A2(
        MULT_mult_6_SUMB_3__6_), .ZN(MULT_mult_6_net84928) );
  NAND2_X1 MULT_mult_6_U2332 ( .A1(MULT_mult_6_CARRYB_3__5_), .A2(
        MULT_mult_6_SUMB_3__6_), .ZN(MULT_mult_6_net84929) );
  NAND2_X2 MULT_mult_6_U2331 ( .A1(MULT_mult_6_CARRYB_4__5_), .A2(
        MULT_mult_6_SUMB_4__6_), .ZN(MULT_mult_6_net88211) );
  XNOR2_X1 MULT_mult_6_U2330 ( .A(MULT_mult_6_ab_5__5_), .B(
        MULT_mult_6_CARRYB_4__5_), .ZN(MULT_mult_6_net89958) );
  NAND2_X1 MULT_mult_6_U2329 ( .A1(MULT_mult_6_ab_5__5_), .A2(
        MULT_mult_6_CARRYB_4__5_), .ZN(MULT_mult_6_net88209) );
  NAND3_X2 MULT_mult_6_U2328 ( .A1(MULT_mult_6_n735), .A2(MULT_mult_6_net84928), .A3(MULT_mult_6_net84929), .ZN(MULT_mult_6_CARRYB_4__5_) );
  NOR2_X2 MULT_mult_6_U2327 ( .A1(MULT_mult_6_net147421), .A2(MULT_mult_6_n357), .ZN(MULT_mult_6_n719) );
  NAND2_X4 MULT_mult_6_U2326 ( .A1(MULT_mult_6_n711), .A2(MULT_mult_6_n712), 
        .ZN(MULT_mult_6_net147421) );
  INV_X2 MULT_mult_6_U2325 ( .A(MULT_mult_6_n716), .ZN(MULT_mult_6_n713) );
  AOI21_X4 MULT_mult_6_U2324 ( .B1(MULT_mult_6_n717), .B2(MULT_mult_6_n718), 
        .A(MULT_mult_6_net147444), .ZN(MULT_mult_6_n716) );
  INV_X1 MULT_mult_6_U2323 ( .A(MULT_mult_6_CARRYB_8__2_), .ZN(
        MULT_mult_6_n715) );
  INV_X8 MULT_mult_6_U2322 ( .A(MULT_mult_6_net147451), .ZN(
        MULT_mult_6_net147444) );
  NAND2_X4 MULT_mult_6_U2321 ( .A1(MULT_mult_6_n722), .A2(MULT_mult_6_n354), 
        .ZN(MULT_mult_6_n718) );
  NAND2_X1 MULT_mult_6_U2320 ( .A1(MULT_mult_6_ab_9__3_), .A2(
        MULT_mult_6_SUMB_8__4_), .ZN(MULT_mult_6_net82849) );
  INV_X2 MULT_mult_6_U2319 ( .A(MULT_mult_6_CARRYB_8__3_), .ZN(
        MULT_mult_6_n729) );
  INV_X4 MULT_mult_6_U2318 ( .A(MULT_mult_6_n729), .ZN(MULT_mult_6_n728) );
  INV_X2 MULT_mult_6_U2317 ( .A(MULT_mult_6_SUMB_8__3_), .ZN(MULT_mult_6_n727)
         );
  INV_X4 MULT_mult_6_U2316 ( .A(MULT_mult_6_n727), .ZN(MULT_mult_6_n726) );
  NAND2_X1 MULT_mult_6_U2315 ( .A1(MULT_mult_6_ab_9__3_), .A2(MULT_mult_6_n728), .ZN(MULT_mult_6_net82848) );
  XNOR2_X1 MULT_mult_6_U2314 ( .A(MULT_mult_6_ab_9__3_), .B(MULT_mult_6_n728), 
        .ZN(MULT_mult_6_n723) );
  OAI211_X1 MULT_mult_6_U2313 ( .C1(MULT_mult_6_net77878), .C2(
        MULT_mult_6_net70475), .A(MULT_mult_6_n711), .B(MULT_mult_6_n712), 
        .ZN(MULT_mult_6_n717) );
  INV_X32 MULT_mult_6_U2312 ( .A(n6005), .ZN(MULT_mult_6_net77878) );
  XNOR2_X2 MULT_mult_6_U2311 ( .A(MULT_mult_6_n726), .B(MULT_mult_6_ab_9__2_), 
        .ZN(MULT_mult_6_n725) );
  MUX2_X2 MULT_mult_6_U2310 ( .A(MULT_mult_6_n723), .B(MULT_mult_6_n356), .S(
        MULT_mult_6_SUMB_8__4_), .Z(MULT_mult_6_n722) );
  INV_X4 MULT_mult_6_U2309 ( .A(MULT_mult_6_n724), .ZN(MULT_mult_6_SUMB_9__2_)
         );
  XNOR2_X2 MULT_mult_6_U2308 ( .A(MULT_mult_6_n725), .B(MULT_mult_6_n715), 
        .ZN(MULT_mult_6_n724) );
  INV_X4 MULT_mult_6_U2307 ( .A(MULT_mult_6_n720), .ZN(MULT_mult_6_n721) );
  NAND2_X2 MULT_mult_6_U2306 ( .A1(MULT_mult_6_n726), .A2(MULT_mult_6_ab_9__2_), .ZN(MULT_mult_6_n711) );
  OAI21_X4 MULT_mult_6_U2305 ( .B1(MULT_mult_6_ab_9__2_), .B2(MULT_mult_6_n726), .A(MULT_mult_6_CARRYB_8__2_), .ZN(MULT_mult_6_n712) );
  XNOR2_X2 MULT_mult_6_U2304 ( .A(MULT_mult_6_n721), .B(MULT_mult_6_n718), 
        .ZN(MULT_mult_6_SUMB_10__2_) );
  XNOR2_X2 MULT_mult_6_U2303 ( .A(MULT_mult_6_n716), .B(MULT_mult_6_net85032), 
        .ZN(MULT_mult_6_net122130) );
  NOR2_X4 MULT_mult_6_U2302 ( .A1(MULT_mult_6_n719), .A2(MULT_mult_6_net147444), .ZN(MULT_mult_6_n720) );
  INV_X4 MULT_mult_6_U2301 ( .A(MULT_mult_6_ab_9__3_), .ZN(MULT_mult_6_n714)
         );
  NAND2_X2 MULT_mult_6_U2300 ( .A1(MULT_mult_6_n713), .A2(
        MULT_mult_6_SUMB_10__3_), .ZN(MULT_mult_6_net81615) );
  NAND2_X2 MULT_mult_6_U2299 ( .A1(MULT_mult_6_n713), .A2(
        MULT_mult_6_ab_11__2_), .ZN(MULT_mult_6_net81617) );
  NAND2_X4 MULT_mult_6_U2298 ( .A1(MULT_mult_6_n210), .A2(
        MULT_mult_6_ab_14__9_), .ZN(MULT_mult_6_n1939) );
  INV_X4 MULT_mult_6_U2297 ( .A(MULT_mult_6_CARRYB_15__12_), .ZN(
        MULT_mult_6_net87004) );
  INV_X4 MULT_mult_6_U2296 ( .A(MULT_mult_6_n1356), .ZN(MULT_mult_6_n1262) );
  INV_X2 MULT_mult_6_U2295 ( .A(MULT_mult_6_n709), .ZN(MULT_mult_6_n710) );
  NAND2_X2 MULT_mult_6_U2294 ( .A1(MULT_mult_6_CARRYB_8__4_), .A2(
        MULT_mult_6_SUMB_8__5_), .ZN(MULT_mult_6_net82101) );
  NAND3_X4 MULT_mult_6_U2293 ( .A1(MULT_mult_6_net81615), .A2(
        MULT_mult_6_net81616), .A3(MULT_mult_6_net81617), .ZN(
        MULT_mult_6_CARRYB_11__2_) );
  BUF_X4 MULT_mult_6_U2292 ( .A(MULT_mult_6_SUMB_7__10_), .Z(MULT_mult_6_n1325) );
  INV_X4 MULT_mult_6_U2291 ( .A(MULT_mult_6_SUMB_5__17_), .ZN(
        MULT_mult_6_n1528) );
  NAND2_X4 MULT_mult_6_U2290 ( .A1(MULT_mult_6_ab_6__18_), .A2(
        MULT_mult_6_SUMB_5__19_), .ZN(MULT_mult_6_n1681) );
  NAND2_X4 MULT_mult_6_U2289 ( .A1(MULT_mult_6_n1601), .A2(MULT_mult_6_n1602), 
        .ZN(MULT_mult_6_n2303) );
  NAND3_X1 MULT_mult_6_U2288 ( .A1(MULT_mult_6_n1714), .A2(MULT_mult_6_n1715), 
        .A3(MULT_mult_6_n1716), .ZN(MULT_mult_6_n861) );
  NAND2_X2 MULT_mult_6_U2287 ( .A1(MULT_mult_6_n1419), .A2(
        MULT_mult_6_SUMB_3__20_), .ZN(MULT_mult_6_n1422) );
  INV_X4 MULT_mult_6_U2286 ( .A(MULT_mult_6_n708), .ZN(MULT_mult_6_n1205) );
  XNOR2_X2 MULT_mult_6_U2285 ( .A(MULT_mult_6_ab_5__18_), .B(
        MULT_mult_6_CARRYB_4__18_), .ZN(MULT_mult_6_n708) );
  NAND2_X1 MULT_mult_6_U2284 ( .A1(MULT_mult_6_CARRYB_16__12_), .A2(
        MULT_mult_6_SUMB_16__13_), .ZN(MULT_mult_6_n892) );
  NAND2_X4 MULT_mult_6_U2283 ( .A1(MULT_mult_6_n1174), .A2(MULT_mult_6_n1175), 
        .ZN(MULT_mult_6_n1618) );
  INV_X1 MULT_mult_6_U2282 ( .A(MULT_mult_6_SUMB_9__9_), .ZN(MULT_mult_6_n705)
         );
  INV_X4 MULT_mult_6_U2281 ( .A(MULT_mult_6_n1773), .ZN(MULT_mult_6_n704) );
  NAND2_X2 MULT_mult_6_U2280 ( .A1(MULT_mult_6_n706), .A2(MULT_mult_6_n707), 
        .ZN(MULT_mult_6_SUMB_10__8_) );
  NAND2_X1 MULT_mult_6_U2279 ( .A1(MULT_mult_6_n1773), .A2(MULT_mult_6_n705), 
        .ZN(MULT_mult_6_n706) );
  NAND3_X4 MULT_mult_6_U2278 ( .A1(MULT_mult_6_n1639), .A2(MULT_mult_6_n1641), 
        .A3(MULT_mult_6_n1640), .ZN(MULT_mult_6_CARRYB_13__4_) );
  NAND2_X1 MULT_mult_6_U2277 ( .A1(MULT_mult_6_SUMB_12__14_), .A2(
        MULT_mult_6_ab_13__13_), .ZN(MULT_mult_6_n1574) );
  NAND2_X2 MULT_mult_6_U2276 ( .A1(MULT_mult_6_n1727), .A2(MULT_mult_6_n1728), 
        .ZN(MULT_mult_6_SUMB_16__11_) );
  INV_X2 MULT_mult_6_U2275 ( .A(MULT_mult_6_n1067), .ZN(MULT_mult_6_n701) );
  NAND2_X4 MULT_mult_6_U2274 ( .A1(MULT_mult_6_n702), .A2(MULT_mult_6_n703), 
        .ZN(MULT_mult_6_SUMB_12__14_) );
  NAND2_X1 MULT_mult_6_U2273 ( .A1(MULT_mult_6_n1067), .A2(
        MULT_mult_6_SUMB_11__15_), .ZN(MULT_mult_6_n702) );
  INV_X4 MULT_mult_6_U2272 ( .A(MULT_mult_6_n2282), .ZN(MULT_mult_6_n696) );
  NAND2_X4 MULT_mult_6_U2271 ( .A1(MULT_mult_6_n698), .A2(MULT_mult_6_n699), 
        .ZN(MULT_mult_6_n1780) );
  NAND2_X4 MULT_mult_6_U2270 ( .A1(MULT_mult_6_n696), .A2(MULT_mult_6_n697), 
        .ZN(MULT_mult_6_n699) );
  NAND2_X2 MULT_mult_6_U2269 ( .A1(MULT_mult_6_n2282), .A2(
        MULT_mult_6_SUMB_22__7_), .ZN(MULT_mult_6_n698) );
  INV_X4 MULT_mult_6_U2268 ( .A(MULT_mult_6_net81113), .ZN(MULT_mult_6_n692)
         );
  INV_X4 MULT_mult_6_U2267 ( .A(MULT_mult_6_SUMB_20__9_), .ZN(MULT_mult_6_n691) );
  NAND2_X4 MULT_mult_6_U2266 ( .A1(MULT_mult_6_n693), .A2(MULT_mult_6_n694), 
        .ZN(MULT_mult_6_SUMB_21__8_) );
  NAND2_X4 MULT_mult_6_U2265 ( .A1(MULT_mult_6_n691), .A2(MULT_mult_6_n692), 
        .ZN(MULT_mult_6_n694) );
  NAND2_X2 MULT_mult_6_U2264 ( .A1(MULT_mult_6_net81113), .A2(
        MULT_mult_6_SUMB_20__9_), .ZN(MULT_mult_6_n693) );
  INV_X4 MULT_mult_6_U2263 ( .A(MULT_mult_6_net92323), .ZN(MULT_mult_6_n688)
         );
  INV_X4 MULT_mult_6_U2262 ( .A(MULT_mult_6_net92322), .ZN(MULT_mult_6_n687)
         );
  NAND2_X4 MULT_mult_6_U2261 ( .A1(MULT_mult_6_n689), .A2(MULT_mult_6_n690), 
        .ZN(MULT_mult_6_net92321) );
  NAND2_X4 MULT_mult_6_U2260 ( .A1(MULT_mult_6_n687), .A2(MULT_mult_6_n688), 
        .ZN(MULT_mult_6_n690) );
  NAND2_X2 MULT_mult_6_U2259 ( .A1(MULT_mult_6_net92322), .A2(
        MULT_mult_6_net92323), .ZN(MULT_mult_6_n689) );
  NAND2_X4 MULT_mult_6_U2258 ( .A1(MULT_mult_6_n685), .A2(MULT_mult_6_n686), 
        .ZN(MULT_mult_6_SUMB_22__7_) );
  NAND2_X4 MULT_mult_6_U2257 ( .A1(MULT_mult_6_n1728), .A2(MULT_mult_6_n1727), 
        .ZN(MULT_mult_6_n682) );
  NAND2_X2 MULT_mult_6_U2256 ( .A1(MULT_mult_6_ab_10__8_), .A2(
        MULT_mult_6_CARRYB_9__8_), .ZN(MULT_mult_6_n1774) );
  INV_X8 MULT_mult_6_U2255 ( .A(MULT_mult_6_net86844), .ZN(
        MULT_mult_6_net120468) );
  NAND2_X4 MULT_mult_6_U2253 ( .A1(MULT_mult_6_n2364), .A2(
        MULT_mult_6_net147938), .ZN(MULT_mult_6_net147940) );
  NAND3_X2 MULT_mult_6_U2251 ( .A1(MULT_mult_6_n1776), .A2(MULT_mult_6_n1775), 
        .A3(MULT_mult_6_n1774), .ZN(MULT_mult_6_net147936) );
  INV_X4 MULT_mult_6_U2250 ( .A(MULT_mult_6_n1120), .ZN(MULT_mult_6_n679) );
  NAND2_X4 MULT_mult_6_U2249 ( .A1(MULT_mult_6_n681), .A2(MULT_mult_6_n680), 
        .ZN(MULT_mult_6_SUMB_3__12_) );
  NAND2_X2 MULT_mult_6_U2248 ( .A1(MULT_mult_6_n1928), .A2(MULT_mult_6_n1120), 
        .ZN(MULT_mult_6_n680) );
  NAND2_X2 MULT_mult_6_U2247 ( .A1(MULT_mult_6_n677), .A2(
        MULT_mult_6_net147922), .ZN(MULT_mult_6_net82757) );
  NAND2_X2 MULT_mult_6_U2246 ( .A1(MULT_mult_6_CARRYB_11__5_), .A2(
        MULT_mult_6_ab_12__5_), .ZN(MULT_mult_6_n1636) );
  INV_X1 MULT_mult_6_U2245 ( .A(MULT_mult_6_net83796), .ZN(
        MULT_mult_6_net84891) );
  INV_X1 MULT_mult_6_U2244 ( .A(MULT_mult_6_SUMB_6__13_), .ZN(
        MULT_mult_6_net88166) );
  XNOR2_X2 MULT_mult_6_U2243 ( .A(MULT_mult_6_n1222), .B(MULT_mult_6_ab_15__3_), .ZN(MULT_mult_6_n1010) );
  XNOR2_X2 MULT_mult_6_U2242 ( .A(MULT_mult_6_CARRYB_8__7_), .B(
        MULT_mult_6_ab_9__7_), .ZN(MULT_mult_6_n1176) );
  CLKBUF_X3 MULT_mult_6_U2241 ( .A(MULT_mult_6_n1261), .Z(MULT_mult_6_n946) );
  INV_X1 MULT_mult_6_U2240 ( .A(MULT_mult_6_n1750), .ZN(MULT_mult_6_n676) );
  NAND2_X2 MULT_mult_6_U2239 ( .A1(MULT_mult_6_SUMB_11__4_), .A2(
        MULT_mult_6_CARRYB_11__3_), .ZN(MULT_mult_6_n1675) );
  XNOR2_X2 MULT_mult_6_U2238 ( .A(MULT_mult_6_CARRYB_15__3_), .B(
        MULT_mult_6_ab_16__3_), .ZN(MULT_mult_6_n862) );
  NAND2_X2 MULT_mult_6_U2237 ( .A1(MULT_mult_6_SUMB_2__6_), .A2(
        MULT_mult_6_CARRYB_2__5_), .ZN(MULT_mult_6_n732) );
  NAND2_X4 MULT_mult_6_U2236 ( .A1(MULT_mult_6_CARRYB_19__0_), .A2(
        MULT_mult_6_SUMB_19__1_), .ZN(MULT_mult_6_n2102) );
  NAND2_X4 MULT_mult_6_U2235 ( .A1(MULT_mult_6_ab_17__1_), .A2(
        MULT_mult_6_CARRYB_16__1_), .ZN(MULT_mult_6_n743) );
  NAND2_X2 MULT_mult_6_U2234 ( .A1(MULT_mult_6_CARRYB_14__0_), .A2(
        MULT_mult_6_SUMB_14__1_), .ZN(MULT_mult_6_n1409) );
  NOR2_X4 MULT_mult_6_U2233 ( .A1(MULT_mult_6_net77906), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__6_) );
  NOR2_X4 MULT_mult_6_U2232 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__4_) );
  INV_X4 MULT_mult_6_U2231 ( .A(MULT_mult_6_ab_9__6_), .ZN(MULT_mult_6_n672)
         );
  INV_X4 MULT_mult_6_U2230 ( .A(MULT_mult_6_CARRYB_8__6_), .ZN(
        MULT_mult_6_n671) );
  NAND2_X1 MULT_mult_6_U2229 ( .A1(MULT_mult_6_CARRYB_8__6_), .A2(
        MULT_mult_6_ab_9__6_), .ZN(MULT_mult_6_n673) );
  INV_X4 MULT_mult_6_U2228 ( .A(MULT_mult_6_net86385), .ZN(
        MULT_mult_6_net147999) );
  INV_X4 MULT_mult_6_U2227 ( .A(MULT_mult_6_net81431), .ZN(
        MULT_mult_6_net147998) );
  NAND2_X4 MULT_mult_6_U2226 ( .A1(MULT_mult_6_n669), .A2(MULT_mult_6_n670), 
        .ZN(multOut[2]) );
  NAND2_X4 MULT_mult_6_U2225 ( .A1(MULT_mult_6_net147998), .A2(
        MULT_mult_6_net147999), .ZN(MULT_mult_6_n670) );
  NAND2_X2 MULT_mult_6_U2224 ( .A1(MULT_mult_6_net81431), .A2(
        MULT_mult_6_net86385), .ZN(MULT_mult_6_n669) );
  INV_X1 MULT_mult_6_U2223 ( .A(MULT_mult_6_ab_12__4_), .ZN(MULT_mult_6_n666)
         );
  INV_X4 MULT_mult_6_U2222 ( .A(MULT_mult_6_CARRYB_11__4_), .ZN(
        MULT_mult_6_n665) );
  NAND2_X4 MULT_mult_6_U2221 ( .A1(MULT_mult_6_n667), .A2(MULT_mult_6_n668), 
        .ZN(MULT_mult_6_n1243) );
  NAND2_X4 MULT_mult_6_U2220 ( .A1(MULT_mult_6_n665), .A2(MULT_mult_6_n666), 
        .ZN(MULT_mult_6_n668) );
  CLKBUF_X2 MULT_mult_6_U2219 ( .A(MULT_mult_6_CARRYB_22__4_), .Z(
        MULT_mult_6_net84213) );
  NAND2_X2 MULT_mult_6_U2218 ( .A1(MULT_mult_6_CARRYB_7__7_), .A2(
        MULT_mult_6_SUMB_7__8_), .ZN(MULT_mult_6_n1861) );
  NAND2_X4 MULT_mult_6_U2217 ( .A1(MULT_mult_6_net88887), .A2(
        MULT_mult_6_ab_20__4_), .ZN(MULT_mult_6_n2229) );
  INV_X4 MULT_mult_6_U2216 ( .A(MULT_mult_6_net83202), .ZN(
        MULT_mult_6_net147928) );
  INV_X8 MULT_mult_6_U2215 ( .A(MULT_mult_6_CARRYB_9__14_), .ZN(
        MULT_mult_6_n1038) );
  INV_X8 MULT_mult_6_U2214 ( .A(MULT_mult_6_CARRYB_11__13_), .ZN(
        MULT_mult_6_n1041) );
  INV_X1 MULT_mult_6_U2213 ( .A(MULT_mult_6_ab_9__13_), .ZN(
        MULT_mult_6_net83438) );
  INV_X2 MULT_mult_6_U2212 ( .A(MULT_mult_6_ab_4__16_), .ZN(MULT_mult_6_n803)
         );
  INV_X4 MULT_mult_6_U2211 ( .A(MULT_mult_6_net83438), .ZN(MULT_mult_6_n662)
         );
  INV_X4 MULT_mult_6_U2210 ( .A(MULT_mult_6_net84447), .ZN(MULT_mult_6_n661)
         );
  NAND2_X4 MULT_mult_6_U2209 ( .A1(MULT_mult_6_n663), .A2(MULT_mult_6_n664), 
        .ZN(MULT_mult_6_net80346) );
  NAND2_X4 MULT_mult_6_U2208 ( .A1(MULT_mult_6_n661), .A2(MULT_mult_6_n662), 
        .ZN(MULT_mult_6_n664) );
  NAND2_X2 MULT_mult_6_U2207 ( .A1(MULT_mult_6_CARRYB_8__13_), .A2(
        MULT_mult_6_net83438), .ZN(MULT_mult_6_n663) );
  INV_X4 MULT_mult_6_U2206 ( .A(MULT_mult_6_net80833), .ZN(
        MULT_mult_6_net148051) );
  NAND2_X2 MULT_mult_6_U2205 ( .A1(MULT_mult_6_net80833), .A2(
        MULT_mult_6_SUMB_3__17_), .ZN(MULT_mult_6_net148053) );
  INV_X1 MULT_mult_6_U2204 ( .A(MULT_mult_6_ab_16__9_), .ZN(MULT_mult_6_n659)
         );
  NAND2_X4 MULT_mult_6_U2203 ( .A1(MULT_mult_6_n658), .A2(MULT_mult_6_n659), 
        .ZN(MULT_mult_6_n660) );
  INV_X4 MULT_mult_6_U2202 ( .A(MULT_mult_6_n803), .ZN(MULT_mult_6_n655) );
  NAND2_X4 MULT_mult_6_U2201 ( .A1(MULT_mult_6_n656), .A2(MULT_mult_6_n657), 
        .ZN(MULT_mult_6_net80833) );
  NAND2_X4 MULT_mult_6_U2200 ( .A1(MULT_mult_6_n654), .A2(MULT_mult_6_n655), 
        .ZN(MULT_mult_6_n657) );
  NAND2_X1 MULT_mult_6_U2199 ( .A1(MULT_mult_6_ab_4__18_), .A2(
        MULT_mult_6_SUMB_3__19_), .ZN(MULT_mult_6_n1724) );
  INV_X8 MULT_mult_6_U2198 ( .A(MULT_mult_6_net89876), .ZN(
        MULT_mult_6_SUMB_20__4_) );
  NAND3_X4 MULT_mult_6_U2197 ( .A1(MULT_mult_6_n766), .A2(MULT_mult_6_net86134), .A3(MULT_mult_6_net86135), .ZN(MULT_mult_6_CARRYB_14__1_) );
  NOR2_X2 MULT_mult_6_U2196 ( .A1(MULT_mult_6_net77868), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__1_) );
  NAND2_X2 MULT_mult_6_U2195 ( .A1(MULT_mult_6_CARRYB_14__1_), .A2(
        MULT_mult_6_SUMB_14__2_), .ZN(MULT_mult_6_n651) );
  NAND3_X4 MULT_mult_6_U2192 ( .A1(MULT_mult_6_n647), .A2(MULT_mult_6_n648), 
        .A3(MULT_mult_6_n649), .ZN(MULT_mult_6_CARRYB_16__1_) );
  NAND2_X2 MULT_mult_6_U2191 ( .A1(MULT_mult_6_ab_16__1_), .A2(
        MULT_mult_6_SUMB_15__2_), .ZN(MULT_mult_6_n649) );
  NAND2_X2 MULT_mult_6_U2190 ( .A1(MULT_mult_6_SUMB_15__2_), .A2(
        MULT_mult_6_CARRYB_15__1_), .ZN(MULT_mult_6_n647) );
  XOR2_X2 MULT_mult_6_U2189 ( .A(MULT_mult_6_CARRYB_15__1_), .B(
        MULT_mult_6_n646), .Z(MULT_mult_6_SUMB_16__1_) );
  NAND2_X4 MULT_mult_6_U2188 ( .A1(MULT_mult_6_SUMB_3__11_), .A2(
        MULT_mult_6_ab_4__10_), .ZN(MULT_mult_6_n1395) );
  NAND2_X2 MULT_mult_6_U2187 ( .A1(MULT_mult_6_net83445), .A2(
        MULT_mult_6_SUMB_13__14_), .ZN(MULT_mult_6_net86630) );
  NAND2_X4 MULT_mult_6_U2186 ( .A1(MULT_mult_6_n1205), .A2(MULT_mult_6_n1576), 
        .ZN(MULT_mult_6_n1578) );
  INV_X8 MULT_mult_6_U2185 ( .A(MULT_mult_6_CARRYB_18__5_), .ZN(
        MULT_mult_6_net84707) );
  NAND2_X2 MULT_mult_6_U2184 ( .A1(MULT_mult_6_net124434), .A2(
        MULT_mult_6_SUMB_11__13_), .ZN(MULT_mult_6_net86158) );
  NAND2_X2 MULT_mult_6_U2183 ( .A1(MULT_mult_6_SUMB_11__13_), .A2(
        MULT_mult_6_ab_12__12_), .ZN(MULT_mult_6_net86159) );
  AND3_X2 MULT_mult_6_U2182 ( .A1(MULT_mult_6_net86158), .A2(
        MULT_mult_6_net86159), .A3(MULT_mult_6_n1019), .ZN(MULT_mult_6_n645)
         );
  INV_X4 MULT_mult_6_U2181 ( .A(MULT_mult_6_net93683), .ZN(MULT_mult_6_n642)
         );
  INV_X1 MULT_mult_6_U2180 ( .A(MULT_mult_6_ab_5__16_), .ZN(MULT_mult_6_n637)
         );
  NAND2_X2 MULT_mult_6_U2179 ( .A1(MULT_mult_6_ab_5__16_), .A2(
        MULT_mult_6_CARRYB_4__16_), .ZN(MULT_mult_6_n639) );
  NAND2_X4 MULT_mult_6_U2178 ( .A1(MULT_mult_6_n678), .A2(
        MULT_mult_6_net147930), .ZN(MULT_mult_6_SUMB_20__5_) );
  NAND2_X4 MULT_mult_6_U2177 ( .A1(MULT_mult_6_net120653), .A2(
        MULT_mult_6_n1011), .ZN(MULT_mult_6_SUMB_10__12_) );
  NAND2_X2 MULT_mult_6_U2176 ( .A1(MULT_mult_6_ab_14__9_), .A2(
        MULT_mult_6_net85043), .ZN(MULT_mult_6_n1938) );
  NAND2_X4 MULT_mult_6_U2175 ( .A1(MULT_mult_6_n830), .A2(MULT_mult_6_n831), 
        .ZN(MULT_mult_6_net84818) );
  INV_X4 MULT_mult_6_U2174 ( .A(MULT_mult_6_n1628), .ZN(MULT_mult_6_n1191) );
  NAND2_X4 MULT_mult_6_U2173 ( .A1(MULT_mult_6_n638), .A2(MULT_mult_6_n637), 
        .ZN(MULT_mult_6_n640) );
  INV_X4 MULT_mult_6_U2172 ( .A(MULT_mult_6_n1504), .ZN(MULT_mult_6_n885) );
  INV_X4 MULT_mult_6_U2171 ( .A(MULT_mult_6_SUMB_2__8_), .ZN(
        MULT_mult_6_net85035) );
  NAND2_X2 MULT_mult_6_U2170 ( .A1(MULT_mult_6_CARRYB_13__4_), .A2(
        MULT_mult_6_ab_14__4_), .ZN(MULT_mult_6_n1633) );
  NAND2_X4 MULT_mult_6_U2169 ( .A1(MULT_mult_6_n1341), .A2(
        MULT_mult_6_net88638), .ZN(MULT_mult_6_n1336) );
  NAND2_X4 MULT_mult_6_U2168 ( .A1(MULT_mult_6_SUMB_18__3_), .A2(
        MULT_mult_6_ab_19__2_), .ZN(MULT_mult_6_n1912) );
  INV_X8 MULT_mult_6_U2167 ( .A(MULT_mult_6_CARRYB_18__4_), .ZN(
        MULT_mult_6_n1858) );
  NAND2_X4 MULT_mult_6_U2166 ( .A1(MULT_mult_6_CARRYB_3__10_), .A2(
        MULT_mult_6_ab_4__10_), .ZN(MULT_mult_6_n1393) );
  XNOR2_X2 MULT_mult_6_U2165 ( .A(MULT_mult_6_n2111), .B(
        MULT_mult_6_SUMB_2__19_), .ZN(MULT_mult_6_n852) );
  NAND2_X2 MULT_mult_6_U2164 ( .A1(MULT_mult_6_ab_9__7_), .A2(
        MULT_mult_6_CARRYB_8__7_), .ZN(MULT_mult_6_n2018) );
  NAND2_X2 MULT_mult_6_U2163 ( .A1(MULT_mult_6_SUMB_18__5_), .A2(
        MULT_mult_6_n2109), .ZN(MULT_mult_6_n1348) );
  BUF_X4 MULT_mult_6_U2162 ( .A(MULT_mult_6_SUMB_15__7_), .Z(
        MULT_mult_6_net84657) );
  BUF_X4 MULT_mult_6_U2161 ( .A(MULT_mult_6_SUMB_13__8_), .Z(MULT_mult_6_n1284) );
  NAND2_X4 MULT_mult_6_U2158 ( .A1(MULT_mult_6_n635), .A2(MULT_mult_6_n636), 
        .ZN(MULT_mult_6_SUMB_18__5_) );
  NAND2_X2 MULT_mult_6_U2157 ( .A1(MULT_mult_6_n634), .A2(
        MULT_mult_6_net148235), .ZN(MULT_mult_6_n636) );
  NAND2_X1 MULT_mult_6_U2156 ( .A1(MULT_mult_6_n1718), .A2(
        MULT_mult_6_net86662), .ZN(MULT_mult_6_n635) );
  INV_X4 MULT_mult_6_U2155 ( .A(MULT_mult_6_net84657), .ZN(
        MULT_mult_6_net148230) );
  INV_X4 MULT_mult_6_U2154 ( .A(MULT_mult_6_n1856), .ZN(MULT_mult_6_n631) );
  NAND2_X4 MULT_mult_6_U2153 ( .A1(MULT_mult_6_n632), .A2(MULT_mult_6_n633), 
        .ZN(MULT_mult_6_SUMB_16__6_) );
  NAND2_X4 MULT_mult_6_U2152 ( .A1(MULT_mult_6_n631), .A2(
        MULT_mult_6_net148230), .ZN(MULT_mult_6_n633) );
  NAND2_X2 MULT_mult_6_U2151 ( .A1(MULT_mult_6_n1856), .A2(
        MULT_mult_6_net84657), .ZN(MULT_mult_6_n632) );
  INV_X8 MULT_mult_6_U2150 ( .A(MULT_mult_6_n1284), .ZN(MULT_mult_6_n627) );
  NAND2_X4 MULT_mult_6_U2149 ( .A1(MULT_mult_6_n630), .A2(MULT_mult_6_n629), 
        .ZN(MULT_mult_6_SUMB_14__7_) );
  NAND2_X4 MULT_mult_6_U2148 ( .A1(MULT_mult_6_n627), .A2(MULT_mult_6_n628), 
        .ZN(MULT_mult_6_n630) );
  NAND2_X2 MULT_mult_6_U2147 ( .A1(MULT_mult_6_n1284), .A2(MULT_mult_6_n1553), 
        .ZN(MULT_mult_6_n629) );
  XNOR2_X2 MULT_mult_6_U2146 ( .A(MULT_mult_6_ab_14__3_), .B(
        MULT_mult_6_CARRYB_13__3_), .ZN(MULT_mult_6_n942) );
  NAND2_X2 MULT_mult_6_U2145 ( .A1(MULT_mult_6_n888), .A2(MULT_mult_6_n889), 
        .ZN(MULT_mult_6_n890) );
  INV_X4 MULT_mult_6_U2144 ( .A(MULT_mult_6_n1218), .ZN(MULT_mult_6_n1219) );
  INV_X2 MULT_mult_6_U2143 ( .A(MULT_mult_6_net90702), .ZN(
        MULT_mult_6_net86601) );
  NAND2_X4 MULT_mult_6_U2142 ( .A1(MULT_mult_6_SUMB_20__5_), .A2(
        MULT_mult_6_ab_21__4_), .ZN(MULT_mult_6_net82407) );
  NAND2_X2 MULT_mult_6_U2141 ( .A1(MULT_mult_6_CARRYB_15__12_), .A2(
        MULT_mult_6_SUMB_15__13_), .ZN(MULT_mult_6_n1087) );
  NAND2_X2 MULT_mult_6_U2140 ( .A1(MULT_mult_6_n704), .A2(
        MULT_mult_6_SUMB_9__9_), .ZN(MULT_mult_6_n707) );
  NAND2_X2 MULT_mult_6_U2139 ( .A1(MULT_mult_6_CARRYB_10__0_), .A2(
        MULT_mult_6_ab_11__0_), .ZN(MULT_mult_6_n1140) );
  XOR2_X1 MULT_mult_6_U2138 ( .A(MULT_mult_6_CARRYB_10__0_), .B(
        MULT_mult_6_ab_11__0_), .Z(MULT_mult_6_n1139) );
  NAND2_X4 MULT_mult_6_U2137 ( .A1(MULT_mult_6_n625), .A2(MULT_mult_6_n626), 
        .ZN(MULT_mult_6_net87411) );
  NAND2_X2 MULT_mult_6_U2136 ( .A1(MULT_mult_6_net92405), .A2(
        MULT_mult_6_net148015), .ZN(MULT_mult_6_n625) );
  INV_X4 MULT_mult_6_U2135 ( .A(MULT_mult_6_net88700), .ZN(MULT_mult_6_n622)
         );
  NAND2_X4 MULT_mult_6_U2134 ( .A1(MULT_mult_6_n623), .A2(MULT_mult_6_n624), 
        .ZN(MULT_mult_6_net90818) );
  NAND2_X4 MULT_mult_6_U2133 ( .A1(MULT_mult_6_n1349), .A2(MULT_mult_6_n1348), 
        .ZN(MULT_mult_6_SUMB_19__4_) );
  NAND2_X2 MULT_mult_6_U2132 ( .A1(MULT_mult_6_ab_4__22_), .A2(
        MULT_mult_6_n843), .ZN(MULT_mult_6_net84313) );
  NOR2_X1 MULT_mult_6_U2131 ( .A1(MULT_mult_6_net70478), .A2(
        MULT_mult_6_net77964), .ZN(MULT_mult_6_ab_3__22_) );
  NAND2_X1 MULT_mult_6_U2130 ( .A1(MULT_mult_6_ab_7__21_), .A2(
        MULT_mult_6_SUMB_6__22_), .ZN(MULT_mult_6_n987) );
  NAND2_X2 MULT_mult_6_U2129 ( .A1(MULT_mult_6_n1766), .A2(
        MULT_mult_6_net90702), .ZN(MULT_mult_6_n1604) );
  NAND2_X2 MULT_mult_6_U2128 ( .A1(MULT_mult_6_ab_7__8_), .A2(
        MULT_mult_6_n1425), .ZN(MULT_mult_6_n2059) );
  NAND3_X2 MULT_mult_6_U2127 ( .A1(MULT_mult_6_n2057), .A2(MULT_mult_6_n2058), 
        .A3(MULT_mult_6_n2059), .ZN(MULT_mult_6_CARRYB_7__8_) );
  NAND3_X4 MULT_mult_6_U2126 ( .A1(MULT_mult_6_n2057), .A2(MULT_mult_6_n2058), 
        .A3(MULT_mult_6_n2059), .ZN(MULT_mult_6_n621) );
  NAND2_X2 MULT_mult_6_U2125 ( .A1(MULT_mult_6_ab_5__22_), .A2(
        MULT_mult_6_SUMB_4__23_), .ZN(MULT_mult_6_net80795) );
  XNOR2_X2 MULT_mult_6_U2124 ( .A(MULT_mult_6_CARRYB_18__12_), .B(
        MULT_mult_6_ab_19__12_), .ZN(MULT_mult_6_n620) );
  XNOR2_X2 MULT_mult_6_U2123 ( .A(MULT_mult_6_SUMB_17__14_), .B(
        MULT_mult_6_n951), .ZN(MULT_mult_6_n619) );
  XNOR2_X2 MULT_mult_6_U2122 ( .A(MULT_mult_6_n619), .B(MULT_mult_6_n620), 
        .ZN(MULT_mult_6_n1413) );
  NAND2_X4 MULT_mult_6_U2121 ( .A1(MULT_mult_6_n1393), .A2(MULT_mult_6_n890), 
        .ZN(MULT_mult_6_n1339) );
  INV_X4 MULT_mult_6_U2120 ( .A(MULT_mult_6_CARRYB_8__15_), .ZN(
        MULT_mult_6_n1366) );
  NAND2_X2 MULT_mult_6_U2119 ( .A1(MULT_mult_6_CARRYB_8__15_), .A2(
        MULT_mult_6_ab_9__15_), .ZN(MULT_mult_6_n1709) );
  NAND2_X4 MULT_mult_6_U2118 ( .A1(MULT_mult_6_SUMB_7__9_), .A2(
        MULT_mult_6_ab_8__8_), .ZN(MULT_mult_6_n2005) );
  INV_X8 MULT_mult_6_U2117 ( .A(MULT_mult_6_CARRYB_4__16_), .ZN(
        MULT_mult_6_n638) );
  NAND3_X4 MULT_mult_6_U2116 ( .A1(MULT_mult_6_n1071), .A2(
        MULT_mult_6_net80267), .A3(MULT_mult_6_net80268), .ZN(
        MULT_mult_6_CARRYB_22__7_) );
  NAND3_X4 MULT_mult_6_U2115 ( .A1(MULT_mult_6_n1870), .A2(MULT_mult_6_n1871), 
        .A3(MULT_mult_6_n1872), .ZN(MULT_mult_6_CARRYB_14__15_) );
  INV_X2 MULT_mult_6_U2114 ( .A(MULT_mult_6_n2188), .ZN(MULT_mult_6_n616) );
  INV_X2 MULT_mult_6_U2113 ( .A(MULT_mult_6_SUMB_13__17_), .ZN(
        MULT_mult_6_n615) );
  NAND2_X4 MULT_mult_6_U2112 ( .A1(MULT_mult_6_n617), .A2(MULT_mult_6_n618), 
        .ZN(MULT_mult_6_n1252) );
  NAND2_X2 MULT_mult_6_U2111 ( .A1(MULT_mult_6_SUMB_13__17_), .A2(
        MULT_mult_6_n2188), .ZN(MULT_mult_6_n617) );
  NAND3_X2 MULT_mult_6_U2110 ( .A1(MULT_mult_6_n612), .A2(MULT_mult_6_n613), 
        .A3(MULT_mult_6_n614), .ZN(MULT_mult_6_CARRYB_15__15_) );
  NAND2_X1 MULT_mult_6_U2109 ( .A1(MULT_mult_6_ab_15__15_), .A2(
        MULT_mult_6_CARRYB_14__15_), .ZN(MULT_mult_6_n614) );
  NAND2_X1 MULT_mult_6_U2108 ( .A1(MULT_mult_6_ab_15__15_), .A2(
        MULT_mult_6_n1252), .ZN(MULT_mult_6_n613) );
  NAND2_X1 MULT_mult_6_U2107 ( .A1(MULT_mult_6_CARRYB_14__15_), .A2(
        MULT_mult_6_n1252), .ZN(MULT_mult_6_n612) );
  XOR2_X2 MULT_mult_6_U2106 ( .A(MULT_mult_6_n1252), .B(MULT_mult_6_n611), .Z(
        MULT_mult_6_SUMB_15__15_) );
  XOR2_X2 MULT_mult_6_U2105 ( .A(MULT_mult_6_CARRYB_14__15_), .B(
        MULT_mult_6_ab_15__15_), .Z(MULT_mult_6_n611) );
  NAND3_X2 MULT_mult_6_U2104 ( .A1(MULT_mult_6_n2206), .A2(MULT_mult_6_n2207), 
        .A3(MULT_mult_6_n2205), .ZN(MULT_mult_6_CARRYB_6__16_) );
  NAND2_X2 MULT_mult_6_U2103 ( .A1(MULT_mult_6_ab_16__12_), .A2(
        MULT_mult_6_SUMB_15__13_), .ZN(MULT_mult_6_n1086) );
  INV_X4 MULT_mult_6_U2102 ( .A(MULT_mult_6_n2197), .ZN(MULT_mult_6_n1788) );
  NAND2_X4 MULT_mult_6_U2101 ( .A1(MULT_mult_6_net120655), .A2(
        MULT_mult_6_net120656), .ZN(MULT_mult_6_n804) );
  NAND2_X2 MULT_mult_6_U2100 ( .A1(MULT_mult_6_net93203), .A2(
        MULT_mult_6_n1901), .ZN(MULT_mult_6_n1128) );
  NAND2_X2 MULT_mult_6_U2099 ( .A1(MULT_mult_6_SUMB_18__9_), .A2(
        MULT_mult_6_net88700), .ZN(MULT_mult_6_n623) );
  NAND3_X2 MULT_mult_6_U2098 ( .A1(MULT_mult_6_n2236), .A2(MULT_mult_6_n2235), 
        .A3(MULT_mult_6_n2234), .ZN(MULT_mult_6_CARRYB_19__4_) );
  NAND2_X4 MULT_mult_6_U2097 ( .A1(MULT_mult_6_CARRYB_17__3_), .A2(
        MULT_mult_6_ab_18__3_), .ZN(MULT_mult_6_n1416) );
  XNOR2_X1 MULT_mult_6_U2096 ( .A(MULT_mult_6_n1268), .B(MULT_mult_6_n1241), 
        .ZN(MULT_mult_6_n868) );
  NAND3_X1 MULT_mult_6_U2095 ( .A1(MULT_mult_6_net86170), .A2(
        MULT_mult_6_net86171), .A3(MULT_mult_6_net86172), .ZN(
        MULT_mult_6_n1186) );
  NAND2_X2 MULT_mult_6_U2094 ( .A1(MULT_mult_6_n1589), .A2(MULT_mult_6_n1456), 
        .ZN(MULT_mult_6_n1591) );
  XOR2_X2 MULT_mult_6_U2092 ( .A(MULT_mult_6_n1470), .B(MULT_mult_6_net124757), 
        .Z(MULT_mult_6_SUMB_10__1_) );
  XNOR2_X2 MULT_mult_6_U2091 ( .A(MULT_mult_6_ab_3__6_), .B(
        MULT_mult_6_CARRYB_2__6_), .ZN(MULT_mult_6_n610) );
  XNOR2_X2 MULT_mult_6_U2090 ( .A(MULT_mult_6_n610), .B(MULT_mult_6_net87962), 
        .ZN(MULT_mult_6_SUMB_3__6_) );
  INV_X4 MULT_mult_6_U2089 ( .A(MULT_mult_6_SUMB_13__14_), .ZN(
        MULT_mult_6_net86629) );
  NAND2_X1 MULT_mult_6_U2088 ( .A1(MULT_mult_6_ab_25__5_), .A2(
        MULT_mult_6_SUMB_24__6_), .ZN(MULT_mult_6_net79867) );
  INV_X2 MULT_mult_6_U2087 ( .A(MULT_mult_6_net84707), .ZN(
        MULT_mult_6_net148582) );
  BUF_X8 MULT_mult_6_U2085 ( .A(MULT_mult_6_SUMB_13__6_), .Z(MULT_mult_6_n1202) );
  BUF_X8 MULT_mult_6_U2084 ( .A(MULT_mult_6_CARRYB_16__9_), .Z(
        MULT_mult_6_net89819) );
  NAND2_X2 MULT_mult_6_U2083 ( .A1(MULT_mult_6_CARRYB_18__8_), .A2(
        MULT_mult_6_ab_19__8_), .ZN(MULT_mult_6_net123293) );
  NAND2_X4 MULT_mult_6_U2082 ( .A1(MULT_mult_6_n609), .A2(MULT_mult_6_n608), 
        .ZN(multOut[0]) );
  NAND2_X4 MULT_mult_6_U2081 ( .A1(MULT_mult_6_n606), .A2(MULT_mult_6_n607), 
        .ZN(MULT_mult_6_n609) );
  INV_X1 MULT_mult_6_U2080 ( .A(MULT_mult_6_ab_8__14_), .ZN(MULT_mult_6_n603)
         );
  XNOR2_X2 MULT_mult_6_U2079 ( .A(MULT_mult_6_n350), .B(MULT_mult_6_ab_2__6_), 
        .ZN(MULT_mult_6_n758) );
  NAND3_X4 MULT_mult_6_U2078 ( .A1(MULT_mult_6_n1471), .A2(MULT_mult_6_n1472), 
        .A3(MULT_mult_6_n1473), .ZN(MULT_mult_6_CARRYB_10__1_) );
  NAND2_X2 MULT_mult_6_U2077 ( .A1(MULT_mult_6_CARRYB_10__0_), .A2(
        MULT_mult_6_SUMB_10__1_), .ZN(MULT_mult_6_n1142) );
  NAND2_X4 MULT_mult_6_U2076 ( .A1(MULT_mult_6_CARRYB_19__0_), .A2(
        MULT_mult_6_ab_20__0_), .ZN(MULT_mult_6_n2100) );
  BUF_X8 MULT_mult_6_U2075 ( .A(MULT_mult_6_SUMB_15__5_), .Z(MULT_mult_6_n1265) );
  INV_X4 MULT_mult_6_U2074 ( .A(MULT_mult_6_n1265), .ZN(MULT_mult_6_n599) );
  INV_X4 MULT_mult_6_U2073 ( .A(MULT_mult_6_n1731), .ZN(MULT_mult_6_n598) );
  NAND2_X4 MULT_mult_6_U2072 ( .A1(MULT_mult_6_n600), .A2(MULT_mult_6_n601), 
        .ZN(MULT_mult_6_SUMB_16__4_) );
  NAND2_X4 MULT_mult_6_U2071 ( .A1(MULT_mult_6_n598), .A2(MULT_mult_6_n599), 
        .ZN(MULT_mult_6_n601) );
  NAND2_X2 MULT_mult_6_U2070 ( .A1(MULT_mult_6_n1731), .A2(MULT_mult_6_n1265), 
        .ZN(MULT_mult_6_n600) );
  NAND3_X2 MULT_mult_6_U2069 ( .A1(MULT_mult_6_n1914), .A2(MULT_mult_6_n1916), 
        .A3(MULT_mult_6_n1915), .ZN(MULT_mult_6_n596) );
  XNOR2_X2 MULT_mult_6_U2068 ( .A(MULT_mult_6_SUMB_11__4_), .B(
        MULT_mult_6_ab_12__3_), .ZN(MULT_mult_6_n985) );
  BUF_X4 MULT_mult_6_U2067 ( .A(MULT_mult_6_SUMB_4__8_), .Z(MULT_mult_6_n1389)
         );
  INV_X4 MULT_mult_6_U2066 ( .A(MULT_mult_6_n947), .ZN(MULT_mult_6_n948) );
  INV_X4 MULT_mult_6_U2065 ( .A(MULT_mult_6_n1276), .ZN(MULT_mult_6_n593) );
  NAND2_X2 MULT_mult_6_U2064 ( .A1(MULT_mult_6_n592), .A2(MULT_mult_6_n593), 
        .ZN(MULT_mult_6_n595) );
  NAND2_X1 MULT_mult_6_U2063 ( .A1(MULT_mult_6_n563), .A2(MULT_mult_6_n1276), 
        .ZN(MULT_mult_6_n594) );
  INV_X4 MULT_mult_6_U2062 ( .A(MULT_mult_6_n1551), .ZN(MULT_mult_6_n589) );
  NAND2_X4 MULT_mult_6_U2061 ( .A1(MULT_mult_6_n590), .A2(MULT_mult_6_n591), 
        .ZN(MULT_mult_6_SUMB_4__8_) );
  NAND2_X4 MULT_mult_6_U2060 ( .A1(MULT_mult_6_n589), .A2(MULT_mult_6_n947), 
        .ZN(MULT_mult_6_n591) );
  NAND2_X2 MULT_mult_6_U2059 ( .A1(MULT_mult_6_n1551), .A2(MULT_mult_6_n948), 
        .ZN(MULT_mult_6_n590) );
  CLKBUF_X3 MULT_mult_6_U2058 ( .A(MULT_mult_6_SUMB_11__8_), .Z(
        MULT_mult_6_n1248) );
  INV_X4 MULT_mult_6_U2057 ( .A(MULT_mult_6_n2337), .ZN(
        MULT_mult_6_SUMB_1__12_) );
  INV_X4 MULT_mult_6_U2056 ( .A(MULT_mult_6_n1044), .ZN(MULT_mult_6_n588) );
  NAND2_X1 MULT_mult_6_U2055 ( .A1(MULT_mult_6_ab_15__12_), .A2(
        MULT_mult_6_CARRYB_14__12_), .ZN(MULT_mult_6_n2200) );
  INV_X2 MULT_mult_6_U2054 ( .A(MULT_mult_6_net148233), .ZN(
        MULT_mult_6_net148754) );
  OR2_X4 MULT_mult_6_U2053 ( .A1(MULT_mult_6_n830), .A2(MULT_mult_6_n831), 
        .ZN(MULT_mult_6_n827) );
  INV_X4 MULT_mult_6_U2052 ( .A(MULT_mult_6_n1118), .ZN(MULT_mult_6_n955) );
  NAND2_X4 MULT_mult_6_U2051 ( .A1(MULT_mult_6_net80021), .A2(
        MULT_mult_6_SUMB_23__5_), .ZN(MULT_mult_6_net86023) );
  INV_X8 MULT_mult_6_U2050 ( .A(MULT_mult_6_n2334), .ZN(
        MULT_mult_6_CARRYB_1__11_) );
  NAND2_X4 MULT_mult_6_U2049 ( .A1(MULT_mult_6_n585), .A2(MULT_mult_6_n586), 
        .ZN(MULT_mult_6_n587) );
  INV_X2 MULT_mult_6_U2048 ( .A(MULT_mult_6_net80927), .ZN(MULT_mult_6_n581)
         );
  NAND2_X1 MULT_mult_6_U2047 ( .A1(MULT_mult_6_net80927), .A2(
        MULT_mult_6_net89104), .ZN(MULT_mult_6_n583) );
  NAND2_X4 MULT_mult_6_U2046 ( .A1(MULT_mult_6_n579), .A2(MULT_mult_6_n580), 
        .ZN(MULT_mult_6_net86884) );
  NAND2_X4 MULT_mult_6_U2045 ( .A1(MULT_mult_6_n577), .A2(MULT_mult_6_n578), 
        .ZN(MULT_mult_6_n580) );
  NAND2_X2 MULT_mult_6_U2044 ( .A1(MULT_mult_6_net83030), .A2(
        MULT_mult_6_net81663), .ZN(MULT_mult_6_n579) );
  NAND2_X4 MULT_mult_6_U2043 ( .A1(MULT_mult_6_SUMB_7__8_), .A2(
        MULT_mult_6_ab_8__7_), .ZN(MULT_mult_6_n1862) );
  NAND2_X2 MULT_mult_6_U2042 ( .A1(MULT_mult_6_CARRYB_5__12_), .A2(
        MULT_mult_6_ab_6__12_), .ZN(MULT_mult_6_n1417) );
  NAND2_X4 MULT_mult_6_U2041 ( .A1(MULT_mult_6_SUMB_5__14_), .A2(
        MULT_mult_6_ab_6__13_), .ZN(MULT_mult_6_n2069) );
  INV_X8 MULT_mult_6_U2040 ( .A(MULT_mult_6_SUMB_18__9_), .ZN(MULT_mult_6_n641) );
  INV_X4 MULT_mult_6_U2039 ( .A(MULT_mult_6_n576), .ZN(MULT_mult_6_SUMB_18__9_) );
  XNOR2_X2 MULT_mult_6_U2038 ( .A(MULT_mult_6_net81782), .B(MULT_mult_6_n825), 
        .ZN(MULT_mult_6_n576) );
  NAND2_X4 MULT_mult_6_U2037 ( .A1(MULT_mult_6_ab_2__11_), .A2(
        MULT_mult_6_CARRYB_1__11_), .ZN(MULT_mult_6_n1642) );
  NAND2_X4 MULT_mult_6_U2036 ( .A1(MULT_mult_6_n1366), .A2(MULT_mult_6_n1708), 
        .ZN(MULT_mult_6_n1710) );
  INV_X2 MULT_mult_6_U2035 ( .A(MULT_mult_6_SUMB_11__15_), .ZN(
        MULT_mult_6_n700) );
  INV_X8 MULT_mult_6_U2034 ( .A(MULT_mult_6_net80392), .ZN(
        MULT_mult_6_net124610) );
  NOR2_X4 MULT_mult_6_U2033 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net77964), .ZN(MULT_mult_6_ab_3__12_) );
  XOR2_X2 MULT_mult_6_U2032 ( .A(MULT_mult_6_n1207), .B(MULT_mult_6_ab_3__12_), 
        .Z(MULT_mult_6_n575) );
  NAND2_X1 MULT_mult_6_U2031 ( .A1(MULT_mult_6_ab_9__8_), .A2(
        MULT_mult_6_CARRYB_8__8_), .ZN(MULT_mult_6_n2086) );
  NAND2_X2 MULT_mult_6_U2030 ( .A1(MULT_mult_6_n1154), .A2(
        MULT_mult_6_CARRYB_1__10_), .ZN(MULT_mult_6_n1156) );
  NAND2_X2 MULT_mult_6_U2029 ( .A1(MULT_mult_6_net92863), .A2(
        MULT_mult_6_net92862), .ZN(MULT_mult_6_n1617) );
  XNOR2_X2 MULT_mult_6_U2028 ( .A(MULT_mult_6_n574), .B(
        MULT_mult_6_SUMB_14__3_), .ZN(MULT_mult_6_SUMB_15__2_) );
  XOR2_X2 MULT_mult_6_U2027 ( .A(MULT_mult_6_SUMB_8__19_), .B(
        MULT_mult_6_net79950), .Z(MULT_mult_6_n573) );
  XNOR2_X2 MULT_mult_6_U2026 ( .A(MULT_mult_6_n1339), .B(MULT_mult_6_n1229), 
        .ZN(MULT_mult_6_n572) );
  BUF_X8 MULT_mult_6_U2025 ( .A(MULT_mult_6_SUMB_15__3_), .Z(MULT_mult_6_n571)
         );
  NAND2_X2 MULT_mult_6_U2024 ( .A1(MULT_mult_6_n1004), .A2(MULT_mult_6_n1683), 
        .ZN(MULT_mult_6_n1685) );
  NAND2_X4 MULT_mult_6_U2023 ( .A1(MULT_mult_6_SUMB_19__5_), .A2(
        MULT_mult_6_CARRYB_19__4_), .ZN(MULT_mult_6_n2230) );
  INV_X4 MULT_mult_6_U2022 ( .A(MULT_mult_6_n37), .ZN(MULT_mult_6_n1593) );
  INV_X4 MULT_mult_6_U2021 ( .A(MULT_mult_6_n1593), .ZN(MULT_mult_6_n570) );
  XNOR2_X2 MULT_mult_6_U2020 ( .A(MULT_mult_6_CARRYB_17__4_), .B(
        MULT_mult_6_ab_18__4_), .ZN(MULT_mult_6_n569) );
  XNOR2_X2 MULT_mult_6_U2019 ( .A(MULT_mult_6_n1204), .B(
        MULT_mult_6_SUMB_19__11_), .ZN(MULT_mult_6_n568) );
  NAND2_X2 MULT_mult_6_U2018 ( .A1(MULT_mult_6_ab_8__7_), .A2(
        MULT_mult_6_CARRYB_7__7_), .ZN(MULT_mult_6_n1863) );
  NAND3_X4 MULT_mult_6_U2017 ( .A1(MULT_mult_6_n1861), .A2(MULT_mult_6_n1862), 
        .A3(MULT_mult_6_n1863), .ZN(MULT_mult_6_CARRYB_8__7_) );
  OR2_X2 MULT_mult_6_U2016 ( .A1(MULT_mult_6_n1037), .A2(MULT_mult_6_n1038), 
        .ZN(MULT_mult_6_n1302) );
  NAND2_X2 MULT_mult_6_U2015 ( .A1(MULT_mult_6_n979), .A2(MULT_mult_6_n980), 
        .ZN(MULT_mult_6_net86557) );
  NOR2_X2 MULT_mult_6_U2014 ( .A1(MULT_mult_6_net70456), .A2(
        MULT_mult_6_net119855), .ZN(MULT_mult_6_ab_4__11_) );
  XNOR2_X2 MULT_mult_6_U2013 ( .A(MULT_mult_6_net81995), .B(MULT_mult_6_n833), 
        .ZN(MULT_mult_6_n565) );
  CLKBUF_X3 MULT_mult_6_U2012 ( .A(MULT_mult_6_SUMB_22__3_), .Z(
        MULT_mult_6_n564) );
  XOR2_X2 MULT_mult_6_U2011 ( .A(MULT_mult_6_n1315), .B(MULT_mult_6_n730), .Z(
        MULT_mult_6_SUMB_11__1_) );
  NAND2_X2 MULT_mult_6_U2010 ( .A1(MULT_mult_6_SUMB_11__1_), .A2(
        MULT_mult_6_CARRYB_11__0_), .ZN(MULT_mult_6_n1146) );
  NAND2_X2 MULT_mult_6_U2009 ( .A1(MULT_mult_6_ab_12__0_), .A2(
        MULT_mult_6_SUMB_11__1_), .ZN(MULT_mult_6_n1144) );
  INV_X4 MULT_mult_6_U2008 ( .A(MULT_mult_6_SUMB_10__5_), .ZN(MULT_mult_6_n592) );
  NAND2_X2 MULT_mult_6_U2007 ( .A1(MULT_mult_6_CARRYB_3__16_), .A2(
        MULT_mult_6_n803), .ZN(MULT_mult_6_n656) );
  INV_X1 MULT_mult_6_U2006 ( .A(MULT_mult_6_n1041), .ZN(MULT_mult_6_n562) );
  XNOR2_X2 MULT_mult_6_U2005 ( .A(MULT_mult_6_SUMB_7__7_), .B(MULT_mult_6_n561), .ZN(MULT_mult_6_SUMB_8__6_) );
  XNOR2_X2 MULT_mult_6_U2004 ( .A(MULT_mult_6_n559), .B(MULT_mult_6_n560), 
        .ZN(MULT_mult_6_SUMB_17__3_) );
  INV_X4 MULT_mult_6_U2003 ( .A(MULT_mult_6_net149605), .ZN(
        MULT_mult_6_net92405) );
  NAND2_X2 MULT_mult_6_U2001 ( .A1(MULT_mult_6_n886), .A2(MULT_mult_6_n887), 
        .ZN(MULT_mult_6_n558) );
  NAND2_X4 MULT_mult_6_U2000 ( .A1(MULT_mult_6_n1709), .A2(MULT_mult_6_n1710), 
        .ZN(MULT_mult_6_n2031) );
  NAND2_X2 MULT_mult_6_U1999 ( .A1(MULT_mult_6_CARRYB_8__15_), .A2(
        MULT_mult_6_n151), .ZN(MULT_mult_6_n2048) );
  NAND3_X4 MULT_mult_6_U1998 ( .A1(MULT_mult_6_n2048), .A2(MULT_mult_6_n2049), 
        .A3(MULT_mult_6_n2050), .ZN(MULT_mult_6_CARRYB_9__15_) );
  NOR2_X2 MULT_mult_6_U1997 ( .A1(MULT_mult_6_net84698), .A2(
        MULT_mult_6_net77926), .ZN(MULT_mult_6_ab_8__14_) );
  NAND2_X2 MULT_mult_6_U1996 ( .A1(MULT_mult_6_net88407), .A2(
        MULT_mult_6_net88408), .ZN(MULT_mult_6_net88410) );
  INV_X8 MULT_mult_6_U1994 ( .A(MULT_mult_6__UDW__112704_net78605), .ZN(
        MULT_mult_6_SUMB_1__13_) );
  XNOR2_X2 MULT_mult_6_U1993 ( .A(MULT_mult_6_ab_3__21_), .B(
        MULT_mult_6_CARRYB_2__21_), .ZN(MULT_mult_6_n557) );
  INV_X4 MULT_mult_6_U1992 ( .A(MULT_mult_6_SUMB_9__16_), .ZN(
        MULT_mult_6_n1220) );
  INV_X4 MULT_mult_6_U1991 ( .A(MULT_mult_6_n554), .ZN(MULT_mult_6_n555) );
  NAND2_X2 MULT_mult_6_U1990 ( .A1(MULT_mult_6_ab_20__2_), .A2(
        MULT_mult_6_SUMB_19__3_), .ZN(MULT_mult_6_n1914) );
  NAND2_X2 MULT_mult_6_U1989 ( .A1(MULT_mult_6_n1699), .A2(MULT_mult_6_n1698), 
        .ZN(MULT_mult_6_n1701) );
  INV_X4 MULT_mult_6_U1988 ( .A(MULT_mult_6_net149916), .ZN(
        MULT_mult_6_net149917) );
  INV_X4 MULT_mult_6_U1987 ( .A(MULT_mult_6_net85096), .ZN(
        MULT_mult_6_net149916) );
  INV_X4 MULT_mult_6_U1986 ( .A(MULT_mult_6_net148015), .ZN(
        MULT_mult_6_net148302) );
  XNOR2_X2 MULT_mult_6_U1985 ( .A(MULT_mult_6_net87619), .B(
        MULT_mult_6_ab_18__7_), .ZN(MULT_mult_6_n549) );
  NAND2_X2 MULT_mult_6_U1984 ( .A1(MULT_mult_6_net83776), .A2(
        MULT_mult_6_CARRYB_16__8_), .ZN(MULT_mult_6_n551) );
  INV_X1 MULT_mult_6_U1983 ( .A(MULT_mult_6_n550), .ZN(MULT_mult_6_net93410)
         );
  INV_X8 MULT_mult_6_U1982 ( .A(MULT_mult_6_CARRYB_16__8_), .ZN(
        MULT_mult_6_n550) );
  NAND2_X4 MULT_mult_6_U1981 ( .A1(MULT_mult_6_n550), .A2(
        MULT_mult_6_ab_17__8_), .ZN(MULT_mult_6_net84374) );
  NAND2_X4 MULT_mult_6_U1980 ( .A1(MULT_mult_6_n551), .A2(MULT_mult_6_net84374), .ZN(MULT_mult_6_n548) );
  XNOR2_X2 MULT_mult_6_U1979 ( .A(MULT_mult_6_n548), .B(
        MULT_mult_6_SUMB_16__9_), .ZN(MULT_mult_6_n552) );
  NAND2_X4 MULT_mult_6_U1978 ( .A1(MULT_mult_6_SUMB_17__8_), .A2(
        MULT_mult_6_ab_18__7_), .ZN(MULT_mult_6_net81065) );
  NAND2_X4 MULT_mult_6_U1977 ( .A1(MULT_mult_6_SUMB_17__8_), .A2(
        MULT_mult_6_net87619), .ZN(MULT_mult_6_net81066) );
  INV_X4 MULT_mult_6_U1976 ( .A(MULT_mult_6_n552), .ZN(MULT_mult_6_SUMB_17__8_) );
  INV_X4 MULT_mult_6_U1975 ( .A(MULT_mult_6_net84348), .ZN(MULT_mult_6_n543)
         );
  NAND2_X4 MULT_mult_6_U1974 ( .A1(MULT_mult_6_n543), .A2(MULT_mult_6_n544), 
        .ZN(MULT_mult_6_n546) );
  NAND2_X2 MULT_mult_6_U1972 ( .A1(MULT_mult_6_net84348), .A2(MULT_mult_6_n547), .ZN(MULT_mult_6_n545) );
  NAND2_X4 MULT_mult_6_U1971 ( .A1(MULT_mult_6_n546), .A2(MULT_mult_6_n545), 
        .ZN(MULT_mult_6_SUMB_20__6_) );
  NAND2_X1 MULT_mult_6_U1970 ( .A1(MULT_mult_6_net83172), .A2(MULT_mult_6_n541), .ZN(MULT_mult_6_net83175) );
  INV_X4 MULT_mult_6_U1969 ( .A(MULT_mult_6_CARRYB_20__3_), .ZN(
        MULT_mult_6_n541) );
  NAND2_X4 MULT_mult_6_U1968 ( .A1(MULT_mult_6_n542), .A2(
        MULT_mult_6_SUMB_20__4_), .ZN(MULT_mult_6_net80511) );
  NOR2_X4 MULT_mult_6_U1967 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70451), .ZN(MULT_mult_6_ab_22__3_) );
  NAND3_X2 MULT_mult_6_U1966 ( .A1(MULT_mult_6_net80509), .A2(
        MULT_mult_6_net80511), .A3(MULT_mult_6_net80510), .ZN(
        MULT_mult_6_net124949) );
  XNOR2_X2 MULT_mult_6_U1965 ( .A(MULT_mult_6_SUMB_21__4_), .B(
        MULT_mult_6_ab_22__3_), .ZN(MULT_mult_6_net81493) );
  INV_X4 MULT_mult_6_U1964 ( .A(WIRE_ALU_A_MUX2TO1_32BIT_7__MUX_N1), .ZN(
        MULT_mult_6_net70447) );
  NOR2_X1 MULT_mult_6_U1963 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70447), .ZN(MULT_mult_6_ab_24__3_) );
  INV_X4 MULT_mult_6_U1962 ( .A(MULT_mult_6_net82024), .ZN(MULT_mult_6_n537)
         );
  NAND2_X4 MULT_mult_6_U1961 ( .A1(MULT_mult_6_SUMB_1__18_), .A2(
        MULT_mult_6_ab_2__17_), .ZN(MULT_mult_6_net82027) );
  INV_X8 MULT_mult_6_U1960 ( .A(MULT_mult_6_n536), .ZN(MULT_mult_6_SUMB_1__18_) );
  NAND2_X4 MULT_mult_6_U1959 ( .A1(MULT_mult_6_n540), .A2(MULT_mult_6_n539), 
        .ZN(MULT_mult_6_net84327) );
  NAND2_X2 MULT_mult_6_U1958 ( .A1(MULT_mult_6_net149526), .A2(
        MULT_mult_6_net88123), .ZN(MULT_mult_6_net123430) );
  NAND2_X4 MULT_mult_6_U1957 ( .A1(MULT_mult_6_ab_0__17_), .A2(
        MULT_mult_6_net88123), .ZN(MULT_mult_6__UDW__112689_net78561) );
  NOR2_X4 MULT_mult_6_U1956 ( .A1(MULT_mult_6_ab_2__16_), .A2(
        MULT_mult_6_CARRYB_1__16_), .ZN(MULT_mult_6_net119901) );
  INV_X8 MULT_mult_6_U1955 ( .A(MULT_mult_6__UDW__112689_net78561), .ZN(
        MULT_mult_6_CARRYB_1__16_) );
  NAND2_X2 MULT_mult_6_U1954 ( .A1(MULT_mult_6_CARRYB_1__16_), .A2(
        MULT_mult_6_ab_2__16_), .ZN(MULT_mult_6_net119899) );
  NAND2_X4 MULT_mult_6_U1953 ( .A1(MULT_mult_6_CARRYB_28__1_), .A2(
        MULT_mult_6_ab_29__1_), .ZN(MULT_mult_6_net85096) );
  INV_X4 MULT_mult_6_U1952 ( .A(MULT_mult_6_net92337), .ZN(
        MULT_mult_6_ab_29__1_) );
  NAND2_X4 MULT_mult_6_U1951 ( .A1(MULT_mult_6_net85094), .A2(
        MULT_mult_6_net92337), .ZN(MULT_mult_6_n532) );
  INV_X4 MULT_mult_6_U1950 ( .A(MULT_mult_6_n402), .ZN(MULT_mult_6_n530) );
  NAND2_X4 MULT_mult_6_U1949 ( .A1(MULT_mult_6_n533), .A2(MULT_mult_6_n530), 
        .ZN(MULT_mult_6_n535) );
  NAND2_X2 MULT_mult_6_U1948 ( .A1(MULT_mult_6_SUMB_28__2_), .A2(
        MULT_mult_6_ab_29__1_), .ZN(MULT_mult_6_net80667) );
  XNOR2_X2 MULT_mult_6_U1947 ( .A(MULT_mult_6_net81158), .B(MULT_mult_6_n4), 
        .ZN(MULT_mult_6_net89453) );
  NAND2_X4 MULT_mult_6_U1946 ( .A1(MULT_mult_6_n535), .A2(MULT_mult_6_n534), 
        .ZN(MULT_mult_6_SUMB_28__2_) );
  XNOR2_X2 MULT_mult_6_U1945 ( .A(MULT_mult_6_n531), .B(MULT_mult_6_n200), 
        .ZN(MULT_mult_6_net86055) );
  INV_X4 MULT_mult_6_U1944 ( .A(WIRE_ALU_A_MUX2TO1_32BIT_4__MUX_N1), .ZN(
        MULT_mult_6_net70441) );
  NAND2_X4 MULT_mult_6_U1943 ( .A1(MULT_mult_6_net119817), .A2(
        MULT_mult_6_ab_4__14_), .ZN(MULT_mult_6_n528) );
  NAND3_X4 MULT_mult_6_U1942 ( .A1(MULT_mult_6_n529), .A2(MULT_mult_6_n528), 
        .A3(MULT_mult_6_net92718), .ZN(MULT_mult_6_CARRYB_4__14_) );
  NOR2_X1 MULT_mult_6_U1941 ( .A1(MULT_mult_6_net36614), .A2(
        MULT_mult_6_net77866), .ZN(MULT_mult_6_net81548) );
  INV_X4 MULT_mult_6_U1940 ( .A(WIRE_ALU_A_MUX2TO1_32BIT_1__MUX_N1), .ZN(
        MULT_mult_6_net36614) );
  NOR2_X1 MULT_mult_6_U1939 ( .A1(MULT_mult_6_net36614), .A2(
        MULT_mult_6_net77858), .ZN(MULT_mult_6_ab_30__0_) );
  XNOR2_X2 MULT_mult_6_U1938 ( .A(MULT_mult_6_net83536), .B(
        MULT_mult_6_net86055), .ZN(multOut[1]) );
  NAND2_X4 MULT_mult_6_U1937 ( .A1(MULT_mult_6_net88856), .A2(
        MULT_mult_6_SUMB_18__7_), .ZN(MULT_mult_6_net81069) );
  INV_X16 MULT_mult_6_U1936 ( .A(WIRE_ALU_A_MUX2TO1_32BIT_10__MUX_N1), .ZN(
        MULT_mult_6_net70453) );
  NOR2_X4 MULT_mult_6_U1935 ( .A1(MULT_mult_6_net77900), .A2(
        MULT_mult_6_net70453), .ZN(MULT_mult_6_ab_21__5_) );
  INV_X4 MULT_mult_6_U1934 ( .A(MULT_mult_6_net124367), .ZN(MULT_mult_6_n526)
         );
  NAND2_X4 MULT_mult_6_U1933 ( .A1(MULT_mult_6_net148051), .A2(
        MULT_mult_6_n526), .ZN(MULT_mult_6_n527) );
  NAND2_X4 MULT_mult_6_U1932 ( .A1(MULT_mult_6_n527), .A2(
        MULT_mult_6_net148053), .ZN(MULT_mult_6_net84856) );
  NAND2_X2 MULT_mult_6_U1931 ( .A1(MULT_mult_6_SUMB_4__16_), .A2(
        MULT_mult_6_n137), .ZN(MULT_mult_6_net80840) );
  NAND2_X2 MULT_mult_6_U1930 ( .A1(MULT_mult_6_SUMB_4__16_), .A2(
        MULT_mult_6_ab_5__15_), .ZN(MULT_mult_6_net80839) );
  INV_X8 MULT_mult_6_U1929 ( .A(MULT_mult_6_net84856), .ZN(
        MULT_mult_6_SUMB_4__16_) );
  NAND2_X4 MULT_mult_6_U1928 ( .A1(MULT_mult_6_net84445), .A2(
        MULT_mult_6_net84446), .ZN(MULT_mult_6_SUMB_5__15_) );
  NOR2_X1 MULT_mult_6_U1927 ( .A1(MULT_mult_6_net84698), .A2(
        MULT_mult_6_net77940), .ZN(MULT_mult_6_ab_6__14_) );
  NAND2_X2 MULT_mult_6_U1926 ( .A1(MULT_mult_6_net83919), .A2(
        MULT_mult_6_CARRYB_4__14_), .ZN(MULT_mult_6_net82297) );
  INV_X2 MULT_mult_6_U1925 ( .A(MULT_mult_6_CARRYB_6__14_), .ZN(
        MULT_mult_6_net88880) );
  INV_X4 MULT_mult_6_U1924 ( .A(MULT_mult_6_SUMB_6__14_), .ZN(
        MULT_mult_6_net88660) );
  NAND2_X4 MULT_mult_6_U1923 ( .A1(MULT_mult_6_net90897), .A2(
        MULT_mult_6_ab_7__13_), .ZN(MULT_mult_6_net80844) );
  NAND2_X4 MULT_mult_6_U1922 ( .A1(MULT_mult_6_net90897), .A2(
        MULT_mult_6_net88444), .ZN(MULT_mult_6_net80845) );
  INV_X8 MULT_mult_6_U1921 ( .A(MULT_mult_6_net88660), .ZN(
        MULT_mult_6_net90897) );
  XNOR2_X2 MULT_mult_6_U1920 ( .A(MULT_mult_6_net90897), .B(
        MULT_mult_6_net81756), .ZN(MULT_mult_6_net90348) );
  XNOR2_X2 MULT_mult_6_U1919 ( .A(MULT_mult_6_CARRYB_24__1_), .B(
        MULT_mult_6_ab_25__1_), .ZN(MULT_mult_6_net124874) );
  NAND2_X4 MULT_mult_6_U1918 ( .A1(MULT_mult_6_SUMB_24__2_), .A2(
        MULT_mult_6_ab_25__1_), .ZN(MULT_mult_6_n524) );
  NAND2_X4 MULT_mult_6_U1917 ( .A1(MULT_mult_6_CARRYB_24__1_), .A2(
        MULT_mult_6_SUMB_24__2_), .ZN(MULT_mult_6_n523) );
  NAND2_X4 MULT_mult_6_U1916 ( .A1(MULT_mult_6_CARRYB_24__1_), .A2(
        MULT_mult_6_ab_25__1_), .ZN(MULT_mult_6_n525) );
  INV_X1 MULT_mult_6_U1915 ( .A(MULT_mult_6_CARRYB_25__1_), .ZN(
        MULT_mult_6_net88655) );
  NAND3_X4 MULT_mult_6_U1914 ( .A1(MULT_mult_6_n523), .A2(MULT_mult_6_n524), 
        .A3(MULT_mult_6_n525), .ZN(MULT_mult_6_CARRYB_25__1_) );
  XNOR2_X2 MULT_mult_6_U1913 ( .A(MULT_mult_6_CARRYB_16__7_), .B(
        MULT_mult_6_ab_17__7_), .ZN(MULT_mult_6_n522) );
  NAND2_X2 MULT_mult_6_U1912 ( .A1(MULT_mult_6_SUMB_17__7_), .A2(
        MULT_mult_6_ab_18__6_), .ZN(MULT_mult_6_net81269) );
  XNOR2_X2 MULT_mult_6_U1911 ( .A(MULT_mult_6_n522), .B(
        MULT_mult_6_SUMB_16__8_), .ZN(MULT_mult_6_SUMB_17__7_) );
  NAND2_X2 MULT_mult_6_U1910 ( .A1(MULT_mult_6_SUMB_15__7_), .A2(
        MULT_mult_6_net90347), .ZN(MULT_mult_6_net80541) );
  NAND2_X2 MULT_mult_6_U1909 ( .A1(MULT_mult_6_SUMB_15__7_), .A2(
        MULT_mult_6_ab_16__6_), .ZN(MULT_mult_6_net80540) );
  NAND2_X2 MULT_mult_6_U1908 ( .A1(MULT_mult_6_net90347), .A2(
        MULT_mult_6_ab_16__6_), .ZN(MULT_mult_6_n521) );
  NAND3_X2 MULT_mult_6_U1907 ( .A1(MULT_mult_6_net80541), .A2(
        MULT_mult_6_net80540), .A3(MULT_mult_6_n521), .ZN(
        MULT_mult_6_CARRYB_16__6_) );
  INV_X16 MULT_mult_6_U1906 ( .A(WIRE_ALU_A_MUX2TO1_32BIT_14__MUX_N1), .ZN(
        MULT_mult_6_net70461) );
  NAND2_X4 MULT_mult_6_U1905 ( .A1(MULT_mult_6_net92790), .A2(
        MULT_mult_6_net93840), .ZN(MULT_mult_6_net80261) );
  XNOR2_X2 MULT_mult_6_U1904 ( .A(MULT_mult_6_SUMB_25__2_), .B(
        MULT_mult_6_ab_26__1_), .ZN(MULT_mult_6_net86427) );
  NAND2_X2 MULT_mult_6_U1903 ( .A1(MULT_mult_6_CARRYB_25__1_), .A2(
        MULT_mult_6_SUMB_25__2_), .ZN(MULT_mult_6_net83975) );
  NAND2_X2 MULT_mult_6_U1902 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_2__MUX_N1), .A2(
        n6005), .ZN(MULT_mult_6_net92341) );
  XNOR2_X2 MULT_mult_6_U1901 ( .A(MULT_mult_6_net90348), .B(
        MULT_mult_6_net85212), .ZN(MULT_mult_6_net90687) );
  NOR2_X2 MULT_mult_6_U1900 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__12_) );
  INV_X16 MULT_mult_6_U1899 ( .A(n10916), .ZN(MULT_mult_6_net123000) );
  NAND2_X2 MULT_mult_6_U1898 ( .A1(MULT_mult_6_net86959), .A2(
        MULT_mult_6_net87050), .ZN(MULT_mult_6_n520) );
  NOR2_X4 MULT_mult_6_U1897 ( .A1(MULT_mult_6_net70470), .A2(
        MULT_mult_6_net82149), .ZN(MULT_mult_6_net85688) );
  NAND2_X4 MULT_mult_6_U1896 ( .A1(MULT_mult_6_net85688), .A2(
        MULT_mult_6_ab_1__17_), .ZN(MULT_mult_6__UDW__112684_net78547) );
  NAND2_X4 MULT_mult_6_U1895 ( .A1(MULT_mult_6_net82286), .A2(MULT_mult_6_n520), .ZN(MULT_mult_6__UDW__112684_net78549) );
  NAND2_X2 MULT_mult_6_U1894 ( .A1(MULT_mult_6_ab_18__6_), .A2(
        MULT_mult_6_net85611), .ZN(MULT_mult_6_net81268) );
  NAND3_X2 MULT_mult_6_U1893 ( .A1(MULT_mult_6_net81270), .A2(
        MULT_mult_6_net81269), .A3(MULT_mult_6_net81268), .ZN(
        MULT_mult_6_net124627) );
  NAND2_X2 MULT_mult_6_U1892 ( .A1(MULT_mult_6_SUMB_17__7_), .A2(
        MULT_mult_6_net85611), .ZN(MULT_mult_6_net81270) );
  INV_X4 MULT_mult_6_U1891 ( .A(n10924), .ZN(MULT_mult_6_net77908) );
  INV_X16 MULT_mult_6_U1890 ( .A(WIRE_ALU_A_MUX2TO1_32BIT_12__MUX_N1), .ZN(
        MULT_mult_6_net70457) );
  NAND2_X4 MULT_mult_6_U1889 ( .A1(MULT_mult_6_SUMB_18__7_), .A2(
        MULT_mult_6_ab_19__6_), .ZN(MULT_mult_6_net81068) );
  NAND2_X2 MULT_mult_6_U1888 ( .A1(MULT_mult_6_ab_19__6_), .A2(
        MULT_mult_6_net124627), .ZN(MULT_mult_6_net81067) );
  NOR2_X4 MULT_mult_6_U1887 ( .A1(MULT_mult_6_net77908), .A2(
        MULT_mult_6_net70457), .ZN(MULT_mult_6_ab_19__6_) );
  NAND3_X2 MULT_mult_6_U1886 ( .A1(MULT_mult_6_net81270), .A2(
        MULT_mult_6_net81269), .A3(MULT_mult_6_net81268), .ZN(
        MULT_mult_6_net93914) );
  NAND2_X4 MULT_mult_6_U1885 ( .A1(MULT_mult_6_n518), .A2(MULT_mult_6_n519), 
        .ZN(MULT_mult_6_net90810) );
  INV_X8 MULT_mult_6_U1884 ( .A(n10925), .ZN(MULT_mult_6_net70444) );
  INV_X16 MULT_mult_6_U1883 ( .A(WIRE_ALU_A_MUX2TO1_32BIT_11__MUX_N1), .ZN(
        MULT_mult_6_net70455) );
  INV_X1 MULT_mult_6_U1882 ( .A(MULT_mult_6_ab_20__5_), .ZN(
        MULT_mult_6_net120626) );
  NOR2_X4 MULT_mult_6_U1881 ( .A1(MULT_mult_6_net77900), .A2(
        MULT_mult_6_net70455), .ZN(MULT_mult_6_ab_20__5_) );
  NAND2_X2 MULT_mult_6_U1880 ( .A1(MULT_mult_6_SUMB_19__6_), .A2(
        MULT_mult_6_ab_20__5_), .ZN(MULT_mult_6_net82405) );
  NAND3_X2 MULT_mult_6_U1879 ( .A1(MULT_mult_6_net81374), .A2(
        MULT_mult_6_net81375), .A3(MULT_mult_6_net81373), .ZN(
        MULT_mult_6_CARRYB_9__12_) );
  NAND2_X4 MULT_mult_6_U1878 ( .A1(MULT_mult_6_net89356), .A2(
        MULT_mult_6_net88943), .ZN(MULT_mult_6_net81372) );
  NAND2_X4 MULT_mult_6_U1877 ( .A1(MULT_mult_6_SUMB_7__14_), .A2(
        MULT_mult_6_ab_8__13_), .ZN(MULT_mult_6_net81371) );
  INV_X2 MULT_mult_6_U1876 ( .A(MULT_mult_6_net84868), .ZN(
        MULT_mult_6_net89149) );
  INV_X1 MULT_mult_6_U1875 ( .A(MULT_mult_6_ab_9__12_), .ZN(
        MULT_mult_6_net84867) );
  NAND2_X4 MULT_mult_6_U1874 ( .A1(MULT_mult_6_net88841), .A2(
        MULT_mult_6_net82837), .ZN(MULT_mult_6_net84671) );
  NAND2_X4 MULT_mult_6_U1873 ( .A1(MULT_mult_6_net84870), .A2(
        MULT_mult_6_net81373), .ZN(MULT_mult_6_net82837) );
  NAND2_X2 MULT_mult_6_U1872 ( .A1(MULT_mult_6_net89356), .A2(
        MULT_mult_6_net81958), .ZN(MULT_mult_6_net85461) );
  INV_X4 MULT_mult_6_U1871 ( .A(MULT_mult_6_net81958), .ZN(
        MULT_mult_6_net85459) );
  NAND2_X4 MULT_mult_6_U1870 ( .A1(MULT_mult_6_net85459), .A2(
        MULT_mult_6_net85460), .ZN(MULT_mult_6_n517) );
  INV_X4 MULT_mult_6_U1868 ( .A(MULT_mult_6_net82837), .ZN(
        MULT_mult_6_net84669) );
  INV_X4 MULT_mult_6_U1867 ( .A(MULT_mult_6_net84670), .ZN(
        MULT_mult_6_net88841) );
  INV_X4 MULT_mult_6_U1866 ( .A(MULT_mult_6_n2360), .ZN(MULT_mult_6_net84670)
         );
  NAND2_X4 MULT_mult_6_U1865 ( .A1(MULT_mult_6_net84669), .A2(
        MULT_mult_6_net84670), .ZN(MULT_mult_6_net84672) );
  NAND2_X1 MULT_mult_6_U1864 ( .A1(MULT_mult_6_ab_10__11_), .A2(
        MULT_mult_6_CARRYB_9__11_), .ZN(MULT_mult_6_net80958) );
  NAND2_X2 MULT_mult_6_U1863 ( .A1(MULT_mult_6_CARRYB_9__11_), .A2(
        MULT_mult_6_ab_10__11_), .ZN(MULT_mult_6_n515) );
  INV_X4 MULT_mult_6_U1862 ( .A(MULT_mult_6_CARRYB_9__11_), .ZN(
        MULT_mult_6_n514) );
  NAND2_X4 MULT_mult_6_U1861 ( .A1(MULT_mult_6_n514), .A2(MULT_mult_6_net83876), .ZN(MULT_mult_6_n516) );
  NAND2_X4 MULT_mult_6_U1860 ( .A1(MULT_mult_6_n516), .A2(MULT_mult_6_n515), 
        .ZN(MULT_mult_6_net82838) );
  NAND2_X4 MULT_mult_6_U1859 ( .A1(MULT_mult_6_net82838), .A2(
        MULT_mult_6_net91003), .ZN(MULT_mult_6_net87366) );
  NAND2_X4 MULT_mult_6_U1858 ( .A1(MULT_mult_6_net84672), .A2(
        MULT_mult_6_net84671), .ZN(MULT_mult_6_net91003) );
  INV_X4 MULT_mult_6_U1857 ( .A(MULT_mult_6_net82838), .ZN(
        MULT_mult_6_net87365) );
  NAND2_X2 MULT_mult_6_U1856 ( .A1(MULT_mult_6_net87366), .A2(
        MULT_mult_6_net87367), .ZN(MULT_mult_6_net91243) );
  NAND2_X4 MULT_mult_6_U1855 ( .A1(MULT_mult_6_net87367), .A2(
        MULT_mult_6_net87366), .ZN(MULT_mult_6_SUMB_10__11_) );
  NAND2_X4 MULT_mult_6_U1854 ( .A1(MULT_mult_6_net87365), .A2(
        MULT_mult_6_net87364), .ZN(MULT_mult_6_net87367) );
  NAND2_X1 MULT_mult_6_U1853 ( .A1(n10928), .A2(MULT_mult_6_net80392), .ZN(
        MULT_mult_6_net70435) );
  NAND2_X1 MULT_mult_6_U1852 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_3__MUX_N1), .A2(
        n10926), .ZN(MULT_mult_6_net92320) );
  INV_X4 MULT_mult_6_U1851 ( .A(n10928), .ZN(MULT_mult_6_net70436) );
  INV_X32 MULT_mult_6_U1850 ( .A(MULT_mult_6_net77864), .ZN(
        MULT_mult_6_net77860) );
  NAND2_X1 MULT_mult_6_U1849 ( .A1(MULT_mult_6_CARRYB_10__10_), .A2(
        MULT_mult_6_ab_11__10_), .ZN(MULT_mult_6_net92862) );
  INV_X2 MULT_mult_6_U1848 ( .A(MULT_mult_6_SUMB_10__11_), .ZN(
        MULT_mult_6_net85373) );
  NAND2_X1 MULT_mult_6_U1847 ( .A1(MULT_mult_6_ab_11__10_), .A2(
        MULT_mult_6_CARRYB_10__10_), .ZN(MULT_mult_6_net83882) );
  NAND2_X2 MULT_mult_6_U1846 ( .A1(MULT_mult_6_SUMB_10__11_), .A2(
        MULT_mult_6_ab_11__10_), .ZN(MULT_mult_6_net83881) );
  NAND2_X2 MULT_mult_6_U1845 ( .A1(MULT_mult_6_n201), .A2(MULT_mult_6_net87045), .ZN(MULT_mult_6_net92863) );
  INV_X1 MULT_mult_6_U1844 ( .A(MULT_mult_6_n201), .ZN(MULT_mult_6_net121898)
         );
  NAND3_X2 MULT_mult_6_U1843 ( .A1(MULT_mult_6_net83880), .A2(
        MULT_mult_6_net83881), .A3(MULT_mult_6_net83882), .ZN(
        MULT_mult_6_CARRYB_11__10_) );
  NAND2_X2 MULT_mult_6_U1842 ( .A1(MULT_mult_6_net121898), .A2(
        MULT_mult_6_SUMB_10__11_), .ZN(MULT_mult_6_net83880) );
  NOR2_X2 MULT_mult_6_U1841 ( .A1(MULT_mult_6_net91660), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__10_) );
  XNOR2_X2 MULT_mult_6_U1840 ( .A(MULT_mult_6_SUMB_27__1_), .B(
        MULT_mult_6_n345), .ZN(MULT_mult_6_net92378) );
  NAND2_X4 MULT_mult_6_U1839 ( .A1(MULT_mult_6_SUMB_27__1_), .A2(
        MULT_mult_6_n345), .ZN(MULT_mult_6_net80771) );
  NAND2_X4 MULT_mult_6_U1838 ( .A1(MULT_mult_6_CARRYB_27__0_), .A2(
        MULT_mult_6_n345), .ZN(MULT_mult_6_n513) );
  NAND3_X4 MULT_mult_6_U1837 ( .A1(MULT_mult_6_net80768), .A2(
        MULT_mult_6_net80769), .A3(MULT_mult_6_net80767), .ZN(
        MULT_mult_6_CARRYB_27__0_) );
  NAND3_X4 MULT_mult_6_U1836 ( .A1(MULT_mult_6_net80773), .A2(MULT_mult_6_n513), .A3(MULT_mult_6_net80771), .ZN(MULT_mult_6_CARRYB_28__0_) );
  NAND2_X4 MULT_mult_6_U1835 ( .A1(MULT_mult_6_SUMB_27__1_), .A2(
        MULT_mult_6_CARRYB_27__0_), .ZN(MULT_mult_6_net80773) );
  INV_X4 MULT_mult_6_U1834 ( .A(MULT_mult_6_SUMB_17__6_), .ZN(
        MULT_mult_6_net86661) );
  INV_X4 MULT_mult_6_U1833 ( .A(MULT_mult_6_net85610), .ZN(
        MULT_mult_6_net85611) );
  XNOR2_X2 MULT_mult_6_U1832 ( .A(MULT_mult_6_net85611), .B(
        MULT_mult_6_net82748), .ZN(MULT_mult_6_net81264) );
  XNOR2_X2 MULT_mult_6_U1831 ( .A(MULT_mult_6_net81264), .B(
        MULT_mult_6_SUMB_17__7_), .ZN(MULT_mult_6_net88878) );
  NAND2_X4 MULT_mult_6_U1830 ( .A1(MULT_mult_6_SUMB_18__6_), .A2(
        MULT_mult_6_net148582), .ZN(MULT_mult_6_n512) );
  XNOR2_X2 MULT_mult_6_U1829 ( .A(MULT_mult_6_SUMB_18__6_), .B(
        MULT_mult_6_net92542), .ZN(MULT_mult_6_net88887) );
  XNOR2_X2 MULT_mult_6_U1828 ( .A(MULT_mult_6_n8), .B(MULT_mult_6_net92542), 
        .ZN(MULT_mult_6_SUMB_19__5_) );
  NAND2_X4 MULT_mult_6_U1827 ( .A1(MULT_mult_6_SUMB_18__6_), .A2(
        MULT_mult_6_ab_19__5_), .ZN(MULT_mult_6_n511) );
  NAND2_X2 MULT_mult_6_U1826 ( .A1(MULT_mult_6_net91377), .A2(
        MULT_mult_6_ab_20__5_), .ZN(MULT_mult_6_net120627) );
  NAND3_X4 MULT_mult_6_U1825 ( .A1(MULT_mult_6_n512), .A2(MULT_mult_6_n511), 
        .A3(MULT_mult_6_net84708), .ZN(MULT_mult_6_net91377) );
  XNOR2_X2 MULT_mult_6_U1824 ( .A(MULT_mult_6_net90810), .B(
        MULT_mult_6_net90576), .ZN(MULT_mult_6_SUMB_19__6_) );
  INV_X2 MULT_mult_6_U1823 ( .A(MULT_mult_6_net124589), .ZN(
        MULT_mult_6_net147929) );
  NAND2_X2 MULT_mult_6_U1822 ( .A1(MULT_mult_6_net83202), .A2(
        MULT_mult_6_net124589), .ZN(MULT_mult_6_net147930) );
  XNOR2_X2 MULT_mult_6_U1821 ( .A(MULT_mult_6_net90810), .B(
        MULT_mult_6_net90576), .ZN(MULT_mult_6_net124589) );
  INV_X8 MULT_mult_6_U1820 ( .A(MULT_mult_6_net91377), .ZN(
        MULT_mult_6_net120625) );
  NAND2_X4 MULT_mult_6_U1819 ( .A1(MULT_mult_6_net86806), .A2(
        MULT_mult_6_ab_20__5_), .ZN(MULT_mult_6_net82403) );
  NAND3_X4 MULT_mult_6_U1818 ( .A1(MULT_mult_6_net82404), .A2(
        MULT_mult_6_net82403), .A3(MULT_mult_6_net82405), .ZN(
        MULT_mult_6_CARRYB_20__5_) );
  NAND2_X4 MULT_mult_6_U1817 ( .A1(MULT_mult_6_net124589), .A2(
        MULT_mult_6_net86806), .ZN(MULT_mult_6_net82404) );
  CLKBUF_X3 MULT_mult_6_U1816 ( .A(MULT_mult_6_net84873), .Z(
        MULT_mult_6_net88455) );
  NAND3_X2 MULT_mult_6_U1815 ( .A1(MULT_mult_6_net88295), .A2(
        MULT_mult_6_net88296), .A3(MULT_mult_6_net88297), .ZN(
        MULT_mult_6_CARRYB_12__9_) );
  NAND2_X1 MULT_mult_6_U1814 ( .A1(MULT_mult_6_ab_13__9_), .A2(
        MULT_mult_6_CARRYB_12__9_), .ZN(MULT_mult_6_net81059) );
  NAND2_X4 MULT_mult_6_U1813 ( .A1(MULT_mult_6_n510), .A2(MULT_mult_6_net86142), .ZN(MULT_mult_6_net86145) );
  INV_X4 MULT_mult_6_U1812 ( .A(MULT_mult_6_net81182), .ZN(
        MULT_mult_6_net86142) );
  INV_X1 MULT_mult_6_U1811 ( .A(MULT_mult_6_ab_13__9_), .ZN(
        MULT_mult_6_net81182) );
  NAND2_X4 MULT_mult_6_U1810 ( .A1(MULT_mult_6_CARRYB_12__9_), .A2(
        MULT_mult_6_net81182), .ZN(MULT_mult_6_net86144) );
  NAND2_X4 MULT_mult_6_U1809 ( .A1(MULT_mult_6_net86145), .A2(
        MULT_mult_6_net86144), .ZN(MULT_mult_6_net92622) );
  NAND2_X2 MULT_mult_6_U1808 ( .A1(MULT_mult_6_SUMB_12__10_), .A2(
        MULT_mult_6_ab_13__9_), .ZN(MULT_mult_6_net81060) );
  INV_X4 MULT_mult_6_U1807 ( .A(MULT_mult_6_net83848), .ZN(
        MULT_mult_6_SUMB_12__10_) );
  INV_X4 MULT_mult_6_U1806 ( .A(MULT_mult_6_net92622), .ZN(
        MULT_mult_6_net82292) );
  NAND2_X4 MULT_mult_6_U1805 ( .A1(MULT_mult_6_SUMB_12__10_), .A2(
        MULT_mult_6_net82292), .ZN(MULT_mult_6_net82295) );
  NAND2_X2 MULT_mult_6_U1804 ( .A1(MULT_mult_6_net92622), .A2(
        MULT_mult_6_net83848), .ZN(MULT_mult_6_net82294) );
  NAND2_X1 MULT_mult_6_U1803 ( .A1(MULT_mult_6_ab_12__10_), .A2(
        MULT_mult_6_CARRYB_11__10_), .ZN(MULT_mult_6_net81056) );
  XNOR2_X2 MULT_mult_6_U1802 ( .A(MULT_mult_6_net89065), .B(
        MULT_mult_6_net80983), .ZN(MULT_mult_6_net89167) );
  NAND3_X2 MULT_mult_6_U1801 ( .A1(MULT_mult_6_net80957), .A2(
        MULT_mult_6_net80956), .A3(MULT_mult_6_net80958), .ZN(
        MULT_mult_6_CARRYB_10__11_) );
  INV_X1 MULT_mult_6_U1800 ( .A(MULT_mult_6_n508), .ZN(MULT_mult_6_net87490)
         );
  INV_X4 MULT_mult_6_U1799 ( .A(MULT_mult_6_CARRYB_10__11_), .ZN(
        MULT_mult_6_n508) );
  NAND2_X4 MULT_mult_6_U1798 ( .A1(MULT_mult_6_n508), .A2(
        MULT_mult_6_ab_11__11_), .ZN(MULT_mult_6_net85539) );
  INV_X1 MULT_mult_6_U1797 ( .A(MULT_mult_6_ab_11__11_), .ZN(
        MULT_mult_6_net85537) );
  NAND2_X2 MULT_mult_6_U1796 ( .A1(MULT_mult_6_net88525), .A2(
        MULT_mult_6_net85537), .ZN(MULT_mult_6_n509) );
  NAND2_X4 MULT_mult_6_U1795 ( .A1(MULT_mult_6_net85539), .A2(MULT_mult_6_n509), .ZN(MULT_mult_6_net81165) );
  NAND3_X2 MULT_mult_6_U1794 ( .A1(MULT_mult_6_net83880), .A2(
        MULT_mult_6_net83882), .A3(MULT_mult_6_net83881), .ZN(
        MULT_mult_6_net89369) );
  INV_X4 MULT_mult_6_U1793 ( .A(MULT_mult_6_net89369), .ZN(
        MULT_mult_6_net92550) );
  INV_X1 MULT_mult_6_U1792 ( .A(MULT_mult_6_ab_12__10_), .ZN(
        MULT_mult_6_net88303) );
  INV_X4 MULT_mult_6_U1791 ( .A(MULT_mult_6_net88303), .ZN(
        MULT_mult_6_net92551) );
  NAND2_X4 MULT_mult_6_U1790 ( .A1(MULT_mult_6_net92552), .A2(
        MULT_mult_6_net92553), .ZN(MULT_mult_6_net88302) );
  NAND2_X2 MULT_mult_6_U1789 ( .A1(MULT_mult_6_net81165), .A2(
        MULT_mult_6_net89167), .ZN(MULT_mult_6_n506) );
  INV_X4 MULT_mult_6_U1788 ( .A(MULT_mult_6_net89167), .ZN(MULT_mult_6_n504)
         );
  INV_X4 MULT_mult_6_U1787 ( .A(MULT_mult_6_net81165), .ZN(MULT_mult_6_n505)
         );
  NAND2_X2 MULT_mult_6_U1786 ( .A1(MULT_mult_6_net88302), .A2(
        MULT_mult_6_SUMB_11__11_), .ZN(MULT_mult_6_net84873) );
  NAND2_X2 MULT_mult_6_U1785 ( .A1(MULT_mult_6_CARRYB_11__10_), .A2(
        MULT_mult_6_SUMB_11__11_), .ZN(MULT_mult_6_net81058) );
  NAND2_X4 MULT_mult_6_U1784 ( .A1(MULT_mult_6_ab_12__10_), .A2(
        MULT_mult_6_SUMB_11__11_), .ZN(MULT_mult_6_net81057) );
  INV_X8 MULT_mult_6_U1783 ( .A(MULT_mult_6_net89447), .ZN(
        MULT_mult_6_SUMB_11__11_) );
  INV_X4 MULT_mult_6_U1782 ( .A(MULT_mult_6_net88302), .ZN(
        MULT_mult_6_net87043) );
  AND2_X2 MULT_mult_6_U1781 ( .A1(MULT_mult_6_net84874), .A2(
        MULT_mult_6_CARRYB_12__9_), .ZN(MULT_mult_6_net85044) );
  NAND2_X4 MULT_mult_6_U1780 ( .A1(MULT_mult_6_net84874), .A2(
        MULT_mult_6_net84873), .ZN(MULT_mult_6_net83848) );
  NAND2_X4 MULT_mult_6_U1779 ( .A1(MULT_mult_6_net89840), .A2(
        MULT_mult_6_net87043), .ZN(MULT_mult_6_net84874) );
  INV_X8 MULT_mult_6_U1778 ( .A(n10926), .ZN(MULT_mult_6_net77882) );
  BUF_X32 MULT_mult_6_U1777 ( .A(MULT_mult_6_net77882), .Z(
        MULT_mult_6_net77886) );
  NAND2_X2 MULT_mult_6_U1776 ( .A1(MULT_mult_6_ab_22__3_), .A2(
        MULT_mult_6_SUMB_21__4_), .ZN(MULT_mult_6_n501) );
  NAND3_X2 MULT_mult_6_U1775 ( .A1(MULT_mult_6_net80511), .A2(
        MULT_mult_6_net80510), .A3(MULT_mult_6_net80509), .ZN(
        MULT_mult_6_CARRYB_21__3_) );
  NAND3_X2 MULT_mult_6_U1773 ( .A1(MULT_mult_6_n503), .A2(MULT_mult_6_n501), 
        .A3(MULT_mult_6_n502), .ZN(MULT_mult_6_CARRYB_22__3_) );
  NAND2_X4 MULT_mult_6_U1771 ( .A1(MULT_mult_6_net86520), .A2(
        MULT_mult_6_ab_24__2_), .ZN(MULT_mult_6_net80257) );
  INV_X8 MULT_mult_6_U1770 ( .A(MULT_mult_6_net86519), .ZN(
        MULT_mult_6_net86520) );
  NAND2_X4 MULT_mult_6_U1769 ( .A1(MULT_mult_6_net86520), .A2(
        MULT_mult_6_CARRYB_23__2_), .ZN(MULT_mult_6_n500) );
  NAND3_X4 MULT_mult_6_U1768 ( .A1(MULT_mult_6_net80257), .A2(MULT_mult_6_n500), .A3(MULT_mult_6_net80258), .ZN(MULT_mult_6_CARRYB_24__2_) );
  INV_X4 MULT_mult_6_U1766 ( .A(MULT_mult_6_net92568), .ZN(
        MULT_mult_6_net92569) );
  NAND2_X4 MULT_mult_6_U1765 ( .A1(MULT_mult_6_n499), .A2(MULT_mult_6_n498), 
        .ZN(MULT_mult_6_SUMB_25__2_) );
  XNOR2_X2 MULT_mult_6_U1764 ( .A(MULT_mult_6_SUMB_7__13_), .B(
        MULT_mult_6_net85212), .ZN(MULT_mult_6_net91118) );
  XNOR2_X2 MULT_mult_6_U1763 ( .A(MULT_mult_6_net90897), .B(
        MULT_mult_6_net81756), .ZN(MULT_mult_6_SUMB_7__13_) );
  NAND2_X4 MULT_mult_6_U1762 ( .A1(MULT_mult_6_n497), .A2(MULT_mult_6_net85251), .ZN(MULT_mult_6_net85254) );
  INV_X8 MULT_mult_6_U1761 ( .A(MULT_mult_6_CARRYB_6__12_), .ZN(
        MULT_mult_6_n497) );
  INV_X2 MULT_mult_6_U1760 ( .A(MULT_mult_6_n497), .ZN(MULT_mult_6_n492) );
  NAND2_X4 MULT_mult_6_U1759 ( .A1(MULT_mult_6_net124104), .A2(
        MULT_mult_6_n492), .ZN(MULT_mult_6_n496) );
  NAND2_X4 MULT_mult_6_U1758 ( .A1(MULT_mult_6_SUMB_6__13_), .A2(
        MULT_mult_6_ab_7__12_), .ZN(MULT_mult_6_n495) );
  INV_X4 MULT_mult_6_U1757 ( .A(MULT_mult_6_CARRYB_7__12_), .ZN(
        MULT_mult_6_net87309) );
  NAND3_X4 MULT_mult_6_U1756 ( .A1(MULT_mult_6_n494), .A2(MULT_mult_6_n496), 
        .A3(MULT_mult_6_n495), .ZN(MULT_mult_6_CARRYB_7__12_) );
  NOR2_X4 MULT_mult_6_U1755 ( .A1(MULT_mult_6_net82247), .A2(
        MULT_mult_6_net70458), .ZN(MULT_mult_6_ab_0__12_) );
  INV_X8 MULT_mult_6_U1754 ( .A(n10918), .ZN(MULT_mult_6_net70458) );
  INV_X4 MULT_mult_6_U1753 ( .A(MULT_mult_6_n491), .ZN(MULT_mult_6_net83784)
         );
  INV_X1 MULT_mult_6_U1752 ( .A(MULT_mult_6_ab_8__12_), .ZN(
        MULT_mult_6_net87308) );
  NOR2_X2 MULT_mult_6_U1751 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net77926), .ZN(MULT_mult_6_ab_8__12_) );
  NAND2_X2 MULT_mult_6_U1750 ( .A1(MULT_mult_6_ab_8__12_), .A2(
        MULT_mult_6_net90348), .ZN(MULT_mult_6_net80847) );
  NAND2_X2 MULT_mult_6_U1749 ( .A1(MULT_mult_6_SUMB_7__13_), .A2(
        MULT_mult_6_CARRYB_7__12_), .ZN(MULT_mult_6_net80848) );
  NAND2_X1 MULT_mult_6_U1748 ( .A1(MULT_mult_6_ab_8__12_), .A2(
        MULT_mult_6_CARRYB_7__12_), .ZN(MULT_mult_6_n493) );
  NAND3_X4 MULT_mult_6_U1747 ( .A1(MULT_mult_6_net80847), .A2(
        MULT_mult_6_net80848), .A3(MULT_mult_6_n493), .ZN(
        MULT_mult_6_CARRYB_8__12_) );
  INV_X16 MULT_mult_6_U1746 ( .A(n5761), .ZN(MULT_mult_6_net119855) );
  INV_X8 MULT_mult_6_U1745 ( .A(n5761), .ZN(MULT_mult_6_net77956) );
  INV_X1 MULT_mult_6_U1744 ( .A(MULT_mult_6_net81424), .ZN(
        MULT_mult_6_net123752) );
  NAND2_X1 MULT_mult_6_U1743 ( .A1(n5761), .A2(MULT_mult_6_net123752), .ZN(
        MULT_mult_6_net119928) );
  XNOR2_X2 MULT_mult_6_U1742 ( .A(MULT_mult_6_net119952), .B(
        MULT_mult_6__UDW__112684_net78549), .ZN(MULT_mult_6_net119949) );
  NAND2_X1 MULT_mult_6_U1741 ( .A1(MULT_mult_6__UDW__112684_net78549), .A2(
        MULT_mult_6_net119899), .ZN(MULT_mult_6_net119920) );
  AOI21_X4 MULT_mult_6_U1740 ( .B1(MULT_mult_6_net119899), .B2(
        MULT_mult_6__UDW__112684_net78549), .A(MULT_mult_6_net119901), .ZN(
        MULT_mult_6_net87363) );
  BUF_X8 MULT_mult_6_U1739 ( .A(MULT_mult_6_net89652), .Z(MULT_mult_6_net88344) );
  INV_X2 MULT_mult_6_U1737 ( .A(MULT_mult_6_n817), .ZN(MULT_mult_6_net148829)
         );
  NAND2_X4 MULT_mult_6_U1736 ( .A1(MULT_mult_6_net82295), .A2(
        MULT_mult_6_net82294), .ZN(MULT_mult_6_SUMB_13__9_) );
  INV_X16 MULT_mult_6_U1735 ( .A(aluA[17]), .ZN(MULT_mult_6_net70467) );
  INV_X1 MULT_mult_6_U1734 ( .A(MULT_mult_6_net86375), .ZN(
        MULT_mult_6_net120517) );
  NAND2_X1 MULT_mult_6_U1733 ( .A1(MULT_mult_6_net83755), .A2(
        MULT_mult_6_net86375), .ZN(MULT_mult_6_net120519) );
  NAND2_X4 MULT_mult_6_U1732 ( .A1(MULT_mult_6_net86375), .A2(
        MULT_mult_6_ab_15__7_), .ZN(MULT_mult_6_net80537) );
  NAND2_X4 MULT_mult_6_U1731 ( .A1(MULT_mult_6_n306), .A2(MULT_mult_6_n346), 
        .ZN(MULT_mult_6_net80538) );
  NAND2_X2 MULT_mult_6_U1730 ( .A1(MULT_mult_6_ab_15__7_), .A2(
        MULT_mult_6_CARRYB_14__7_), .ZN(MULT_mult_6_net80536) );
  NAND3_X4 MULT_mult_6_U1729 ( .A1(MULT_mult_6_net80537), .A2(
        MULT_mult_6_net80538), .A3(MULT_mult_6_net80536), .ZN(
        MULT_mult_6_CARRYB_15__7_) );
  INV_X8 MULT_mult_6_U1728 ( .A(n10923), .ZN(MULT_mult_6_net70448) );
  INV_X16 MULT_mult_6_U1727 ( .A(MULT_mult_6_net77916), .ZN(
        MULT_mult_6_net77912) );
  INV_X16 MULT_mult_6_U1726 ( .A(MULT_mult_6_net70448), .ZN(
        MULT_mult_6_net77916) );
  INV_X32 MULT_mult_6_U1725 ( .A(MULT_mult_6_net77916), .ZN(
        MULT_mult_6_net77914) );
  INV_X16 MULT_mult_6_U1724 ( .A(WIRE_ALU_A_MUX2TO1_32BIT_15__MUX_N1), .ZN(
        MULT_mult_6_net70463) );
  NAND2_X2 MULT_mult_6_U1723 ( .A1(MULT_mult_6_CARRYB_15__7_), .A2(
        MULT_mult_6_ab_16__7_), .ZN(MULT_mult_6_net80564) );
  NOR2_X2 MULT_mult_6_U1722 ( .A1(MULT_mult_6_net77914), .A2(
        MULT_mult_6_net70463), .ZN(MULT_mult_6_ab_16__7_) );
  INV_X2 MULT_mult_6_U1721 ( .A(MULT_mult_6_net119928), .ZN(
        MULT_mult_6_net123267) );
  NAND2_X2 MULT_mult_6_U1720 ( .A1(MULT_mult_6_net123266), .A2(
        MULT_mult_6_net123267), .ZN(MULT_mult_6_net123269) );
  INV_X4 MULT_mult_6_U1719 ( .A(MULT_mult_6_net119960), .ZN(
        MULT_mult_6_net119909) );
  BUF_X8 MULT_mult_6_U1718 ( .A(MULT_mult_6_CARRYB_2__15_), .Z(
        MULT_mult_6_net119974) );
  INV_X16 MULT_mult_6_U1717 ( .A(MULT_mult_6_net70444), .ZN(
        MULT_mult_6_net77904) );
  INV_X32 MULT_mult_6_U1716 ( .A(MULT_mult_6_net77904), .ZN(
        MULT_mult_6_net77900) );
  INV_X16 MULT_mult_6_U1715 ( .A(WIRE_ALU_A_MUX2TO1_32BIT_9__MUX_N1), .ZN(
        MULT_mult_6_net70451) );
  NOR2_X4 MULT_mult_6_U1714 ( .A1(MULT_mult_6_net77900), .A2(
        MULT_mult_6_net70451), .ZN(MULT_mult_6_ab_22__5_) );
  INV_X4 MULT_mult_6_U1713 ( .A(MULT_mult_6_net149530), .ZN(
        MULT_mult_6_net84666) );
  NAND2_X4 MULT_mult_6_U1712 ( .A1(MULT_mult_6_net84666), .A2(
        MULT_mult_6_net87681), .ZN(MULT_mult_6_net84668) );
  NAND2_X4 MULT_mult_6_U1711 ( .A1(MULT_mult_6_net83101), .A2(MULT_mult_6_n311), .ZN(MULT_mult_6_net84667) );
  NAND2_X4 MULT_mult_6_U1710 ( .A1(MULT_mult_6_net84668), .A2(
        MULT_mult_6_net84667), .ZN(MULT_mult_6_SUMB_21__6_) );
  NAND2_X1 MULT_mult_6_U1709 ( .A1(MULT_mult_6_ab_23__5_), .A2(
        MULT_mult_6_CARRYB_22__5_), .ZN(MULT_mult_6_net79904) );
  XNOR2_X2 MULT_mult_6_U1708 ( .A(MULT_mult_6_CARRYB_22__5_), .B(
        MULT_mult_6_ab_23__5_), .ZN(MULT_mult_6_net81983) );
  INV_X1 MULT_mult_6_U1707 ( .A(MULT_mult_6_CARRYB_22__5_), .ZN(
        MULT_mult_6_net88859) );
  INV_X4 MULT_mult_6_U1706 ( .A(MULT_mult_6_net88648), .ZN(
        MULT_mult_6_net124635) );
  NAND2_X4 MULT_mult_6_U1705 ( .A1(MULT_mult_6_n102), .A2(MULT_mult_6_net84213), .ZN(MULT_mult_6_net80290) );
  XNOR2_X2 MULT_mult_6_U1704 ( .A(MULT_mult_6_CARRYB_22__4_), .B(
        MULT_mult_6_ab_23__4_), .ZN(MULT_mult_6_net86109) );
  NAND2_X2 MULT_mult_6_U1703 ( .A1(MULT_mult_6_SUMB_23__4_), .A2(
        MULT_mult_6_ab_24__3_), .ZN(MULT_mult_6_net84679) );
  XNOR2_X2 MULT_mult_6_U1702 ( .A(MULT_mult_6_n102), .B(MULT_mult_6_net86109), 
        .ZN(MULT_mult_6_SUMB_23__4_) );
  NAND2_X2 MULT_mult_6_U1701 ( .A1(MULT_mult_6_n364), .A2(MULT_mult_6_net89455), .ZN(MULT_mult_6_net120366) );
  INV_X2 MULT_mult_6_U1700 ( .A(MULT_mult_6_SUMB_23__4_), .ZN(
        MULT_mult_6_net89455) );
  INV_X4 MULT_mult_6_U1699 ( .A(MULT_mult_6_net89455), .ZN(
        MULT_mult_6_net120364) );
  NAND2_X4 MULT_mult_6_U1698 ( .A1(MULT_mult_6_net120366), .A2(
        MULT_mult_6_n489), .ZN(MULT_mult_6_net92790) );
  NAND2_X4 MULT_mult_6_U1697 ( .A1(MULT_mult_6_net120364), .A2(
        MULT_mult_6_n285), .ZN(MULT_mult_6_n489) );
  INV_X1 MULT_mult_6_U1696 ( .A(MULT_mult_6_net82289), .ZN(
        MULT_mult_6_net85372) );
  INV_X8 MULT_mult_6_U1695 ( .A(MULT_mult_6_CARRYB_15__7_), .ZN(
        MULT_mult_6_net82289) );
  INV_X2 MULT_mult_6_U1694 ( .A(MULT_mult_6_ab_16__7_), .ZN(
        MULT_mult_6_net82288) );
  NAND2_X4 MULT_mult_6_U1693 ( .A1(MULT_mult_6_net82289), .A2(
        MULT_mult_6_net82288), .ZN(MULT_mult_6_n488) );
  NAND2_X4 MULT_mult_6_U1692 ( .A1(MULT_mult_6_net80564), .A2(MULT_mult_6_n488), .ZN(MULT_mult_6_net80906) );
  NAND2_X4 MULT_mult_6_U1691 ( .A1(MULT_mult_6_net93791), .A2(
        MULT_mult_6_net121814), .ZN(MULT_mult_6_n487) );
  NAND2_X2 MULT_mult_6_U1690 ( .A1(MULT_mult_6_n486), .A2(MULT_mult_6_n487), 
        .ZN(MULT_mult_6_SUMB_26__2_) );
  NAND3_X2 MULT_mult_6_U1689 ( .A1(MULT_mult_6_net83975), .A2(
        MULT_mult_6_net83977), .A3(MULT_mult_6_net83976), .ZN(
        MULT_mult_6_CARRYB_26__1_) );
  NAND2_X4 MULT_mult_6_U1688 ( .A1(MULT_mult_6_CARRYB_26__1_), .A2(
        MULT_mult_6_ab_27__1_), .ZN(MULT_mult_6_net80990) );
  NAND2_X4 MULT_mult_6_U1687 ( .A1(MULT_mult_6_net123365), .A2(
        MULT_mult_6_ab_27__1_), .ZN(MULT_mult_6_net80991) );
  NAND2_X4 MULT_mult_6_U1686 ( .A1(MULT_mult_6_n486), .A2(MULT_mult_6_n487), 
        .ZN(MULT_mult_6_net123365) );
  NAND3_X2 MULT_mult_6_U1685 ( .A1(MULT_mult_6_net83975), .A2(
        MULT_mult_6_net83977), .A3(MULT_mult_6_net83976), .ZN(
        MULT_mult_6_net89460) );
  XNOR2_X2 MULT_mult_6_U1684 ( .A(MULT_mult_6_net89460), .B(
        MULT_mult_6_net81867), .ZN(MULT_mult_6_net80986) );
  NAND2_X1 MULT_mult_6_U1683 ( .A1(MULT_mult_6_net80986), .A2(
        MULT_mult_6_net83623), .ZN(MULT_mult_6_net83624) );
  NAND2_X4 MULT_mult_6_U1682 ( .A1(MULT_mult_6_net83625), .A2(
        MULT_mult_6_net83624), .ZN(MULT_mult_6_SUMB_27__1_) );
  OR2_X2 MULT_mult_6_U1681 ( .A1(MULT_mult_6_net80986), .A2(
        MULT_mult_6_net83623), .ZN(MULT_mult_6_net83625) );
  XNOR2_X2 MULT_mult_6_U1680 ( .A(MULT_mult_6_CARRYB_20__5_), .B(
        MULT_mult_6_ab_21__5_), .ZN(MULT_mult_6_net83705) );
  NAND2_X2 MULT_mult_6_U1679 ( .A1(MULT_mult_6_SUMB_20__6_), .A2(
        MULT_mult_6_CARRYB_20__5_), .ZN(MULT_mult_6_net79991) );
  XNOR2_X2 MULT_mult_6_U1678 ( .A(MULT_mult_6_CARRYB_20__5_), .B(
        MULT_mult_6_ab_21__5_), .ZN(MULT_mult_6_net149133) );
  XNOR2_X2 MULT_mult_6_U1677 ( .A(MULT_mult_6_net149133), .B(MULT_mult_6_n71), 
        .ZN(MULT_mult_6_SUMB_21__5_) );
  INV_X4 MULT_mult_6_U1676 ( .A(MULT_mult_6_net80862), .ZN(
        MULT_mult_6_net147924) );
  INV_X4 MULT_mult_6_U1675 ( .A(MULT_mult_6_SUMB_21__5_), .ZN(
        MULT_mult_6_net147925) );
  NAND2_X4 MULT_mult_6_U1674 ( .A1(MULT_mult_6_n485), .A2(
        MULT_mult_6_net147926), .ZN(MULT_mult_6_SUMB_22__4_) );
  NAND2_X4 MULT_mult_6_U1673 ( .A1(MULT_mult_6_net147924), .A2(
        MULT_mult_6_net147925), .ZN(MULT_mult_6_n485) );
  INV_X4 MULT_mult_6_U1672 ( .A(MULT_mult_6_SUMB_14__8_), .ZN(
        MULT_mult_6_net86374) );
  INV_X2 MULT_mult_6_U1671 ( .A(MULT_mult_6_CARRYB_14__8_), .ZN(
        MULT_mult_6_net86536) );
  XNOR2_X2 MULT_mult_6_U1670 ( .A(MULT_mult_6_ab_15__8_), .B(
        MULT_mult_6_net86537), .ZN(MULT_mult_6_net93878) );
  NAND2_X2 MULT_mult_6_U1669 ( .A1(MULT_mult_6_ab_15__8_), .A2(
        MULT_mult_6_net86537), .ZN(MULT_mult_6_net80561) );
  INV_X4 MULT_mult_6_U1668 ( .A(MULT_mult_6_net86536), .ZN(
        MULT_mult_6_net86537) );
  XNOR2_X2 MULT_mult_6_U1667 ( .A(MULT_mult_6_ab_15__8_), .B(
        MULT_mult_6_net86537), .ZN(MULT_mult_6_net83273) );
  INV_X4 MULT_mult_6_U1666 ( .A(MULT_mult_6_ab_14__9_), .ZN(MULT_mult_6_n483)
         );
  XNOR2_X2 MULT_mult_6_U1665 ( .A(MULT_mult_6_n483), .B(MULT_mult_6_net85043), 
        .ZN(MULT_mult_6_n482) );
  XNOR2_X2 MULT_mult_6_U1664 ( .A(MULT_mult_6_n482), .B(MULT_mult_6_n210), 
        .ZN(MULT_mult_6_net88904) );
  NAND2_X4 MULT_mult_6_U1663 ( .A1(MULT_mult_6_net86537), .A2(
        MULT_mult_6_SUMB_14__9_), .ZN(MULT_mult_6_net80563) );
  NAND2_X4 MULT_mult_6_U1662 ( .A1(MULT_mult_6_SUMB_14__9_), .A2(
        MULT_mult_6_ab_15__8_), .ZN(MULT_mult_6_net80562) );
  INV_X8 MULT_mult_6_U1661 ( .A(MULT_mult_6_net88904), .ZN(
        MULT_mult_6_SUMB_14__9_) );
  NAND2_X4 MULT_mult_6_U1660 ( .A1(MULT_mult_6_net83273), .A2(
        MULT_mult_6_SUMB_14__9_), .ZN(MULT_mult_6_n484) );
  NAND2_X2 MULT_mult_6_U1659 ( .A1(MULT_mult_6_ab_16__7_), .A2(
        MULT_mult_6_SUMB_15__8_), .ZN(MULT_mult_6_net80565) );
  NAND2_X2 MULT_mult_6_U1658 ( .A1(MULT_mult_6_net80906), .A2(MULT_mult_6_n104), .ZN(MULT_mult_6_net81668) );
  NAND2_X2 MULT_mult_6_U1657 ( .A1(MULT_mult_6_SUMB_15__8_), .A2(
        MULT_mult_6_net85372), .ZN(MULT_mult_6_net80566) );
  NAND2_X4 MULT_mult_6_U1656 ( .A1(MULT_mult_6_net85543), .A2(MULT_mult_6_n484), .ZN(MULT_mult_6_SUMB_15__8_) );
  INV_X4 MULT_mult_6_U1655 ( .A(MULT_mult_6_net80906), .ZN(
        MULT_mult_6_net81666) );
  INV_X4 MULT_mult_6_U1654 ( .A(MULT_mult_6_n104), .ZN(MULT_mult_6_net81667)
         );
  NAND2_X4 MULT_mult_6_U1653 ( .A1(MULT_mult_6_n481), .A2(MULT_mult_6_net81668), .ZN(MULT_mult_6_SUMB_16__7_) );
  NAND2_X4 MULT_mult_6_U1652 ( .A1(MULT_mult_6_net81666), .A2(
        MULT_mult_6_net81667), .ZN(MULT_mult_6_n481) );
  NAND2_X2 MULT_mult_6_U1651 ( .A1(MULT_mult_6_n353), .A2(
        MULT_mult_6_net119949), .ZN(MULT_mult_6_net119960) );
  XNOR2_X2 MULT_mult_6_U1650 ( .A(MULT_mult_6_CARRYB_2__15_), .B(
        MULT_mult_6_n353), .ZN(MULT_mult_6_net121859) );
  NOR2_X2 MULT_mult_6_U1649 ( .A1(MULT_mult_6_net119949), .A2(MULT_mult_6_n353), .ZN(MULT_mult_6_net119948) );
  OAI21_X4 MULT_mult_6_U1648 ( .B1(MULT_mult_6_net119908), .B2(
        MULT_mult_6_net123267), .A(MULT_mult_6_net123266), .ZN(
        MULT_mult_6_net124908) );
  OAI21_X4 MULT_mult_6_U1647 ( .B1(MULT_mult_6_net119909), .B2(
        MULT_mult_6_net119910), .A(MULT_mult_6_n477), .ZN(
        MULT_mult_6_net119908) );
  INV_X1 MULT_mult_6_U1646 ( .A(MULT_mult_6_ab_5__14_), .ZN(
        MULT_mult_6_net84946) );
  NOR2_X4 MULT_mult_6_U1645 ( .A1(MULT_mult_6_net84698), .A2(
        MULT_mult_6_net77948), .ZN(MULT_mult_6_ab_5__14_) );
  INV_X4 MULT_mult_6_U1644 ( .A(MULT_mult_6_net119927), .ZN(
        MULT_mult_6_net148837) );
  NAND2_X4 MULT_mult_6_U1643 ( .A1(MULT_mult_6_net148836), .A2(
        MULT_mult_6_net148837), .ZN(MULT_mult_6_n478) );
  NAND2_X4 MULT_mult_6_U1642 ( .A1(MULT_mult_6_n478), .A2(
        MULT_mult_6_net148838), .ZN(MULT_mult_6_net83918) );
  INV_X8 MULT_mult_6_U1641 ( .A(MULT_mult_6_net83918), .ZN(
        MULT_mult_6_net83919) );
  NAND3_X2 MULT_mult_6_U1640 ( .A1(MULT_mult_6_net82297), .A2(MULT_mult_6_n479), .A3(MULT_mult_6_n480), .ZN(MULT_mult_6_CARRYB_5__14_) );
  NAND2_X4 MULT_mult_6_U1639 ( .A1(MULT_mult_6_net87411), .A2(MULT_mult_6_n344), .ZN(MULT_mult_6_net79884) );
  INV_X32 MULT_mult_6_U1638 ( .A(net78051), .ZN(MULT_mult_6_net77868) );
  INV_X4 MULT_mult_6_U1637 ( .A(MULT_mult_6_net77866), .ZN(
        MULT_mult_6_net92331) );
  NAND2_X4 MULT_mult_6_U1636 ( .A1(MULT_mult_6_net89110), .A2(
        MULT_mult_6_ab_28__1_), .ZN(MULT_mult_6_net79881) );
  XNOR2_X2 MULT_mult_6_U1635 ( .A(MULT_mult_6_CARRYB_27__1_), .B(
        MULT_mult_6_ab_28__1_), .ZN(MULT_mult_6_net149605) );
  INV_X4 MULT_mult_6_U1634 ( .A(MULT_mult_6_net92330), .ZN(
        MULT_mult_6_ab_28__1_) );
  XNOR2_X2 MULT_mult_6_U1633 ( .A(MULT_mult_6_CARRYB_27__1_), .B(
        MULT_mult_6_net92330), .ZN(MULT_mult_6_n476) );
  NAND2_X4 MULT_mult_6_U1632 ( .A1(MULT_mult_6_CARRYB_28__0_), .A2(
        MULT_mult_6_net86792), .ZN(MULT_mult_6_net79885) );
  XNOR2_X2 MULT_mult_6_U1631 ( .A(MULT_mult_6_net87798), .B(
        MULT_mult_6_ab_30__0_), .ZN(MULT_mult_6_net83536) );
  NAND3_X4 MULT_mult_6_U1630 ( .A1(MULT_mult_6_net79885), .A2(
        MULT_mult_6_net79884), .A3(MULT_mult_6_net79883), .ZN(
        MULT_mult_6_net87798) );
  NOR2_X4 MULT_mult_6_U1628 ( .A1(MULT_mult_6_net87396), .A2(
        MULT_mult_6_net80409), .ZN(MULT_mult_6_ab_1__15_) );
  INV_X4 MULT_mult_6_U1627 ( .A(n10931), .ZN(MULT_mult_6_net77926) );
  NAND2_X2 MULT_mult_6_U1626 ( .A1(MULT_mult_6_net123072), .A2(n10931), .ZN(
        MULT_mult_6_net123019) );
  NOR2_X2 MULT_mult_6_U1625 ( .A1(MULT_mult_6_net91660), .A2(
        MULT_mult_6_net77924), .ZN(MULT_mult_6_ab_8__10_) );
  NAND2_X4 MULT_mult_6_U1624 ( .A1(MULT_mult_6_net119982), .A2(
        MULT_mult_6_net88297), .ZN(MULT_mult_6_net89168) );
  NAND2_X1 MULT_mult_6_U1623 ( .A1(MULT_mult_6_net122062), .A2(
        MULT_mult_6_net89168), .ZN(MULT_mult_6_net123143) );
  XNOR2_X2 MULT_mult_6_U1622 ( .A(MULT_mult_6_CARRYB_6__10_), .B(
        MULT_mult_6_ab_7__10_), .ZN(MULT_mult_6_net81586) );
  NAND2_X2 MULT_mult_6_U1621 ( .A1(MULT_mult_6_SUMB_6__11_), .A2(
        MULT_mult_6_ab_7__10_), .ZN(MULT_mult_6_n474) );
  NAND2_X1 MULT_mult_6_U1620 ( .A1(MULT_mult_6_ab_7__10_), .A2(
        MULT_mult_6_CARRYB_6__10_), .ZN(MULT_mult_6_n475) );
  NAND3_X2 MULT_mult_6_U1619 ( .A1(MULT_mult_6_n473), .A2(MULT_mult_6_n474), 
        .A3(MULT_mult_6_n475), .ZN(MULT_mult_6_CARRYB_7__10_) );
  INV_X32 MULT_mult_6_U1618 ( .A(n6007), .ZN(MULT_mult_6_net77966) );
  INV_X16 MULT_mult_6_U1617 ( .A(n6007), .ZN(MULT_mult_6_net77964) );
  NAND2_X4 MULT_mult_6_U1616 ( .A1(MULT_mult_6_ab_3__13_), .A2(
        MULT_mult_6_SUMB_2__14_), .ZN(MULT_mult_6_net81514) );
  NOR2_X2 MULT_mult_6_U1615 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net77964), .ZN(MULT_mult_6_ab_3__13_) );
  NOR2_X4 MULT_mult_6_U1614 ( .A1(MULT_mult_6_net87396), .A2(
        MULT_mult_6_net82149), .ZN(MULT_mult_6_ab_0__15_) );
  AND2_X2 MULT_mult_6_U1613 ( .A1(n10924), .A2(MULT_mult_6_n341), .ZN(
        MULT_mult_6_ab_1__6_) );
  INV_X1 MULT_mult_6_U1612 ( .A(MULT_mult_6_ab_11__8_), .ZN(
        MULT_mult_6_net120464) );
  NAND2_X4 MULT_mult_6_U1611 ( .A1(MULT_mult_6_net147936), .A2(
        MULT_mult_6_ab_11__8_), .ZN(MULT_mult_6_net84656) );
  NAND2_X4 MULT_mult_6_U1610 ( .A1(MULT_mult_6_net120466), .A2(
        MULT_mult_6_net84656), .ZN(MULT_mult_6_net86844) );
  NAND2_X4 MULT_mult_6_U1609 ( .A1(MULT_mult_6_CARRYB_10__8_), .A2(
        MULT_mult_6_SUMB_10__9_), .ZN(MULT_mult_6_net84654) );
  INV_X4 MULT_mult_6_U1608 ( .A(MULT_mult_6_net91419), .ZN(
        MULT_mult_6_net120514) );
  INV_X16 MULT_mult_6_U1607 ( .A(n10921), .ZN(MULT_mult_6_net70452) );
  NAND3_X4 MULT_mult_6_U1606 ( .A1(MULT_mult_6_net84267), .A2(
        MULT_mult_6_net84268), .A3(MULT_mult_6_net93306), .ZN(
        MULT_mult_6_CARRYB_11__9_) );
  NAND3_X2 MULT_mult_6_U1605 ( .A1(MULT_mult_6_n471), .A2(MULT_mult_6_n325), 
        .A3(MULT_mult_6_n472), .ZN(MULT_mult_6_CARRYB_10__9_) );
  NAND2_X4 MULT_mult_6_U1604 ( .A1(MULT_mult_6_net93304), .A2(
        MULT_mult_6_net93305), .ZN(MULT_mult_6_net93307) );
  NAND2_X4 MULT_mult_6_U1603 ( .A1(MULT_mult_6_net93306), .A2(
        MULT_mult_6_net93307), .ZN(MULT_mult_6_net90735) );
  NAND2_X2 MULT_mult_6_U1602 ( .A1(MULT_mult_6_net91118), .A2(
        MULT_mult_6_ab_9__11_), .ZN(MULT_mult_6_net81258) );
  XNOR2_X2 MULT_mult_6_U1601 ( .A(MULT_mult_6_net91118), .B(
        MULT_mult_6_net83042), .ZN(MULT_mult_6_SUMB_9__11_) );
  NAND2_X4 MULT_mult_6_U1600 ( .A1(MULT_mult_6_net84069), .A2(MULT_mult_6_n70), 
        .ZN(MULT_mult_6_net84072) );
  NAND2_X4 MULT_mult_6_U1599 ( .A1(MULT_mult_6_SUMB_10__10_), .A2(
        MULT_mult_6_ab_11__9_), .ZN(MULT_mult_6_net93306) );
  INV_X4 MULT_mult_6_U1598 ( .A(MULT_mult_6_SUMB_10__10_), .ZN(
        MULT_mult_6_net93304) );
  NAND2_X4 MULT_mult_6_U1597 ( .A1(MULT_mult_6_net86895), .A2(
        MULT_mult_6_net86896), .ZN(MULT_mult_6_net83042) );
  NAND2_X2 MULT_mult_6_U1596 ( .A1(MULT_mult_6_net90687), .A2(MULT_mult_6_n229), .ZN(MULT_mult_6_net81259) );
  NAND2_X2 MULT_mult_6_U1595 ( .A1(MULT_mult_6_net86896), .A2(
        MULT_mult_6_net86895), .ZN(MULT_mult_6_n470) );
  XNOR2_X2 MULT_mult_6_U1594 ( .A(MULT_mult_6_n470), .B(MULT_mult_6_net90687), 
        .ZN(MULT_mult_6_net91259) );
  INV_X1 MULT_mult_6_U1593 ( .A(MULT_mult_6_net91259), .ZN(
        MULT_mult_6_net84070) );
  NAND2_X4 MULT_mult_6_U1592 ( .A1(MULT_mult_6_net84072), .A2(
        MULT_mult_6_net84071), .ZN(MULT_mult_6_SUMB_10__10_) );
  INV_X8 MULT_mult_6_U1591 ( .A(net36463), .ZN(MULT_mult_6_net84698) );
  NAND2_X4 MULT_mult_6_U1590 ( .A1(n10916), .A2(MULT_mult_6_net77984), .ZN(
        MULT_mult_6_net87050) );
  INV_X16 MULT_mult_6_U1589 ( .A(MULT_mult_6_net70493), .ZN(
        MULT_mult_6_net77984) );
  INV_X16 MULT_mult_6_U1588 ( .A(MULT_mult_6_net77984), .ZN(
        MULT_mult_6_net86101) );
  NAND2_X4 MULT_mult_6_U1587 ( .A1(MULT_mult_6_net87465), .A2(
        MULT_mult_6_net87464), .ZN(MULT_mult_6_n469) );
  NAND2_X4 MULT_mult_6_U1586 ( .A1(MULT_mult_6_n469), .A2(MULT_mult_6_net81204), .ZN(MULT_mult_6_net86151) );
  INV_X32 MULT_mult_6_U1585 ( .A(n10930), .ZN(MULT_mult_6_net77938) );
  NOR2_X1 MULT_mult_6_U1584 ( .A1(MULT_mult_6_net70456), .A2(
        MULT_mult_6_net77938), .ZN(MULT_mult_6_ab_6__11_) );
  NAND2_X2 MULT_mult_6_U1583 ( .A1(MULT_mult_6_net91419), .A2(
        MULT_mult_6_net82723), .ZN(MULT_mult_6_net120515) );
  XNOR2_X2 MULT_mult_6_U1582 ( .A(MULT_mult_6_net82723), .B(
        MULT_mult_6_net91419), .ZN(MULT_mult_6_n468) );
  NAND2_X4 MULT_mult_6_U1581 ( .A1(MULT_mult_6_n468), .A2(
        MULT_mult_6_ab_11__8_), .ZN(MULT_mult_6_n467) );
  NAND3_X4 MULT_mult_6_U1580 ( .A1(MULT_mult_6_net84654), .A2(MULT_mult_6_n467), .A3(MULT_mult_6_net84656), .ZN(MULT_mult_6_CARRYB_11__8_) );
  INV_X16 MULT_mult_6_U1579 ( .A(aluA[19]), .ZN(MULT_mult_6_net70471) );
  NOR2_X2 MULT_mult_6_U1578 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__8_) );
  NAND2_X2 MULT_mult_6_U1577 ( .A1(MULT_mult_6_net123072), .A2(n10932), .ZN(
        MULT_mult_6_net123055) );
  NAND3_X2 MULT_mult_6_U1576 ( .A1(MULT_mult_6_net81216), .A2(MULT_mult_6_n461), .A3(MULT_mult_6_net81215), .ZN(MULT_mult_6_CARRYB_8__10_) );
  INV_X4 MULT_mult_6_U1575 ( .A(MULT_mult_6_net80993), .ZN(MULT_mult_6_n462)
         );
  NAND2_X2 MULT_mult_6_U1574 ( .A1(MULT_mult_6_n463), .A2(MULT_mult_6_net80993), .ZN(MULT_mult_6_n464) );
  INV_X2 MULT_mult_6_U1573 ( .A(MULT_mult_6_SUMB_7__12_), .ZN(MULT_mult_6_n463) );
  INV_X2 MULT_mult_6_U1572 ( .A(MULT_mult_6_n463), .ZN(MULT_mult_6_n460) );
  NAND2_X4 MULT_mult_6_U1571 ( .A1(MULT_mult_6_n462), .A2(MULT_mult_6_n460), 
        .ZN(MULT_mult_6_n465) );
  NAND2_X4 MULT_mult_6_U1570 ( .A1(MULT_mult_6_n464), .A2(MULT_mult_6_n465), 
        .ZN(MULT_mult_6_SUMB_8__11_) );
  INV_X4 MULT_mult_6_U1569 ( .A(n10932), .ZN(MULT_mult_6_net70477) );
  NAND2_X2 MULT_mult_6_U1568 ( .A1(MULT_mult_6_SUMB_10__10_), .A2(
        MULT_mult_6_CARRYB_10__9_), .ZN(MULT_mult_6_net84267) );
  NAND2_X2 MULT_mult_6_U1567 ( .A1(MULT_mult_6_CARRYB_10__9_), .A2(
        MULT_mult_6_ab_11__9_), .ZN(MULT_mult_6_net84268) );
  XNOR2_X2 MULT_mult_6_U1566 ( .A(MULT_mult_6_CARRYB_11__8_), .B(
        MULT_mult_6_ab_12__8_), .ZN(MULT_mult_6_net82548) );
  INV_X1 MULT_mult_6_U1565 ( .A(MULT_mult_6_net89537), .ZN(
        MULT_mult_6_net93309) );
  NOR2_X2 MULT_mult_6_U1564 ( .A1(MULT_mult_6_net124610), .A2(
        MULT_mult_6_net70450), .ZN(MULT_mult_6_ab_0__8_) );
  INV_X8 MULT_mult_6_U1563 ( .A(n10922), .ZN(MULT_mult_6_net70450) );
  INV_X4 MULT_mult_6_U1562 ( .A(MULT_mult_6_net70450), .ZN(
        MULT_mult_6_net77922) );
  INV_X32 MULT_mult_6_U1561 ( .A(MULT_mult_6_net77922), .ZN(
        MULT_mult_6_net77920) );
  INV_X16 MULT_mult_6_U1560 ( .A(aluA[18]), .ZN(MULT_mult_6_net70469) );
  XNOR2_X1 MULT_mult_6_U1559 ( .A(MULT_mult_6_n183), .B(MULT_mult_6_net88104), 
        .ZN(MULT_mult_6_net149580) );
  NAND2_X1 MULT_mult_6_U1558 ( .A1(MULT_mult_6_net90735), .A2(
        MULT_mult_6_net88104), .ZN(MULT_mult_6_net121447) );
  INV_X2 MULT_mult_6_U1557 ( .A(MULT_mult_6_net88104), .ZN(
        MULT_mult_6_net121446) );
  BUF_X4 MULT_mult_6_U1556 ( .A(MULT_mult_6_CARRYB_10__9_), .Z(
        MULT_mult_6_net88104) );
  XNOR2_X2 MULT_mult_6_U1555 ( .A(MULT_mult_6_net90735), .B(
        MULT_mult_6_net88104), .ZN(MULT_mult_6_SUMB_11__9_) );
  NAND2_X2 MULT_mult_6_U1554 ( .A1(MULT_mult_6_SUMB_11__9_), .A2(
        MULT_mult_6_CARRYB_11__8_), .ZN(MULT_mult_6_net81115) );
  NAND2_X2 MULT_mult_6_U1553 ( .A1(MULT_mult_6_ab_12__8_), .A2(
        MULT_mult_6_CARRYB_11__8_), .ZN(MULT_mult_6_n459) );
  NAND2_X4 MULT_mult_6_U1552 ( .A1(MULT_mult_6_net89537), .A2(
        MULT_mult_6_ab_12__8_), .ZN(MULT_mult_6_net81116) );
  NAND2_X2 MULT_mult_6_U1551 ( .A1(MULT_mult_6_SUMB_12__9_), .A2(
        MULT_mult_6_CARRYB_12__8_), .ZN(MULT_mult_6_net80505) );
  INV_X4 MULT_mult_6_U1550 ( .A(MULT_mult_6_CARRYB_12__8_), .ZN(
        MULT_mult_6_net84710) );
  NAND2_X2 MULT_mult_6_U1549 ( .A1(MULT_mult_6_net80694), .A2(
        MULT_mult_6_CARRYB_12__8_), .ZN(MULT_mult_6_net84712) );
  NAND3_X4 MULT_mult_6_U1548 ( .A1(MULT_mult_6_net81115), .A2(MULT_mult_6_n459), .A3(MULT_mult_6_net81116), .ZN(MULT_mult_6_CARRYB_12__8_) );
  NAND3_X2 MULT_mult_6_U1547 ( .A1(MULT_mult_6_net80506), .A2(
        MULT_mult_6_net80505), .A3(MULT_mult_6_net80507), .ZN(
        MULT_mult_6_CARRYB_13__8_) );
  NAND2_X2 MULT_mult_6_U1546 ( .A1(MULT_mult_6_CARRYB_12__8_), .A2(
        MULT_mult_6_ab_13__8_), .ZN(MULT_mult_6_net80507) );
  NAND2_X2 MULT_mult_6_U1545 ( .A1(MULT_mult_6_net81630), .A2(n10920), .ZN(
        MULT_mult_6_net90174) );
  NAND3_X4 MULT_mult_6_U1544 ( .A1(n10933), .A2(n6005), .A3(
        MULT_mult_6_net147421), .ZN(MULT_mult_6_net147451) );
  INV_X1 MULT_mult_6_U1543 ( .A(MULT_mult_6_ab_9__10_), .ZN(
        MULT_mult_6_net87456) );
  NAND2_X2 MULT_mult_6_U1542 ( .A1(MULT_mult_6_CARRYB_8__10_), .A2(
        MULT_mult_6_ab_9__10_), .ZN(MULT_mult_6_net87458) );
  NAND2_X4 MULT_mult_6_U1541 ( .A1(MULT_mult_6_net87458), .A2(
        MULT_mult_6_net87459), .ZN(MULT_mult_6_net83736) );
  INV_X8 MULT_mult_6_U1540 ( .A(n10920), .ZN(MULT_mult_6_net70454) );
  INV_X4 MULT_mult_6_U1539 ( .A(n10933), .ZN(MULT_mult_6_net70475) );
  NAND2_X4 MULT_mult_6_U1538 ( .A1(MULT_mult_6_net91259), .A2(
        MULT_mult_6_ab_10__10_), .ZN(MULT_mult_6_net81261) );
  INV_X4 MULT_mult_6_U1537 ( .A(MULT_mult_6_n2378), .ZN(MULT_mult_6_net87457)
         );
  INV_X4 MULT_mult_6_U1536 ( .A(MULT_mult_6_net87457), .ZN(
        MULT_mult_6_net91298) );
  NAND2_X4 MULT_mult_6_U1535 ( .A1(MULT_mult_6_net91298), .A2(
        MULT_mult_6_SUMB_8__11_), .ZN(MULT_mult_6_net81001) );
  NAND2_X4 MULT_mult_6_U1534 ( .A1(MULT_mult_6_SUMB_8__11_), .A2(
        MULT_mult_6_ab_9__10_), .ZN(MULT_mult_6_n457) );
  NAND2_X2 MULT_mult_6_U1533 ( .A1(MULT_mult_6_SUMB_9__11_), .A2(
        MULT_mult_6_CARRYB_9__10_), .ZN(MULT_mult_6_net81262) );
  NAND2_X2 MULT_mult_6_U1532 ( .A1(MULT_mult_6_CARRYB_9__10_), .A2(
        MULT_mult_6_ab_10__10_), .ZN(MULT_mult_6_net81260) );
  NAND3_X4 MULT_mult_6_U1531 ( .A1(MULT_mult_6_net81001), .A2(MULT_mult_6_n457), .A3(MULT_mult_6_net87458), .ZN(MULT_mult_6_CARRYB_9__10_) );
  INV_X4 MULT_mult_6_U1530 ( .A(MULT_mult_6_CARRYB_9__10_), .ZN(
        MULT_mult_6_net83061) );
  NAND2_X2 MULT_mult_6_U1529 ( .A1(MULT_mult_6_CARRYB_9__10_), .A2(
        MULT_mult_6_net81643), .ZN(MULT_mult_6_net83062) );
  INV_X4 MULT_mult_6_U1528 ( .A(MULT_mult_6_net81256), .ZN(
        MULT_mult_6_net84069) );
  NAND2_X4 MULT_mult_6_U1526 ( .A1(MULT_mult_6_n458), .A2(MULT_mult_6_net83062), .ZN(MULT_mult_6_net81256) );
  NOR2_X4 MULT_mult_6_U1525 ( .A1(MULT_mult_6_net70462), .A2(
        MULT_mult_6_net86101), .ZN(MULT_mult_6_ab_1__14_) );
  INV_X8 MULT_mult_6_U1524 ( .A(net36463), .ZN(MULT_mult_6_net70462) );
  XNOR2_X2 MULT_mult_6_U1523 ( .A(MULT_mult_6_ab_0__14_), .B(
        MULT_mult_6_ab_1__13_), .ZN(MULT_mult_6__UDW__112704_net78605) );
  INV_X4 MULT_mult_6_U1522 ( .A(MULT_mult_6_net120391), .ZN(
        MULT_mult_6_net120392) );
  INV_X16 MULT_mult_6_U1521 ( .A(MULT_mult_6_net120392), .ZN(
        MULT_mult_6_net70460) );
  INV_X16 MULT_mult_6_U1520 ( .A(aluA[29]), .ZN(MULT_mult_6_net70491) );
  NOR2_X4 MULT_mult_6_U1519 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net70491), .ZN(MULT_mult_6_ab_2__13_) );
  NOR2_X4 MULT_mult_6_U1518 ( .A1(MULT_mult_6_net80727), .A2(MULT_mult_6_n175), 
        .ZN(MULT_mult_6_ab_2__20_) );
  XNOR2_X2 MULT_mult_6_U1517 ( .A(MULT_mult_6_ab_1__14_), .B(
        MULT_mult_6_ab_0__15_), .ZN(MULT_mult_6__UDW__112699_net78591) );
  XNOR2_X2 MULT_mult_6_U1516 ( .A(MULT_mult_6_n456), .B(
        MULT_mult_6_SUMB_1__14_), .ZN(MULT_mult_6_SUMB_2__13_) );
  INV_X8 MULT_mult_6_U1515 ( .A(MULT_mult_6__UDW__112699_net78591), .ZN(
        MULT_mult_6_SUMB_1__14_) );
  NAND2_X2 MULT_mult_6_U1514 ( .A1(MULT_mult_6_ab_0__14_), .A2(
        MULT_mult_6_ab_1__13_), .ZN(MULT_mult_6_n452) );
  XNOR2_X2 MULT_mult_6_U1513 ( .A(MULT_mult_6_CARRYB_1__13_), .B(
        MULT_mult_6_ab_2__13_), .ZN(MULT_mult_6_n456) );
  NAND2_X2 MULT_mult_6_U1512 ( .A1(MULT_mult_6_net124833), .A2(
        MULT_mult_6_CARRYB_1__13_), .ZN(MULT_mult_6_n455) );
  NAND2_X2 MULT_mult_6_U1511 ( .A1(MULT_mult_6_n99), .A2(MULT_mult_6_ab_3__13_), .ZN(MULT_mult_6_net81515) );
  NAND3_X4 MULT_mult_6_U1510 ( .A1(MULT_mult_6_n454), .A2(MULT_mult_6_n453), 
        .A3(MULT_mult_6_n455), .ZN(MULT_mult_6_CARRYB_2__13_) );
  NAND2_X4 MULT_mult_6_U1509 ( .A1(MULT_mult_6_SUMB_3__12_), .A2(
        MULT_mult_6_ab_4__11_), .ZN(MULT_mult_6_net88085) );
  NAND2_X2 MULT_mult_6_U1508 ( .A1(MULT_mult_6_SUMB_3__12_), .A2(
        MULT_mult_6_CARRYB_3__11_), .ZN(MULT_mult_6_net88084) );
  INV_X2 MULT_mult_6_U1507 ( .A(MULT_mult_6_SUMB_4__12_), .ZN(
        MULT_mult_6_net123898) );
  NAND2_X1 MULT_mult_6_U1506 ( .A1(MULT_mult_6_net82757), .A2(
        MULT_mult_6_SUMB_4__12_), .ZN(MULT_mult_6_net123899) );
  INV_X8 MULT_mult_6_U1505 ( .A(aluA[26]), .ZN(MULT_mult_6_n449) );
  NOR2_X4 MULT_mult_6_U1504 ( .A1(MULT_mult_6_net70456), .A2(
        MULT_mult_6_net77946), .ZN(MULT_mult_6_ab_5__11_) );
  NAND2_X1 MULT_mult_6_U1503 ( .A1(MULT_mult_6_CARRYB_4__11_), .A2(
        MULT_mult_6_net83351), .ZN(MULT_mult_6_net147922) );
  NAND3_X2 MULT_mult_6_U1502 ( .A1(MULT_mult_6_net88084), .A2(
        MULT_mult_6_net88085), .A3(MULT_mult_6_net88086), .ZN(
        MULT_mult_6_CARRYB_4__11_) );
  NAND3_X1 MULT_mult_6_U1501 ( .A1(MULT_mult_6_net88084), .A2(
        MULT_mult_6_net88085), .A3(MULT_mult_6_net88086), .ZN(
        MULT_mult_6_net124527) );
  NAND2_X4 MULT_mult_6_U1500 ( .A1(MULT_mult_6_SUMB_4__12_), .A2(
        MULT_mult_6_net124527), .ZN(MULT_mult_6_net82762) );
  NAND2_X4 MULT_mult_6_U1499 ( .A1(MULT_mult_6_SUMB_4__12_), .A2(
        MULT_mult_6_ab_5__11_), .ZN(MULT_mult_6_net82763) );
  NAND2_X1 MULT_mult_6_U1498 ( .A1(MULT_mult_6_ab_5__11_), .A2(
        MULT_mult_6_CARRYB_4__11_), .ZN(MULT_mult_6_n451) );
  NAND3_X4 MULT_mult_6_U1497 ( .A1(MULT_mult_6_net82762), .A2(
        MULT_mult_6_net82763), .A3(MULT_mult_6_n451), .ZN(
        MULT_mult_6_CARRYB_5__11_) );
  NAND2_X2 MULT_mult_6_U1496 ( .A1(MULT_mult_6_ab_5__12_), .A2(
        MULT_mult_6_SUMB_4__13_), .ZN(MULT_mult_6_net81205) );
  NAND2_X2 MULT_mult_6_U1495 ( .A1(MULT_mult_6_SUMB_4__13_), .A2(
        MULT_mult_6_CARRYB_4__12_), .ZN(MULT_mult_6_net81206) );
  INV_X2 MULT_mult_6_U1494 ( .A(MULT_mult_6_net86151), .ZN(
        MULT_mult_6_net121453) );
  INV_X2 MULT_mult_6_U1493 ( .A(MULT_mult_6_n448), .ZN(MULT_mult_6_net121454)
         );
  NAND2_X2 MULT_mult_6_U1492 ( .A1(MULT_mult_6_net86151), .A2(MULT_mult_6_n448), .ZN(MULT_mult_6_net121455) );
  XNOR2_X2 MULT_mult_6_U1491 ( .A(MULT_mult_6_net86151), .B(MULT_mult_6_n448), 
        .ZN(MULT_mult_6_SUMB_5__12_) );
  NAND2_X4 MULT_mult_6_U1490 ( .A1(MULT_mult_6_SUMB_5__12_), .A2(
        MULT_mult_6_ab_6__11_), .ZN(MULT_mult_6_n446) );
  NAND2_X4 MULT_mult_6_U1489 ( .A1(MULT_mult_6_net90731), .A2(
        MULT_mult_6_net84652), .ZN(MULT_mult_6_n445) );
  INV_X4 MULT_mult_6_U1488 ( .A(MULT_mult_6_n146), .ZN(MULT_mult_6_net84652)
         );
  NAND2_X4 MULT_mult_6_U1487 ( .A1(MULT_mult_6_net84652), .A2(
        MULT_mult_6_ab_6__11_), .ZN(MULT_mult_6_n447) );
  NAND3_X4 MULT_mult_6_U1486 ( .A1(MULT_mult_6_n445), .A2(MULT_mult_6_n447), 
        .A3(MULT_mult_6_n446), .ZN(MULT_mult_6_CARRYB_6__11_) );
  INV_X16 MULT_mult_6_U1485 ( .A(n10919), .ZN(MULT_mult_6_net70456) );
  INV_X4 MULT_mult_6_U1484 ( .A(net36391), .ZN(MULT_mult_6_n443) );
  NOR2_X1 MULT_mult_6_U1483 ( .A1(MULT_mult_6_net70456), .A2(
        MULT_mult_6_net77930), .ZN(MULT_mult_6_ab_7__11_) );
  INV_X8 MULT_mult_6_U1482 ( .A(aluA[31]), .ZN(MULT_mult_6_net77988) );
  XNOR2_X2 MULT_mult_6_U1481 ( .A(MULT_mult_6_CARRYB_2__13_), .B(
        MULT_mult_6_ab_3__13_), .ZN(MULT_mult_6_net81694) );
  XNOR2_X2 MULT_mult_6_U1480 ( .A(MULT_mult_6_ab_2__14_), .B(
        MULT_mult_6_CARRYB_1__14_), .ZN(MULT_mult_6_net86864) );
  XNOR2_X1 MULT_mult_6_U1479 ( .A(MULT_mult_6_CARRYB_1__14_), .B(
        MULT_mult_6_ab_2__14_), .ZN(MULT_mult_6_n438) );
  NOR2_X4 MULT_mult_6_U1478 ( .A1(MULT_mult_6_net70466), .A2(
        MULT_mult_6_net80409), .ZN(MULT_mult_6_net88123) );
  INV_X16 MULT_mult_6_U1477 ( .A(aluA[31]), .ZN(MULT_mult_6_net82149) );
  NOR2_X4 MULT_mult_6_U1476 ( .A1(MULT_mult_6_net70466), .A2(
        MULT_mult_6_net82149), .ZN(MULT_mult_6_ab_0__16_) );
  NAND2_X2 MULT_mult_6_U1475 ( .A1(MULT_mult_6_SUMB_1__15_), .A2(
        MULT_mult_6_ab_2__14_), .ZN(MULT_mult_6_net86170) );
  CLKBUF_X3 MULT_mult_6_U1474 ( .A(MULT_mult_6_SUMB_1__15_), .Z(
        MULT_mult_6_n440) );
  XNOR2_X2 MULT_mult_6_U1473 ( .A(MULT_mult_6_n438), .B(MULT_mult_6_n440), 
        .ZN(MULT_mult_6_net84270) );
  NAND2_X1 MULT_mult_6_U1472 ( .A1(MULT_mult_6_SUMB_3__13_), .A2(
        MULT_mult_6_n89), .ZN(MULT_mult_6_net82760) );
  INV_X4 MULT_mult_6_U1471 ( .A(MULT_mult_6_net89227), .ZN(MULT_mult_6_n439)
         );
  NAND2_X2 MULT_mult_6_U1470 ( .A1(MULT_mult_6_net89227), .A2(
        MULT_mult_6_net85493), .ZN(MULT_mult_6_n441) );
  INV_X4 MULT_mult_6_U1469 ( .A(MULT_mult_6_net85493), .ZN(
        MULT_mult_6_net88010) );
  NAND2_X4 MULT_mult_6_U1468 ( .A1(MULT_mult_6_n441), .A2(MULT_mult_6_n442), 
        .ZN(MULT_mult_6_SUMB_4__12_) );
  NAND2_X4 MULT_mult_6_U1467 ( .A1(MULT_mult_6_n439), .A2(MULT_mult_6_net88010), .ZN(MULT_mult_6_n442) );
  NAND2_X2 MULT_mult_6_U1466 ( .A1(MULT_mult_6_ab_7__11_), .A2(
        MULT_mult_6_CARRYB_6__11_), .ZN(MULT_mult_6_net81211) );
  NAND2_X2 MULT_mult_6_U1465 ( .A1(MULT_mult_6_SUMB_5__13_), .A2(
        MULT_mult_6_ab_6__12_), .ZN(MULT_mult_6_net81713) );
  NAND2_X2 MULT_mult_6_U1464 ( .A1(MULT_mult_6_SUMB_5__13_), .A2(
        MULT_mult_6_n1439), .ZN(MULT_mult_6_net81714) );
  INV_X4 MULT_mult_6_U1463 ( .A(MULT_mult_6_CARRYB_6__11_), .ZN(
        MULT_mult_6_net87460) );
  NAND2_X2 MULT_mult_6_U1462 ( .A1(MULT_mult_6_net83045), .A2(
        MULT_mult_6_CARRYB_6__11_), .ZN(MULT_mult_6_net87462) );
  INV_X1 MULT_mult_6_U1461 ( .A(MULT_mult_6_ab_7__11_), .ZN(
        MULT_mult_6_net83045) );
  INV_X4 MULT_mult_6_U1460 ( .A(MULT_mult_6_net83045), .ZN(
        MULT_mult_6_net87461) );
  NAND2_X4 MULT_mult_6_U1459 ( .A1(MULT_mult_6_net87460), .A2(
        MULT_mult_6_net87461), .ZN(MULT_mult_6_n435) );
  NAND2_X4 MULT_mult_6_U1458 ( .A1(MULT_mult_6_net87462), .A2(MULT_mult_6_n435), .ZN(MULT_mult_6_net81209) );
  NAND2_X2 MULT_mult_6_U1457 ( .A1(MULT_mult_6_net82089), .A2(MULT_mult_6_n434), .ZN(MULT_mult_6_n432) );
  INV_X4 MULT_mult_6_U1456 ( .A(MULT_mult_6_net82089), .ZN(MULT_mult_6_n430)
         );
  INV_X2 MULT_mult_6_U1455 ( .A(MULT_mult_6_n431), .ZN(MULT_mult_6_n434) );
  INV_X2 MULT_mult_6_U1454 ( .A(MULT_mult_6_SUMB_5__13_), .ZN(MULT_mult_6_n431) );
  NAND2_X4 MULT_mult_6_U1453 ( .A1(MULT_mult_6_n430), .A2(MULT_mult_6_n431), 
        .ZN(MULT_mult_6_n433) );
  NAND2_X2 MULT_mult_6_U1452 ( .A1(MULT_mult_6_SUMB_6__12_), .A2(
        MULT_mult_6_CARRYB_6__11_), .ZN(MULT_mult_6_net81213) );
  NAND2_X2 MULT_mult_6_U1451 ( .A1(MULT_mult_6_ab_7__11_), .A2(
        MULT_mult_6_SUMB_6__12_), .ZN(MULT_mult_6_net81212) );
  NAND2_X4 MULT_mult_6_U1450 ( .A1(MULT_mult_6_n432), .A2(MULT_mult_6_n433), 
        .ZN(MULT_mult_6_SUMB_6__12_) );
  INV_X4 MULT_mult_6_U1449 ( .A(MULT_mult_6_net81209), .ZN(
        MULT_mult_6_net88105) );
  NAND2_X2 MULT_mult_6_U1448 ( .A1(MULT_mult_6_net88106), .A2(
        MULT_mult_6_net81209), .ZN(MULT_mult_6_net88107) );
  INV_X4 MULT_mult_6_U1447 ( .A(MULT_mult_6_net88106), .ZN(
        MULT_mult_6_net89021) );
  NAND2_X4 MULT_mult_6_U1446 ( .A1(MULT_mult_6_net88107), .A2(MULT_mult_6_n436), .ZN(MULT_mult_6_SUMB_7__11_) );
  NAND2_X4 MULT_mult_6_U1445 ( .A1(MULT_mult_6_net88105), .A2(
        MULT_mult_6_net89021), .ZN(MULT_mult_6_n436) );
  NAND2_X2 MULT_mult_6_U1444 ( .A1(MULT_mult_6_CARRYB_24__3_), .A2(
        MULT_mult_6_SUMB_24__4_), .ZN(MULT_mult_6_net81006) );
  NAND3_X2 MULT_mult_6_U1443 ( .A1(MULT_mult_6_n1528), .A2(MULT_mult_6_n1892), 
        .A3(MULT_mult_6_n2205), .ZN(MULT_mult_6_n1497) );
  XNOR2_X2 MULT_mult_6_U1442 ( .A(MULT_mult_6_n926), .B(
        MULT_mult_6_CARRYB_7__17_), .ZN(MULT_mult_6_net88703) );
  XNOR2_X2 MULT_mult_6_U1441 ( .A(MULT_mult_6_n1094), .B(
        MULT_mult_6_SUMB_10__16_), .ZN(MULT_mult_6_SUMB_11__15_) );
  INV_X1 MULT_mult_6_U1440 ( .A(MULT_mult_6_ab_8__16_), .ZN(MULT_mult_6_n429)
         );
  OAI211_X4 MULT_mult_6_U1439 ( .C1(MULT_mult_6_n428), .C2(MULT_mult_6_n429), 
        .A(MULT_mult_6_n2298), .B(MULT_mult_6_n2297), .ZN(
        MULT_mult_6_CARRYB_8__16_) );
  NAND2_X2 MULT_mult_6_U1438 ( .A1(MULT_mult_6_n584), .A2(MULT_mult_6_n583), 
        .ZN(MULT_mult_6_net89110) );
  NAND3_X2 MULT_mult_6_U1437 ( .A1(MULT_mult_6_net81157), .A2(MULT_mult_6_n690), .A3(MULT_mult_6_n689), .ZN(MULT_mult_6_n835) );
  NAND3_X2 MULT_mult_6_U1436 ( .A1(MULT_mult_6_n250), .A2(MULT_mult_6_net79885), .A3(MULT_mult_6_net79884), .ZN(MULT_mult_6_net87797) );
  NAND3_X2 MULT_mult_6_U1435 ( .A1(MULT_mult_6_net86022), .A2(
        MULT_mult_6_net79907), .A3(MULT_mult_6_n784), .ZN(MULT_mult_6_net86024) );
  INV_X8 MULT_mult_6_U1434 ( .A(MULT_mult_6_n427), .ZN(MULT_mult_6_net92318)
         );
  NAND3_X4 MULT_mult_6_U1433 ( .A1(MULT_mult_6_net80472), .A2(
        MULT_mult_6_net80473), .A3(MULT_mult_6_net80474), .ZN(MULT_mult_6_n427) );
  NAND2_X4 MULT_mult_6_U1432 ( .A1(MULT_mult_6_n4), .A2(MULT_mult_6_net148179), 
        .ZN(MULT_mult_6_net80668) );
  NAND2_X4 MULT_mult_6_U1431 ( .A1(MULT_mult_6_net82009), .A2(
        MULT_mult_6_ab_19__6_), .ZN(MULT_mult_6_n519) );
  INV_X4 MULT_mult_6_U1430 ( .A(MULT_mult_6_net92317), .ZN(MULT_mult_6_n606)
         );
  NAND2_X2 MULT_mult_6_U1429 ( .A1(MULT_mult_6_ab_14__2_), .A2(
        MULT_mult_6_SUMB_13__3_), .ZN(MULT_mult_6_net81779) );
  XNOR2_X2 MULT_mult_6_U1428 ( .A(MULT_mult_6_CARRYB_18__2_), .B(
        MULT_mult_6_ab_19__2_), .ZN(MULT_mult_6_n1254) );
  INV_X4 MULT_mult_6_U1427 ( .A(MULT_mult_6_ab_17__3_), .ZN(MULT_mult_6_n2013)
         );
  NAND2_X4 MULT_mult_6_U1426 ( .A1(MULT_mult_6_SUMB_16__4_), .A2(
        MULT_mult_6_ab_17__3_), .ZN(MULT_mult_6_n2107) );
  BUF_X8 MULT_mult_6_U1425 ( .A(MULT_mult_6_n424), .Z(MULT_mult_6_n1241) );
  NOR2_X2 MULT_mult_6_U1424 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__9_) );
  INV_X4 MULT_mult_6_U1423 ( .A(MULT_mult_6_ab_11__9_), .ZN(
        MULT_mult_6_net93305) );
  NAND2_X2 MULT_mult_6_U1422 ( .A1(MULT_mult_6_SUMB_4__10_), .A2(
        MULT_mult_6_n943), .ZN(MULT_mult_6_n1398) );
  NAND2_X2 MULT_mult_6_U1421 ( .A1(MULT_mult_6_net124627), .A2(
        MULT_mult_6_net81947), .ZN(MULT_mult_6_n518) );
  INV_X4 MULT_mult_6_U1420 ( .A(MULT_mult_6_ab_24__2_), .ZN(
        MULT_mult_6_net121380) );
  NAND2_X4 MULT_mult_6_U1419 ( .A1(MULT_mult_6_net119976), .A2(
        MULT_mult_6_SUMB_4__16_), .ZN(MULT_mult_6_net84446) );
  INV_X4 MULT_mult_6_U1418 ( .A(MULT_mult_6_SUMB_9__13_), .ZN(
        MULT_mult_6_net120652) );
  NAND2_X4 MULT_mult_6_U1417 ( .A1(MULT_mult_6_SUMB_10__12_), .A2(
        MULT_mult_6_ab_11__11_), .ZN(MULT_mult_6_net81167) );
  NAND2_X4 MULT_mult_6_U1416 ( .A1(MULT_mult_6_n895), .A2(
        MULT_mult_6_net123430), .ZN(MULT_mult_6_n2338) );
  INV_X2 MULT_mult_6_U1415 ( .A(MULT_mult_6_ab_7__12_), .ZN(
        MULT_mult_6_net85251) );
  NOR2_X1 MULT_mult_6_U1414 ( .A1(MULT_mult_6_net83784), .A2(
        MULT_mult_6_net77932), .ZN(MULT_mult_6_ab_7__12_) );
  NAND2_X4 MULT_mult_6_U1413 ( .A1(MULT_mult_6_SUMB_1__14_), .A2(
        MULT_mult_6_CARRYB_1__13_), .ZN(MULT_mult_6_n453) );
  XNOR2_X2 MULT_mult_6_U1412 ( .A(MULT_mult_6_ab_20__2_), .B(
        MULT_mult_6_SUMB_19__3_), .ZN(MULT_mult_6_n1232) );
  XNOR2_X2 MULT_mult_6_U1411 ( .A(MULT_mult_6_SUMB_13__2_), .B(
        MULT_mult_6_ab_14__1_), .ZN(MULT_mult_6_n426) );
  XNOR2_X2 MULT_mult_6_U1410 ( .A(MULT_mult_6_n35), .B(MULT_mult_6_n426), .ZN(
        MULT_mult_6_SUMB_14__1_) );
  NAND2_X2 MULT_mult_6_U1409 ( .A1(MULT_mult_6_CARRYB_3__13_), .A2(
        MULT_mult_6_SUMB_3__14_), .ZN(MULT_mult_6_n2091) );
  INV_X4 MULT_mult_6_U1408 ( .A(MULT_mult_6_net82009), .ZN(
        MULT_mult_6_net88856) );
  NAND2_X4 MULT_mult_6_U1407 ( .A1(MULT_mult_6_SUMB_20__5_), .A2(
        MULT_mult_6_CARRYB_20__4_), .ZN(MULT_mult_6_net82408) );
  INV_X2 MULT_mult_6_U1406 ( .A(MULT_mult_6_n1190), .ZN(MULT_mult_6_n544) );
  NOR2_X4 MULT_mult_6_U1405 ( .A1(MULT_mult_6_net82247), .A2(
        MULT_mult_6_net120391), .ZN(MULT_mult_6_ab_0__13_) );
  INV_X4 MULT_mult_6_U1404 ( .A(MULT_mult_6_net86884), .ZN(
        MULT_mult_6_net89103) );
  NAND2_X4 MULT_mult_6_U1403 ( .A1(MULT_mult_6_SUMB_18__5_), .A2(
        MULT_mult_6_ab_19__4_), .ZN(MULT_mult_6_n2235) );
  NAND2_X4 MULT_mult_6_U1402 ( .A1(MULT_mult_6_ab_4__13_), .A2(
        MULT_mult_6_SUMB_3__14_), .ZN(MULT_mult_6_n2090) );
  NAND2_X2 MULT_mult_6_U1401 ( .A1(MULT_mult_6_n1023), .A2(
        MULT_mult_6_net120501), .ZN(MULT_mult_6_n1025) );
  INV_X4 MULT_mult_6_U1400 ( .A(MULT_mult_6_ab_27__1_), .ZN(
        MULT_mult_6_net81867) );
  NAND2_X2 MULT_mult_6_U1399 ( .A1(MULT_mult_6_CARRYB_20__0_), .A2(
        MULT_mult_6_SUMB_20__1_), .ZN(MULT_mult_6_n1805) );
  NAND2_X4 MULT_mult_6_U1398 ( .A1(MULT_mult_6_n1642), .A2(MULT_mult_6_n587), 
        .ZN(MULT_mult_6_n1485) );
  NAND2_X2 MULT_mult_6_U1397 ( .A1(MULT_mult_6_ab_21__8_), .A2(
        MULT_mult_6_SUMB_20__9_), .ZN(MULT_mult_6_net81037) );
  XNOR2_X2 MULT_mult_6_U1396 ( .A(MULT_mult_6_CARRYB_19__1_), .B(
        MULT_mult_6_net89997), .ZN(MULT_mult_6_n425) );
  NAND2_X4 MULT_mult_6_U1395 ( .A1(MULT_mult_6_net92321), .A2(
        MULT_mult_6_net92325), .ZN(MULT_mult_6_n834) );
  NAND2_X2 MULT_mult_6_U1394 ( .A1(MULT_mult_6_ab_2__10_), .A2(
        MULT_mult_6_CARRYB_1__10_), .ZN(MULT_mult_6_n1652) );
  INV_X2 MULT_mult_6_U1393 ( .A(MULT_mult_6_SUMB_20__5_), .ZN(
        MULT_mult_6_net87874) );
  INV_X4 MULT_mult_6_U1392 ( .A(MULT_mult_6_net87874), .ZN(
        MULT_mult_6_net88638) );
  NOR2_X2 MULT_mult_6_U1391 ( .A1(MULT_mult_6_net70456), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__11_) );
  INV_X2 MULT_mult_6_U1390 ( .A(MULT_mult_6_ab_9__11_), .ZN(
        MULT_mult_6_net86894) );
  XNOR2_X2 MULT_mult_6_U1389 ( .A(MULT_mult_6_n1936), .B(MULT_mult_6_n863), 
        .ZN(MULT_mult_6_n424) );
  BUF_X4 MULT_mult_6_U1388 ( .A(MULT_mult_6_n864), .Z(MULT_mult_6_n1228) );
  INV_X4 MULT_mult_6_U1387 ( .A(MULT_mult_6_n1228), .ZN(MULT_mult_6_n1151) );
  NAND2_X4 MULT_mult_6_U1386 ( .A1(MULT_mult_6_n1721), .A2(MULT_mult_6_n1228), 
        .ZN(MULT_mult_6_n1152) );
  NAND2_X4 MULT_mult_6_U1385 ( .A1(MULT_mult_6_SUMB_17__4_), .A2(
        MULT_mult_6_ab_18__3_), .ZN(MULT_mult_6_n1415) );
  NOR2_X1 MULT_mult_6_U1384 ( .A1(MULT_mult_6_net77906), .A2(
        MULT_mult_6_net77924), .ZN(MULT_mult_6_ab_8__6_) );
  INV_X2 MULT_mult_6_U1383 ( .A(MULT_mult_6_ab_8__6_), .ZN(MULT_mult_6_n1650)
         );
  NAND2_X4 MULT_mult_6_U1382 ( .A1(MULT_mult_6_ab_8__6_), .A2(
        MULT_mult_6_SUMB_7__7_), .ZN(MULT_mult_6_n1826) );
  XNOR2_X2 MULT_mult_6_U1381 ( .A(MULT_mult_6_n423), .B(MULT_mult_6_n571), 
        .ZN(MULT_mult_6_SUMB_16__2_) );
  XNOR2_X1 MULT_mult_6_U1380 ( .A(MULT_mult_6_n1902), .B(MULT_mult_6_n1248), 
        .ZN(MULT_mult_6_n553) );
  INV_X4 MULT_mult_6_U1379 ( .A(MULT_mult_6_ab_12__9_), .ZN(MULT_mult_6_n1054)
         );
  NAND2_X2 MULT_mult_6_U1378 ( .A1(MULT_mult_6_SUMB_17__2_), .A2(
        MULT_mult_6_ab_18__1_), .ZN(MULT_mult_6_n745) );
  NAND3_X4 MULT_mult_6_U1377 ( .A1(MULT_mult_6_n747), .A2(MULT_mult_6_n746), 
        .A3(MULT_mult_6_n745), .ZN(MULT_mult_6_CARRYB_18__1_) );
  NAND2_X1 MULT_mult_6_U1376 ( .A1(MULT_mult_6_SUMB_2__20_), .A2(
        MULT_mult_6_CARRYB_2__19_), .ZN(MULT_mult_6_n2056) );
  NOR2_X4 MULT_mult_6_U1375 ( .A1(MULT_mult_6_net85716), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__11_) );
  INV_X4 MULT_mult_6_U1374 ( .A(MULT_mult_6_ab_10__11_), .ZN(
        MULT_mult_6_net83876) );
  AND3_X4 MULT_mult_6_U1373 ( .A1(MULT_mult_6_net88295), .A2(
        MULT_mult_6_net88296), .A3(MULT_mult_6_net88297), .ZN(MULT_mult_6_n510) );
  NAND2_X4 MULT_mult_6_U1372 ( .A1(MULT_mult_6_n641), .A2(MULT_mult_6_n642), 
        .ZN(MULT_mult_6_n644) );
  NAND2_X4 MULT_mult_6_U1371 ( .A1(MULT_mult_6_SUMB_1__18_), .A2(
        MULT_mult_6_net87683), .ZN(MULT_mult_6_net82028) );
  NAND2_X4 MULT_mult_6_U1370 ( .A1(MULT_mult_6_net123143), .A2(
        MULT_mult_6_n909), .ZN(MULT_mult_6_net91301) );
  NAND2_X4 MULT_mult_6_U1369 ( .A1(MULT_mult_6_SUMB_9__12_), .A2(
        MULT_mult_6_ab_10__11_), .ZN(MULT_mult_6_net80957) );
  INV_X4 MULT_mult_6_U1368 ( .A(MULT_mult_6_net91003), .ZN(
        MULT_mult_6_net87364) );
  NAND2_X2 MULT_mult_6_U1367 ( .A1(MULT_mult_6_CARRYB_15__3_), .A2(
        MULT_mult_6_SUMB_15__4_), .ZN(MULT_mult_6_n1129) );
  NOR2_X1 MULT_mult_6_U1366 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70449), .ZN(MULT_mult_6_ab_23__3_) );
  NAND2_X4 MULT_mult_6_U1365 ( .A1(MULT_mult_6_n418), .A2(MULT_mult_6_n413), 
        .ZN(MULT_mult_6_n417) );
  NOR2_X2 MULT_mult_6_U1364 ( .A1(MULT_mult_6_n422), .A2(MULT_mult_6_n404), 
        .ZN(MULT_mult_6_n411) );
  NOR2_X4 MULT_mult_6_U1363 ( .A1(MULT_mult_6_n404), .A2(MULT_mult_6_n406), 
        .ZN(MULT_mult_6_n408) );
  INV_X4 MULT_mult_6_U1362 ( .A(MULT_mult_6_ab_23__3_), .ZN(MULT_mult_6_n406)
         );
  NAND2_X4 MULT_mult_6_U1361 ( .A1(MULT_mult_6_SUMB_25__3_), .A2(
        MULT_mult_6_n30), .ZN(MULT_mult_6_net80989) );
  XNOR2_X2 MULT_mult_6_U1360 ( .A(MULT_mult_6_CARRYB_2__4_), .B(
        MULT_mult_6_ab_3__4_), .ZN(MULT_mult_6_n403) );
  XNOR2_X2 MULT_mult_6_U1359 ( .A(MULT_mult_6_SUMB_2__5_), .B(MULT_mult_6_n403), .ZN(MULT_mult_6_SUMB_3__4_) );
  NAND2_X2 MULT_mult_6_U1358 ( .A1(MULT_mult_6_net93747), .A2(MULT_mult_6_n826), .ZN(MULT_mult_6_net80879) );
  NAND3_X4 MULT_mult_6_U1357 ( .A1(MULT_mult_6_n1130), .A2(MULT_mult_6_n1129), 
        .A3(MULT_mult_6_n1131), .ZN(MULT_mult_6_CARRYB_16__3_) );
  XNOR2_X2 MULT_mult_6_U1356 ( .A(MULT_mult_6_CARRYB_16__3_), .B(
        MULT_mult_6_n2013), .ZN(MULT_mult_6_n559) );
  NAND2_X4 MULT_mult_6_U1355 ( .A1(MULT_mult_6_SUMB_16__4_), .A2(
        MULT_mult_6_CARRYB_16__3_), .ZN(MULT_mult_6_n2108) );
  NAND2_X4 MULT_mult_6_U1354 ( .A1(MULT_mult_6_CARRYB_17__3_), .A2(
        MULT_mult_6_n424), .ZN(MULT_mult_6_n1414) );
  INV_X4 MULT_mult_6_U1353 ( .A(MULT_mult_6_ab_21__4_), .ZN(MULT_mult_6_n945)
         );
  NAND2_X4 MULT_mult_6_U1352 ( .A1(MULT_mult_6_CARRYB_20__4_), .A2(
        MULT_mult_6_ab_21__4_), .ZN(MULT_mult_6_n1882) );
  NAND2_X2 MULT_mult_6_U1351 ( .A1(MULT_mult_6_net92317), .A2(
        MULT_mult_6_net92318), .ZN(MULT_mult_6_n608) );
  NAND2_X4 MULT_mult_6_U1350 ( .A1(MULT_mult_6_n1363), .A2(
        MULT_mult_6_net148754), .ZN(MULT_mult_6_n1365) );
  NAND2_X4 MULT_mult_6_U1349 ( .A1(MULT_mult_6_CARRYB_25__1_), .A2(
        MULT_mult_6_ab_26__1_), .ZN(MULT_mult_6_net83976) );
  XNOR2_X2 MULT_mult_6_U1348 ( .A(MULT_mult_6_SUMB_13__3_), .B(
        MULT_mult_6_ab_14__2_), .ZN(MULT_mult_6_n765) );
  NAND3_X4 MULT_mult_6_U1347 ( .A1(MULT_mult_6_n1414), .A2(MULT_mult_6_n1415), 
        .A3(MULT_mult_6_n1416), .ZN(MULT_mult_6_CARRYB_18__3_) );
  NOR2_X2 MULT_mult_6_U1346 ( .A1(MULT_mult_6_net77908), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__6_) );
  INV_X4 MULT_mult_6_U1345 ( .A(MULT_mult_6_ab_14__6_), .ZN(MULT_mult_6_n1607)
         );
  NAND2_X2 MULT_mult_6_U1344 ( .A1(MULT_mult_6_net80862), .A2(
        MULT_mult_6_SUMB_21__5_), .ZN(MULT_mult_6_net147926) );
  NAND2_X2 MULT_mult_6_U1343 ( .A1(MULT_mult_6_ab_2__21_), .A2(
        MULT_mult_6_CARRYB_1__21_), .ZN(MULT_mult_6_n2189) );
  NAND2_X2 MULT_mult_6_U1342 ( .A1(MULT_mult_6_ab_3__19_), .A2(
        MULT_mult_6_SUMB_2__20_), .ZN(MULT_mult_6_n2055) );
  NOR2_X4 MULT_mult_6_U1341 ( .A1(MULT_mult_6_net85716), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__11_) );
  NAND2_X1 MULT_mult_6_U1340 ( .A1(MULT_mult_6_ab_12__11_), .A2(
        MULT_mult_6_net90604), .ZN(MULT_mult_6_n806) );
  NAND2_X2 MULT_mult_6_U1339 ( .A1(MULT_mult_6_net90604), .A2(
        MULT_mult_6_ab_12__11_), .ZN(MULT_mult_6_net84825) );
  INV_X4 MULT_mult_6_U1338 ( .A(MULT_mult_6_ab_12__11_), .ZN(
        MULT_mult_6_net84824) );
  NAND2_X2 MULT_mult_6_U1337 ( .A1(MULT_mult_6_CARRYB_20__5_), .A2(
        MULT_mult_6_ab_21__5_), .ZN(MULT_mult_6_net79989) );
  NOR2_X4 MULT_mult_6_U1336 ( .A1(MULT_mult_6_net85716), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__11_) );
  NOR2_X1 MULT_mult_6_U1335 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__2_) );
  NAND2_X2 MULT_mult_6_U1334 ( .A1(MULT_mult_6_ab_13__2_), .A2(MULT_mult_6_n19), .ZN(MULT_mult_6_n762) );
  NAND2_X2 MULT_mult_6_U1333 ( .A1(MULT_mult_6_ab_15__3_), .A2(
        MULT_mult_6_SUMB_14__4_), .ZN(MULT_mult_6_n1992) );
  INV_X8 MULT_mult_6_U1332 ( .A(MULT_mult_6_net80264), .ZN(MULT_mult_6_n683)
         );
  XNOR2_X2 MULT_mult_6_U1331 ( .A(MULT_mult_6_n683), .B(MULT_mult_6_net89461), 
        .ZN(MULT_mult_6_net89402) );
  INV_X8 MULT_mult_6_U1330 ( .A(MULT_mult_6_n1486), .ZN(MULT_mult_6_n1345) );
  NAND2_X4 MULT_mult_6_U1329 ( .A1(MULT_mult_6_n1529), .A2(MULT_mult_6_n2064), 
        .ZN(MULT_mult_6_n1496) );
  XNOR2_X2 MULT_mult_6_U1328 ( .A(MULT_mult_6_ab_15__2_), .B(
        MULT_mult_6_CARRYB_14__2_), .ZN(MULT_mult_6_n574) );
  XNOR2_X2 MULT_mult_6_U1327 ( .A(MULT_mult_6_SUMB_26__4_), .B(
        MULT_mult_6_n1758), .ZN(MULT_mult_6_n402) );
  NAND3_X2 MULT_mult_6_U1326 ( .A1(MULT_mult_6_net81110), .A2(
        MULT_mult_6_net81111), .A3(MULT_mult_6_net81112), .ZN(
        MULT_mult_6_CARRYB_18__2_) );
  XNOR2_X2 MULT_mult_6_U1325 ( .A(MULT_mult_6_n736), .B(
        MULT_mult_6_SUMB_12__2_), .ZN(MULT_mult_6_SUMB_13__1_) );
  INV_X4 MULT_mult_6_U1324 ( .A(MULT_mult_6_n399), .ZN(MULT_mult_6_net83445)
         );
  XNOR2_X2 MULT_mult_6_U1323 ( .A(MULT_mult_6_CARRYB_13__13_), .B(
        MULT_mult_6_n400), .ZN(MULT_mult_6_n399) );
  NAND3_X2 MULT_mult_6_U1322 ( .A1(MULT_mult_6_n750), .A2(MULT_mult_6_n751), 
        .A3(MULT_mult_6_n752), .ZN(MULT_mult_6_n398) );
  NAND2_X1 MULT_mult_6_U1321 ( .A1(MULT_mult_6_CARRYB_4__20_), .A2(
        MULT_mult_6_SUMB_4__21_), .ZN(MULT_mult_6_n1883) );
  NOR2_X1 MULT_mult_6_U1320 ( .A1(MULT_mult_6_net77868), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__1_) );
  NOR2_X1 MULT_mult_6_U1319 ( .A1(MULT_mult_6_net77868), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__1_) );
  NAND2_X2 MULT_mult_6_U1318 ( .A1(MULT_mult_6_net84209), .A2(MULT_mult_6_n795), .ZN(MULT_mult_6_net84212) );
  INV_X1 MULT_mult_6_U1317 ( .A(MULT_mult_6_n795), .ZN(MULT_mult_6_n796) );
  NAND2_X4 MULT_mult_6_U1316 ( .A1(MULT_mult_6_net147928), .A2(
        MULT_mult_6_net147929), .ZN(MULT_mult_6_n678) );
  NOR2_X1 MULT_mult_6_U1315 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net77970), .ZN(MULT_mult_6_ab_2__2_) );
  INV_X2 MULT_mult_6_U1314 ( .A(MULT_mult_6_net124949), .ZN(
        MULT_mult_6_net88867) );
  NOR2_X4 MULT_mult_6_U1313 ( .A1(MULT_mult_6_n409), .A2(MULT_mult_6_n410), 
        .ZN(MULT_mult_6_n414) );
  NAND2_X4 MULT_mult_6_U1312 ( .A1(MULT_mult_6_n414), .A2(MULT_mult_6_n415), 
        .ZN(MULT_mult_6_n416) );
  NOR2_X4 MULT_mult_6_U1311 ( .A1(MULT_mult_6_net70470), .A2(
        MULT_mult_6_net70491), .ZN(MULT_mult_6_ab_2__18_) );
  NAND2_X4 MULT_mult_6_U1310 ( .A1(MULT_mult_6_net86162), .A2(
        MULT_mult_6_net80834), .ZN(MULT_mult_6_net84445) );
  NAND2_X4 MULT_mult_6_U1309 ( .A1(MULT_mult_6_n1592), .A2(MULT_mult_6_n570), 
        .ZN(MULT_mult_6_n1595) );
  NOR2_X4 MULT_mult_6_U1308 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net70465), .ZN(MULT_mult_6_ab_15__9_) );
  INV_X4 MULT_mult_6_U1307 ( .A(MULT_mult_6_ab_15__9_), .ZN(MULT_mult_6_n830)
         );
  NAND2_X4 MULT_mult_6_U1306 ( .A1(MULT_mult_6_ab_15__9_), .A2(
        MULT_mult_6_SUMB_14__10_), .ZN(MULT_mult_6_n828) );
  INV_X2 MULT_mult_6_U1305 ( .A(MULT_mult_6_net87935), .ZN(
        MULT_mult_6_net121285) );
  NAND2_X4 MULT_mult_6_U1304 ( .A1(MULT_mult_6_SUMB_1__14_), .A2(
        MULT_mult_6_net124833), .ZN(MULT_mult_6_n454) );
  INV_X8 MULT_mult_6_U1303 ( .A(MULT_mult_6_n2340), .ZN(
        MULT_mult_6_SUMB_1__19_) );
  INV_X2 MULT_mult_6_U1302 ( .A(MULT_mult_6_SUMB_1__19_), .ZN(
        MULT_mult_6_n1498) );
  NAND2_X4 MULT_mult_6_U1301 ( .A1(MULT_mult_6_SUMB_1__19_), .A2(
        MULT_mult_6_ab_2__18_), .ZN(MULT_mult_6_n1712) );
  NAND2_X4 MULT_mult_6_U1300 ( .A1(MULT_mult_6_n710), .A2(
        MULT_mult_6_SUMB_1__19_), .ZN(MULT_mult_6_n1713) );
  NOR2_X2 MULT_mult_6_U1299 ( .A1(MULT_mult_6_net84698), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__14_) );
  INV_X4 MULT_mult_6_U1298 ( .A(MULT_mult_6_ab_10__14_), .ZN(MULT_mult_6_n1037) );
  NAND2_X4 MULT_mult_6_U1297 ( .A1(MULT_mult_6_net120585), .A2(
        MULT_mult_6_net120586), .ZN(MULT_mult_6_n1020) );
  INV_X2 MULT_mult_6_U1296 ( .A(MULT_mult_6_net120585), .ZN(
        MULT_mult_6_net124434) );
  NOR2_X4 MULT_mult_6_U1295 ( .A1(MULT_mult_6_net123000), .A2(
        MULT_mult_6_net77940), .ZN(MULT_mult_6_ab_6__17_) );
  NAND2_X2 MULT_mult_6_U1294 ( .A1(MULT_mult_6_ab_6__17_), .A2(
        MULT_mult_6_n1490), .ZN(MULT_mult_6_n2247) );
  NAND2_X4 MULT_mult_6_U1293 ( .A1(MULT_mult_6_n1490), .A2(
        MULT_mult_6_ab_6__17_), .ZN(MULT_mult_6_n2046) );
  INV_X4 MULT_mult_6_U1292 ( .A(MULT_mult_6_ab_6__17_), .ZN(MULT_mult_6_n2045)
         );
  NOR2_X4 MULT_mult_6_U1291 ( .A1(MULT_mult_6_net77866), .A2(
        MULT_mult_6_net70445), .ZN(MULT_mult_6_ab_25__1_) );
  NAND3_X2 MULT_mult_6_U1290 ( .A1(MULT_mult_6_n1406), .A2(
        MULT_mult_6_net86651), .A3(MULT_mult_6_net86652), .ZN(
        MULT_mult_6_CARRYB_16__0_) );
  NAND2_X4 MULT_mult_6_U1289 ( .A1(MULT_mult_6_n366), .A2(
        MULT_mult_6_ab_22__4_), .ZN(MULT_mult_6_net79993) );
  INV_X4 MULT_mult_6_U1288 ( .A(MULT_mult_6_net92318), .ZN(MULT_mult_6_n607)
         );
  NAND2_X4 MULT_mult_6_U1287 ( .A1(MULT_mult_6_n1536), .A2(MULT_mult_6_n1535), 
        .ZN(MULT_mult_6_n1758) );
  NAND2_X4 MULT_mult_6_U1286 ( .A1(MULT_mult_6_net148828), .A2(
        MULT_mult_6_net148829), .ZN(MULT_mult_6_n490) );
  NAND3_X4 MULT_mult_6_U1285 ( .A1(MULT_mult_6_net82030), .A2(
        MULT_mult_6_net82029), .A3(MULT_mult_6_net82031), .ZN(
        MULT_mult_6_CARRYB_3__16_) );
  INV_X1 MULT_mult_6_U1284 ( .A(MULT_mult_6_SUMB_1__21_), .ZN(
        MULT_mult_6_n1683) );
  NAND2_X2 MULT_mult_6_U1283 ( .A1(MULT_mult_6_SUMB_1__21_), .A2(
        MULT_mult_6_CARRYB_1__20_), .ZN(MULT_mult_6_n2053) );
  NOR2_X2 MULT_mult_6_U1282 ( .A1(MULT_mult_6_n411), .A2(MULT_mult_6_n412), 
        .ZN(MULT_mult_6_n415) );
  NAND2_X4 MULT_mult_6_U1281 ( .A1(MULT_mult_6_n395), .A2(
        MULT_mult_6_ab_15__4_), .ZN(MULT_mult_6_n1706) );
  XNOR2_X2 MULT_mult_6_U1280 ( .A(MULT_mult_6_n1584), .B(MULT_mult_6_n1202), 
        .ZN(MULT_mult_6_n395) );
  NAND2_X4 MULT_mult_6_U1279 ( .A1(MULT_mult_6_n2248), .A2(MULT_mult_6_n1593), 
        .ZN(MULT_mult_6_n1594) );
  NAND2_X4 MULT_mult_6_U1278 ( .A1(MULT_mult_6_n504), .A2(MULT_mult_6_n505), 
        .ZN(MULT_mult_6_n507) );
  NAND2_X4 MULT_mult_6_U1277 ( .A1(MULT_mult_6_n506), .A2(MULT_mult_6_n507), 
        .ZN(MULT_mult_6_net89447) );
  INV_X8 MULT_mult_6_U1276 ( .A(MULT_mult_6_net89103), .ZN(
        MULT_mult_6_net89104) );
  NAND2_X4 MULT_mult_6_U1274 ( .A1(MULT_mult_6_n1159), .A2(MULT_mult_6_n1160), 
        .ZN(MULT_mult_6_n1162) );
  NOR2_X4 MULT_mult_6_U1273 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net70471), .ZN(MULT_mult_6_ab_12__9_) );
  NOR2_X4 MULT_mult_6_U1272 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__8_) );
  INV_X4 MULT_mult_6_U1271 ( .A(MULT_mult_6_ab_13__8_), .ZN(
        MULT_mult_6_net80694) );
  XNOR2_X2 MULT_mult_6_U1270 ( .A(MULT_mult_6_SUMB_13__17_), .B(
        MULT_mult_6_n2188), .ZN(MULT_mult_6_SUMB_14__16_) );
  NAND2_X2 MULT_mult_6_U1269 ( .A1(MULT_mult_6_SUMB_7__15_), .A2(
        MULT_mult_6_ab_8__14_), .ZN(MULT_mult_6_n604) );
  INV_X4 MULT_mult_6_U1268 ( .A(MULT_mult_6_SUMB_7__15_), .ZN(MULT_mult_6_n602) );
  INV_X1 MULT_mult_6_U1267 ( .A(MULT_mult_6_n1160), .ZN(MULT_mult_6_n972) );
  NAND2_X4 MULT_mult_6_U1266 ( .A1(MULT_mult_6_n972), .A2(MULT_mult_6_n1256), 
        .ZN(MULT_mult_6_n2070) );
  NAND3_X2 MULT_mult_6_U1265 ( .A1(MULT_mult_6_net80925), .A2(
        MULT_mult_6_net80924), .A3(MULT_mult_6_net80926), .ZN(MULT_mult_6_n394) );
  INV_X2 MULT_mult_6_U1264 ( .A(MULT_mult_6_SUMB_1__20_), .ZN(
        MULT_mult_6_n1012) );
  INV_X4 MULT_mult_6_U1263 ( .A(MULT_mult_6_net85902), .ZN(
        MULT_mult_6_net85903) );
  XNOR2_X2 MULT_mult_6_U1262 ( .A(MULT_mult_6_CARRYB_25__5_), .B(
        MULT_mult_6_ab_26__5_), .ZN(MULT_mult_6_n393) );
  NAND2_X1 MULT_mult_6_U1261 ( .A1(MULT_mult_6_ab_6__6_), .A2(
        MULT_mult_6_SUMB_5__7_), .ZN(MULT_mult_6_n1950) );
  NAND3_X4 MULT_mult_6_U1260 ( .A1(MULT_mult_6_n1330), .A2(MULT_mult_6_n1331), 
        .A3(MULT_mult_6_n1332), .ZN(MULT_mult_6_CARRYB_6__7_) );
  OAI21_X2 MULT_mult_6_U1259 ( .B1(MULT_mult_6_n1499), .B2(
        MULT_mult_6_CARRYB_6__7_), .A(MULT_mult_6_n1443), .ZN(
        MULT_mult_6_n1821) );
  NAND2_X2 MULT_mult_6_U1258 ( .A1(MULT_mult_6_ab_19__2_), .A2(
        MULT_mult_6_n2373), .ZN(MULT_mult_6_n1911) );
  INV_X4 MULT_mult_6_U1257 ( .A(MULT_mult_6_ab_21__3_), .ZN(
        MULT_mult_6_net82834) );
  NAND2_X4 MULT_mult_6_U1256 ( .A1(MULT_mult_6_SUMB_20__4_), .A2(
        MULT_mult_6_ab_21__3_), .ZN(MULT_mult_6_net80510) );
  NAND2_X4 MULT_mult_6_U1255 ( .A1(MULT_mult_6_CARRYB_23__1_), .A2(
        MULT_mult_6_ab_24__1_), .ZN(MULT_mult_6_net80922) );
  INV_X8 MULT_mult_6_U1254 ( .A(MULT_mult_6_n416), .ZN(MULT_mult_6_net86519)
         );
  AND2_X2 MULT_mult_6_U1253 ( .A1(MULT_mult_6_n247), .A2(
        MULT_mult_6_SUMB_22__4_), .ZN(MULT_mult_6_n407) );
  INV_X2 MULT_mult_6_U1252 ( .A(MULT_mult_6_n279), .ZN(MULT_mult_6_net119927)
         );
  XNOR2_X2 MULT_mult_6_U1251 ( .A(MULT_mult_6_ab_18__2_), .B(
        MULT_mult_6_CARRYB_17__2_), .ZN(MULT_mult_6_n754) );
  NAND2_X4 MULT_mult_6_U1250 ( .A1(MULT_mult_6_ab_22__7_), .A2(
        MULT_mult_6_net89461), .ZN(MULT_mult_6_net80267) );
  AND2_X2 MULT_mult_6_U1249 ( .A1(MULT_mult_6_n105), .A2(MULT_mult_6_n385), 
        .ZN(MULT_mult_6_n381) );
  OR2_X4 MULT_mult_6_U1248 ( .A1(MULT_mult_6_n375), .A2(MULT_mult_6_n376), 
        .ZN(MULT_mult_6_n391) );
  NAND2_X4 MULT_mult_6_U1247 ( .A1(MULT_mult_6_n387), .A2(MULT_mult_6_n388), 
        .ZN(MULT_mult_6_n389) );
  NOR2_X4 MULT_mult_6_U1246 ( .A1(MULT_mult_6_n381), .A2(MULT_mult_6_n382), 
        .ZN(MULT_mult_6_n388) );
  NOR2_X4 MULT_mult_6_U1245 ( .A1(MULT_mult_6_n379), .A2(MULT_mult_6_n380), 
        .ZN(MULT_mult_6_n387) );
  INV_X4 MULT_mult_6_U1244 ( .A(MULT_mult_6_n386), .ZN(MULT_mult_6_n383) );
  NOR2_X4 MULT_mult_6_U1243 ( .A1(MULT_mult_6_n374), .A2(MULT_mult_6_n375), 
        .ZN(MULT_mult_6_n386) );
  NOR2_X2 MULT_mult_6_U1242 ( .A1(MULT_mult_6_SUMB_15__11_), .A2(
        MULT_mult_6_ab_16__10_), .ZN(MULT_mult_6_n385) );
  NOR2_X2 MULT_mult_6_U1241 ( .A1(MULT_mult_6_n377), .A2(MULT_mult_6_n378), 
        .ZN(MULT_mult_6_n384) );
  NOR2_X4 MULT_mult_6_U1240 ( .A1(MULT_mult_6_n383), .A2(MULT_mult_6_n376), 
        .ZN(MULT_mult_6_n382) );
  NOR2_X4 MULT_mult_6_U1239 ( .A1(MULT_mult_6_n333), .A2(MULT_mult_6_n352), 
        .ZN(MULT_mult_6_n380) );
  NOR2_X4 MULT_mult_6_U1238 ( .A1(MULT_mult_6_n376), .A2(MULT_mult_6_n339), 
        .ZN(MULT_mult_6_n379) );
  NOR2_X2 MULT_mult_6_U1237 ( .A1(MULT_mult_6_n374), .A2(MULT_mult_6_n376), 
        .ZN(MULT_mult_6_n378) );
  NOR2_X2 MULT_mult_6_U1236 ( .A1(MULT_mult_6_n374), .A2(MULT_mult_6_n375), 
        .ZN(MULT_mult_6_n377) );
  INV_X1 MULT_mult_6_U1235 ( .A(MULT_mult_6_ab_16__10_), .ZN(MULT_mult_6_n376)
         );
  INV_X8 MULT_mult_6_U1234 ( .A(MULT_mult_6_SUMB_15__11_), .ZN(
        MULT_mult_6_n375) );
  INV_X4 MULT_mult_6_U1233 ( .A(MULT_mult_6_n105), .ZN(MULT_mult_6_n374) );
  XNOR2_X2 MULT_mult_6_U1232 ( .A(MULT_mult_6_net88776), .B(
        MULT_mult_6_net85903), .ZN(MULT_mult_6_n597) );
  NAND2_X2 MULT_mult_6_U1231 ( .A1(MULT_mult_6_n1035), .A2(MULT_mult_6_n1036), 
        .ZN(MULT_mult_6_SUMB_26__5_) );
  NAND2_X4 MULT_mult_6_U1230 ( .A1(MULT_mult_6_n1590), .A2(MULT_mult_6_n1591), 
        .ZN(MULT_mult_6_n1694) );
  INV_X1 MULT_mult_6_U1229 ( .A(MULT_mult_6_ab_7__20_), .ZN(
        MULT_mult_6_net81340) );
  NOR2_X4 MULT_mult_6_U1228 ( .A1(MULT_mult_6_net91660), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__10_) );
  INV_X2 MULT_mult_6_U1227 ( .A(MULT_mult_6_ab_10__10_), .ZN(
        MULT_mult_6_net81643) );
  XNOR2_X2 MULT_mult_6_U1226 ( .A(MULT_mult_6_ab_10__18_), .B(
        MULT_mult_6_CARRYB_9__18_), .ZN(MULT_mult_6_n373) );
  XNOR2_X2 MULT_mult_6_U1225 ( .A(MULT_mult_6_n373), .B(
        MULT_mult_6_SUMB_9__19_), .ZN(MULT_mult_6_SUMB_10__18_) );
  NOR2_X4 MULT_mult_6_U1224 ( .A1(MULT_mult_6_net124723), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__16_) );
  INV_X2 MULT_mult_6_U1223 ( .A(MULT_mult_6_ab_9__16_), .ZN(MULT_mult_6_n1600)
         );
  INV_X16 MULT_mult_6_U1222 ( .A(MULT_mult_6_net82149), .ZN(
        MULT_mult_6_net80392) );
  NAND3_X2 MULT_mult_6_U1221 ( .A1(MULT_mult_6_n2186), .A2(MULT_mult_6_n2185), 
        .A3(MULT_mult_6_n2187), .ZN(MULT_mult_6_n372) );
  NAND2_X4 MULT_mult_6_U1220 ( .A1(MULT_mult_6_ab_1__14_), .A2(
        MULT_mult_6_ab_0__15_), .ZN(MULT_mult_6__UDW__112699_net78589) );
  INV_X8 MULT_mult_6_U1219 ( .A(MULT_mult_6__UDW__112699_net78589), .ZN(
        MULT_mult_6_CARRYB_1__14_) );
  NAND2_X4 MULT_mult_6_U1218 ( .A1(MULT_mult_6_net122156), .A2(
        MULT_mult_6_CARRYB_23__1_), .ZN(MULT_mult_6_net80920) );
  INV_X2 MULT_mult_6_U1217 ( .A(MULT_mult_6_net122156), .ZN(
        MULT_mult_6_net85902) );
  INV_X2 MULT_mult_6_U1216 ( .A(MULT_mult_6_SUMB_7__14_), .ZN(
        MULT_mult_6_net85460) );
  NAND2_X4 MULT_mult_6_U1213 ( .A1(MULT_mult_6_n604), .A2(MULT_mult_6_n605), 
        .ZN(MULT_mult_6_net81995) );
  NAND2_X4 MULT_mult_6_U1212 ( .A1(MULT_mult_6_SUMB_3__11_), .A2(
        MULT_mult_6_CARRYB_3__10_), .ZN(MULT_mult_6_n1394) );
  INV_X2 MULT_mult_6_U1211 ( .A(MULT_mult_6_n369), .ZN(MULT_mult_6_n370) );
  INV_X1 MULT_mult_6_U1210 ( .A(MULT_mult_6_CARRYB_20__9_), .ZN(
        MULT_mult_6_n369) );
  NAND2_X4 MULT_mult_6_U1209 ( .A1(MULT_mult_6_SUMB_25__3_), .A2(
        MULT_mult_6_ab_26__2_), .ZN(MULT_mult_6_net80988) );
  BUF_X4 MULT_mult_6_U1208 ( .A(MULT_mult_6_n1195), .Z(MULT_mult_6_n863) );
  NAND2_X4 MULT_mult_6_U1207 ( .A1(MULT_mult_6_n602), .A2(MULT_mult_6_n603), 
        .ZN(MULT_mult_6_n605) );
  XNOR2_X2 MULT_mult_6_U1206 ( .A(MULT_mult_6_net88881), .B(
        MULT_mult_6_ab_7__14_), .ZN(MULT_mult_6_n797) );
  CLKBUF_X3 MULT_mult_6_U1205 ( .A(MULT_mult_6_SUMB_20__3_), .Z(
        MULT_mult_6_net122087) );
  NAND2_X1 MULT_mult_6_U1204 ( .A1(MULT_mult_6_CARRYB_12__14_), .A2(
        MULT_mult_6_net88756), .ZN(MULT_mult_6_net82658) );
  NAND2_X1 MULT_mult_6_U1203 ( .A1(MULT_mult_6_ab_13__14_), .A2(
        MULT_mult_6_net88756), .ZN(MULT_mult_6_net82657) );
  CLKBUF_X3 MULT_mult_6_U1202 ( .A(MULT_mult_6_n1185), .Z(MULT_mult_6_n844) );
  CLKBUF_X3 MULT_mult_6_U1201 ( .A(MULT_mult_6_CARRYB_7__14_), .Z(
        MULT_mult_6_n833) );
  NOR2_X4 MULT_mult_6_U1200 ( .A1(MULT_mult_6_net70472), .A2(
        MULT_mult_6_net82149), .ZN(MULT_mult_6_n365) );
  INV_X4 MULT_mult_6_U1199 ( .A(MULT_mult_6_net87067), .ZN(MULT_mult_6_n554)
         );
  NAND2_X2 MULT_mult_6_U1198 ( .A1(MULT_mult_6_ab_7__7_), .A2(
        MULT_mult_6_CARRYB_6__7_), .ZN(MULT_mult_6_n1822) );
  NAND2_X4 MULT_mult_6_U1197 ( .A1(MULT_mult_6_CARRYB_19__2_), .A2(
        MULT_mult_6_ab_20__2_), .ZN(MULT_mult_6_n1915) );
  INV_X8 MULT_mult_6_U1196 ( .A(MULT_mult_6__UDW__112684_net78547), .ZN(
        MULT_mult_6_net87683) );
  NAND3_X1 MULT_mult_6_U1195 ( .A1(MULT_mult_6_n2209), .A2(MULT_mult_6_n2208), 
        .A3(MULT_mult_6_n2210), .ZN(MULT_mult_6_n858) );
  NAND2_X4 MULT_mult_6_U1194 ( .A1(MULT_mult_6_CARRYB_21__7_), .A2(
        MULT_mult_6_SUMB_21__8_), .ZN(MULT_mult_6_net80268) );
  XNOR2_X2 MULT_mult_6_U1193 ( .A(MULT_mult_6_CARRYB_7__6_), .B(
        MULT_mult_6_n363), .ZN(MULT_mult_6_n561) );
  INV_X8 MULT_mult_6_U1192 ( .A(MULT_mult_6__UDW__112679_net78533), .ZN(
        MULT_mult_6_CARRYB_1__18_) );
  NAND2_X4 MULT_mult_6_U1191 ( .A1(MULT_mult_6_n401), .A2(MULT_mult_6_n365), 
        .ZN(MULT_mult_6__UDW__112679_net78533) );
  XNOR2_X2 MULT_mult_6_U1190 ( .A(MULT_mult_6_n1266), .B(
        MULT_mult_6_CARRYB_20__1_), .ZN(MULT_mult_6_SUMB_21__1_) );
  INV_X4 MULT_mult_6_U1189 ( .A(MULT_mult_6_n1224), .ZN(MULT_mult_6_n1225) );
  NAND2_X4 MULT_mult_6_U1188 ( .A1(MULT_mult_6_SUMB_13__11_), .A2(
        MULT_mult_6_ab_14__10_), .ZN(MULT_mult_6_net82161) );
  INV_X8 MULT_mult_6_U1187 ( .A(MULT_mult_6_n389), .ZN(MULT_mult_6_net85807)
         );
  NAND3_X4 MULT_mult_6_U1186 ( .A1(MULT_mult_6_net81779), .A2(
        MULT_mult_6_net81780), .A3(MULT_mult_6_net81781), .ZN(
        MULT_mult_6_CARRYB_14__2_) );
  NAND2_X2 MULT_mult_6_U1185 ( .A1(MULT_mult_6_ab_15__2_), .A2(
        MULT_mult_6_CARRYB_14__2_), .ZN(MULT_mult_6_n1970) );
  INV_X8 MULT_mult_6_U1184 ( .A(MULT_mult_6_CARRYB_15__9_), .ZN(
        MULT_mult_6_n658) );
  BUF_X8 MULT_mult_6_U1183 ( .A(MULT_mult_6_net86101), .Z(MULT_mult_6_net83263) );
  INV_X2 MULT_mult_6_U1182 ( .A(MULT_mult_6_n566), .ZN(MULT_mult_6_n567) );
  NAND2_X4 MULT_mult_6_U1180 ( .A1(MULT_mult_6_net92550), .A2(
        MULT_mult_6_net92551), .ZN(MULT_mult_6_net92553) );
  INV_X2 MULT_mult_6_U1179 ( .A(MULT_mult_6_CARRYB_17__6_), .ZN(
        MULT_mult_6_net85610) );
  NAND2_X2 MULT_mult_6_U1177 ( .A1(MULT_mult_6_ab_8__15_), .A2(
        MULT_mult_6_n858), .ZN(MULT_mult_6_n2252) );
  INV_X2 MULT_mult_6_U1176 ( .A(MULT_mult_6_n395), .ZN(MULT_mult_6_n1224) );
  XNOR2_X2 MULT_mult_6_U1175 ( .A(MULT_mult_6_n765), .B(
        MULT_mult_6_CARRYB_13__2_), .ZN(MULT_mult_6_SUMB_14__2_) );
  XNOR2_X2 MULT_mult_6_U1174 ( .A(MULT_mult_6_CARRYB_2__5_), .B(
        MULT_mult_6_ab_3__5_), .ZN(MULT_mult_6_n361) );
  XNOR2_X1 MULT_mult_6_U1173 ( .A(MULT_mult_6_SUMB_2__6_), .B(MULT_mult_6_n361), .ZN(MULT_mult_6_SUMB_3__5_) );
  NAND2_X4 MULT_mult_6_U1172 ( .A1(MULT_mult_6_n1631), .A2(MULT_mult_6_n1632), 
        .ZN(MULT_mult_6_n1634) );
  NAND2_X4 MULT_mult_6_U1171 ( .A1(MULT_mult_6_n1633), .A2(MULT_mult_6_n1634), 
        .ZN(MULT_mult_6_n1993) );
  NAND2_X2 MULT_mult_6_U1170 ( .A1(MULT_mult_6_ab_4__6_), .A2(
        MULT_mult_6_CARRYB_3__6_), .ZN(MULT_mult_6_net88206) );
  NAND2_X4 MULT_mult_6_U1169 ( .A1(MULT_mult_6_ab_0__6_), .A2(
        MULT_mult_6_ab_1__5_), .ZN(MULT_mult_6_n2329) );
  NAND2_X1 MULT_mult_6_U1168 ( .A1(MULT_mult_6_ab_1__11_), .A2(
        MULT_mult_6_ab_0__12_), .ZN(MULT_mult_6_n1024) );
  NAND3_X2 MULT_mult_6_U1167 ( .A1(MULT_mult_6_n1972), .A2(MULT_mult_6_n1971), 
        .A3(MULT_mult_6_n1970), .ZN(MULT_mult_6_CARRYB_15__2_) );
  XNOR2_X2 MULT_mult_6_U1166 ( .A(MULT_mult_6_ab_1__4_), .B(
        MULT_mult_6_ab_0__5_), .ZN(MULT_mult_6_n2328) );
  INV_X8 MULT_mult_6_U1164 ( .A(MULT_mult_6_CARRYB_11__7_), .ZN(
        MULT_mult_6_n1286) );
  OR2_X2 MULT_mult_6_U1163 ( .A1(MULT_mult_6_n405), .A2(MULT_mult_6_n406), 
        .ZN(MULT_mult_6_n418) );
  NAND2_X4 MULT_mult_6_U1162 ( .A1(MULT_mult_6_n1458), .A2(
        MULT_mult_6_SUMB_10__6_), .ZN(MULT_mult_6_n1460) );
  NAND2_X2 MULT_mult_6_U1161 ( .A1(MULT_mult_6_n1271), .A2(MULT_mult_6_n1835), 
        .ZN(MULT_mult_6_n1783) );
  INV_X4 MULT_mult_6_U1160 ( .A(MULT_mult_6_CARRYB_2__7_), .ZN(
        MULT_mult_6_n566) );
  XNOR2_X2 MULT_mult_6_U1159 ( .A(MULT_mult_6_ab_17__2_), .B(
        MULT_mult_6_SUMB_16__3_), .ZN(MULT_mult_6_n742) );
  XNOR2_X2 MULT_mult_6_U1158 ( .A(MULT_mult_6_ab_16__2_), .B(
        MULT_mult_6_CARRYB_15__2_), .ZN(MULT_mult_6_n423) );
  XNOR2_X1 MULT_mult_6_U1157 ( .A(MULT_mult_6_CARRYB_20__0_), .B(
        MULT_mult_6_ab_21__0_), .ZN(MULT_mult_6_n360) );
  NAND2_X2 MULT_mult_6_U1155 ( .A1(MULT_mult_6_n2377), .A2(
        MULT_mult_6_ab_6__8_), .ZN(MULT_mult_6_n2079) );
  NAND2_X2 MULT_mult_6_U1154 ( .A1(MULT_mult_6_SUMB_5__9_), .A2(
        MULT_mult_6_CARRYB_5__8_), .ZN(MULT_mult_6_n2077) );
  XOR2_X1 MULT_mult_6_U1152 ( .A(MULT_mult_6_ab_1__0_), .B(
        MULT_mult_6_ab_0__1_), .Z(multOut[30]) );
  NAND2_X1 MULT_mult_6_U1151 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_3__MUX_N1), .A2(
        MULT_mult_6_net92331), .ZN(MULT_mult_6_net92330) );
  NAND2_X1 MULT_mult_6_U1150 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_2__MUX_N1), .A2(
        MULT_mult_6_net92331), .ZN(MULT_mult_6_net92337) );
  INV_X2 MULT_mult_6_U1149 ( .A(MULT_mult_6_ab_22__6_), .ZN(MULT_mult_6_n824)
         );
  INV_X8 MULT_mult_6_U1148 ( .A(MULT_mult_6_net70436), .ZN(
        MULT_mult_6_net77864) );
  INV_X16 MULT_mult_6_U1147 ( .A(MULT_mult_6_net77864), .ZN(
        MULT_mult_6_net77858) );
  INV_X2 MULT_mult_6_U1146 ( .A(MULT_mult_6_ab_17__8_), .ZN(
        MULT_mult_6_net83776) );
  INV_X2 MULT_mult_6_U1145 ( .A(MULT_mult_6_ab_19__6_), .ZN(
        MULT_mult_6_net81947) );
  INV_X4 MULT_mult_6_U1144 ( .A(MULT_mult_6_ab_26__2_), .ZN(
        MULT_mult_6_net93792) );
  INV_X16 MULT_mult_6_U1143 ( .A(MULT_mult_6_n444), .ZN(MULT_mult_6_net77930)
         );
  INV_X16 MULT_mult_6_U1142 ( .A(MULT_mult_6_n443), .ZN(MULT_mult_6_n444) );
  INV_X16 MULT_mult_6_U1141 ( .A(n10930), .ZN(MULT_mult_6_net77940) );
  AND2_X2 MULT_mult_6_U1140 ( .A1(n6005), .A2(n10933), .ZN(MULT_mult_6_n357)
         );
  NOR2_X2 MULT_mult_6_U1139 ( .A1(MULT_mult_6_net91660), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__10_) );
  INV_X8 MULT_mult_6_U1138 ( .A(MULT_mult_6_n450), .ZN(MULT_mult_6_net77946)
         );
  INV_X8 MULT_mult_6_U1137 ( .A(MULT_mult_6_n450), .ZN(MULT_mult_6_net77948)
         );
  INV_X8 MULT_mult_6_U1136 ( .A(MULT_mult_6_n449), .ZN(MULT_mult_6_n450) );
  INV_X2 MULT_mult_6_U1135 ( .A(MULT_mult_6_ab_5__11_), .ZN(
        MULT_mult_6_net83351) );
  INV_X4 MULT_mult_6_U1134 ( .A(MULT_mult_6_net82238), .ZN(
        MULT_mult_6_net82239) );
  INV_X1 MULT_mult_6_U1133 ( .A(MULT_mult_6_n1111), .ZN(MULT_mult_6_net82238)
         );
  OR2_X2 MULT_mult_6_U1132 ( .A1(MULT_mult_6_ab_9__3_), .A2(MULT_mult_6_n728), 
        .ZN(MULT_mult_6_n356) );
  XOR2_X2 MULT_mult_6_U1131 ( .A(MULT_mult_6_ab_1__30_), .B(
        MULT_mult_6_ab_0__31_), .Z(MULT_mult_6_n355) );
  INV_X4 MULT_mult_6_U1130 ( .A(MULT_mult_6_n2346), .ZN(MULT_mult_6_n1692) );
  OR2_X4 MULT_mult_6_U1129 ( .A1(MULT_mult_6_net82850), .A2(MULT_mult_6_n714), 
        .ZN(MULT_mult_6_n354) );
  INV_X4 MULT_mult_6_U1128 ( .A(MULT_mult_6_n2332), .ZN(
        MULT_mult_6_CARRYB_1__10_) );
  INV_X4 MULT_mult_6_U1127 ( .A(MULT_mult_6_net90174), .ZN(
        MULT_mult_6_net88177) );
  OR2_X2 MULT_mult_6_U1125 ( .A1(MULT_mult_6_ab_16__10_), .A2(
        MULT_mult_6_CARRYB_15__10_), .ZN(MULT_mult_6_n352) );
  NAND3_X1 MULT_mult_6_U1124 ( .A1(MULT_mult_6_net80942), .A2(
        MULT_mult_6_net80941), .A3(MULT_mult_6_net80940), .ZN(MULT_mult_6_n351) );
  AND2_X2 MULT_mult_6_U1123 ( .A1(MULT_mult_6_ab_0__7_), .A2(
        MULT_mult_6_ab_1__6_), .ZN(MULT_mult_6_n350) );
  AND2_X2 MULT_mult_6_U1122 ( .A1(MULT_mult_6_ab_0__26_), .A2(
        MULT_mult_6_ab_1__25_), .ZN(MULT_mult_6_n349) );
  INV_X4 MULT_mult_6_U1121 ( .A(MULT_mult_6_CARRYB_4__10_), .ZN(
        MULT_mult_6_n1029) );
  AND3_X4 MULT_mult_6_U1120 ( .A1(MULT_mult_6_n809), .A2(MULT_mult_6_net80686), 
        .A3(MULT_mult_6_net93918), .ZN(MULT_mult_6_n348) );
  AND2_X2 MULT_mult_6_U1119 ( .A1(MULT_mult_6_ab_0__29_), .A2(
        MULT_mult_6_ab_1__28_), .ZN(MULT_mult_6_n347) );
  NAND3_X1 MULT_mult_6_U1118 ( .A1(MULT_mult_6_net84998), .A2(
        MULT_mult_6_net84999), .A3(MULT_mult_6_net85000), .ZN(MULT_mult_6_n346) );
  INV_X4 MULT_mult_6_U1117 ( .A(MULT_mult_6_n215), .ZN(MULT_mult_6_n428) );
  INV_X16 MULT_mult_6_U1116 ( .A(net78051), .ZN(MULT_mult_6_net77866) );
  AND2_X2 MULT_mult_6_U1115 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_3__MUX_N1), .A2(
        MULT_mult_6_net77864), .ZN(MULT_mult_6_n345) );
  AND2_X2 MULT_mult_6_U1114 ( .A1(WIRE_ALU_A_MUX2TO1_32BIT_2__MUX_N1), .A2(
        MULT_mult_6_net77864), .ZN(MULT_mult_6_n344) );
  NOR2_X1 MULT_mult_6_U1113 ( .A1(MULT_mult_6_net77858), .A2(
        MULT_mult_6_net70443), .ZN(MULT_mult_6_ab_26__0_) );
  NOR2_X2 MULT_mult_6_U1112 ( .A1(MULT_mult_6_net77866), .A2(
        MULT_mult_6_net77956), .ZN(MULT_mult_6_ab_4__1_) );
  NOR2_X1 MULT_mult_6_U1111 ( .A1(MULT_mult_6_net77858), .A2(
        MULT_mult_6_net70441), .ZN(MULT_mult_6_ab_27__0_) );
  INV_X4 MULT_mult_6_U1110 ( .A(MULT_mult_6_ab_20__1_), .ZN(
        MULT_mult_6_net89997) );
  NAND2_X2 MULT_mult_6_U1109 ( .A1(MULT_mult_6_CARRYB_16__1_), .A2(
        MULT_mult_6_SUMB_16__2_), .ZN(MULT_mult_6_n744) );
  NAND3_X2 MULT_mult_6_U1108 ( .A1(MULT_mult_6_n744), .A2(MULT_mult_6_net82534), .A3(MULT_mult_6_n743), .ZN(MULT_mult_6_CARRYB_17__1_) );
  NOR2_X1 MULT_mult_6_U1107 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net77946), .ZN(MULT_mult_6_ab_5__4_) );
  NOR2_X2 MULT_mult_6_U1106 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net77946), .ZN(MULT_mult_6_ab_5__3_) );
  INV_X4 MULT_mult_6_U1105 ( .A(MULT_mult_6_n2325), .ZN(
        MULT_mult_6_CARRYB_1__3_) );
  INV_X8 MULT_mult_6_U1104 ( .A(WIRE_ALU_A_MUX2TO1_32BIT_8__MUX_N1), .ZN(
        MULT_mult_6_net70449) );
  NOR2_X2 MULT_mult_6_U1103 ( .A1(MULT_mult_6_net81673), .A2(
        MULT_mult_6_net77882), .ZN(MULT_mult_6_ab_0__3_) );
  NOR2_X1 MULT_mult_6_U1102 ( .A1(MULT_mult_6_n1078), .A2(MULT_mult_6_net77858), .ZN(MULT_mult_6_ab_31__0_) );
  NOR2_X1 MULT_mult_6_U1101 ( .A1(MULT_mult_6_net77866), .A2(
        MULT_mult_6_net70441), .ZN(MULT_mult_6_ab_27__1_) );
  NOR2_X2 MULT_mult_6_U1100 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net70455), .ZN(MULT_mult_6_ab_20__3_) );
  NOR2_X1 MULT_mult_6_U1099 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70441), .ZN(MULT_mult_6_ab_27__2_) );
  INV_X4 MULT_mult_6_U1098 ( .A(MULT_mult_6_ab_13__4_), .ZN(MULT_mult_6_n1530)
         );
  INV_X4 MULT_mult_6_U1097 ( .A(MULT_mult_6_n1650), .ZN(MULT_mult_6_n363) );
  NOR2_X2 MULT_mult_6_U1096 ( .A1(MULT_mult_6_net77914), .A2(
        MULT_mult_6_net86101), .ZN(MULT_mult_6_ab_1__7_) );
  INV_X4 MULT_mult_6_U1095 ( .A(MULT_mult_6_ab_24__3_), .ZN(
        MULT_mult_6_net85109) );
  NAND2_X2 MULT_mult_6_U1094 ( .A1(MULT_mult_6_ab_22__2_), .A2(
        MULT_mult_6_SUMB_21__3_), .ZN(MULT_mult_6_net80925) );
  INV_X4 MULT_mult_6_U1093 ( .A(MULT_mult_6_ab_18__6_), .ZN(
        MULT_mult_6_net82748) );
  NAND2_X2 MULT_mult_6_U1092 ( .A1(MULT_mult_6_n683), .A2(
        MULT_mult_6_SUMB_21__8_), .ZN(MULT_mult_6_n686) );
  INV_X4 MULT_mult_6_U1091 ( .A(MULT_mult_6_ab_23__6_), .ZN(MULT_mult_6_n1234)
         );
  NAND2_X2 MULT_mult_6_U1090 ( .A1(MULT_mult_6_CARRYB_14__5_), .A2(
        MULT_mult_6_ab_15__5_), .ZN(MULT_mult_6_n1977) );
  CLKBUF_X3 MULT_mult_6_U1089 ( .A(MULT_mult_6_SUMB_14__7_), .Z(
        MULT_mult_6_n1123) );
  NOR2_X1 MULT_mult_6_U1088 ( .A1(MULT_mult_6_net77906), .A2(
        MULT_mult_6_net70473), .ZN(MULT_mult_6_ab_11__6_) );
  INV_X4 MULT_mult_6_U1087 ( .A(MULT_mult_6_n1429), .ZN(MULT_mult_6_n1430) );
  BUF_X8 MULT_mult_6_U1086 ( .A(MULT_mult_6_net70456), .Z(MULT_mult_6_net85716) );
  NOR2_X2 MULT_mult_6_U1085 ( .A1(MULT_mult_6_net77908), .A2(
        MULT_mult_6_net70453), .ZN(MULT_mult_6_ab_21__6_) );
  INV_X8 MULT_mult_6_U1084 ( .A(MULT_mult_6_net77988), .ZN(
        MULT_mult_6_net81630) );
  NAND2_X2 MULT_mult_6_U1083 ( .A1(MULT_mult_6_n615), .A2(MULT_mult_6_n616), 
        .ZN(MULT_mult_6_n618) );
  NAND2_X2 MULT_mult_6_U1082 ( .A1(MULT_mult_6_ab_14__13_), .A2(
        MULT_mult_6_SUMB_13__14_), .ZN(MULT_mult_6_n1060) );
  NAND3_X2 MULT_mult_6_U1081 ( .A1(MULT_mult_6_net79891), .A2(
        MULT_mult_6_net79892), .A3(MULT_mult_6_net79893), .ZN(
        MULT_mult_6_CARRYB_13__15_) );
  INV_X2 MULT_mult_6_U1080 ( .A(MULT_mult_6_ab_14__13_), .ZN(MULT_mult_6_n400)
         );
  INV_X4 MULT_mult_6_U1079 ( .A(MULT_mult_6_net84007), .ZN(
        MULT_mult_6_net84209) );
  NOR2_X2 MULT_mult_6_U1078 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__8_) );
  INV_X4 MULT_mult_6_U1077 ( .A(MULT_mult_6_ab_10__19_), .ZN(MULT_mult_6_n1886) );
  NAND2_X2 MULT_mult_6_U1076 ( .A1(MULT_mult_6_net121447), .A2(
        MULT_mult_6_n466), .ZN(MULT_mult_6_net89537) );
  NAND3_X2 MULT_mult_6_U1075 ( .A1(MULT_mult_6_n1843), .A2(MULT_mult_6_n1842), 
        .A3(MULT_mult_6_n1844), .ZN(MULT_mult_6_CARRYB_11__14_) );
  NOR2_X2 MULT_mult_6_U1074 ( .A1(MULT_mult_6_net124723), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__16_) );
  NAND2_X2 MULT_mult_6_U1073 ( .A1(MULT_mult_6_n1040), .A2(MULT_mult_6_n1039), 
        .ZN(MULT_mult_6_n1227) );
  NAND2_X2 MULT_mult_6_U1072 ( .A1(MULT_mult_6_SUMB_9__14_), .A2(
        MULT_mult_6_CARRYB_9__13_), .ZN(MULT_mult_6_net80248) );
  NOR2_X2 MULT_mult_6_U1071 ( .A1(MULT_mult_6_net91660), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__10_) );
  INV_X4 MULT_mult_6_U1070 ( .A(MULT_mult_6_CARRYB_4__12_), .ZN(
        MULT_mult_6_net87465) );
  INV_X16 MULT_mult_6_U1069 ( .A(MULT_mult_6_n444), .ZN(MULT_mult_6_net77932)
         );
  NAND2_X2 MULT_mult_6_U1068 ( .A1(MULT_mult_6_n957), .A2(MULT_mult_6_n958), 
        .ZN(MULT_mult_6_n960) );
  CLKBUF_X3 MULT_mult_6_U1067 ( .A(MULT_mult_6_SUMB_3__24_), .Z(
        MULT_mult_6_n1089) );
  NAND2_X2 MULT_mult_6_U1066 ( .A1(MULT_mult_6_n2360), .A2(
        MULT_mult_6_ab_9__12_), .ZN(MULT_mult_6_net81374) );
  NOR2_X2 MULT_mult_6_U1065 ( .A1(MULT_mult_6_net81424), .A2(
        MULT_mult_6_net77932), .ZN(MULT_mult_6_ab_7__15_) );
  INV_X4 MULT_mult_6_U1064 ( .A(MULT_mult_6_n2043), .ZN(MULT_mult_6_n1749) );
  NOR2_X2 MULT_mult_6_U1063 ( .A1(MULT_mult_6_net84358), .A2(MULT_mult_6_n331), 
        .ZN(MULT_mult_6_ab_2__23_) );
  NAND2_X2 MULT_mult_6_U1062 ( .A1(MULT_mult_6_ab_4__13_), .A2(
        MULT_mult_6_CARRYB_3__13_), .ZN(MULT_mult_6_n2089) );
  NAND3_X2 MULT_mult_6_U1061 ( .A1(MULT_mult_6_n2146), .A2(MULT_mult_6_n2147), 
        .A3(MULT_mult_6_n1548), .ZN(MULT_mult_6_CARRYB_3__18_) );
  NOR2_X2 MULT_mult_6_U1060 ( .A1(MULT_mult_6_net86565), .A2(
        MULT_mult_6_net77964), .ZN(MULT_mult_6_ab_3__19_) );
  NAND2_X2 MULT_mult_6_U1059 ( .A1(MULT_mult_6_n95), .A2(
        MULT_mult_6_SUMB_2__18_), .ZN(MULT_mult_6_n1716) );
  NAND2_X2 MULT_mult_6_U1058 ( .A1(MULT_mult_6_net82024), .A2(
        MULT_mult_6_SUMB_1__18_), .ZN(MULT_mult_6_n539) );
  NOR2_X1 MULT_mult_6_U1057 ( .A1(MULT_mult_6_net77860), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__0_) );
  NOR2_X2 MULT_mult_6_U1056 ( .A1(MULT_mult_6_net77860), .A2(
        MULT_mult_6_net77924), .ZN(MULT_mult_6_ab_8__0_) );
  NOR2_X1 MULT_mult_6_U1055 ( .A1(MULT_mult_6_net77858), .A2(
        MULT_mult_6_net77966), .ZN(MULT_mult_6_ab_3__0_) );
  INV_X4 MULT_mult_6_U1054 ( .A(MULT_mult_6_ab_17__1_), .ZN(
        MULT_mult_6_net88712) );
  NOR2_X1 MULT_mult_6_U1053 ( .A1(MULT_mult_6_net77866), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__1_) );
  NOR2_X1 MULT_mult_6_U1052 ( .A1(MULT_mult_6_net77866), .A2(
        MULT_mult_6_net77966), .ZN(MULT_mult_6_ab_3__1_) );
  NOR2_X1 MULT_mult_6_U1051 ( .A1(MULT_mult_6_net77858), .A2(
        MULT_mult_6_net70445), .ZN(MULT_mult_6_ab_25__0_) );
  NOR2_X2 MULT_mult_6_U1050 ( .A1(MULT_mult_6_net77898), .A2(
        MULT_mult_6_net77956), .ZN(MULT_mult_6_ab_4__5_) );
  NOR2_X2 MULT_mult_6_U1049 ( .A1(MULT_mult_6_net77886), .A2(
        MULT_mult_6_net77924), .ZN(MULT_mult_6_ab_8__3_) );
  NAND2_X2 MULT_mult_6_U1048 ( .A1(MULT_mult_6_ab_2__6_), .A2(
        MULT_mult_6_SUMB_1__7_), .ZN(MULT_mult_6_n760) );
  INV_X4 MULT_mult_6_U1047 ( .A(MULT_mult_6_net87961), .ZN(
        MULT_mult_6_net87962) );
  INV_X4 MULT_mult_6_U1046 ( .A(MULT_mult_6_n592), .ZN(MULT_mult_6_n563) );
  NOR2_X1 MULT_mult_6_U1045 ( .A1(MULT_mult_6_net77898), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__5_) );
  NOR2_X2 MULT_mult_6_U1044 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__4_) );
  NAND3_X2 MULT_mult_6_U1043 ( .A1(MULT_mult_6_n1948), .A2(MULT_mult_6_n1947), 
        .A3(MULT_mult_6_n143), .ZN(MULT_mult_6_CARRYB_5__7_) );
  NOR2_X2 MULT_mult_6_U1042 ( .A1(MULT_mult_6_net77908), .A2(
        MULT_mult_6_net70459), .ZN(MULT_mult_6_ab_18__6_) );
  INV_X4 MULT_mult_6_U1041 ( .A(MULT_mult_6_n1588), .ZN(MULT_mult_6_n1445) );
  INV_X2 MULT_mult_6_U1040 ( .A(MULT_mult_6_ab_18__10_), .ZN(MULT_mult_6_n897)
         );
  INV_X4 MULT_mult_6_U1039 ( .A(MULT_mult_6_n1553), .ZN(MULT_mult_6_n628) );
  INV_X4 MULT_mult_6_U1038 ( .A(MULT_mult_6_n1830), .ZN(MULT_mult_6_n1760) );
  NOR2_X2 MULT_mult_6_U1037 ( .A1(MULT_mult_6_net81424), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__15_) );
  INV_X4 MULT_mult_6_U1036 ( .A(MULT_mult_6_ab_9__20_), .ZN(MULT_mult_6_n1889)
         );
  NAND3_X2 MULT_mult_6_U1035 ( .A1(MULT_mult_6_n2260), .A2(MULT_mult_6_n2261), 
        .A3(MULT_mult_6_n2262), .ZN(MULT_mult_6_CARRYB_2__28_) );
  INV_X4 MULT_mult_6_U1034 ( .A(MULT_mult_6_ab_10__15_), .ZN(MULT_mult_6_n1624) );
  NAND3_X2 MULT_mult_6_U1033 ( .A1(MULT_mult_6_n2165), .A2(MULT_mult_6_n2166), 
        .A3(MULT_mult_6_n2167), .ZN(MULT_mult_6_CARRYB_2__25_) );
  NOR2_X2 MULT_mult_6_U1032 ( .A1(MULT_mult_6_net80727), .A2(
        MULT_mult_6_net77956), .ZN(MULT_mult_6_ab_4__20_) );
  NAND3_X2 MULT_mult_6_U1031 ( .A1(MULT_mult_6_n1931), .A2(MULT_mult_6_n1930), 
        .A3(MULT_mult_6_n1932), .ZN(MULT_mult_6_CARRYB_2__22_) );
  INV_X4 MULT_mult_6_U1030 ( .A(MULT_mult_6__UDW__112694_net78575), .ZN(
        MULT_mult_6_CARRYB_1__15_) );
  INV_X4 MULT_mult_6_U1029 ( .A(MULT_mult_6_n2344), .ZN(
        MULT_mult_6_SUMB_1__21_) );
  NOR2_X1 MULT_mult_6_U1028 ( .A1(MULT_mult_6_net77860), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__0_) );
  NOR2_X1 MULT_mult_6_U1027 ( .A1(MULT_mult_6_net77858), .A2(
        MULT_mult_6_net77946), .ZN(MULT_mult_6_ab_5__0_) );
  NOR2_X1 MULT_mult_6_U1026 ( .A1(MULT_mult_6_net81673), .A2(
        MULT_mult_6_net77866), .ZN(MULT_mult_6_ab_0__1_) );
  INV_X4 MULT_mult_6_U1025 ( .A(n10931), .ZN(MULT_mult_6_net77924) );
  NOR2_X1 MULT_mult_6_U1024 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net77946), .ZN(MULT_mult_6_ab_5__2_) );
  INV_X4 MULT_mult_6_U1023 ( .A(MULT_mult_6_ab_11__2_), .ZN(
        MULT_mult_6_net85032) );
  NOR2_X1 MULT_mult_6_U1022 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net77956), .ZN(MULT_mult_6_ab_4__4_) );
  NOR2_X1 MULT_mult_6_U1021 ( .A1(MULT_mult_6_net77906), .A2(
        MULT_mult_6_net77946), .ZN(MULT_mult_6_ab_5__6_) );
  NAND2_X2 MULT_mult_6_U1020 ( .A1(MULT_mult_6_n671), .A2(MULT_mult_6_n672), 
        .ZN(MULT_mult_6_n674) );
  NAND2_X2 MULT_mult_6_U1019 ( .A1(MULT_mult_6_n673), .A2(MULT_mult_6_n674), 
        .ZN(MULT_mult_6_n1198) );
  NOR2_X1 MULT_mult_6_U1018 ( .A1(MULT_mult_6_net77908), .A2(
        MULT_mult_6_net70461), .ZN(MULT_mult_6_ab_17__6_) );
  NOR2_X2 MULT_mult_6_U1017 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__8_) );
  NOR2_X2 MULT_mult_6_U1016 ( .A1(MULT_mult_6_net81673), .A2(MULT_mult_6_n2353), .ZN(MULT_mult_6_ab_0__30_) );
  INV_X4 MULT_mult_6_U1015 ( .A(net36466), .ZN(MULT_mult_6_n2353) );
  NOR2_X2 MULT_mult_6_U1014 ( .A1(MULT_mult_6_net81424), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__15_) );
  NOR2_X1 MULT_mult_6_U1013 ( .A1(MULT_mult_6_net77860), .A2(
        MULT_mult_6_net70477), .ZN(MULT_mult_6_ab_9__0_) );
  NOR2_X1 MULT_mult_6_U1012 ( .A1(MULT_mult_6_net77858), .A2(
        MULT_mult_6_net119855), .ZN(MULT_mult_6_ab_4__0_) );
  NOR2_X1 MULT_mult_6_U1011 ( .A1(MULT_mult_6_net77860), .A2(
        MULT_mult_6_net70467), .ZN(MULT_mult_6_ab_14__0_) );
  NOR2_X1 MULT_mult_6_U1010 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net77966), .ZN(MULT_mult_6_ab_3__2_) );
  INV_X8 MULT_mult_6_U1009 ( .A(aluA[20]), .ZN(MULT_mult_6_net70473) );
  NOR2_X2 MULT_mult_6_U1008 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net77924), .ZN(MULT_mult_6_ab_8__2_) );
  NOR2_X1 MULT_mult_6_U1007 ( .A1(MULT_mult_6_net77882), .A2(
        MULT_mult_6_net77966), .ZN(MULT_mult_6_ab_3__3_) );
  NOR2_X2 MULT_mult_6_U1006 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net77930), .ZN(MULT_mult_6_ab_7__4_) );
  NAND2_X2 MULT_mult_6_U1005 ( .A1(MULT_mult_6_ab_12__4_), .A2(
        MULT_mult_6_SUMB_11__5_), .ZN(MULT_mult_6_n1296) );
  NOR2_X2 MULT_mult_6_U1004 ( .A1(MULT_mult_6_net77860), .A2(
        MULT_mult_6_net77930), .ZN(MULT_mult_6_ab_7__0_) );
  NOR2_X1 MULT_mult_6_U1003 ( .A1(MULT_mult_6_net77860), .A2(
        MULT_mult_6_net77970), .ZN(MULT_mult_6_ab_2__0_) );
  NOR2_X2 MULT_mult_6_U1002 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net77930), .ZN(MULT_mult_6_ab_7__2_) );
  NOR2_X2 MULT_mult_6_U1001 ( .A1(MULT_mult_6_net77866), .A2(
        MULT_mult_6_net77970), .ZN(MULT_mult_6_ab_2__1_) );
  INV_X16 MULT_mult_6_U1000 ( .A(MULT_mult_6_net81630), .ZN(
        MULT_mult_6_net82247) );
  NOR2_X4 MULT_mult_6_U999 ( .A1(MULT_mult_6_net82247), .A2(
        MULT_mult_6_net70480), .ZN(MULT_mult_6_ab_0__23_) );
  NOR2_X4 MULT_mult_6_U998 ( .A1(MULT_mult_6_net123000), .A2(
        MULT_mult_6_net82247), .ZN(MULT_mult_6_ab_0__17_) );
  NAND2_X1 MULT_mult_6_U996 ( .A1(MULT_mult_6_SUMB_4__22_), .A2(
        MULT_mult_6_ab_5__21_), .ZN(MULT_mult_6_n1116) );
  INV_X1 MULT_mult_6_U994 ( .A(MULT_mult_6_SUMB_28__2_), .ZN(MULT_mult_6_n531)
         );
  NOR2_X4 MULT_mult_6_U993 ( .A1(MULT_mult_6_net89652), .A2(
        MULT_mult_6_net70491), .ZN(MULT_mult_6_ab_2__16_) );
  NOR2_X4 MULT_mult_6_U992 ( .A1(MULT_mult_6_n407), .A2(MULT_mult_6_n408), 
        .ZN(MULT_mult_6_n413) );
  INV_X1 MULT_mult_6_U991 ( .A(MULT_mult_6_SUMB_18__5_), .ZN(MULT_mult_6_n1347) );
  NOR2_X2 MULT_mult_6_U990 ( .A1(MULT_mult_6_n404), .A2(MULT_mult_6_n419), 
        .ZN(MULT_mult_6_n412) );
  NOR2_X4 MULT_mult_6_U989 ( .A1(MULT_mult_6_net70462), .A2(
        MULT_mult_6_net82149), .ZN(MULT_mult_6_ab_0__14_) );
  NOR2_X4 MULT_mult_6_U988 ( .A1(MULT_mult_6_net70474), .A2(
        MULT_mult_6_net80409), .ZN(MULT_mult_6_ab_1__20_) );
  NAND2_X4 MULT_mult_6_U987 ( .A1(MULT_mult_6_net82544), .A2(
        MULT_mult_6_net121770), .ZN(MULT_mult_6_net121451) );
  NAND2_X4 MULT_mult_6_U986 ( .A1(MULT_mult_6_n1155), .A2(MULT_mult_6_n1156), 
        .ZN(MULT_mult_6_n1651) );
  NAND2_X2 MULT_mult_6_U985 ( .A1(MULT_mult_6_CARRYB_5__3_), .A2(
        MULT_mult_6_SUMB_5__4_), .ZN(MULT_mult_6_n1564) );
  BUF_X16 MULT_mult_6_U984 ( .A(MULT_mult_6_SUMB_10__2_), .Z(MULT_mult_6_n730)
         );
  INV_X2 MULT_mult_6_U983 ( .A(MULT_mult_6_net123365), .ZN(
        MULT_mult_6_net83623) );
  NAND2_X2 MULT_mult_6_U982 ( .A1(MULT_mult_6_CARRYB_11__4_), .A2(
        MULT_mult_6_SUMB_11__5_), .ZN(MULT_mult_6_n1295) );
  NAND3_X4 MULT_mult_6_U981 ( .A1(MULT_mult_6_n1295), .A2(MULT_mult_6_n1296), 
        .A3(MULT_mult_6_n667), .ZN(MULT_mult_6_CARRYB_12__4_) );
  INV_X4 MULT_mult_6_U980 ( .A(MULT_mult_6_n342), .ZN(MULT_mult_6_n343) );
  INV_X2 MULT_mult_6_U979 ( .A(MULT_mult_6_CARRYB_5__4_), .ZN(MULT_mult_6_n342) );
  NAND2_X4 MULT_mult_6_U978 ( .A1(MULT_mult_6_n542), .A2(MULT_mult_6_ab_21__3_), .ZN(MULT_mult_6_net80509) );
  NAND2_X4 MULT_mult_6_U977 ( .A1(MULT_mult_6_ab_5__8_), .A2(
        MULT_mult_6_CARRYB_4__8_), .ZN(MULT_mult_6_n1964) );
  NAND2_X2 MULT_mult_6_U976 ( .A1(MULT_mult_6_CARRYB_5__20_), .A2(
        MULT_mult_6_SUMB_5__21_), .ZN(MULT_mult_6_net79935) );
  NAND2_X4 MULT_mult_6_U975 ( .A1(MULT_mult_6_net88692), .A2(
        MULT_mult_6_ab_19__8_), .ZN(MULT_mult_6_n1391) );
  NAND3_X4 MULT_mult_6_U974 ( .A1(MULT_mult_6_n1390), .A2(MULT_mult_6_n1391), 
        .A3(MULT_mult_6_n1392), .ZN(MULT_mult_6_CARRYB_19__8_) );
  INV_X16 MULT_mult_6_U973 ( .A(MULT_mult_6_net80392), .ZN(MULT_mult_6_n392)
         );
  NOR2_X4 MULT_mult_6_U972 ( .A1(MULT_mult_6_n392), .A2(MULT_mult_6_net70482), 
        .ZN(MULT_mult_6_ab_0__24_) );
  INV_X8 MULT_mult_6_U971 ( .A(MULT_mult_6_CARRYB_14__9_), .ZN(
        MULT_mult_6_n831) );
  NAND3_X4 MULT_mult_6_U970 ( .A1(MULT_mult_6_n1579), .A2(MULT_mult_6_n1580), 
        .A3(MULT_mult_6_net84746), .ZN(MULT_mult_6_CARRYB_17__10_) );
  NOR2_X4 MULT_mult_6_U969 ( .A1(MULT_mult_6_net70482), .A2(
        MULT_mult_6_net80409), .ZN(MULT_mult_6_ab_1__24_) );
  INV_X4 MULT_mult_6_U968 ( .A(MULT_mult_6_n825), .ZN(MULT_mult_6_n826) );
  BUF_X4 MULT_mult_6_U967 ( .A(MULT_mult_6_CARRYB_19__8_), .Z(
        MULT_mult_6_net89467) );
  INV_X2 MULT_mult_6_U966 ( .A(MULT_mult_6_net81663), .ZN(MULT_mult_6_n577) );
  NAND2_X4 MULT_mult_6_U965 ( .A1(MULT_mult_6_net92790), .A2(
        MULT_mult_6_ab_25__2_), .ZN(MULT_mult_6_net80262) );
  NAND2_X1 MULT_mult_6_U964 ( .A1(MULT_mult_6_SUMB_16__13_), .A2(
        MULT_mult_6_ab_17__12_), .ZN(MULT_mult_6_n893) );
  NAND2_X4 MULT_mult_6_U963 ( .A1(MULT_mult_6_ab_3__14_), .A2(
        MULT_mult_6_SUMB_2__15_), .ZN(MULT_mult_6_n1988) );
  NOR2_X4 MULT_mult_6_U962 ( .A1(MULT_mult_6_n392), .A2(MULT_mult_6_net70456), 
        .ZN(MULT_mult_6_ab_0__11_) );
  INV_X8 MULT_mult_6_U960 ( .A(MULT_mult_6__UDW__112644_net78437), .ZN(
        MULT_mult_6_SUMB_1__25_) );
  BUF_X4 MULT_mult_6_U959 ( .A(MULT_mult_6_net80564), .Z(MULT_mult_6_net83296)
         );
  NAND2_X4 MULT_mult_6_U958 ( .A1(MULT_mult_6_SUMB_4__14_), .A2(
        MULT_mult_6_ab_5__13_), .ZN(MULT_mult_6_n1981) );
  NAND2_X4 MULT_mult_6_U957 ( .A1(MULT_mult_6_SUMB_20__6_), .A2(
        MULT_mult_6_ab_21__5_), .ZN(MULT_mult_6_net79990) );
  XNOR2_X2 MULT_mult_6_U956 ( .A(MULT_mult_6_n343), .B(MULT_mult_6_ab_6__4_), 
        .ZN(MULT_mult_6_net92884) );
  NOR2_X4 MULT_mult_6_U955 ( .A1(MULT_mult_6_net124610), .A2(
        MULT_mult_6_net77912), .ZN(MULT_mult_6_ab_0__7_) );
  INV_X2 MULT_mult_6_U954 ( .A(MULT_mult_6_SUMB_6__12_), .ZN(
        MULT_mult_6_net88106) );
  NAND2_X4 MULT_mult_6_U953 ( .A1(MULT_mult_6_net84945), .A2(
        MULT_mult_6_ab_5__14_), .ZN(MULT_mult_6_net84948) );
  NAND2_X4 MULT_mult_6_U952 ( .A1(MULT_mult_6_n1855), .A2(MULT_mult_6_n1854), 
        .ZN(MULT_mult_6_n675) );
  INV_X4 MULT_mult_6_U951 ( .A(MULT_mult_6_n675), .ZN(MULT_mult_6_n340) );
  INV_X2 MULT_mult_6_U950 ( .A(MULT_mult_6_n929), .ZN(MULT_mult_6_n918) );
  NAND2_X2 MULT_mult_6_U949 ( .A1(MULT_mult_6_ab_8__14_), .A2(
        MULT_mult_6_SUMB_7__15_), .ZN(MULT_mult_6_n2272) );
  INV_X8 MULT_mult_6_U948 ( .A(MULT_mult_6_n2248), .ZN(MULT_mult_6_n1592) );
  OR2_X2 MULT_mult_6_U947 ( .A1(MULT_mult_6_SUMB_15__11_), .A2(
        MULT_mult_6_CARRYB_15__10_), .ZN(MULT_mult_6_n339) );
  BUF_X4 MULT_mult_6_U946 ( .A(MULT_mult_6_SUMB_10__13_), .Z(
        MULT_mult_6_net90262) );
  INV_X2 MULT_mult_6_U945 ( .A(MULT_mult_6_net90262), .ZN(MULT_mult_6_n336) );
  INV_X2 MULT_mult_6_U944 ( .A(MULT_mult_6_net81087), .ZN(MULT_mult_6_n335) );
  NAND2_X4 MULT_mult_6_U943 ( .A1(MULT_mult_6_n337), .A2(MULT_mult_6_n338), 
        .ZN(MULT_mult_6_net89670) );
  NAND2_X4 MULT_mult_6_U942 ( .A1(MULT_mult_6_n335), .A2(MULT_mult_6_n336), 
        .ZN(MULT_mult_6_n338) );
  NAND2_X2 MULT_mult_6_U941 ( .A1(MULT_mult_6_net81087), .A2(
        MULT_mult_6_net90262), .ZN(MULT_mult_6_n337) );
  NAND2_X4 MULT_mult_6_U940 ( .A1(MULT_mult_6_CARRYB_17__4_), .A2(
        MULT_mult_6_ab_18__4_), .ZN(MULT_mult_6_n2040) );
  NAND2_X4 MULT_mult_6_U939 ( .A1(MULT_mult_6_n915), .A2(MULT_mult_6_n916), 
        .ZN(MULT_mult_6_n1199) );
  NAND2_X4 MULT_mult_6_U937 ( .A1(MULT_mult_6_n404), .A2(MULT_mult_6_n406), 
        .ZN(MULT_mult_6_n421) );
  INV_X2 MULT_mult_6_U936 ( .A(MULT_mult_6_net147938), .ZN(MULT_mult_6_n334)
         );
  INV_X4 MULT_mult_6_U935 ( .A(MULT_mult_6_n332), .ZN(MULT_mult_6_n333) );
  INV_X1 MULT_mult_6_U934 ( .A(MULT_mult_6_n375), .ZN(MULT_mult_6_n332) );
  NAND2_X4 MULT_mult_6_U933 ( .A1(MULT_mult_6_n542), .A2(MULT_mult_6_net82834), 
        .ZN(MULT_mult_6_net83174) );
  NAND2_X4 MULT_mult_6_U932 ( .A1(MULT_mult_6_net83175), .A2(
        MULT_mult_6_net83174), .ZN(MULT_mult_6_n2244) );
  NOR2_X2 MULT_mult_6_U931 ( .A1(MULT_mult_6_net81424), .A2(
        MULT_mult_6_net77926), .ZN(MULT_mult_6_ab_8__15_) );
  INV_X1 MULT_mult_6_U930 ( .A(MULT_mult_6_ab_8__15_), .ZN(MULT_mult_6_n328)
         );
  INV_X4 MULT_mult_6_U929 ( .A(MULT_mult_6_CARRYB_7__15_), .ZN(
        MULT_mult_6_n327) );
  NAND2_X2 MULT_mult_6_U928 ( .A1(MULT_mult_6_n329), .A2(MULT_mult_6_n330), 
        .ZN(MULT_mult_6_n1736) );
  NAND2_X2 MULT_mult_6_U927 ( .A1(MULT_mult_6_n327), .A2(MULT_mult_6_n328), 
        .ZN(MULT_mult_6_n330) );
  NAND2_X1 MULT_mult_6_U926 ( .A1(MULT_mult_6_CARRYB_7__15_), .A2(
        MULT_mult_6_ab_8__15_), .ZN(MULT_mult_6_n329) );
  NAND2_X4 MULT_mult_6_U925 ( .A1(MULT_mult_6_n639), .A2(MULT_mult_6_n640), 
        .ZN(MULT_mult_6_n1741) );
  NAND2_X2 MULT_mult_6_U924 ( .A1(MULT_mult_6_CARRYB_3__7_), .A2(
        MULT_mult_6_SUMB_3__8_), .ZN(MULT_mult_6_n1910) );
  NOR2_X4 MULT_mult_6_U923 ( .A1(MULT_mult_6_net70454), .A2(
        MULT_mult_6_net86101), .ZN(MULT_mult_6_ab_1__10_) );
  NAND2_X2 MULT_mult_6_U922 ( .A1(MULT_mult_6_n1376), .A2(
        MULT_mult_6_SUMB_6__16_), .ZN(MULT_mult_6_n1377) );
  NAND2_X4 MULT_mult_6_U921 ( .A1(MULT_mult_6_SUMB_16__8_), .A2(
        MULT_mult_6_ab_17__7_), .ZN(MULT_mult_6_net81266) );
  INV_X8 MULT_mult_6_U920 ( .A(MULT_mult_6_n2329), .ZN(
        MULT_mult_6_CARRYB_1__5_) );
  NAND2_X4 MULT_mult_6_U919 ( .A1(MULT_mult_6_net93840), .A2(
        MULT_mult_6_ab_25__2_), .ZN(MULT_mult_6_net80263) );
  NOR2_X4 MULT_mult_6_U918 ( .A1(MULT_mult_6_net70474), .A2(
        MULT_mult_6_net82149), .ZN(MULT_mult_6_ab_0__20_) );
  NAND2_X2 MULT_mult_6_U917 ( .A1(MULT_mult_6_ab_23__6_), .A2(
        MULT_mult_6_net89402), .ZN(MULT_mult_6_n2284) );
  NAND2_X2 MULT_mult_6_U916 ( .A1(MULT_mult_6_n351), .A2(MULT_mult_6_net89402), 
        .ZN(MULT_mult_6_n2285) );
  NAND2_X4 MULT_mult_6_U915 ( .A1(MULT_mult_6_net80302), .A2(
        MULT_mult_6_net80660), .ZN(MULT_mult_6_net80366) );
  NOR2_X4 MULT_mult_6_U914 ( .A1(MULT_mult_6_net70476), .A2(
        MULT_mult_6_net86101), .ZN(MULT_mult_6_ab_1__21_) );
  CLKBUF_X3 MULT_mult_6_U913 ( .A(MULT_mult_6_SUMB_4__13_), .Z(
        MULT_mult_6_n448) );
  INV_X4 MULT_mult_6_U912 ( .A(MULT_mult_6_net82723), .ZN(
        MULT_mult_6_net120513) );
  NOR2_X2 MULT_mult_6_U911 ( .A1(MULT_mult_6_net70452), .A2(
        MULT_mult_6_net70475), .ZN(MULT_mult_6_ab_10__9_) );
  NAND2_X2 MULT_mult_6_U910 ( .A1(MULT_mult_6_net81581), .A2(
        MULT_mult_6_net120922), .ZN(MULT_mult_6_n873) );
  NOR2_X1 MULT_mult_6_U909 ( .A1(MULT_mult_6_net77914), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__7_) );
  INV_X1 MULT_mult_6_U908 ( .A(MULT_mult_6_ab_10__9_), .ZN(MULT_mult_6_n324)
         );
  NAND2_X4 MULT_mult_6_U907 ( .A1(MULT_mult_6_n325), .A2(MULT_mult_6_n326), 
        .ZN(MULT_mult_6_net82723) );
  INV_X1 MULT_mult_6_U906 ( .A(MULT_mult_6_ab_8__10_), .ZN(MULT_mult_6_n320)
         );
  INV_X2 MULT_mult_6_U905 ( .A(MULT_mult_6_CARRYB_7__10_), .ZN(
        MULT_mult_6_n319) );
  NAND2_X4 MULT_mult_6_U904 ( .A1(MULT_mult_6_n321), .A2(MULT_mult_6_n322), 
        .ZN(MULT_mult_6_net81581) );
  NAND2_X1 MULT_mult_6_U903 ( .A1(MULT_mult_6_CARRYB_7__10_), .A2(
        MULT_mult_6_ab_8__10_), .ZN(MULT_mult_6_n321) );
  NAND2_X4 MULT_mult_6_U902 ( .A1(MULT_mult_6_n317), .A2(MULT_mult_6_n318), 
        .ZN(MULT_mult_6_net89227) );
  NAND2_X1 MULT_mult_6_U901 ( .A1(MULT_mult_6_n89), .A2(MULT_mult_6_ab_4__12_), 
        .ZN(MULT_mult_6_n317) );
  INV_X1 MULT_mult_6_U900 ( .A(MULT_mult_6_ab_13__7_), .ZN(MULT_mult_6_n314)
         );
  NAND2_X4 MULT_mult_6_U898 ( .A1(MULT_mult_6_n2022), .A2(MULT_mult_6_n315), 
        .ZN(MULT_mult_6_n1732) );
  NAND2_X4 MULT_mult_6_U897 ( .A1(MULT_mult_6_n313), .A2(MULT_mult_6_n314), 
        .ZN(MULT_mult_6_n315) );
  NOR2_X1 MULT_mult_6_U896 ( .A1(MULT_mult_6_net70486), .A2(
        MULT_mult_6_net77966), .ZN(MULT_mult_6_ab_3__26_) );
  NAND2_X4 MULT_mult_6_U895 ( .A1(MULT_mult_6_SUMB_1__13_), .A2(
        MULT_mult_6_ab_2__12_), .ZN(MULT_mult_6_n2080) );
  NAND2_X2 MULT_mult_6_U894 ( .A1(net36470), .A2(MULT_mult_6_net81630), .ZN(
        MULT_mult_6_net86959) );
  INV_X16 MULT_mult_6_U893 ( .A(net36470), .ZN(MULT_mult_6_net70470) );
  INV_X8 MULT_mult_6_U892 ( .A(MULT_mult_6_net93914), .ZN(MULT_mult_6_net82009) );
  BUF_X8 MULT_mult_6_U891 ( .A(MULT_mult_6_net88344), .Z(MULT_mult_6_net124723) );
  NOR2_X2 MULT_mult_6_U890 ( .A1(MULT_mult_6_net88344), .A2(
        MULT_mult_6_net77948), .ZN(MULT_mult_6_ab_5__16_) );
  NAND2_X2 MULT_mult_6_U889 ( .A1(MULT_mult_6_net81416), .A2(MULT_mult_6_n112), 
        .ZN(MULT_mult_6__UDW__112694_net78575) );
  NOR2_X1 MULT_mult_6_U888 ( .A1(MULT_mult_6_n2355), .A2(MULT_mult_6_n175), 
        .ZN(MULT_mult_6_ab_2__27_) );
  NOR2_X1 MULT_mult_6_U887 ( .A1(MULT_mult_6_n2354), .A2(MULT_mult_6_n175), 
        .ZN(MULT_mult_6_ab_2__28_) );
  NAND2_X2 MULT_mult_6_U885 ( .A1(MULT_mult_6_ab_22__0_), .A2(
        MULT_mult_6_SUMB_21__1_), .ZN(MULT_mult_6_n1797) );
  INV_X2 MULT_mult_6_U883 ( .A(MULT_mult_6_SUMB_17__8_), .ZN(MULT_mult_6_n308)
         );
  NAND2_X4 MULT_mult_6_U882 ( .A1(MULT_mult_6_n309), .A2(MULT_mult_6_n310), 
        .ZN(MULT_mult_6_SUMB_18__7_) );
  NAND2_X4 MULT_mult_6_U881 ( .A1(MULT_mult_6_n307), .A2(MULT_mult_6_n308), 
        .ZN(MULT_mult_6_n310) );
  NAND2_X2 MULT_mult_6_U880 ( .A1(MULT_mult_6_ab_8__10_), .A2(
        MULT_mult_6_CARRYB_7__10_), .ZN(MULT_mult_6_n461) );
  INV_X4 MULT_mult_6_U879 ( .A(MULT_mult_6_net86374), .ZN(MULT_mult_6_net86375) );
  INV_X4 MULT_mult_6_U878 ( .A(MULT_mult_6_net86374), .ZN(MULT_mult_6_n306) );
  NAND2_X4 MULT_mult_6_U877 ( .A1(MULT_mult_6_net85808), .A2(
        MULT_mult_6_ab_17__9_), .ZN(MULT_mult_6_net80813) );
  NAND2_X4 MULT_mult_6_U876 ( .A1(MULT_mult_6_n575), .A2(MULT_mult_6_n679), 
        .ZN(MULT_mult_6_n681) );
  NAND2_X2 MULT_mult_6_U875 ( .A1(MULT_mult_6_SUMB_18__9_), .A2(
        MULT_mult_6_net93683), .ZN(MULT_mult_6_n643) );
  NAND2_X4 MULT_mult_6_U874 ( .A1(MULT_mult_6_n819), .A2(MULT_mult_6_n820), 
        .ZN(MULT_mult_6_n822) );
  NAND2_X1 MULT_mult_6_U873 ( .A1(MULT_mult_6_net88916), .A2(
        MULT_mult_6_net86696), .ZN(MULT_mult_6_net79868) );
  NAND2_X2 MULT_mult_6_U872 ( .A1(MULT_mult_6_ab_4__12_), .A2(MULT_mult_6_n89), 
        .ZN(MULT_mult_6_n1829) );
  NAND2_X4 MULT_mult_6_U871 ( .A1(MULT_mult_6_n1615), .A2(MULT_mult_6_n1614), 
        .ZN(MULT_mult_6_n1616) );
  NAND2_X2 MULT_mult_6_U870 ( .A1(MULT_mult_6_SUMB_6__6_), .A2(
        MULT_mult_6_CARRYB_6__5_), .ZN(MULT_mult_6_n1519) );
  NAND2_X2 MULT_mult_6_U869 ( .A1(MULT_mult_6_SUMB_22__2_), .A2(
        MULT_mult_6_ab_23__1_), .ZN(MULT_mult_6_n751) );
  NAND3_X4 MULT_mult_6_U868 ( .A1(MULT_mult_6_n1954), .A2(MULT_mult_6_n1953), 
        .A3(MULT_mult_6_n1952), .ZN(MULT_mult_6_CARRYB_16__14_) );
  NAND2_X4 MULT_mult_6_U867 ( .A1(MULT_mult_6_net123269), .A2(
        MULT_mult_6_net123268), .ZN(MULT_mult_6_net119955) );
  XNOR2_X2 MULT_mult_6_U866 ( .A(MULT_mult_6_SUMB_14__15_), .B(
        MULT_mult_6_net86054), .ZN(MULT_mult_6_net90525) );
  NOR2_X4 MULT_mult_6_U865 ( .A1(MULT_mult_6_net82043), .A2(
        MULT_mult_6_net82044), .ZN(MULT_mult_6_net82124) );
  XNOR2_X2 MULT_mult_6_U864 ( .A(MULT_mult_6_ab_4__6_), .B(
        MULT_mult_6_CARRYB_3__6_), .ZN(MULT_mult_6_n774) );
  INV_X8 MULT_mult_6_U863 ( .A(MULT_mult_6_ab_0__16_), .ZN(MULT_mult_6_n303)
         );
  INV_X4 MULT_mult_6_U862 ( .A(MULT_mult_6_ab_1__15_), .ZN(MULT_mult_6_n302)
         );
  NAND2_X4 MULT_mult_6_U861 ( .A1(MULT_mult_6_n304), .A2(MULT_mult_6_n305), 
        .ZN(MULT_mult_6_n437) );
  NAND2_X4 MULT_mult_6_U860 ( .A1(MULT_mult_6_n302), .A2(MULT_mult_6_n303), 
        .ZN(MULT_mult_6_n305) );
  NAND2_X2 MULT_mult_6_U859 ( .A1(MULT_mult_6_n112), .A2(MULT_mult_6_ab_0__16_), .ZN(MULT_mult_6_n304) );
  NAND2_X2 MULT_mult_6_U858 ( .A1(MULT_mult_6_SUMB_10__16_), .A2(
        MULT_mult_6_CARRYB_10__15_), .ZN(MULT_mult_6_n1091) );
  INV_X1 MULT_mult_6_U857 ( .A(MULT_mult_6_n393), .ZN(MULT_mult_6_net84979) );
  NAND2_X4 MULT_mult_6_U856 ( .A1(MULT_mult_6_net82759), .A2(MULT_mult_6_n1829), .ZN(MULT_mult_6_n1734) );
  NAND2_X4 MULT_mult_6_U855 ( .A1(MULT_mult_6_net84672), .A2(
        MULT_mult_6_net84671), .ZN(MULT_mult_6_SUMB_9__12_) );
  INV_X8 MULT_mult_6_U854 ( .A(MULT_mult_6_net84327), .ZN(
        MULT_mult_6_net119921) );
  NAND2_X1 MULT_mult_6_U853 ( .A1(MULT_mult_6_net89168), .A2(
        MULT_mult_6_net122062), .ZN(MULT_mult_6_n300) );
  NAND3_X4 MULT_mult_6_U852 ( .A1(MULT_mult_6_n296), .A2(MULT_mult_6_n297), 
        .A3(MULT_mult_6_n298), .ZN(MULT_mult_6_CARRYB_14__0_) );
  NAND2_X2 MULT_mult_6_U851 ( .A1(MULT_mult_6_SUMB_13__1_), .A2(
        MULT_mult_6_CARRYB_13__0_), .ZN(MULT_mult_6_n298) );
  NAND2_X1 MULT_mult_6_U850 ( .A1(MULT_mult_6_ab_14__0_), .A2(
        MULT_mult_6_CARRYB_13__0_), .ZN(MULT_mult_6_n297) );
  NAND2_X2 MULT_mult_6_U849 ( .A1(MULT_mult_6_ab_14__0_), .A2(
        MULT_mult_6_SUMB_13__1_), .ZN(MULT_mult_6_n296) );
  XOR2_X1 MULT_mult_6_U848 ( .A(MULT_mult_6_n295), .B(
        MULT_mult_6_CARRYB_13__0_), .Z(multOut[17]) );
  XOR2_X1 MULT_mult_6_U847 ( .A(MULT_mult_6_ab_14__0_), .B(
        MULT_mult_6_SUMB_13__1_), .Z(MULT_mult_6_n295) );
  NAND3_X4 MULT_mult_6_U846 ( .A1(MULT_mult_6_n292), .A2(MULT_mult_6_n293), 
        .A3(MULT_mult_6_n294), .ZN(MULT_mult_6_CARRYB_13__0_) );
  NAND2_X2 MULT_mult_6_U845 ( .A1(MULT_mult_6_SUMB_12__1_), .A2(
        MULT_mult_6_CARRYB_12__0_), .ZN(MULT_mult_6_n294) );
  NAND2_X2 MULT_mult_6_U844 ( .A1(MULT_mult_6_ab_13__0_), .A2(
        MULT_mult_6_CARRYB_12__0_), .ZN(MULT_mult_6_n293) );
  NAND2_X2 MULT_mult_6_U843 ( .A1(MULT_mult_6_ab_13__0_), .A2(
        MULT_mult_6_SUMB_12__1_), .ZN(MULT_mult_6_n292) );
  XOR2_X2 MULT_mult_6_U842 ( .A(MULT_mult_6_n291), .B(
        MULT_mult_6_CARRYB_12__0_), .Z(multOut[18]) );
  XOR2_X2 MULT_mult_6_U841 ( .A(MULT_mult_6_ab_13__0_), .B(
        MULT_mult_6_SUMB_12__1_), .Z(MULT_mult_6_n291) );
  NOR2_X4 MULT_mult_6_U840 ( .A1(MULT_mult_6_n405), .A2(MULT_mult_6_n421), 
        .ZN(MULT_mult_6_n410) );
  INV_X8 MULT_mult_6_U839 ( .A(MULT_mult_6_ab_2__11_), .ZN(MULT_mult_6_n585)
         );
  INV_X4 MULT_mult_6_U838 ( .A(MULT_mult_6_SUMB_6__9_), .ZN(MULT_mult_6_n1429)
         );
  XNOR2_X2 MULT_mult_6_U836 ( .A(MULT_mult_6_n1216), .B(MULT_mult_6_n1220), 
        .ZN(MULT_mult_6_n556) );
  XNOR2_X2 MULT_mult_6_U835 ( .A(MULT_mult_6_ab_8__16_), .B(
        MULT_mult_6_CARRYB_7__16_), .ZN(MULT_mult_6_n849) );
  INV_X2 MULT_mult_6_U834 ( .A(MULT_mult_6_SUMB_1__13_), .ZN(
        MULT_mult_6_net123509) );
  NAND2_X2 MULT_mult_6_U833 ( .A1(MULT_mult_6_SUMB_7__11_), .A2(
        MULT_mult_6_CARRYB_7__10_), .ZN(MULT_mult_6_net81216) );
  INV_X2 MULT_mult_6_U831 ( .A(MULT_mult_6_net83755), .ZN(
        MULT_mult_6_net120518) );
  NAND2_X2 MULT_mult_6_U830 ( .A1(MULT_mult_6_SUMB_9__10_), .A2(
        MULT_mult_6_CARRYB_9__9_), .ZN(MULT_mult_6_n472) );
  NAND2_X2 MULT_mult_6_U829 ( .A1(MULT_mult_6_CARRYB_1__15_), .A2(
        MULT_mult_6_SUMB_1__16_), .ZN(MULT_mult_6_n1986) );
  INV_X8 MULT_mult_6_U827 ( .A(MULT_mult_6_CARRYB_18__7_), .ZN(
        MULT_mult_6_n1615) );
  INV_X2 MULT_mult_6_U826 ( .A(MULT_mult_6_n1118), .ZN(MULT_mult_6_net80643)
         );
  NAND3_X4 MULT_mult_6_U825 ( .A1(MULT_mult_6_n1106), .A2(MULT_mult_6_n1105), 
        .A3(MULT_mult_6_n1107), .ZN(MULT_mult_6_CARRYB_8__18_) );
  NAND2_X4 MULT_mult_6_U824 ( .A1(MULT_mult_6_SUMB_10__15_), .A2(
        MULT_mult_6_CARRYB_10__14_), .ZN(MULT_mult_6_n1844) );
  INV_X8 MULT_mult_6_U823 ( .A(MULT_mult_6_n933), .ZN(MULT_mult_6_n936) );
  CLKBUF_X3 MULT_mult_6_U822 ( .A(MULT_mult_6_CARRYB_13__13_), .Z(
        MULT_mult_6_n695) );
  NAND2_X1 MULT_mult_6_U821 ( .A1(MULT_mult_6_ab_15__12_), .A2(
        MULT_mult_6_SUMB_14__13_), .ZN(MULT_mult_6_n2199) );
  NAND2_X1 MULT_mult_6_U820 ( .A1(MULT_mult_6_ab_3__12_), .A2(
        MULT_mult_6_n1207), .ZN(MULT_mult_6_n2009) );
  BUF_X4 MULT_mult_6_U819 ( .A(MULT_mult_6_SUMB_8__11_), .Z(
        MULT_mult_6_net125375) );
  NAND2_X2 MULT_mult_6_U818 ( .A1(MULT_mult_6_n300), .A2(MULT_mult_6_n301), 
        .ZN(MULT_mult_6_SUMB_12__9_) );
  INV_X4 MULT_mult_6_U817 ( .A(MULT_mult_6_SUMB_24__4_), .ZN(
        MULT_mult_6_net87938) );
  INV_X32 MULT_mult_6_U816 ( .A(MULT_mult_6_net85109), .ZN(MULT_mult_6_n286)
         );
  XNOR2_X2 MULT_mult_6_U815 ( .A(MULT_mult_6_n417), .B(MULT_mult_6_n286), .ZN(
        MULT_mult_6_n285) );
  NAND2_X2 MULT_mult_6_U814 ( .A1(MULT_mult_6_n944), .A2(MULT_mult_6_net87874), 
        .ZN(MULT_mult_6_n1337) );
  NAND2_X4 MULT_mult_6_U813 ( .A1(MULT_mult_6_SUMB_25__2_), .A2(
        MULT_mult_6_ab_26__1_), .ZN(MULT_mult_6_net83977) );
  NAND2_X4 MULT_mult_6_U812 ( .A1(MULT_mult_6_CARRYB_28__0_), .A2(
        MULT_mult_6_n344), .ZN(MULT_mult_6_net79883) );
  NAND2_X2 MULT_mult_6_U811 ( .A1(MULT_mult_6_n728), .A2(
        MULT_mult_6_SUMB_8__4_), .ZN(MULT_mult_6_net82850) );
  XNOR2_X2 MULT_mult_6_U810 ( .A(MULT_mult_6_net119952), .B(
        MULT_mult_6__UDW__112684_net78549), .ZN(MULT_mult_6_net149611) );
  INV_X4 MULT_mult_6_U809 ( .A(MULT_mult_6_CARRYB_1__16_), .ZN(
        MULT_mult_6_n281) );
  NAND2_X4 MULT_mult_6_U807 ( .A1(MULT_mult_6_n283), .A2(MULT_mult_6_n282), 
        .ZN(MULT_mult_6_net119952) );
  NAND2_X2 MULT_mult_6_U806 ( .A1(MULT_mult_6_ab_2__16_), .A2(
        MULT_mult_6_CARRYB_1__16_), .ZN(MULT_mult_6_n282) );
  OAI21_X4 MULT_mult_6_U805 ( .B1(MULT_mult_6_net119909), .B2(
        MULT_mult_6_net119910), .A(MULT_mult_6_n477), .ZN(MULT_mult_6_n279) );
  INV_X4 MULT_mult_6_U803 ( .A(MULT_mult_6_n38), .ZN(MULT_mult_6_n1628) );
  NAND2_X4 MULT_mult_6_U802 ( .A1(MULT_mult_6_ab_10__8_), .A2(
        MULT_mult_6_SUMB_9__9_), .ZN(MULT_mult_6_n1775) );
  NAND2_X2 MULT_mult_6_U801 ( .A1(MULT_mult_6_net120625), .A2(
        MULT_mult_6_net120626), .ZN(MULT_mult_6_net120628) );
  NAND2_X2 MULT_mult_6_U800 ( .A1(MULT_mult_6_n1233), .A2(
        MULT_mult_6_ab_4__20_), .ZN(MULT_mult_6_n2238) );
  NAND2_X2 MULT_mult_6_U799 ( .A1(MULT_mult_6_ab_6__19_), .A2(
        MULT_mult_6_SUMB_5__20_), .ZN(MULT_mult_6_n2280) );
  NAND2_X2 MULT_mult_6_U798 ( .A1(MULT_mult_6_n56), .A2(
        MULT_mult_6_SUMB_5__20_), .ZN(MULT_mult_6_n2281) );
  NAND2_X1 MULT_mult_6_U797 ( .A1(n6005), .A2(
        WIRE_ALU_A_MUX2TO1_32BIT_3__MUX_N1), .ZN(MULT_mult_6_net92311) );
  INV_X4 MULT_mult_6_U796 ( .A(MULT_mult_6_net93107), .ZN(MULT_mult_6_n276) );
  INV_X2 MULT_mult_6_U795 ( .A(MULT_mult_6_SUMB_14__14_), .ZN(MULT_mult_6_n275) );
  NAND2_X4 MULT_mult_6_U794 ( .A1(MULT_mult_6_n277), .A2(MULT_mult_6_n278), 
        .ZN(MULT_mult_6_SUMB_15__13_) );
  NAND2_X4 MULT_mult_6_U793 ( .A1(MULT_mult_6_n275), .A2(MULT_mult_6_n276), 
        .ZN(MULT_mult_6_n278) );
  NAND2_X2 MULT_mult_6_U792 ( .A1(MULT_mult_6_SUMB_14__14_), .A2(
        MULT_mult_6_net93107), .ZN(MULT_mult_6_n277) );
  INV_X2 MULT_mult_6_U791 ( .A(MULT_mult_6_SUMB_13__15_), .ZN(MULT_mult_6_n272) );
  INV_X4 MULT_mult_6_U790 ( .A(MULT_mult_6_net85119), .ZN(MULT_mult_6_n271) );
  NAND2_X4 MULT_mult_6_U789 ( .A1(MULT_mult_6_n273), .A2(MULT_mult_6_n274), 
        .ZN(MULT_mult_6_SUMB_14__14_) );
  NAND2_X4 MULT_mult_6_U788 ( .A1(MULT_mult_6_n271), .A2(MULT_mult_6_n272), 
        .ZN(MULT_mult_6_n274) );
  NAND2_X2 MULT_mult_6_U787 ( .A1(MULT_mult_6_net85119), .A2(
        MULT_mult_6_SUMB_13__15_), .ZN(MULT_mult_6_n273) );
  INV_X4 MULT_mult_6_U786 ( .A(MULT_mult_6_net90801), .ZN(MULT_mult_6_n268) );
  INV_X4 MULT_mult_6_U785 ( .A(MULT_mult_6_n859), .ZN(MULT_mult_6_n267) );
  NAND2_X4 MULT_mult_6_U784 ( .A1(MULT_mult_6_n269), .A2(MULT_mult_6_n270), 
        .ZN(MULT_mult_6_net89461) );
  NAND2_X4 MULT_mult_6_U783 ( .A1(MULT_mult_6_n267), .A2(MULT_mult_6_n268), 
        .ZN(MULT_mult_6_n270) );
  NAND2_X2 MULT_mult_6_U782 ( .A1(MULT_mult_6_n859), .A2(MULT_mult_6_net90801), 
        .ZN(MULT_mult_6_n269) );
  INV_X2 MULT_mult_6_U781 ( .A(MULT_mult_6_n866), .ZN(MULT_mult_6_n264) );
  INV_X4 MULT_mult_6_U780 ( .A(MULT_mult_6_n1609), .ZN(MULT_mult_6_n263) );
  NAND2_X4 MULT_mult_6_U779 ( .A1(MULT_mult_6_n265), .A2(MULT_mult_6_n266), 
        .ZN(MULT_mult_6_n1233) );
  NAND2_X4 MULT_mult_6_U778 ( .A1(MULT_mult_6_n263), .A2(MULT_mult_6_n264), 
        .ZN(MULT_mult_6_n266) );
  NAND2_X2 MULT_mult_6_U777 ( .A1(MULT_mult_6_n1609), .A2(MULT_mult_6_n866), 
        .ZN(MULT_mult_6_n265) );
  INV_X1 MULT_mult_6_U776 ( .A(MULT_mult_6_net83116), .ZN(MULT_mult_6_n262) );
  INV_X4 MULT_mult_6_U775 ( .A(MULT_mult_6_n348), .ZN(MULT_mult_6_n260) );
  NOR2_X2 MULT_mult_6_U774 ( .A1(MULT_mult_6_n530), .A2(MULT_mult_6_n261), 
        .ZN(MULT_mult_6_net92314) );
  NOR2_X4 MULT_mult_6_U773 ( .A1(MULT_mult_6_ab_28__2_), .A2(MULT_mult_6_n260), 
        .ZN(MULT_mult_6_n261) );
  NAND2_X4 MULT_mult_6_U772 ( .A1(MULT_mult_6_net88692), .A2(
        MULT_mult_6_net121150), .ZN(MULT_mult_6_n1390) );
  NOR2_X1 MULT_mult_6_U771 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net86101), .ZN(MULT_mult_6_ab_1__2_) );
  NOR2_X2 MULT_mult_6_U770 ( .A1(MULT_mult_6_net77908), .A2(
        MULT_mult_6_net70469), .ZN(MULT_mult_6_ab_13__6_) );
  INV_X1 MULT_mult_6_U769 ( .A(MULT_mult_6_ab_13__6_), .ZN(MULT_mult_6_n257)
         );
  INV_X4 MULT_mult_6_U768 ( .A(MULT_mult_6_SUMB_12__7_), .ZN(MULT_mult_6_n256)
         );
  NAND2_X2 MULT_mult_6_U767 ( .A1(MULT_mult_6_n258), .A2(MULT_mult_6_n259), 
        .ZN(MULT_mult_6_n1899) );
  NAND2_X2 MULT_mult_6_U766 ( .A1(MULT_mult_6_SUMB_12__7_), .A2(
        MULT_mult_6_ab_13__6_), .ZN(MULT_mult_6_n258) );
  BUF_X4 MULT_mult_6_U765 ( .A(MULT_mult_6_SUMB_12__6_), .Z(MULT_mult_6_n1260)
         );
  INV_X4 MULT_mult_6_U764 ( .A(MULT_mult_6_n371), .ZN(MULT_mult_6_n253) );
  INV_X4 MULT_mult_6_U763 ( .A(MULT_mult_6_n1764), .ZN(MULT_mult_6_n252) );
  NAND2_X4 MULT_mult_6_U762 ( .A1(MULT_mult_6_n255), .A2(MULT_mult_6_n254), 
        .ZN(MULT_mult_6_SUMB_12__6_) );
  NAND2_X4 MULT_mult_6_U761 ( .A1(MULT_mult_6_n252), .A2(MULT_mult_6_n253), 
        .ZN(MULT_mult_6_n255) );
  INV_X4 MULT_mult_6_U760 ( .A(MULT_mult_6_n344), .ZN(MULT_mult_6_n249) );
  INV_X2 MULT_mult_6_U759 ( .A(MULT_mult_6_CARRYB_28__0_), .ZN(
        MULT_mult_6_n248) );
  NAND2_X4 MULT_mult_6_U758 ( .A1(MULT_mult_6_n250), .A2(MULT_mult_6_n251), 
        .ZN(MULT_mult_6_net81431) );
  NAND3_X2 MULT_mult_6_U757 ( .A1(MULT_mult_6_n503), .A2(MULT_mult_6_n501), 
        .A3(MULT_mult_6_n502), .ZN(MULT_mult_6_n247) );
  XNOR2_X2 MULT_mult_6_U756 ( .A(MULT_mult_6_CARRYB_19__8_), .B(
        MULT_mult_6_ab_20__8_), .ZN(MULT_mult_6_n368) );
  NAND2_X4 MULT_mult_6_U755 ( .A1(MULT_mult_6_CARRYB_11__7_), .A2(
        MULT_mult_6_ab_12__7_), .ZN(MULT_mult_6_n2019) );
  NAND2_X4 MULT_mult_6_U754 ( .A1(MULT_mult_6_net124367), .A2(
        MULT_mult_6_net123303), .ZN(MULT_mult_6_n2158) );
  INV_X2 MULT_mult_6_U753 ( .A(MULT_mult_6_net121859), .ZN(MULT_mult_6_n244)
         );
  INV_X1 MULT_mult_6_U752 ( .A(MULT_mult_6_net149611), .ZN(MULT_mult_6_n243)
         );
  NAND2_X4 MULT_mult_6_U751 ( .A1(MULT_mult_6_n245), .A2(MULT_mult_6_n246), 
        .ZN(MULT_mult_6_SUMB_3__15_) );
  NAND2_X1 MULT_mult_6_U750 ( .A1(MULT_mult_6_net149611), .A2(
        MULT_mult_6_net121859), .ZN(MULT_mult_6_n245) );
  INV_X4 MULT_mult_6_U749 ( .A(MULT_mult_6_net81581), .ZN(
        MULT_mult_6_net123842) );
  NAND2_X4 MULT_mult_6_U748 ( .A1(MULT_mult_6_SUMB_2__15_), .A2(
        MULT_mult_6_n1186), .ZN(MULT_mult_6_n1989) );
  INV_X2 MULT_mult_6_U747 ( .A(MULT_mult_6_net80409), .ZN(MULT_mult_6_n341) );
  INV_X4 MULT_mult_6_U746 ( .A(MULT_mult_6_n341), .ZN(MULT_mult_6_n242) );
  INV_X1 MULT_mult_6_U745 ( .A(MULT_mult_6_n852), .ZN(MULT_mult_6_n239) );
  NAND2_X2 MULT_mult_6_U744 ( .A1(MULT_mult_6_n240), .A2(MULT_mult_6_n241), 
        .ZN(MULT_mult_6_SUMB_4__17_) );
  NAND2_X2 MULT_mult_6_U743 ( .A1(MULT_mult_6_n238), .A2(MULT_mult_6_n239), 
        .ZN(MULT_mult_6_n241) );
  NAND2_X1 MULT_mult_6_U742 ( .A1(MULT_mult_6_SUMB_5__18_), .A2(
        MULT_mult_6_n1490), .ZN(MULT_mult_6_n2245) );
  CLKBUF_X3 MULT_mult_6_U741 ( .A(MULT_mult_6_SUMB_1__15_), .Z(
        MULT_mult_6_net93243) );
  INV_X16 MULT_mult_6_U740 ( .A(n10917), .ZN(MULT_mult_6_net87396) );
  INV_X16 MULT_mult_6_U739 ( .A(MULT_mult_6_net80392), .ZN(
        MULT_mult_6_net81673) );
  NAND2_X4 MULT_mult_6_U738 ( .A1(MULT_mult_6_n1211), .A2(
        MULT_mult_6_SUMB_14__5_), .ZN(MULT_mult_6_n1707) );
  NAND2_X2 MULT_mult_6_U737 ( .A1(MULT_mult_6_ab_4__7_), .A2(
        MULT_mult_6_SUMB_3__8_), .ZN(MULT_mult_6_n1909) );
  NAND2_X4 MULT_mult_6_U736 ( .A1(MULT_mult_6_CARRYB_23__0_), .A2(
        MULT_mult_6_ab_24__0_), .ZN(MULT_mult_6_n1569) );
  NAND2_X4 MULT_mult_6_U735 ( .A1(MULT_mult_6_n940), .A2(MULT_mult_6_ab_26__0_), .ZN(MULT_mult_6_net81533) );
  NAND2_X4 MULT_mult_6_U734 ( .A1(MULT_mult_6_ab_22__4_), .A2(
        MULT_mult_6_net86464), .ZN(MULT_mult_6_net79992) );
  INV_X2 MULT_mult_6_U733 ( .A(n5851), .ZN(MULT_mult_6_net89652) );
  NAND2_X2 MULT_mult_6_U732 ( .A1(MULT_mult_6_ab_10__9_), .A2(
        MULT_mult_6_SUMB_9__10_), .ZN(MULT_mult_6_n471) );
  INV_X2 MULT_mult_6_U731 ( .A(MULT_mult_6_net88123), .ZN(
        MULT_mult_6_net123429) );
  NAND2_X2 MULT_mult_6_U730 ( .A1(MULT_mult_6_n869), .A2(MULT_mult_6_net83134), 
        .ZN(MULT_mult_6_net86704) );
  NAND2_X4 MULT_mult_6_U729 ( .A1(MULT_mult_6_SUMB_11__10_), .A2(
        MULT_mult_6_ab_12__9_), .ZN(MULT_mult_6_net88296) );
  NAND2_X4 MULT_mult_6_U728 ( .A1(MULT_mult_6_net91301), .A2(
        MULT_mult_6_ab_13__8_), .ZN(MULT_mult_6_net80506) );
  INV_X8 MULT_mult_6_U727 ( .A(MULT_mult_6_n1230), .ZN(MULT_mult_6_SUMB_9__9_)
         );
  XNOR2_X1 MULT_mult_6_U726 ( .A(MULT_mult_6_net81581), .B(
        MULT_mult_6_net120922), .ZN(MULT_mult_6_n941) );
  INV_X4 MULT_mult_6_U725 ( .A(MULT_mult_6_n1618), .ZN(MULT_mult_6_n234) );
  INV_X4 MULT_mult_6_U724 ( .A(MULT_mult_6_n941), .ZN(MULT_mult_6_n233) );
  NAND2_X4 MULT_mult_6_U723 ( .A1(MULT_mult_6_n235), .A2(MULT_mult_6_n236), 
        .ZN(MULT_mult_6_n1230) );
  NAND2_X4 MULT_mult_6_U722 ( .A1(MULT_mult_6_n233), .A2(MULT_mult_6_n234), 
        .ZN(MULT_mult_6_n236) );
  NAND2_X2 MULT_mult_6_U721 ( .A1(MULT_mult_6_n941), .A2(MULT_mult_6_n1618), 
        .ZN(MULT_mult_6_n235) );
  INV_X2 MULT_mult_6_U720 ( .A(MULT_mult_6_net93800), .ZN(MULT_mult_6_n230) );
  NAND2_X2 MULT_mult_6_U719 ( .A1(MULT_mult_6_n231), .A2(MULT_mult_6_n232), 
        .ZN(MULT_mult_6_SUMB_7__14_) );
  NAND2_X1 MULT_mult_6_U718 ( .A1(MULT_mult_6_n797), .A2(MULT_mult_6_net93800), 
        .ZN(MULT_mult_6_n231) );
  INV_X8 MULT_mult_6_U717 ( .A(MULT_mult_6_CARRYB_8__11_), .ZN(
        MULT_mult_6_net86893) );
  NAND2_X4 MULT_mult_6_U715 ( .A1(MULT_mult_6_n1684), .A2(MULT_mult_6_n1685), 
        .ZN(MULT_mult_6_SUMB_2__20_) );
  NAND2_X4 MULT_mult_6_U714 ( .A1(MULT_mult_6_net83061), .A2(
        MULT_mult_6_ab_10__10_), .ZN(MULT_mult_6_n458) );
  NOR2_X2 MULT_mult_6_U713 ( .A1(MULT_mult_6_net82239), .A2(MULT_mult_6_n175), 
        .ZN(MULT_mult_6_ab_2__25_) );
  NAND2_X4 MULT_mult_6_U712 ( .A1(MULT_mult_6_n1343), .A2(MULT_mult_6_n1344), 
        .ZN(MULT_mult_6_net82024) );
  NAND2_X4 MULT_mult_6_U711 ( .A1(MULT_mult_6_net87682), .A2(
        MULT_mult_6_net87683), .ZN(MULT_mult_6_n1344) );
  INV_X4 MULT_mult_6_U710 ( .A(MULT_mult_6_n2095), .ZN(MULT_mult_6_n1725) );
  NOR2_X2 MULT_mult_6_U709 ( .A1(MULT_mult_6_net70470), .A2(
        MULT_mult_6_net86101), .ZN(MULT_mult_6_n401) );
  INV_X4 MULT_mult_6_U708 ( .A(MULT_mult_6_SUMB_13__7_), .ZN(MULT_mult_6_n1308) );
  INV_X1 MULT_mult_6_U707 ( .A(MULT_mult_6_n1308), .ZN(MULT_mult_6_n225) );
  INV_X2 MULT_mult_6_U706 ( .A(MULT_mult_6_n1973), .ZN(MULT_mult_6_n224) );
  NAND2_X4 MULT_mult_6_U705 ( .A1(MULT_mult_6_n226), .A2(MULT_mult_6_n227), 
        .ZN(MULT_mult_6_n864) );
  INV_X1 MULT_mult_6_U702 ( .A(MULT_mult_6_n2001), .ZN(MULT_mult_6_n220) );
  NAND2_X2 MULT_mult_6_U701 ( .A1(MULT_mult_6_n222), .A2(MULT_mult_6_n223), 
        .ZN(MULT_mult_6_SUMB_8__8_) );
  NAND2_X2 MULT_mult_6_U700 ( .A1(MULT_mult_6_n220), .A2(MULT_mult_6_n939), 
        .ZN(MULT_mult_6_n223) );
  NAND2_X1 MULT_mult_6_U699 ( .A1(MULT_mult_6_n221), .A2(MULT_mult_6_n2001), 
        .ZN(MULT_mult_6_n222) );
  XNOR2_X2 MULT_mult_6_U698 ( .A(MULT_mult_6_n11), .B(MULT_mult_6_n1270), .ZN(
        MULT_mult_6_n1189) );
  NAND2_X4 MULT_mult_6_U697 ( .A1(MULT_mult_6_SUMB_12__6_), .A2(
        MULT_mult_6_ab_13__5_), .ZN(MULT_mult_6_n1921) );
  INV_X1 MULT_mult_6_U696 ( .A(MULT_mult_6_n1189), .ZN(MULT_mult_6_n217) );
  INV_X4 MULT_mult_6_U695 ( .A(MULT_mult_6_n569), .ZN(MULT_mult_6_n216) );
  NAND2_X4 MULT_mult_6_U694 ( .A1(MULT_mult_6_n218), .A2(MULT_mult_6_n219), 
        .ZN(MULT_mult_6_n1209) );
  NAND2_X2 MULT_mult_6_U692 ( .A1(MULT_mult_6_net92724), .A2(
        MULT_mult_6__UDW__112694_net78575), .ZN(MULT_mult_6_n1163) );
  NAND2_X2 MULT_mult_6_U691 ( .A1(MULT_mult_6_n1604), .A2(MULT_mult_6_n1605), 
        .ZN(MULT_mult_6_SUMB_7__17_) );
  NAND2_X4 MULT_mult_6_U690 ( .A1(MULT_mult_6_n1604), .A2(MULT_mult_6_n1605), 
        .ZN(MULT_mult_6_n215) );
  NAND2_X2 MULT_mult_6_U689 ( .A1(MULT_mult_6_n857), .A2(MULT_mult_6_n910), 
        .ZN(MULT_mult_6_n912) );
  NOR2_X4 MULT_mult_6_U688 ( .A1(MULT_mult_6_net70460), .A2(
        MULT_mult_6_net119855), .ZN(MULT_mult_6_ab_4__13_) );
  NAND2_X2 MULT_mult_6_U687 ( .A1(MULT_mult_6_n1507), .A2(MULT_mult_6_n1508), 
        .ZN(MULT_mult_6_SUMB_13__10_) );
  INV_X1 MULT_mult_6_U686 ( .A(MULT_mult_6_ab_4__13_), .ZN(MULT_mult_6_n212)
         );
  INV_X2 MULT_mult_6_U685 ( .A(MULT_mult_6_CARRYB_3__13_), .ZN(
        MULT_mult_6_n211) );
  NAND2_X2 MULT_mult_6_U683 ( .A1(MULT_mult_6_n211), .A2(MULT_mult_6_ab_4__13_), .ZN(MULT_mult_6_n214) );
  NAND2_X4 MULT_mult_6_U681 ( .A1(MULT_mult_6_n1507), .A2(MULT_mult_6_n1508), 
        .ZN(MULT_mult_6_n210) );
  NAND2_X4 MULT_mult_6_U680 ( .A1(MULT_mult_6_n45), .A2(MULT_mult_6_n316), 
        .ZN(MULT_mult_6_n318) );
  OR2_X2 MULT_mult_6_U679 ( .A1(MULT_mult_6_n2361), .A2(MULT_mult_6_n2359), 
        .ZN(MULT_mult_6_n209) );
  NAND3_X2 MULT_mult_6_U678 ( .A1(MULT_mult_6_n2115), .A2(MULT_mult_6_n2114), 
        .A3(MULT_mult_6_n2113), .ZN(MULT_mult_6_CARRYB_25__4_) );
  BUF_X4 MULT_mult_6_U677 ( .A(MULT_mult_6_SUMB_3__13_), .Z(
        MULT_mult_6_net85493) );
  NAND2_X4 MULT_mult_6_U676 ( .A1(MULT_mult_6_SUMB_3__13_), .A2(
        MULT_mult_6_ab_4__12_), .ZN(MULT_mult_6_net82759) );
  INV_X2 MULT_mult_6_U675 ( .A(MULT_mult_6_ab_11__10_), .ZN(
        MULT_mult_6_net87045) );
  INV_X8 MULT_mult_6_U674 ( .A(MULT_mult_6_net122062), .ZN(MULT_mult_6_n299)
         );
  INV_X4 MULT_mult_6_U673 ( .A(MULT_mult_6_net84270), .ZN(MULT_mult_6_n206) );
  NAND2_X4 MULT_mult_6_U671 ( .A1(MULT_mult_6_n208), .A2(MULT_mult_6_n207), 
        .ZN(MULT_mult_6_SUMB_3__13_) );
  NAND2_X4 MULT_mult_6_U670 ( .A1(MULT_mult_6_n2366), .A2(MULT_mult_6_n206), 
        .ZN(MULT_mult_6_n208) );
  NAND2_X2 MULT_mult_6_U669 ( .A1(MULT_mult_6_net81694), .A2(
        MULT_mult_6_net84270), .ZN(MULT_mult_6_n207) );
  INV_X1 MULT_mult_6_U668 ( .A(MULT_mult_6_net87045), .ZN(MULT_mult_6_n202) );
  NAND2_X2 MULT_mult_6_U667 ( .A1(MULT_mult_6_n203), .A2(MULT_mult_6_n204), 
        .ZN(MULT_mult_6_net85732) );
  NAND2_X2 MULT_mult_6_U666 ( .A1(MULT_mult_6_n201), .A2(MULT_mult_6_n202), 
        .ZN(MULT_mult_6_n204) );
  NAND2_X2 MULT_mult_6_U665 ( .A1(MULT_mult_6_CARRYB_10__10_), .A2(
        MULT_mult_6_net87045), .ZN(MULT_mult_6_n203) );
  INV_X2 MULT_mult_6_U664 ( .A(MULT_mult_6_SUMB_1__18_), .ZN(MULT_mult_6_n538)
         );
  NAND2_X4 MULT_mult_6_U663 ( .A1(MULT_mult_6_n537), .A2(MULT_mult_6_n538), 
        .ZN(MULT_mult_6_n540) );
  NAND2_X4 MULT_mult_6_U662 ( .A1(MULT_mult_6_n1193), .A2(
        MULT_mult_6_ab_12__6_), .ZN(MULT_mult_6_n1917) );
  XNOR2_X1 MULT_mult_6_U661 ( .A(MULT_mult_6_CARRYB_1__13_), .B(
        MULT_mult_6_ab_2__13_), .ZN(MULT_mult_6_net124618) );
  INV_X2 MULT_mult_6_U660 ( .A(MULT_mult_6_CARRYB_4__11_), .ZN(
        MULT_mult_6_net147920) );
  INV_X8 MULT_mult_6_U659 ( .A(MULT_mult_6_CARRYB_8__8_), .ZN(
        MULT_mult_6_n1177) );
  NAND2_X4 MULT_mult_6_U657 ( .A1(MULT_mult_6_n532), .A2(MULT_mult_6_net85096), 
        .ZN(MULT_mult_6_net81158) );
  INV_X8 MULT_mult_6_U656 ( .A(MULT_mult_6_net82544), .ZN(
        MULT_mult_6_net121449) );
  NAND2_X2 MULT_mult_6_U655 ( .A1(MULT_mult_6_net121450), .A2(
        MULT_mult_6_net121449), .ZN(MULT_mult_6_net121452) );
  NAND2_X4 MULT_mult_6_U654 ( .A1(MULT_mult_6_net121449), .A2(
        MULT_mult_6_net121450), .ZN(MULT_mult_6_n199) );
  NAND2_X2 MULT_mult_6_U653 ( .A1(MULT_mult_6_n549), .A2(
        MULT_mult_6_SUMB_17__8_), .ZN(MULT_mult_6_n309) );
  NAND2_X4 MULT_mult_6_U652 ( .A1(MULT_mult_6_n643), .A2(MULT_mult_6_n644), 
        .ZN(MULT_mult_6_net88699) );
  NAND2_X2 MULT_mult_6_U651 ( .A1(MULT_mult_6_CARRYB_20__8_), .A2(
        MULT_mult_6_n859), .ZN(MULT_mult_6_net81038) );
  NAND3_X4 MULT_mult_6_U650 ( .A1(MULT_mult_6_net81038), .A2(
        MULT_mult_6_net81037), .A3(MULT_mult_6_net81036), .ZN(
        MULT_mult_6_CARRYB_21__8_) );
  NAND2_X1 MULT_mult_6_U649 ( .A1(MULT_mult_6_ab_12__17_), .A2(
        MULT_mult_6_SUMB_11__18_), .ZN(MULT_mult_6_n1468) );
  NAND2_X2 MULT_mult_6_U648 ( .A1(MULT_mult_6_net123142), .A2(MULT_mult_6_n299), .ZN(MULT_mult_6_n301) );
  INV_X4 MULT_mult_6_U647 ( .A(MULT_mult_6_n950), .ZN(MULT_mult_6_n196) );
  INV_X4 MULT_mult_6_U646 ( .A(MULT_mult_6_n2015), .ZN(MULT_mult_6_n195) );
  NAND2_X2 MULT_mult_6_U645 ( .A1(MULT_mult_6_n2015), .A2(MULT_mult_6_n950), 
        .ZN(MULT_mult_6_n197) );
  NAND2_X4 MULT_mult_6_U644 ( .A1(MULT_mult_6_n594), .A2(MULT_mult_6_n595), 
        .ZN(MULT_mult_6_SUMB_11__4_) );
  XNOR2_X2 MULT_mult_6_U643 ( .A(MULT_mult_6_net88776), .B(
        MULT_mult_6_net85903), .ZN(MULT_mult_6_SUMB_24__1_) );
  BUF_X8 MULT_mult_6_U642 ( .A(MULT_mult_6_SUMB_10__8_), .Z(MULT_mult_6_n1249)
         );
  XNOR2_X2 MULT_mult_6_U641 ( .A(MULT_mult_6_SUMB_9__7_), .B(MULT_mult_6_n996), 
        .ZN(MULT_mult_6_n194) );
  INV_X4 MULT_mult_6_U640 ( .A(MULT_mult_6_net121450), .ZN(
        MULT_mult_6_net121770) );
  INV_X4 MULT_mult_6_U638 ( .A(MULT_mult_6_n193), .ZN(MULT_mult_6_net121814)
         );
  INV_X4 MULT_mult_6_U636 ( .A(MULT_mult_6_n1429), .ZN(MULT_mult_6_n288) );
  XNOR2_X2 MULT_mult_6_U635 ( .A(MULT_mult_6_n192), .B(MULT_mult_6_SUMB_26__1_), .ZN(multOut[4]) );
  XNOR2_X2 MULT_mult_6_U634 ( .A(MULT_mult_6_n417), .B(MULT_mult_6_net85109), 
        .ZN(MULT_mult_6_n364) );
  NAND2_X4 MULT_mult_6_U632 ( .A1(MULT_mult_6_net87938), .A2(
        MULT_mult_6_net87939), .ZN(MULT_mult_6_net87941) );
  NAND2_X2 MULT_mult_6_U631 ( .A1(MULT_mult_6_SUMB_9__9_), .A2(
        MULT_mult_6_CARRYB_9__8_), .ZN(MULT_mult_6_n1776) );
  INV_X2 MULT_mult_6_U630 ( .A(MULT_mult_6_SUMB_11__11_), .ZN(
        MULT_mult_6_net89840) );
  INV_X4 MULT_mult_6_U629 ( .A(MULT_mult_6_n290), .ZN(MULT_mult_6_n1134) );
  INV_X2 MULT_mult_6_U627 ( .A(MULT_mult_6_SUMB_15__10_), .ZN(MULT_mult_6_n189) );
  INV_X4 MULT_mult_6_U626 ( .A(MULT_mult_6_net81992), .ZN(MULT_mult_6_n188) );
  NAND2_X4 MULT_mult_6_U625 ( .A1(MULT_mult_6_n190), .A2(MULT_mult_6_n191), 
        .ZN(MULT_mult_6_SUMB_16__9_) );
  NAND2_X2 MULT_mult_6_U624 ( .A1(MULT_mult_6_n188), .A2(MULT_mult_6_n189), 
        .ZN(MULT_mult_6_n191) );
  NAND2_X1 MULT_mult_6_U623 ( .A1(MULT_mult_6_net81992), .A2(
        MULT_mult_6_SUMB_15__10_), .ZN(MULT_mult_6_n190) );
  NAND2_X4 MULT_mult_6_U622 ( .A1(MULT_mult_6_net90022), .A2(
        MULT_mult_6_net90818), .ZN(MULT_mult_6_net87950) );
  INV_X1 MULT_mult_6_U621 ( .A(MULT_mult_6_ab_3__10_), .ZN(MULT_mult_6_n185)
         );
  INV_X4 MULT_mult_6_U620 ( .A(MULT_mult_6_CARRYB_2__10_), .ZN(
        MULT_mult_6_n184) );
  NAND2_X4 MULT_mult_6_U619 ( .A1(MULT_mult_6_n186), .A2(MULT_mult_6_n187), 
        .ZN(MULT_mult_6_n1399) );
  NAND2_X2 MULT_mult_6_U618 ( .A1(MULT_mult_6_n184), .A2(MULT_mult_6_n185), 
        .ZN(MULT_mult_6_n187) );
  NAND2_X4 MULT_mult_6_U616 ( .A1(MULT_mult_6_net147939), .A2(
        MULT_mult_6_net147940), .ZN(MULT_mult_6_SUMB_24__2_) );
  NAND2_X4 MULT_mult_6_U615 ( .A1(MULT_mult_6_net123293), .A2(MULT_mult_6_n776), .ZN(MULT_mult_6_net93683) );
  NAND2_X4 MULT_mult_6_U614 ( .A1(MULT_mult_6_ab_14__4_), .A2(
        MULT_mult_6_CARRYB_13__4_), .ZN(MULT_mult_6_n2152) );
  NAND2_X4 MULT_mult_6_U613 ( .A1(MULT_mult_6_net85808), .A2(
        MULT_mult_6_net84208), .ZN(MULT_mult_6_net87945) );
  NAND2_X2 MULT_mult_6_U612 ( .A1(MULT_mult_6_n1486), .A2(MULT_mult_6_n1487), 
        .ZN(MULT_mult_6_n1489) );
  NAND2_X4 MULT_mult_6_U611 ( .A1(MULT_mult_6_n1768), .A2(
        MULT_mult_6_SUMB_4__19_), .ZN(MULT_mult_6_n2141) );
  INV_X1 MULT_mult_6_U610 ( .A(MULT_mult_6_SUMB_3__20_), .ZN(MULT_mult_6_n1420) );
  NAND2_X1 MULT_mult_6_U609 ( .A1(MULT_mult_6_CARRYB_17__11_), .A2(
        MULT_mult_6_net88647), .ZN(MULT_mult_6_net82666) );
  INV_X8 MULT_mult_6_U608 ( .A(MULT_mult_6_net90735), .ZN(
        MULT_mult_6_net121445) );
  INV_X2 MULT_mult_6_U607 ( .A(MULT_mult_6_net121445), .ZN(MULT_mult_6_n183)
         );
  BUF_X8 MULT_mult_6_U606 ( .A(MULT_mult_6_net70470), .Z(MULT_mult_6_n182) );
  BUF_X4 MULT_mult_6_U605 ( .A(MULT_mult_6_SUMB_3__12_), .Z(
        MULT_mult_6_net121785) );
  BUF_X8 MULT_mult_6_U604 ( .A(MULT_mult_6_SUMB_11__7_), .Z(MULT_mult_6_n371)
         );
  XNOR2_X2 MULT_mult_6_U603 ( .A(MULT_mult_6_net121785), .B(MULT_mult_6_n1311), 
        .ZN(MULT_mult_6_n181) );
  INV_X2 MULT_mult_6_U602 ( .A(MULT_mult_6_n558), .ZN(MULT_mult_6_n178) );
  INV_X4 MULT_mult_6_U601 ( .A(MULT_mult_6_n1199), .ZN(MULT_mult_6_n177) );
  NAND2_X4 MULT_mult_6_U600 ( .A1(MULT_mult_6_n179), .A2(MULT_mult_6_n180), 
        .ZN(MULT_mult_6_SUMB_3__11_) );
  NAND2_X4 MULT_mult_6_U599 ( .A1(MULT_mult_6_n177), .A2(MULT_mult_6_n178), 
        .ZN(MULT_mult_6_n180) );
  NAND2_X2 MULT_mult_6_U598 ( .A1(MULT_mult_6_n1199), .A2(MULT_mult_6_n558), 
        .ZN(MULT_mult_6_n179) );
  NAND2_X2 MULT_mult_6_U597 ( .A1(MULT_mult_6_CARRYB_16__9_), .A2(
        MULT_mult_6_ab_17__9_), .ZN(MULT_mult_6_net120657) );
  NAND2_X4 MULT_mult_6_U596 ( .A1(MULT_mult_6_net123291), .A2(MULT_mult_6_n775), .ZN(MULT_mult_6_n776) );
  XNOR2_X2 MULT_mult_6_U595 ( .A(MULT_mult_6_CARRYB_13__11_), .B(
        MULT_mult_6_ab_14__11_), .ZN(MULT_mult_6_net125934) );
  NAND2_X4 MULT_mult_6_U594 ( .A1(MULT_mult_6_ab_9__9_), .A2(
        MULT_mult_6_CARRYB_8__9_), .ZN(MULT_mult_6_n1621) );
  NOR2_X4 MULT_mult_6_U593 ( .A1(MULT_mult_6_n392), .A2(MULT_mult_6_n2354), 
        .ZN(MULT_mult_6_ab_0__28_) );
  NOR2_X4 MULT_mult_6_U592 ( .A1(MULT_mult_6_n2355), .A2(MULT_mult_6_n242), 
        .ZN(MULT_mult_6_ab_1__27_) );
  NAND2_X2 MULT_mult_6_U591 ( .A1(MULT_mult_6_n319), .A2(MULT_mult_6_n320), 
        .ZN(MULT_mult_6_n322) );
  NAND2_X2 MULT_mult_6_U590 ( .A1(MULT_mult_6_ab_2__23_), .A2(
        MULT_mult_6_n2357), .ZN(MULT_mult_6_net83575) );
  NAND2_X2 MULT_mult_6_U589 ( .A1(MULT_mult_6_net82124), .A2(
        MULT_mult_6_net83044), .ZN(MULT_mult_6_net83576) );
  INV_X8 MULT_mult_6_U588 ( .A(MULT_mult_6_ab_0__24_), .ZN(
        MULT_mult_6_net82044) );
  INV_X4 MULT_mult_6_U587 ( .A(MULT_mult_6_net83919), .ZN(MULT_mult_6_net93203) );
  INV_X4 MULT_mult_6_U586 ( .A(MULT_mult_6_net93203), .ZN(MULT_mult_6_n174) );
  NAND2_X4 MULT_mult_6_U585 ( .A1(MULT_mult_6_net84868), .A2(
        MULT_mult_6_net84867), .ZN(MULT_mult_6_net84870) );
  BUF_X4 MULT_mult_6_U584 ( .A(MULT_mult_6_CARRYB_27__0_), .Z(MULT_mult_6_n284) );
  INV_X2 MULT_mult_6_U583 ( .A(MULT_mult_6_ab_0__12_), .ZN(
        MULT_mult_6_net120501) );
  AND2_X2 MULT_mult_6_U582 ( .A1(n10920), .A2(n6007), .ZN(
        MULT_mult_6_ab_3__10_) );
  NAND2_X4 MULT_mult_6_U581 ( .A1(MULT_mult_6_CARRYB_7__6_), .A2(
        MULT_mult_6_SUMB_7__7_), .ZN(MULT_mult_6_n1827) );
  NAND2_X2 MULT_mult_6_U580 ( .A1(MULT_mult_6_n569), .A2(MULT_mult_6_n1189), 
        .ZN(MULT_mult_6_n218) );
  NAND2_X4 MULT_mult_6_U578 ( .A1(MULT_mult_6_n195), .A2(MULT_mult_6_n196), 
        .ZN(MULT_mult_6_n198) );
  NAND2_X4 MULT_mult_6_U577 ( .A1(MULT_mult_6_n198), .A2(MULT_mult_6_n197), 
        .ZN(MULT_mult_6_SUMB_9__8_) );
  NAND2_X2 MULT_mult_6_U576 ( .A1(MULT_mult_6_ab_30__0_), .A2(
        MULT_mult_6_net87797), .ZN(MULT_mult_6_net80474) );
  NAND2_X4 MULT_mult_6_U575 ( .A1(MULT_mult_6_ab_9__13_), .A2(
        MULT_mult_6_SUMB_8__14_), .ZN(MULT_mult_6_net80349) );
  NOR2_X2 MULT_mult_6_U574 ( .A1(MULT_mult_6_net123000), .A2(
        MULT_mult_6_net82247), .ZN(MULT_mult_6_net88449) );
  INV_X1 MULT_mult_6_U573 ( .A(MULT_mult_6_n1611), .ZN(MULT_mult_6_n1368) );
  XNOR2_X2 MULT_mult_6_U572 ( .A(MULT_mult_6_CARRYB_3__13_), .B(
        MULT_mult_6_ab_4__13_), .ZN(MULT_mult_6_n1562) );
  NAND2_X4 MULT_mult_6_U571 ( .A1(MULT_mult_6_n1362), .A2(MULT_mult_6_net86440), .ZN(MULT_mult_6_n1418) );
  INV_X4 MULT_mult_6_U570 ( .A(MULT_mult_6_n91), .ZN(MULT_mult_6_n578) );
  NOR2_X4 MULT_mult_6_U568 ( .A1(MULT_mult_6_net70470), .A2(
        MULT_mult_6_net86101), .ZN(MULT_mult_6_ab_1__18_) );
  INV_X4 MULT_mult_6_U567 ( .A(MULT_mult_6_net87363), .ZN(
        MULT_mult_6_net148828) );
  INV_X8 MULT_mult_6_U566 ( .A(MULT_mult_6_net85035), .ZN(MULT_mult_6_net85036) );
  INV_X4 MULT_mult_6_U565 ( .A(MULT_mult_6_n172), .ZN(MULT_mult_6_n173) );
  INV_X2 MULT_mult_6_U564 ( .A(MULT_mult_6_CARRYB_10__7_), .ZN(
        MULT_mult_6_n172) );
  NAND3_X2 MULT_mult_6_U563 ( .A1(MULT_mult_6_n651), .A2(MULT_mult_6_n652), 
        .A3(MULT_mult_6_n653), .ZN(MULT_mult_6_CARRYB_15__1_) );
  BUF_X16 MULT_mult_6_U562 ( .A(MULT_mult_6_net70454), .Z(MULT_mult_6_net91660) );
  NOR2_X1 MULT_mult_6_U561 ( .A1(MULT_mult_6_net70454), .A2(
        MULT_mult_6_net77938), .ZN(MULT_mult_6_ab_6__10_) );
  INV_X2 MULT_mult_6_U560 ( .A(MULT_mult_6_SUMB_16__4_), .ZN(MULT_mult_6_n560)
         );
  NAND2_X4 MULT_mult_6_U559 ( .A1(MULT_mult_6_SUMB_23__2_), .A2(
        MULT_mult_6_ab_24__1_), .ZN(MULT_mult_6_net80921) );
  INV_X2 MULT_mult_6_U558 ( .A(MULT_mult_6_CARRYB_2__9_), .ZN(
        MULT_mult_6_n1245) );
  NAND2_X4 MULT_mult_6_U557 ( .A1(MULT_mult_6_CARRYB_14__9_), .A2(
        MULT_mult_6_ab_15__9_), .ZN(MULT_mult_6_net84817) );
  NOR2_X2 MULT_mult_6_U556 ( .A1(MULT_mult_6_net70456), .A2(
        MULT_mult_6_net77966), .ZN(MULT_mult_6_ab_3__11_) );
  INV_X4 MULT_mult_6_U555 ( .A(MULT_mult_6_net81158), .ZN(MULT_mult_6_n200) );
  XNOR2_X2 MULT_mult_6_U554 ( .A(MULT_mult_6_SUMB_23__8_), .B(
        MULT_mult_6_n1084), .ZN(MULT_mult_6_n171) );
  XNOR2_X2 MULT_mult_6_U553 ( .A(MULT_mult_6_n171), .B(MULT_mult_6_n1083), 
        .ZN(MULT_mult_6_n170) );
  NAND2_X2 MULT_mult_6_U552 ( .A1(MULT_mult_6_net121445), .A2(
        MULT_mult_6_net121446), .ZN(MULT_mult_6_n466) );
  NAND3_X4 MULT_mult_6_U551 ( .A1(MULT_mult_6_net84312), .A2(
        MULT_mult_6_net84313), .A3(MULT_mult_6_n1057), .ZN(
        MULT_mult_6_CARRYB_4__22_) );
  NAND2_X2 MULT_mult_6_U550 ( .A1(MULT_mult_6_SUMB_25__5_), .A2(
        MULT_mult_6_ab_26__4_), .ZN(MULT_mult_6_n1080) );
  INV_X4 MULT_mult_6_U549 ( .A(MULT_mult_6_net89109), .ZN(MULT_mult_6_net85287) );
  NAND3_X2 MULT_mult_6_U548 ( .A1(MULT_mult_6_net80925), .A2(
        MULT_mult_6_net80924), .A3(MULT_mult_6_net80926), .ZN(
        MULT_mult_6_CARRYB_22__2_) );
  NOR2_X2 MULT_mult_6_U547 ( .A1(MULT_mult_6_net77866), .A2(
        MULT_mult_6_net70447), .ZN(MULT_mult_6_ab_24__1_) );
  INV_X8 MULT_mult_6_U546 ( .A(MULT_mult_6_n1994), .ZN(MULT_mult_6_n1001) );
  NOR2_X4 MULT_mult_6_U545 ( .A1(MULT_mult_6_net77920), .A2(
        MULT_mult_6_net77938), .ZN(MULT_mult_6_ab_6__8_) );
  INV_X1 MULT_mult_6_U544 ( .A(MULT_mult_6_ab_24__1_), .ZN(MULT_mult_6_n167)
         );
  INV_X4 MULT_mult_6_U543 ( .A(MULT_mult_6_n398), .ZN(MULT_mult_6_n166) );
  NAND2_X4 MULT_mult_6_U542 ( .A1(MULT_mult_6_n168), .A2(MULT_mult_6_n169), 
        .ZN(MULT_mult_6_net88776) );
  NAND2_X4 MULT_mult_6_U541 ( .A1(MULT_mult_6_n166), .A2(MULT_mult_6_n167), 
        .ZN(MULT_mult_6_n169) );
  NAND2_X1 MULT_mult_6_U540 ( .A1(MULT_mult_6_n398), .A2(MULT_mult_6_ab_24__1_), .ZN(MULT_mult_6_n168) );
  NAND3_X2 MULT_mult_6_U539 ( .A1(MULT_mult_6_n1822), .A2(MULT_mult_6_n1823), 
        .A3(MULT_mult_6_n1824), .ZN(MULT_mult_6_n165) );
  INV_X4 MULT_mult_6_U538 ( .A(MULT_mult_6_ab_6__8_), .ZN(MULT_mult_6_n162) );
  INV_X2 MULT_mult_6_U537 ( .A(MULT_mult_6_CARRYB_5__8_), .ZN(MULT_mult_6_n161) );
  NAND2_X4 MULT_mult_6_U536 ( .A1(MULT_mult_6_n163), .A2(MULT_mult_6_n164), 
        .ZN(MULT_mult_6_n1994) );
  NAND2_X4 MULT_mult_6_U535 ( .A1(MULT_mult_6_n161), .A2(MULT_mult_6_n162), 
        .ZN(MULT_mult_6_n164) );
  NAND2_X1 MULT_mult_6_U534 ( .A1(MULT_mult_6_n2377), .A2(MULT_mult_6_ab_6__8_), .ZN(MULT_mult_6_n163) );
  NAND2_X4 MULT_mult_6_U533 ( .A1(MULT_mult_6_n256), .A2(MULT_mult_6_n257), 
        .ZN(MULT_mult_6_n259) );
  NAND2_X4 MULT_mult_6_U532 ( .A1(MULT_mult_6_ab_2__10_), .A2(
        MULT_mult_6_SUMB_1__11_), .ZN(MULT_mult_6_n1653) );
  INV_X4 MULT_mult_6_U531 ( .A(MULT_mult_6_n549), .ZN(MULT_mult_6_n307) );
  INV_X8 MULT_mult_6_U530 ( .A(MULT_mult_6_net119955), .ZN(
        MULT_mult_6_net148836) );
  NAND2_X4 MULT_mult_6_U529 ( .A1(MULT_mult_6_n243), .A2(MULT_mult_6_n244), 
        .ZN(MULT_mult_6_n246) );
  NAND2_X2 MULT_mult_6_U528 ( .A1(MULT_mult_6_SUMB_6__6_), .A2(
        MULT_mult_6_ab_7__5_), .ZN(MULT_mult_6_n1521) );
  NAND2_X2 MULT_mult_6_U527 ( .A1(MULT_mult_6_ab_9__4_), .A2(
        MULT_mult_6_CARRYB_8__4_), .ZN(MULT_mult_6_net82099) );
  NOR2_X1 MULT_mult_6_U526 ( .A1(MULT_mult_6_net77892), .A2(
        MULT_mult_6_net77924), .ZN(MULT_mult_6_ab_8__4_) );
  INV_X1 MULT_mult_6_U525 ( .A(MULT_mult_6_SUMB_5__7_), .ZN(MULT_mult_6_n158)
         );
  INV_X4 MULT_mult_6_U524 ( .A(MULT_mult_6_n1552), .ZN(MULT_mult_6_n157) );
  NAND2_X4 MULT_mult_6_U523 ( .A1(MULT_mult_6_n159), .A2(MULT_mult_6_n160), 
        .ZN(MULT_mult_6_SUMB_6__6_) );
  NAND2_X4 MULT_mult_6_U522 ( .A1(MULT_mult_6_n157), .A2(MULT_mult_6_n158), 
        .ZN(MULT_mult_6_n160) );
  NAND2_X2 MULT_mult_6_U521 ( .A1(MULT_mult_6_n1552), .A2(
        MULT_mult_6_SUMB_5__7_), .ZN(MULT_mult_6_n159) );
  NAND3_X4 MULT_mult_6_U520 ( .A1(MULT_mult_6_n154), .A2(MULT_mult_6_n155), 
        .A3(MULT_mult_6_n156), .ZN(MULT_mult_6_CARRYB_8__4_) );
  NAND2_X2 MULT_mult_6_U519 ( .A1(MULT_mult_6_ab_8__4_), .A2(
        MULT_mult_6_CARRYB_7__4_), .ZN(MULT_mult_6_n156) );
  NAND2_X2 MULT_mult_6_U518 ( .A1(MULT_mult_6_ab_8__4_), .A2(
        MULT_mult_6_SUMB_7__5_), .ZN(MULT_mult_6_n155) );
  NAND2_X2 MULT_mult_6_U517 ( .A1(MULT_mult_6_CARRYB_7__4_), .A2(
        MULT_mult_6_SUMB_7__5_), .ZN(MULT_mult_6_n154) );
  XOR2_X2 MULT_mult_6_U516 ( .A(MULT_mult_6_SUMB_7__5_), .B(MULT_mult_6_n153), 
        .Z(MULT_mult_6_SUMB_8__4_) );
  XOR2_X2 MULT_mult_6_U515 ( .A(MULT_mult_6_CARRYB_7__4_), .B(
        MULT_mult_6_ab_8__4_), .Z(MULT_mult_6_n153) );
  NAND3_X2 MULT_mult_6_U514 ( .A1(MULT_mult_6_n2025), .A2(MULT_mult_6_net81530), .A3(MULT_mult_6_net81531), .ZN(MULT_mult_6_n152) );
  NAND3_X4 MULT_mult_6_U513 ( .A1(MULT_mult_6_n1564), .A2(MULT_mult_6_n1565), 
        .A3(MULT_mult_6_n1566), .ZN(MULT_mult_6_CARRYB_6__3_) );
  INV_X8 MULT_mult_6_U512 ( .A(MULT_mult_6_net77904), .ZN(MULT_mult_6_net77898) );
  INV_X8 MULT_mult_6_U511 ( .A(MULT_mult_6_CARRYB_22__3_), .ZN(
        MULT_mult_6_n404) );
  NAND2_X2 MULT_mult_6_U510 ( .A1(MULT_mult_6_n1387), .A2(MULT_mult_6_n1388), 
        .ZN(MULT_mult_6_SUMB_8__16_) );
  NAND2_X4 MULT_mult_6_U509 ( .A1(MULT_mult_6_n1387), .A2(MULT_mult_6_n1388), 
        .ZN(MULT_mult_6_n151) );
  INV_X4 MULT_mult_6_U508 ( .A(MULT_mult_6_SUMB_6__16_), .ZN(MULT_mult_6_n1375) );
  NOR2_X2 MULT_mult_6_U507 ( .A1(MULT_mult_6_net77988), .A2(
        MULT_mult_6_net70466), .ZN(MULT_mult_6_net81416) );
  INV_X8 MULT_mult_6_U506 ( .A(MULT_mult_6_CARRYB_4__14_), .ZN(
        MULT_mult_6_net84945) );
  NAND2_X4 MULT_mult_6_U504 ( .A1(MULT_mult_6_net87457), .A2(
        MULT_mult_6_net87456), .ZN(MULT_mult_6_net87459) );
  NAND2_X2 MULT_mult_6_U503 ( .A1(MULT_mult_6_CARRYB_7__12_), .A2(
        MULT_mult_6_ab_8__12_), .ZN(MULT_mult_6_net87310) );
  INV_X1 MULT_mult_6_U502 ( .A(MULT_mult_6_ab_6__11_), .ZN(MULT_mult_6_n147)
         );
  NAND2_X4 MULT_mult_6_U501 ( .A1(MULT_mult_6_n146), .A2(MULT_mult_6_n147), 
        .ZN(MULT_mult_6_n149) );
  NAND2_X1 MULT_mult_6_U500 ( .A1(MULT_mult_6_CARRYB_5__11_), .A2(
        MULT_mult_6_ab_6__11_), .ZN(MULT_mult_6_n148) );
  NAND2_X2 MULT_mult_6_U499 ( .A1(MULT_mult_6_n1855), .A2(MULT_mult_6_n1854), 
        .ZN(MULT_mult_6_n145) );
  NAND2_X4 MULT_mult_6_U498 ( .A1(MULT_mult_6_SUMB_25__1_), .A2(
        MULT_mult_6_CARRYB_25__0_), .ZN(MULT_mult_6_net81535) );
  NOR2_X4 MULT_mult_6_U497 ( .A1(MULT_mult_6_net77912), .A2(
        MULT_mult_6_net77946), .ZN(MULT_mult_6_ab_5__7_) );
  INV_X4 MULT_mult_6_U496 ( .A(MULT_mult_6_CARRYB_4__7_), .ZN(MULT_mult_6_n142) );
  INV_X2 MULT_mult_6_U495 ( .A(MULT_mult_6_ab_5__7_), .ZN(MULT_mult_6_n141) );
  NAND2_X2 MULT_mult_6_U494 ( .A1(MULT_mult_6_n143), .A2(MULT_mult_6_n144), 
        .ZN(MULT_mult_6_n1122) );
  NAND2_X2 MULT_mult_6_U493 ( .A1(MULT_mult_6_n141), .A2(MULT_mult_6_n142), 
        .ZN(MULT_mult_6_n144) );
  BUF_X4 MULT_mult_6_U492 ( .A(MULT_mult_6_n312), .Z(MULT_mult_6_n1206) );
  NOR2_X1 MULT_mult_6_U491 ( .A1(MULT_mult_6_net77898), .A2(
        MULT_mult_6_net77924), .ZN(MULT_mult_6_ab_8__5_) );
  NAND3_X2 MULT_mult_6_U490 ( .A1(MULT_mult_6_n138), .A2(MULT_mult_6_n139), 
        .A3(MULT_mult_6_n140), .ZN(MULT_mult_6_n312) );
  NAND2_X1 MULT_mult_6_U489 ( .A1(MULT_mult_6_ab_8__5_), .A2(
        MULT_mult_6_CARRYB_7__5_), .ZN(MULT_mult_6_n140) );
  NAND2_X1 MULT_mult_6_U488 ( .A1(MULT_mult_6_ab_8__5_), .A2(MULT_mult_6_n2375), .ZN(MULT_mult_6_n139) );
  NAND2_X1 MULT_mult_6_U487 ( .A1(MULT_mult_6_CARRYB_7__5_), .A2(
        MULT_mult_6_n2375), .ZN(MULT_mult_6_n138) );
  INV_X8 MULT_mult_6_U486 ( .A(MULT_mult_6_net83866), .ZN(MULT_mult_6_net85455) );
  INV_X8 MULT_mult_6_U484 ( .A(MULT_mult_6_CARRYB_2__17_), .ZN(
        MULT_mult_6_n799) );
  INV_X8 MULT_mult_6_U483 ( .A(MULT_mult_6_n1937), .ZN(MULT_mult_6_n1506) );
  INV_X4 MULT_mult_6_U482 ( .A(MULT_mult_6_SUMB_4__16_), .ZN(
        MULT_mult_6_net86162) );
  NAND2_X4 MULT_mult_6_U481 ( .A1(MULT_mult_6_net80264), .A2(MULT_mult_6_n684), 
        .ZN(MULT_mult_6_n685) );
  NAND2_X4 MULT_mult_6_U480 ( .A1(MULT_mult_6_n72), .A2(MULT_mult_6_net87950), 
        .ZN(MULT_mult_6_net149530) );
  INV_X1 MULT_mult_6_U479 ( .A(MULT_mult_6_net83535), .ZN(MULT_mult_6_n134) );
  NAND2_X2 MULT_mult_6_U478 ( .A1(MULT_mult_6_n135), .A2(MULT_mult_6_n136), 
        .ZN(MULT_mult_6_n816) );
  NAND2_X1 MULT_mult_6_U477 ( .A1(MULT_mult_6_n133), .A2(MULT_mult_6_net83535), 
        .ZN(MULT_mult_6_n136) );
  INV_X2 MULT_mult_6_U476 ( .A(MULT_mult_6_SUMB_1__16_), .ZN(MULT_mult_6_n1352) );
  NAND2_X2 MULT_mult_6_U475 ( .A1(MULT_mult_6_CARRYB_16__11_), .A2(
        MULT_mult_6_SUMB_16__12_), .ZN(MULT_mult_6_net87011) );
  INV_X2 MULT_mult_6_U474 ( .A(MULT_mult_6_n170), .ZN(MULT_mult_6_net84978) );
  NAND2_X4 MULT_mult_6_U473 ( .A1(MULT_mult_6_ab_26__0_), .A2(MULT_mult_6_n152), .ZN(MULT_mult_6_n2027) );
  XNOR2_X2 MULT_mult_6_U472 ( .A(MULT_mult_6_n2031), .B(MULT_mult_6_n151), 
        .ZN(MULT_mult_6_n367) );
  CLKBUF_X3 MULT_mult_6_U471 ( .A(MULT_mult_6_CARRYB_9__11_), .Z(
        MULT_mult_6_net82678) );
  INV_X8 MULT_mult_6_U470 ( .A(MULT_mult_6_CARRYB_5__11_), .ZN(
        MULT_mult_6_n146) );
  NOR2_X4 MULT_mult_6_U469 ( .A1(MULT_mult_6_net77878), .A2(
        MULT_mult_6_net70445), .ZN(MULT_mult_6_ab_25__2_) );
  INV_X1 MULT_mult_6_U468 ( .A(MULT_mult_6_ab_25__2_), .ZN(MULT_mult_6_n130)
         );
  NAND2_X2 MULT_mult_6_U466 ( .A1(MULT_mult_6_n129), .A2(MULT_mult_6_n130), 
        .ZN(MULT_mult_6_n132) );
  CLKBUF_X3 MULT_mult_6_U464 ( .A(MULT_mult_6_SUMB_2__11_), .Z(
        MULT_mult_6_n128) );
  INV_X8 MULT_mult_6_U463 ( .A(MULT_mult_6_CARRYB_9__8_), .ZN(
        MULT_mult_6_n1289) );
  NAND2_X4 MULT_mult_6_U462 ( .A1(MULT_mult_6_SUMB_5__11_), .A2(
        MULT_mult_6_CARRYB_5__10_), .ZN(MULT_mult_6_n1748) );
  NAND2_X2 MULT_mult_6_U461 ( .A1(MULT_mult_6_CARRYB_2__10_), .A2(
        MULT_mult_6_ab_3__10_), .ZN(MULT_mult_6_n186) );
  NOR2_X4 MULT_mult_6_U460 ( .A1(MULT_mult_6_n955), .A2(MULT_mult_6_net70491), 
        .ZN(MULT_mult_6_ab_2__21_) );
  INV_X8 MULT_mult_6_U459 ( .A(MULT_mult_6_CARRYB_28__1_), .ZN(
        MULT_mult_6_net85094) );
  NAND2_X2 MULT_mult_6_U458 ( .A1(MULT_mult_6_SUMB_2__23_), .A2(
        MULT_mult_6_CARRYB_2__22_), .ZN(MULT_mult_6_n1070) );
  NAND2_X4 MULT_mult_6_U457 ( .A1(MULT_mult_6_net123428), .A2(
        MULT_mult_6_net123429), .ZN(MULT_mult_6_n895) );
  CLKBUF_X3 MULT_mult_6_U456 ( .A(MULT_mult_6_CARRYB_4__10_), .Z(
        MULT_mult_6_n228) );
  NAND2_X4 MULT_mult_6_U454 ( .A1(MULT_mult_6_n1533), .A2(MULT_mult_6_n1534), 
        .ZN(MULT_mult_6_n1536) );
  INV_X4 MULT_mult_6_U453 ( .A(MULT_mult_6_CARRYB_13__10_), .ZN(
        MULT_mult_6_net88408) );
  INV_X8 MULT_mult_6_U452 ( .A(MULT_mult_6_net77976), .ZN(MULT_mult_6_n175) );
  NAND2_X4 MULT_mult_6_U451 ( .A1(MULT_mult_6_n25), .A2(MULT_mult_6_ab_22__1_), 
        .ZN(MULT_mult_6_net82543) );
  INV_X4 MULT_mult_6_U450 ( .A(MULT_mult_6_CARRYB_15__5_), .ZN(
        MULT_mult_6_n1454) );
  XNOR2_X1 MULT_mult_6_U449 ( .A(MULT_mult_6_ab_1__2_), .B(
        MULT_mult_6_ab_0__3_), .ZN(MULT_mult_6_n2324) );
  XNOR2_X1 MULT_mult_6_U447 ( .A(MULT_mult_6_ab_13__1_), .B(
        MULT_mult_6_CARRYB_12__1_), .ZN(MULT_mult_6_n736) );
  NAND2_X4 MULT_mult_6_U445 ( .A1(MULT_mult_6_CARRYB_17__1_), .A2(
        MULT_mult_6_ab_18__1_), .ZN(MULT_mult_6_n746) );
  NAND2_X2 MULT_mult_6_U442 ( .A1(MULT_mult_6_net92569), .A2(
        MULT_mult_6_net88665), .ZN(MULT_mult_6_n498) );
  NAND2_X2 MULT_mult_6_U441 ( .A1(MULT_mult_6_n131), .A2(MULT_mult_6_n132), 
        .ZN(MULT_mult_6_net88665) );
  NAND2_X2 MULT_mult_6_U440 ( .A1(MULT_mult_6_CARRYB_12__12_), .A2(
        MULT_mult_6_ab_13__12_), .ZN(MULT_mult_6_n1373) );
  NAND2_X2 MULT_mult_6_U439 ( .A1(MULT_mult_6_SUMB_13__12_), .A2(
        MULT_mult_6_CARRYB_13__11_), .ZN(MULT_mult_6_net82558) );
  INV_X4 MULT_mult_6_U438 ( .A(MULT_mult_6_net87681), .ZN(MULT_mult_6_net83101) );
  INV_X8 MULT_mult_6_U437 ( .A(MULT_mult_6_net119951), .ZN(
        MULT_mult_6_net123266) );
  NAND2_X2 MULT_mult_6_U436 ( .A1(MULT_mult_6_net119928), .A2(
        MULT_mult_6_net119951), .ZN(MULT_mult_6_net123268) );
  INV_X8 MULT_mult_6_U435 ( .A(MULT_mult_6_net81354), .ZN(MULT_mult_6_n125) );
  INV_X8 MULT_mult_6_U434 ( .A(MULT_mult_6_ab_1__18_), .ZN(MULT_mult_6_n124)
         );
  NAND2_X4 MULT_mult_6_U433 ( .A1(MULT_mult_6_n127), .A2(MULT_mult_6_n126), 
        .ZN(MULT_mult_6_n536) );
  NAND2_X4 MULT_mult_6_U432 ( .A1(MULT_mult_6_n124), .A2(MULT_mult_6_n125), 
        .ZN(MULT_mult_6_n127) );
  NAND2_X2 MULT_mult_6_U431 ( .A1(MULT_mult_6_ab_1__18_), .A2(MULT_mult_6_n365), .ZN(MULT_mult_6_n126) );
  NAND2_X4 MULT_mult_6_U429 ( .A1(MULT_mult_6_n123), .A2(MULT_mult_6_n122), 
        .ZN(MULT_mult_6_net119951) );
  NAND2_X2 MULT_mult_6_U427 ( .A1(MULT_mult_6_net82152), .A2(
        MULT_mult_6_net84327), .ZN(MULT_mult_6_n122) );
  INV_X4 MULT_mult_6_U426 ( .A(MULT_mult_6_CARRYB_16__9_), .ZN(
        MULT_mult_6_net120655) );
  NAND2_X2 MULT_mult_6_U425 ( .A1(MULT_mult_6_SUMB_12__13_), .A2(
        MULT_mult_6_CARRYB_12__12_), .ZN(MULT_mult_6_n2123) );
  NAND2_X4 MULT_mult_6_U424 ( .A1(MULT_mult_6_n1242), .A2(
        MULT_mult_6_ab_5__16_), .ZN(MULT_mult_6_n1897) );
  NAND3_X4 MULT_mult_6_U423 ( .A1(MULT_mult_6_n2123), .A2(MULT_mult_6_n2124), 
        .A3(MULT_mult_6_n2125), .ZN(MULT_mult_6_CARRYB_13__12_) );
  INV_X8 MULT_mult_6_U422 ( .A(MULT_mult_6_CARRYB_13__12_), .ZN(
        MULT_mult_6_n1486) );
  NAND2_X1 MULT_mult_6_U421 ( .A1(MULT_mult_6_SUMB_6__19_), .A2(
        MULT_mult_6_ab_7__18_), .ZN(MULT_mult_6_net80303) );
  INV_X2 MULT_mult_6_U420 ( .A(MULT_mult_6_SUMB_21__8_), .ZN(MULT_mult_6_n684)
         );
  INV_X8 MULT_mult_6_U419 ( .A(MULT_mult_6_n437), .ZN(MULT_mult_6_SUMB_1__15_)
         );
  NAND2_X4 MULT_mult_6_U418 ( .A1(MULT_mult_6_n46), .A2(MULT_mult_6_n230), 
        .ZN(MULT_mult_6_n232) );
  INV_X4 MULT_mult_6_U417 ( .A(MULT_mult_6_net84902), .ZN(MULT_mult_6_n533) );
  NAND2_X2 MULT_mult_6_U416 ( .A1(MULT_mult_6_net84902), .A2(MULT_mult_6_n402), 
        .ZN(MULT_mult_6_n534) );
  INV_X4 MULT_mult_6_U415 ( .A(MULT_mult_6_SUMB_4__11_), .ZN(MULT_mult_6_n118)
         );
  INV_X4 MULT_mult_6_U414 ( .A(MULT_mult_6_n1658), .ZN(MULT_mult_6_n117) );
  NAND2_X4 MULT_mult_6_U413 ( .A1(MULT_mult_6_n119), .A2(MULT_mult_6_n120), 
        .ZN(MULT_mult_6_SUMB_5__10_) );
  NAND2_X4 MULT_mult_6_U412 ( .A1(MULT_mult_6_n117), .A2(MULT_mult_6_n118), 
        .ZN(MULT_mult_6_n120) );
  NAND2_X2 MULT_mult_6_U411 ( .A1(MULT_mult_6_n1658), .A2(
        MULT_mult_6_SUMB_4__11_), .ZN(MULT_mult_6_n119) );
  INV_X4 MULT_mult_6_U410 ( .A(MULT_mult_6_ab_28__2_), .ZN(MULT_mult_6_n114)
         );
  INV_X4 MULT_mult_6_U409 ( .A(MULT_mult_6_CARRYB_27__2_), .ZN(
        MULT_mult_6_n113) );
  NAND2_X4 MULT_mult_6_U408 ( .A1(MULT_mult_6_n115), .A2(MULT_mult_6_n116), 
        .ZN(MULT_mult_6_net84902) );
  NAND2_X4 MULT_mult_6_U407 ( .A1(MULT_mult_6_n113), .A2(MULT_mult_6_n114), 
        .ZN(MULT_mult_6_n116) );
  INV_X2 MULT_mult_6_U406 ( .A(MULT_mult_6_SUMB_24__5_), .ZN(MULT_mult_6_n1596) );
  INV_X4 MULT_mult_6_U405 ( .A(MULT_mult_6_CARRYB_13__4_), .ZN(
        MULT_mult_6_n1631) );
  NAND2_X1 MULT_mult_6_U404 ( .A1(MULT_mult_6_ab_24__3_), .A2(MULT_mult_6_n417), .ZN(MULT_mult_6_net84680) );
  NAND2_X4 MULT_mult_6_U403 ( .A1(MULT_mult_6_n700), .A2(MULT_mult_6_n701), 
        .ZN(MULT_mult_6_n703) );
  INV_X32 MULT_mult_6_U401 ( .A(MULT_mult_6_net77984), .ZN(
        MULT_mult_6_net80409) );
  NOR2_X4 MULT_mult_6_U400 ( .A1(MULT_mult_6_net87396), .A2(
        MULT_mult_6_net80409), .ZN(MULT_mult_6_n112) );
  NAND3_X2 MULT_mult_6_U399 ( .A1(MULT_mult_6_n1091), .A2(MULT_mult_6_n1092), 
        .A3(MULT_mult_6_n1093), .ZN(MULT_mult_6_n111) );
  NAND2_X2 MULT_mult_6_U398 ( .A1(MULT_mult_6_CARRYB_7__11_), .A2(
        MULT_mult_6_ab_8__11_), .ZN(MULT_mult_6_n2128) );
  NAND2_X4 MULT_mult_6_U397 ( .A1(MULT_mult_6_n1599), .A2(
        MULT_mult_6_ab_9__16_), .ZN(MULT_mult_6_n1602) );
  NAND2_X2 MULT_mult_6_U396 ( .A1(MULT_mult_6_n814), .A2(
        MULT_mult_6_SUMB_14__12_), .ZN(MULT_mult_6_n815) );
  INV_X2 MULT_mult_6_U395 ( .A(MULT_mult_6_CARRYB_15__11_), .ZN(
        MULT_mult_6_n1733) );
  NAND2_X2 MULT_mult_6_U394 ( .A1(MULT_mult_6_ab_16__11_), .A2(
        MULT_mult_6_CARRYB_15__11_), .ZN(MULT_mult_6_n2097) );
  NAND2_X2 MULT_mult_6_U393 ( .A1(MULT_mult_6_net119955), .A2(
        MULT_mult_6_net119927), .ZN(MULT_mult_6_net148838) );
  XOR2_X2 MULT_mult_6_U392 ( .A(MULT_mult_6_CARRYB_6__20_), .B(
        MULT_mult_6_net81340), .Z(MULT_mult_6_n110) );
  XNOR2_X2 MULT_mult_6_U391 ( .A(MULT_mult_6_SUMB_6__21_), .B(MULT_mult_6_n110), .ZN(MULT_mult_6_SUMB_7__20_) );
  CLKBUF_X3 MULT_mult_6_U390 ( .A(MULT_mult_6_net91088), .Z(
        MULT_mult_6_net122062) );
  INV_X2 MULT_mult_6_U389 ( .A(MULT_mult_6_ab_4__17_), .ZN(MULT_mult_6_n107)
         );
  INV_X4 MULT_mult_6_U388 ( .A(MULT_mult_6_CARRYB_3__17_), .ZN(
        MULT_mult_6_n106) );
  NAND2_X4 MULT_mult_6_U387 ( .A1(MULT_mult_6_n108), .A2(MULT_mult_6_n109), 
        .ZN(MULT_mult_6_n1742) );
  NAND2_X4 MULT_mult_6_U386 ( .A1(MULT_mult_6_n106), .A2(MULT_mult_6_n107), 
        .ZN(MULT_mult_6_n109) );
  NAND2_X2 MULT_mult_6_U385 ( .A1(MULT_mult_6_CARRYB_3__17_), .A2(
        MULT_mult_6_ab_4__17_), .ZN(MULT_mult_6_n108) );
  NAND3_X2 MULT_mult_6_U384 ( .A1(MULT_mult_6_net82561), .A2(
        MULT_mult_6_net82560), .A3(MULT_mult_6_net82559), .ZN(MULT_mult_6_n105) );
  NAND2_X4 MULT_mult_6_U383 ( .A1(MULT_mult_6_net85543), .A2(MULT_mult_6_n484), 
        .ZN(MULT_mult_6_n104) );
  NAND3_X4 MULT_mult_6_U382 ( .A1(MULT_mult_6_n1070), .A2(MULT_mult_6_n1069), 
        .A3(MULT_mult_6_n1068), .ZN(MULT_mult_6_CARRYB_3__22_) );
  NAND2_X4 MULT_mult_6_U381 ( .A1(MULT_mult_6_n279), .A2(MULT_mult_6_net123267), .ZN(MULT_mult_6_net120511) );
  BUF_X8 MULT_mult_6_U380 ( .A(MULT_mult_6_net88079), .Z(MULT_mult_6_n137) );
  NAND2_X2 MULT_mult_6_U379 ( .A1(MULT_mult_6_CARRYB_6__19_), .A2(
        MULT_mult_6_SUMB_6__20_), .ZN(MULT_mult_6_n1103) );
  INV_X4 MULT_mult_6_U378 ( .A(MULT_mult_6_CARRYB_2__11_), .ZN(
        MULT_mult_6_n913) );
  NAND2_X4 MULT_mult_6_U377 ( .A1(MULT_mult_6_SUMB_16__3_), .A2(
        MULT_mult_6_CARRYB_16__2_), .ZN(MULT_mult_6_n1669) );
  NAND2_X4 MULT_mult_6_U376 ( .A1(MULT_mult_6_n1944), .A2(MULT_mult_6_n1328), 
        .ZN(MULT_mult_6_n1551) );
  NAND2_X2 MULT_mult_6_U375 ( .A1(MULT_mult_6_SUMB_3__9_), .A2(
        MULT_mult_6_ab_4__8_), .ZN(MULT_mult_6_n1945) );
  OR2_X2 MULT_mult_6_U374 ( .A1(MULT_mult_6_SUMB_22__4_), .A2(
        MULT_mult_6_ab_23__3_), .ZN(MULT_mult_6_n422) );
  NAND2_X2 MULT_mult_6_U373 ( .A1(MULT_mult_6_SUMB_22__4_), .A2(
        MULT_mult_6_n420), .ZN(MULT_mult_6_n419) );
  INV_X4 MULT_mult_6_U372 ( .A(MULT_mult_6_SUMB_22__4_), .ZN(MULT_mult_6_n405)
         );
  NAND2_X2 MULT_mult_6_U371 ( .A1(MULT_mult_6_n405), .A2(MULT_mult_6_n420), 
        .ZN(MULT_mult_6_n103) );
  NOR2_X2 MULT_mult_6_U370 ( .A1(MULT_mult_6_n247), .A2(MULT_mult_6_n103), 
        .ZN(MULT_mult_6_n409) );
  NAND2_X2 MULT_mult_6_U369 ( .A1(MULT_mult_6_ab_21__0_), .A2(
        MULT_mult_6_SUMB_20__1_), .ZN(MULT_mult_6_n1806) );
  NAND2_X4 MULT_mult_6_U368 ( .A1(MULT_mult_6_net88177), .A2(
        MULT_mult_6_ab_1__9_), .ZN(MULT_mult_6_n1517) );
  NAND2_X4 MULT_mult_6_U367 ( .A1(MULT_mult_6_ab_16__3_), .A2(
        MULT_mult_6_CARRYB_15__3_), .ZN(MULT_mult_6_n1131) );
  NAND2_X1 MULT_mult_6_U366 ( .A1(MULT_mult_6_CARRYB_3__6_), .A2(
        MULT_mult_6_SUMB_3__7_), .ZN(MULT_mult_6_net88208) );
  NAND2_X4 MULT_mult_6_U365 ( .A1(MULT_mult_6_n1031), .A2(MULT_mult_6_n1032), 
        .ZN(MULT_mult_6_n1658) );
  NAND2_X2 MULT_mult_6_U364 ( .A1(MULT_mult_6_n1272), .A2(
        MULT_mult_6_SUMB_26__4_), .ZN(MULT_mult_6_net80816) );
  NAND2_X2 MULT_mult_6_U363 ( .A1(MULT_mult_6_n56), .A2(MULT_mult_6_ab_6__19_), 
        .ZN(MULT_mult_6_n979) );
  NAND2_X1 MULT_mult_6_U362 ( .A1(MULT_mult_6_SUMB_13__12_), .A2(
        MULT_mult_6_ab_14__11_), .ZN(MULT_mult_6_net82557) );
  XNOR2_X1 MULT_mult_6_U361 ( .A(MULT_mult_6_net125934), .B(
        MULT_mult_6_net86801), .ZN(MULT_mult_6_SUMB_14__11_) );
  INV_X4 MULT_mult_6_U360 ( .A(MULT_mult_6_n869), .ZN(MULT_mult_6_net86703) );
  NAND2_X4 MULT_mult_6_U359 ( .A1(MULT_mult_6_net86702), .A2(
        MULT_mult_6_net86703), .ZN(MULT_mult_6_n1401) );
  INV_X4 MULT_mult_6_U358 ( .A(MULT_mult_6_SUMB_22__5_), .ZN(
        MULT_mult_6_net88648) );
  INV_X4 MULT_mult_6_U357 ( .A(MULT_mult_6_net88648), .ZN(MULT_mult_6_n102) );
  NAND2_X4 MULT_mult_6_U356 ( .A1(MULT_mult_6_n280), .A2(MULT_mult_6_n281), 
        .ZN(MULT_mult_6_n283) );
  NAND2_X4 MULT_mult_6_U355 ( .A1(MULT_mult_6_ab_8__10_), .A2(
        MULT_mult_6_SUMB_7__11_), .ZN(MULT_mult_6_net81215) );
  INV_X4 MULT_mult_6_U354 ( .A(MULT_mult_6_n100), .ZN(MULT_mult_6_n101) );
  NAND2_X2 MULT_mult_6_U353 ( .A1(MULT_mult_6_n101), .A2(MULT_mult_6_net82407), 
        .ZN(MULT_mult_6_net86464) );
  NAND2_X2 MULT_mult_6_U352 ( .A1(MULT_mult_6_n1882), .A2(MULT_mult_6_net82408), .ZN(MULT_mult_6_n100) );
  NAND2_X2 MULT_mult_6_U351 ( .A1(MULT_mult_6_ab_2__17_), .A2(
        MULT_mult_6__UDW__112684_net78547), .ZN(MULT_mult_6_n1343) );
  NAND2_X4 MULT_mult_6_U349 ( .A1(MULT_mult_6_n818), .A2(MULT_mult_6_ab_22__6_), .ZN(MULT_mult_6_n820) );
  INV_X8 MULT_mult_6_U348 ( .A(aluA[30]), .ZN(MULT_mult_6_net70493) );
  NAND3_X2 MULT_mult_6_U347 ( .A1(MULT_mult_6_n454), .A2(MULT_mult_6_n453), 
        .A3(MULT_mult_6_n455), .ZN(MULT_mult_6_n99) );
  NAND2_X4 MULT_mult_6_U346 ( .A1(MULT_mult_6_CARRYB_20__6_), .A2(
        MULT_mult_6_net81042), .ZN(MULT_mult_6_n781) );
  XNOR2_X1 MULT_mult_6_U345 ( .A(MULT_mult_6_CARRYB_24__1_), .B(
        MULT_mult_6_ab_25__1_), .ZN(MULT_mult_6_net93880) );
  INV_X8 MULT_mult_6_U344 ( .A(n10924), .ZN(MULT_mult_6_net77906) );
  NOR2_X4 MULT_mult_6_U343 ( .A1(MULT_mult_6_net124610), .A2(
        MULT_mult_6_net77906), .ZN(MULT_mult_6_ab_0__6_) );
  NAND2_X2 MULT_mult_6_U342 ( .A1(MULT_mult_6_ab_17__0_), .A2(
        MULT_mult_6_SUMB_16__1_), .ZN(MULT_mult_6_net86654) );
  NAND2_X2 MULT_mult_6_U341 ( .A1(MULT_mult_6_CARRYB_25__2_), .A2(
        MULT_mult_6_ab_26__2_), .ZN(MULT_mult_6_n1033) );
  INV_X32 MULT_mult_6_U340 ( .A(MULT_mult_6_ab_16__1_), .ZN(MULT_mult_6_n98)
         );
  XNOR2_X2 MULT_mult_6_U339 ( .A(MULT_mult_6_SUMB_15__2_), .B(MULT_mult_6_n98), 
        .ZN(MULT_mult_6_n646) );
  NAND2_X4 MULT_mult_6_U338 ( .A1(MULT_mult_6_ab_9__15_), .A2(MULT_mult_6_n151), .ZN(MULT_mult_6_n2049) );
  INV_X8 MULT_mult_6_U337 ( .A(MULT_mult_6_SUMB_22__7_), .ZN(MULT_mult_6_n697)
         );
  INV_X8 MULT_mult_6_U336 ( .A(MULT_mult_6_n96), .ZN(MULT_mult_6_n97) );
  INV_X4 MULT_mult_6_U335 ( .A(MULT_mult_6_net87936), .ZN(MULT_mult_6_n96) );
  INV_X1 MULT_mult_6_U334 ( .A(MULT_mult_6_n799), .ZN(MULT_mult_6_n95) );
  INV_X2 MULT_mult_6_U333 ( .A(MULT_mult_6_SUMB_2__15_), .ZN(MULT_mult_6_n1557) );
  NAND2_X4 MULT_mult_6_U332 ( .A1(MULT_mult_6_net147920), .A2(
        MULT_mult_6_ab_5__11_), .ZN(MULT_mult_6_n677) );
  INV_X8 MULT_mult_6_U331 ( .A(MULT_mult_6_n917), .ZN(MULT_mult_6_n927) );
  INV_X2 MULT_mult_6_U329 ( .A(MULT_mult_6_n910), .ZN(MULT_mult_6_n94) );
  NAND2_X4 MULT_mult_6_U328 ( .A1(MULT_mult_6_n1126), .A2(MULT_mult_6_n174), 
        .ZN(MULT_mult_6_n1127) );
  INV_X2 MULT_mult_6_U327 ( .A(MULT_mult_6_n92), .ZN(MULT_mult_6_n93) );
  INV_X1 MULT_mult_6_U326 ( .A(MULT_mult_6_net88079), .ZN(MULT_mult_6_n92) );
  NAND2_X2 MULT_mult_6_U325 ( .A1(MULT_mult_6_CARRYB_4__10_), .A2(
        MULT_mult_6_ab_5__10_), .ZN(MULT_mult_6_n1031) );
  NAND2_X2 MULT_mult_6_U324 ( .A1(MULT_mult_6_n181), .A2(MULT_mult_6_n228), 
        .ZN(MULT_mult_6_n1745) );
  NAND2_X2 MULT_mult_6_U323 ( .A1(MULT_mult_6_ab_5__10_), .A2(MULT_mult_6_n181), .ZN(MULT_mult_6_n1746) );
  NAND2_X2 MULT_mult_6_U322 ( .A1(MULT_mult_6_CARRYB_28__0_), .A2(
        MULT_mult_6_n344), .ZN(MULT_mult_6_n250) );
  NAND2_X1 MULT_mult_6_U321 ( .A1(MULT_mult_6_ab_13__16_), .A2(
        MULT_mult_6_SUMB_12__17_), .ZN(MULT_mult_6_n2317) );
  NAND2_X4 MULT_mult_6_U320 ( .A1(MULT_mult_6_SUMB_16__9_), .A2(
        MULT_mult_6_ab_17__8_), .ZN(MULT_mult_6_n811) );
  INV_X2 MULT_mult_6_U319 ( .A(MULT_mult_6_SUMB_7__8_), .ZN(MULT_mult_6_n1864)
         );
  NOR2_X4 MULT_mult_6_U318 ( .A1(MULT_mult_6_net70458), .A2(
        MULT_mult_6_net80409), .ZN(MULT_mult_6_n237) );
  NAND2_X4 MULT_mult_6_U317 ( .A1(MULT_mult_6_n1516), .A2(MULT_mult_6_net90174), .ZN(MULT_mult_6_n1518) );
  NAND2_X1 MULT_mult_6_U316 ( .A1(MULT_mult_6_CARRYB_3__21_), .A2(
        MULT_mult_6_SUMB_3__22_), .ZN(MULT_mult_6_n2276) );
  NOR2_X2 MULT_mult_6_U315 ( .A1(MULT_mult_6_net123000), .A2(
        MULT_mult_6_net82247), .ZN(MULT_mult_6_net149526) );
  INV_X4 MULT_mult_6_U314 ( .A(MULT_mult_6_net87050), .ZN(
        MULT_mult_6_ab_1__17_) );
  INV_X2 MULT_mult_6_U313 ( .A(MULT_mult_6_net87396), .ZN(MULT_mult_6_n90) );
  NAND2_X4 MULT_mult_6_U312 ( .A1(MULT_mult_6_ab_17__2_), .A2(
        MULT_mult_6_CARRYB_16__2_), .ZN(MULT_mult_6_n1668) );
  NOR2_X4 MULT_mult_6_U311 ( .A1(MULT_mult_6_n68), .A2(MULT_mult_6_net70491), 
        .ZN(MULT_mult_6_ab_2__12_) );
  INV_X2 MULT_mult_6_U310 ( .A(MULT_mult_6_SUMB_18__7_), .ZN(
        MULT_mult_6_net90576) );
  NOR2_X2 MULT_mult_6_U308 ( .A1(MULT_mult_6_net84698), .A2(
        MULT_mult_6_net77932), .ZN(MULT_mult_6_ab_7__14_) );
  NAND2_X2 MULT_mult_6_U307 ( .A1(MULT_mult_6_ab_10__15_), .A2(
        MULT_mult_6_SUMB_9__16_), .ZN(MULT_mult_6_n1840) );
  NAND2_X2 MULT_mult_6_U306 ( .A1(MULT_mult_6_SUMB_9__16_), .A2(
        MULT_mult_6_CARRYB_9__15_), .ZN(MULT_mult_6_n1841) );
  NAND2_X4 MULT_mult_6_U305 ( .A1(MULT_mult_6_ab_17__10_), .A2(
        MULT_mult_6_SUMB_16__11_), .ZN(MULT_mult_6_n1580) );
  NOR2_X2 MULT_mult_6_U304 ( .A1(MULT_mult_6_net70486), .A2(
        MULT_mult_6_net80409), .ZN(MULT_mult_6_ab_1__26_) );
  NAND2_X4 MULT_mult_6_U303 ( .A1(MULT_mult_6_net84817), .A2(
        MULT_mult_6_net84818), .ZN(MULT_mult_6_n1743) );
  INV_X8 MULT_mult_6_U302 ( .A(MULT_mult_6_net119974), .ZN(
        MULT_mult_6_net119910) );
  INV_X4 MULT_mult_6_U301 ( .A(MULT_mult_6_net119948), .ZN(MULT_mult_6_n477)
         );
  INV_X4 MULT_mult_6_U300 ( .A(MULT_mult_6_n1901), .ZN(MULT_mult_6_n1126) );
  NAND2_X4 MULT_mult_6_U299 ( .A1(MULT_mult_6_CARRYB_4__14_), .A2(
        MULT_mult_6_net84946), .ZN(MULT_mult_6_net84947) );
  INV_X4 MULT_mult_6_U298 ( .A(MULT_mult_6_n1742), .ZN(MULT_mult_6_n238) );
  NAND2_X4 MULT_mult_6_U297 ( .A1(MULT_mult_6_ab_5__18_), .A2(
        MULT_mult_6_SUMB_4__19_), .ZN(MULT_mult_6_n2140) );
  NOR2_X4 MULT_mult_6_U296 ( .A1(MULT_mult_6_net92314), .A2(MULT_mult_6_n1181), 
        .ZN(MULT_mult_6_n1182) );
  NAND2_X4 MULT_mult_6_U295 ( .A1(MULT_mult_6_CARRYB_18__3_), .A2(
        MULT_mult_6_ab_19__3_), .ZN(MULT_mult_6_n2275) );
  CLKBUF_X3 MULT_mult_6_U294 ( .A(MULT_mult_6_n1425), .Z(MULT_mult_6_n1157) );
  NAND3_X4 MULT_mult_6_U293 ( .A1(MULT_mult_6_n1590), .A2(MULT_mult_6_n1747), 
        .A3(MULT_mult_6_n1748), .ZN(MULT_mult_6_CARRYB_6__10_) );
  NAND2_X4 MULT_mult_6_U292 ( .A1(MULT_mult_6_ab_21__2_), .A2(MULT_mult_6_n596), .ZN(MULT_mult_6_n2187) );
  NAND2_X4 MULT_mult_6_U291 ( .A1(MULT_mult_6_n641), .A2(MULT_mult_6_n622), 
        .ZN(MULT_mult_6_n624) );
  NAND3_X2 MULT_mult_6_U289 ( .A1(MULT_mult_6_n2007), .A2(MULT_mult_6_n2008), 
        .A3(MULT_mult_6_n2009), .ZN(MULT_mult_6_n89) );
  NAND2_X4 MULT_mult_6_U288 ( .A1(MULT_mult_6_net82029), .A2(MULT_mult_6_n490), 
        .ZN(MULT_mult_6_net82152) );
  NAND3_X4 MULT_mult_6_U286 ( .A1(MULT_mult_6_n2104), .A2(MULT_mult_6_n2103), 
        .A3(MULT_mult_6_n2105), .ZN(MULT_mult_6_n176) );
  NAND2_X4 MULT_mult_6_U285 ( .A1(MULT_mult_6_ab_11__4_), .A2(MULT_mult_6_n563), .ZN(MULT_mult_6_n1833) );
  INV_X8 MULT_mult_6_U284 ( .A(MULT_mult_6_CARRYB_1__11_), .ZN(
        MULT_mult_6_n586) );
  INV_X2 MULT_mult_6_U283 ( .A(MULT_mult_6_SUMB_13__13_), .ZN(MULT_mult_6_n133) );
  NAND2_X2 MULT_mult_6_U282 ( .A1(MULT_mult_6_SUMB_13__13_), .A2(
        MULT_mult_6_n134), .ZN(MULT_mult_6_n135) );
  NAND2_X4 MULT_mult_6_U281 ( .A1(MULT_mult_6_SUMB_13__13_), .A2(
        MULT_mult_6_n1345), .ZN(MULT_mult_6_n2120) );
  NAND2_X4 MULT_mult_6_U280 ( .A1(MULT_mult_6_n562), .A2(
        MULT_mult_6_SUMB_11__14_), .ZN(MULT_mult_6_n1793) );
  INV_X8 MULT_mult_6_U279 ( .A(MULT_mult_6_SUMB_17__10_), .ZN(MULT_mult_6_n825) );
  INV_X2 MULT_mult_6_U278 ( .A(MULT_mult_6_SUMB_12__14_), .ZN(MULT_mult_6_n86)
         );
  INV_X4 MULT_mult_6_U277 ( .A(MULT_mult_6_n1323), .ZN(MULT_mult_6_n85) );
  NAND2_X4 MULT_mult_6_U276 ( .A1(MULT_mult_6_n87), .A2(MULT_mult_6_n88), .ZN(
        MULT_mult_6_SUMB_13__13_) );
  NAND2_X2 MULT_mult_6_U275 ( .A1(MULT_mult_6_n85), .A2(MULT_mult_6_n86), .ZN(
        MULT_mult_6_n88) );
  INV_X4 MULT_mult_6_U274 ( .A(MULT_mult_6_n556), .ZN(MULT_mult_6_n82) );
  INV_X4 MULT_mult_6_U273 ( .A(MULT_mult_6_n1226), .ZN(MULT_mult_6_n81) );
  NAND2_X4 MULT_mult_6_U272 ( .A1(MULT_mult_6_n83), .A2(MULT_mult_6_n84), .ZN(
        MULT_mult_6_SUMB_11__14_) );
  NAND2_X4 MULT_mult_6_U271 ( .A1(MULT_mult_6_n81), .A2(MULT_mult_6_n82), .ZN(
        MULT_mult_6_n84) );
  NAND2_X2 MULT_mult_6_U270 ( .A1(MULT_mult_6_n1226), .A2(MULT_mult_6_n556), 
        .ZN(MULT_mult_6_n83) );
  INV_X4 MULT_mult_6_U269 ( .A(MULT_mult_6_n682), .ZN(MULT_mult_6_n78) );
  INV_X4 MULT_mult_6_U268 ( .A(MULT_mult_6_net85325), .ZN(MULT_mult_6_n77) );
  NAND2_X4 MULT_mult_6_U267 ( .A1(MULT_mult_6_n79), .A2(MULT_mult_6_n80), .ZN(
        MULT_mult_6_SUMB_17__10_) );
  NAND2_X4 MULT_mult_6_U266 ( .A1(MULT_mult_6_n77), .A2(MULT_mult_6_n78), .ZN(
        MULT_mult_6_n80) );
  NAND2_X2 MULT_mult_6_U265 ( .A1(MULT_mult_6_net85325), .A2(MULT_mult_6_n682), 
        .ZN(MULT_mult_6_n79) );
  INV_X2 MULT_mult_6_U264 ( .A(MULT_mult_6_SUMB_11__13_), .ZN(MULT_mult_6_n785) );
  CLKBUF_X3 MULT_mult_6_U263 ( .A(MULT_mult_6_n1207), .Z(MULT_mult_6_n1324) );
  INV_X4 MULT_mult_6_U261 ( .A(MULT_mult_6_CARRYB_9__9_), .ZN(MULT_mult_6_n323) );
  NAND2_X4 MULT_mult_6_U260 ( .A1(MULT_mult_6_n323), .A2(MULT_mult_6_n324), 
        .ZN(MULT_mult_6_n326) );
  AND2_X4 MULT_mult_6_U259 ( .A1(n10917), .A2(aluA[29]), .ZN(
        MULT_mult_6_ab_2__15_) );
  XNOR2_X2 MULT_mult_6_U258 ( .A(MULT_mult_6_ab_2__18_), .B(
        MULT_mult_6__UDW__112679_net78533), .ZN(MULT_mult_6_n287) );
  NAND2_X2 MULT_mult_6_U257 ( .A1(MULT_mult_6_n1845), .A2(MULT_mult_6_n1255), 
        .ZN(MULT_mult_6_n1542) );
  NAND2_X4 MULT_mult_6_U256 ( .A1(MULT_mult_6_n1543), .A2(MULT_mult_6_n1542), 
        .ZN(MULT_mult_6_n362) );
  NAND2_X2 MULT_mult_6_U255 ( .A1(MULT_mult_6_CARRYB_3__11_), .A2(
        MULT_mult_6_ab_4__11_), .ZN(MULT_mult_6_net88086) );
  INV_X4 MULT_mult_6_U254 ( .A(MULT_mult_6_ab_22__4_), .ZN(MULT_mult_6_n74) );
  NAND2_X4 MULT_mult_6_U252 ( .A1(MULT_mult_6_n76), .A2(MULT_mult_6_n75), .ZN(
        MULT_mult_6_net80862) );
  NAND2_X4 MULT_mult_6_U251 ( .A1(MULT_mult_6_n73), .A2(MULT_mult_6_n74), .ZN(
        MULT_mult_6_n76) );
  NAND2_X2 MULT_mult_6_U250 ( .A1(MULT_mult_6_CARRYB_21__4_), .A2(
        MULT_mult_6_ab_22__4_), .ZN(MULT_mult_6_n75) );
  INV_X4 MULT_mult_6_U249 ( .A(MULT_mult_6_CARRYB_6__22_), .ZN(
        MULT_mult_6_n876) );
  BUF_X8 MULT_mult_6_U248 ( .A(MULT_mult_6_SUMB_12__18_), .Z(MULT_mult_6_n1240) );
  INV_X8 MULT_mult_6_U247 ( .A(MULT_mult_6_net120625), .ZN(
        MULT_mult_6_net86806) );
  INV_X8 MULT_mult_6_U246 ( .A(MULT_mult_6_net90022), .ZN(MULT_mult_6_n777) );
  NAND2_X2 MULT_mult_6_U245 ( .A1(MULT_mult_6_n777), .A2(MULT_mult_6_net87391), 
        .ZN(MULT_mult_6_net87949) );
  NAND2_X4 MULT_mult_6_U244 ( .A1(MULT_mult_6_n777), .A2(MULT_mult_6_net87391), 
        .ZN(MULT_mult_6_n72) );
  XNOR2_X2 MULT_mult_6_U243 ( .A(MULT_mult_6_CARRYB_22__7_), .B(
        MULT_mult_6_ab_23__7_), .ZN(MULT_mult_6_n867) );
  NAND2_X2 MULT_mult_6_U242 ( .A1(MULT_mult_6_ab_15__13_), .A2(
        MULT_mult_6_SUMB_14__14_), .ZN(MULT_mult_6_net80484) );
  NAND2_X2 MULT_mult_6_U241 ( .A1(MULT_mult_6_CARRYB_14__6_), .A2(
        MULT_mult_6_ab_15__6_), .ZN(MULT_mult_6_n1438) );
  NAND2_X4 MULT_mult_6_U240 ( .A1(MULT_mult_6_SUMB_14__14_), .A2(
        MULT_mult_6_CARRYB_14__13_), .ZN(MULT_mult_6_net80485) );
  NAND3_X4 MULT_mult_6_U239 ( .A1(MULT_mult_6_net80484), .A2(
        MULT_mult_6_net80485), .A3(MULT_mult_6_n1058), .ZN(
        MULT_mult_6_CARRYB_15__13_) );
  NAND2_X2 MULT_mult_6_U238 ( .A1(MULT_mult_6_CARRYB_12__5_), .A2(
        MULT_mult_6_ab_13__5_), .ZN(MULT_mult_6_n1920) );
  NAND2_X2 MULT_mult_6_U237 ( .A1(MULT_mult_6_CARRYB_24__0_), .A2(
        MULT_mult_6_SUMB_24__1_), .ZN(MULT_mult_6_net81530) );
  NAND2_X2 MULT_mult_6_U235 ( .A1(MULT_mult_6_SUMB_23__4_), .A2(
        MULT_mult_6_n417), .ZN(MULT_mult_6_net84678) );
  NAND2_X2 MULT_mult_6_U234 ( .A1(MULT_mult_6_SUMB_26__3_), .A2(
        MULT_mult_6_ab_27__2_), .ZN(MULT_mult_6_n809) );
  INV_X8 MULT_mult_6_U233 ( .A(MULT_mult_6_CARRYB_10__10_), .ZN(
        MULT_mult_6_n201) );
  XNOR2_X2 MULT_mult_6_U232 ( .A(MULT_mult_6_ab_2__18_), .B(
        MULT_mult_6_CARRYB_1__18_), .ZN(MULT_mult_6_n397) );
  NAND2_X2 MULT_mult_6_U231 ( .A1(MULT_mult_6_n1742), .A2(MULT_mult_6_n852), 
        .ZN(MULT_mult_6_n240) );
  CLKBUF_X3 MULT_mult_6_U230 ( .A(MULT_mult_6_SUMB_9__11_), .Z(MULT_mult_6_n70) );
  INV_X8 MULT_mult_6_U229 ( .A(n5759), .ZN(MULT_mult_6_net120391) );
  NOR2_X4 MULT_mult_6_U228 ( .A1(MULT_mult_6_net120391), .A2(
        MULT_mult_6_net80409), .ZN(MULT_mult_6_ab_1__13_) );
  INV_X8 MULT_mult_6_U227 ( .A(MULT_mult_6_CARRYB_20__6_), .ZN(
        MULT_mult_6_net81553) );
  INV_X1 MULT_mult_6_U226 ( .A(MULT_mult_6_net81553), .ZN(MULT_mult_6_n69) );
  OR2_X4 MULT_mult_6_U225 ( .A1(MULT_mult_6_net85251), .A2(MULT_mult_6_n497), 
        .ZN(MULT_mult_6_n494) );
  INV_X2 MULT_mult_6_U224 ( .A(MULT_mult_6_net86893), .ZN(MULT_mult_6_n229) );
  INV_X4 MULT_mult_6_U223 ( .A(MULT_mult_6_net82551), .ZN(MULT_mult_6_net90433) );
  NAND2_X4 MULT_mult_6_U222 ( .A1(MULT_mult_6_n1385), .A2(MULT_mult_6_net87005), .ZN(MULT_mult_6_net82641) );
  NOR2_X4 MULT_mult_6_U221 ( .A1(MULT_mult_6_net70478), .A2(
        MULT_mult_6_net86101), .ZN(MULT_mult_6_n2196) );
  INV_X4 MULT_mult_6_U220 ( .A(MULT_mult_6_n491), .ZN(MULT_mult_6_n68) );
  INV_X2 MULT_mult_6_U219 ( .A(MULT_mult_6_n1699), .ZN(MULT_mult_6_n67) );
  NAND2_X2 MULT_mult_6_U218 ( .A1(MULT_mult_6_SUMB_6__11_), .A2(
        MULT_mult_6_CARRYB_6__10_), .ZN(MULT_mult_6_n473) );
  NAND3_X4 MULT_mult_6_U216 ( .A1(MULT_mult_6_n1874), .A2(MULT_mult_6_n1875), 
        .A3(MULT_mult_6_n1876), .ZN(MULT_mult_6_CARRYB_10__18_) );
  CLKBUF_X2 MULT_mult_6_U215 ( .A(MULT_mult_6_SUMB_6__11_), .Z(
        MULT_mult_6_net149004) );
  XNOR2_X2 MULT_mult_6_U214 ( .A(MULT_mult_6_CARRYB_20__4_), .B(
        MULT_mult_6_n945), .ZN(MULT_mult_6_n66) );
  NAND2_X2 MULT_mult_6_U213 ( .A1(MULT_mult_6_SUMB_13__5_), .A2(
        MULT_mult_6_ab_14__4_), .ZN(MULT_mult_6_n2151) );
  NAND2_X4 MULT_mult_6_U212 ( .A1(MULT_mult_6_n1271), .A2(
        MULT_mult_6_SUMB_10__6_), .ZN(MULT_mult_6_n2061) );
  NAND2_X2 MULT_mult_6_U211 ( .A1(MULT_mult_6_SUMB_25__4_), .A2(
        MULT_mult_6_ab_26__3_), .ZN(MULT_mult_6_net81052) );
  CLKBUF_X2 MULT_mult_6_U210 ( .A(MULT_mult_6_SUMB_25__4_), .Z(
        MULT_mult_6_net83030) );
  NAND2_X2 MULT_mult_6_U209 ( .A1(MULT_mult_6_n1598), .A2(MULT_mult_6_n1597), 
        .ZN(MULT_mult_6_n91) );
  NOR2_X4 MULT_mult_6_U208 ( .A1(MULT_mult_6_n392), .A2(MULT_mult_6_n2355), 
        .ZN(MULT_mult_6_ab_0__27_) );
  NAND2_X4 MULT_mult_6_U207 ( .A1(MULT_mult_6_n148), .A2(MULT_mult_6_n149), 
        .ZN(MULT_mult_6_net82154) );
  NAND2_X2 MULT_mult_6_U206 ( .A1(MULT_mult_6_n366), .A2(MULT_mult_6_net86464), 
        .ZN(MULT_mult_6_n2302) );
  BUF_X4 MULT_mult_6_U205 ( .A(MULT_mult_6_SUMB_20__6_), .Z(MULT_mult_6_n71)
         );
  INV_X4 MULT_mult_6_U204 ( .A(MULT_mult_6_n71), .ZN(MULT_mult_6_n63) );
  INV_X4 MULT_mult_6_U203 ( .A(MULT_mult_6_net83705), .ZN(MULT_mult_6_n62) );
  NAND2_X4 MULT_mult_6_U202 ( .A1(MULT_mult_6_n64), .A2(MULT_mult_6_n65), .ZN(
        MULT_mult_6_n366) );
  NAND2_X4 MULT_mult_6_U201 ( .A1(MULT_mult_6_n62), .A2(MULT_mult_6_n63), .ZN(
        MULT_mult_6_n65) );
  NAND2_X2 MULT_mult_6_U200 ( .A1(MULT_mult_6_net83705), .A2(MULT_mult_6_n71), 
        .ZN(MULT_mult_6_n64) );
  NAND2_X4 MULT_mult_6_U199 ( .A1(MULT_mult_6_n1562), .A2(MULT_mult_6_n94), 
        .ZN(MULT_mult_6_n911) );
  BUF_X8 MULT_mult_6_U198 ( .A(MULT_mult_6_SUMB_7__11_), .Z(
        MULT_mult_6_net120922) );
  INV_X8 MULT_mult_6_U197 ( .A(MULT_mult_6_net83736), .ZN(
        MULT_mult_6_net121606) );
  NAND2_X2 MULT_mult_6_U196 ( .A1(MULT_mult_6_ab_1__17_), .A2(
        MULT_mult_6_net85688), .ZN(MULT_mult_6_net82286) );
  NAND2_X4 MULT_mult_6_U195 ( .A1(MULT_mult_6_SUMB_14__6_), .A2(
        MULT_mult_6_ab_15__5_), .ZN(MULT_mult_6_n1978) );
  NAND2_X4 MULT_mult_6_U194 ( .A1(MULT_mult_6_n216), .A2(MULT_mult_6_n217), 
        .ZN(MULT_mult_6_n219) );
  INV_X4 MULT_mult_6_U193 ( .A(MULT_mult_6_n1927), .ZN(MULT_mult_6_n1524) );
  INV_X2 MULT_mult_6_U192 ( .A(MULT_mult_6_CARRYB_4__18_), .ZN(
        MULT_mult_6_n1767) );
  NAND2_X1 MULT_mult_6_U191 ( .A1(MULT_mult_6_net90702), .A2(
        MULT_mult_6_CARRYB_6__17_), .ZN(MULT_mult_6_n932) );
  INV_X4 MULT_mult_6_U190 ( .A(MULT_mult_6_CARRYB_8__16_), .ZN(
        MULT_mult_6_n1599) );
  NAND2_X4 MULT_mult_6_U189 ( .A1(MULT_mult_6_SUMB_1__15_), .A2(
        MULT_mult_6_CARRYB_1__14_), .ZN(MULT_mult_6_net86171) );
  NAND2_X2 MULT_mult_6_U188 ( .A1(MULT_mult_6_ab_14__15_), .A2(
        MULT_mult_6_SUMB_13__16_), .ZN(MULT_mult_6_n1871) );
  NAND2_X2 MULT_mult_6_U187 ( .A1(MULT_mult_6_ab_8__18_), .A2(
        MULT_mult_6_n1109), .ZN(MULT_mult_6_n1105) );
  NAND2_X4 MULT_mult_6_U186 ( .A1(MULT_mult_6_net123055), .A2(MULT_mult_6_n927), .ZN(MULT_mult_6_n928) );
  NAND2_X4 MULT_mult_6_U185 ( .A1(MULT_mult_6_net80657), .A2(
        MULT_mult_6_net80658), .ZN(MULT_mult_6_net80660) );
  NAND3_X2 MULT_mult_6_U184 ( .A1(MULT_mult_6_net82667), .A2(
        MULT_mult_6_net82668), .A3(MULT_mult_6_net82669), .ZN(
        MULT_mult_6_CARRYB_19__10_) );
  NAND2_X4 MULT_mult_6_U183 ( .A1(MULT_mult_6_SUMB_2__14_), .A2(
        MULT_mult_6_n99), .ZN(MULT_mult_6_net81513) );
  NAND2_X2 MULT_mult_6_U182 ( .A1(MULT_mult_6_SUMB_4__20_), .A2(
        MULT_mult_6_ab_5__19_), .ZN(MULT_mult_6_n2241) );
  NOR2_X2 MULT_mult_6_U181 ( .A1(MULT_mult_6_net77912), .A2(
        MULT_mult_6_net70449), .ZN(MULT_mult_6_ab_23__7_) );
  INV_X4 MULT_mult_6_U180 ( .A(MULT_mult_6_SUMB_17__11_), .ZN(MULT_mult_6_n59)
         );
  INV_X4 MULT_mult_6_U179 ( .A(MULT_mult_6_net87009), .ZN(MULT_mult_6_n58) );
  NAND2_X2 MULT_mult_6_U176 ( .A1(MULT_mult_6_net87009), .A2(
        MULT_mult_6_SUMB_17__11_), .ZN(MULT_mult_6_n60) );
  XNOR2_X2 MULT_mult_6_U175 ( .A(MULT_mult_6_ab_2__21_), .B(
        MULT_mult_6_CARRYB_1__21_), .ZN(MULT_mult_6_n57) );
  NAND3_X2 MULT_mult_6_U174 ( .A1(MULT_mult_6_n2241), .A2(MULT_mult_6_n2240), 
        .A3(MULT_mult_6_n2242), .ZN(MULT_mult_6_n56) );
  INV_X1 MULT_mult_6_U173 ( .A(MULT_mult_6_ab_23__7_), .ZN(MULT_mult_6_n53) );
  INV_X1 MULT_mult_6_U172 ( .A(MULT_mult_6_CARRYB_22__7_), .ZN(MULT_mult_6_n52) );
  NAND2_X2 MULT_mult_6_U171 ( .A1(MULT_mult_6_n54), .A2(MULT_mult_6_n55), .ZN(
        MULT_mult_6_net88961) );
  NAND2_X2 MULT_mult_6_U170 ( .A1(MULT_mult_6_n52), .A2(MULT_mult_6_n53), .ZN(
        MULT_mult_6_n55) );
  NAND2_X1 MULT_mult_6_U169 ( .A1(MULT_mult_6_CARRYB_22__7_), .A2(
        MULT_mult_6_ab_23__7_), .ZN(MULT_mult_6_n54) );
  NAND2_X2 MULT_mult_6_U168 ( .A1(MULT_mult_6_SUMB_3__10_), .A2(
        MULT_mult_6_CARRYB_3__9_), .ZN(MULT_mult_6_n1963) );
  NAND3_X2 MULT_mult_6_U167 ( .A1(MULT_mult_6_n1673), .A2(MULT_mult_6_n1674), 
        .A3(MULT_mult_6_n1675), .ZN(MULT_mult_6_n51) );
  INV_X4 MULT_mult_6_U166 ( .A(MULT_mult_6_n1313), .ZN(MULT_mult_6_n48) );
  INV_X4 MULT_mult_6_U165 ( .A(MULT_mult_6_CARRYB_5__7_), .ZN(MULT_mult_6_n47)
         );
  NAND2_X2 MULT_mult_6_U164 ( .A1(MULT_mult_6_n49), .A2(MULT_mult_6_n50), .ZN(
        MULT_mult_6_n1329) );
  NAND2_X4 MULT_mult_6_U163 ( .A1(MULT_mult_6_n47), .A2(MULT_mult_6_n48), .ZN(
        MULT_mult_6_n50) );
  NAND2_X1 MULT_mult_6_U162 ( .A1(MULT_mult_6_CARRYB_5__7_), .A2(
        MULT_mult_6_n1313), .ZN(MULT_mult_6_n49) );
  NAND2_X2 MULT_mult_6_U161 ( .A1(MULT_mult_6_SUMB_23__5_), .A2(
        MULT_mult_6_net84434), .ZN(MULT_mult_6_net79909) );
  NAND2_X2 MULT_mult_6_U159 ( .A1(MULT_mult_6_ab_14__3_), .A2(
        MULT_mult_6_SUMB_13__4_), .ZN(MULT_mult_6_n1968) );
  BUF_X8 MULT_mult_6_U158 ( .A(MULT_mult_6_SUMB_3__10_), .Z(MULT_mult_6_n1259)
         );
  BUF_X4 MULT_mult_6_U157 ( .A(MULT_mult_6_SUMB_4__10_), .Z(MULT_mult_6_n1258)
         );
  NAND2_X1 MULT_mult_6_U156 ( .A1(MULT_mult_6_ab_15__1_), .A2(
        MULT_mult_6_SUMB_14__2_), .ZN(MULT_mult_6_n652) );
  NAND3_X2 MULT_mult_6_U155 ( .A1(MULT_mult_6_n738), .A2(MULT_mult_6_n739), 
        .A3(MULT_mult_6_n740), .ZN(MULT_mult_6_CARRYB_11__1_) );
  INV_X1 MULT_mult_6_U154 ( .A(MULT_mult_6_net84000), .ZN(MULT_mult_6_net84434) );
  INV_X2 MULT_mult_6_U153 ( .A(MULT_mult_6_CARRYB_4__8_), .ZN(
        MULT_mult_6_n1514) );
  NAND2_X2 MULT_mult_6_U152 ( .A1(MULT_mult_6_CARRYB_1__14_), .A2(
        MULT_mult_6_ab_2__14_), .ZN(MULT_mult_6_net86172) );
  NAND2_X2 MULT_mult_6_U151 ( .A1(MULT_mult_6_ab_25__4_), .A2(
        MULT_mult_6_net90433), .ZN(MULT_mult_6_n2113) );
  INV_X8 MULT_mult_6_U150 ( .A(n5943), .ZN(MULT_mult_6_net70472) );
  XNOR2_X2 MULT_mult_6_U149 ( .A(MULT_mult_6_net93203), .B(MULT_mult_6_n1901), 
        .ZN(MULT_mult_6_SUMB_5__14_) );
  NAND2_X2 MULT_mult_6_U147 ( .A1(MULT_mult_6_n1765), .A2(
        MULT_mult_6_SUMB_2__21_), .ZN(MULT_mult_6_n1433) );
  NAND2_X4 MULT_mult_6_U146 ( .A1(MULT_mult_6_SUMB_16__9_), .A2(
        MULT_mult_6_net93410), .ZN(MULT_mult_6_n812) );
  NAND2_X4 MULT_mult_6_U145 ( .A1(MULT_mult_6_net87949), .A2(
        MULT_mult_6_net87950), .ZN(MULT_mult_6_n311) );
  INV_X4 MULT_mult_6_U144 ( .A(MULT_mult_6_CARRYB_1__18_), .ZN(
        MULT_mult_6_n709) );
  NAND2_X2 MULT_mult_6_U143 ( .A1(MULT_mult_6_n312), .A2(MULT_mult_6_ab_9__5_), 
        .ZN(MULT_mult_6_n1786) );
  NAND2_X2 MULT_mult_6_U142 ( .A1(MULT_mult_6_net93813), .A2(
        MULT_mult_6_ab_24__4_), .ZN(MULT_mult_6_net79908) );
  NAND2_X4 MULT_mult_6_U141 ( .A1(MULT_mult_6_ab_12__13_), .A2(
        MULT_mult_6_CARRYB_11__13_), .ZN(MULT_mult_6_n1795) );
  NAND2_X4 MULT_mult_6_U139 ( .A1(MULT_mult_6_n2156), .A2(MULT_mult_6_n2157), 
        .ZN(MULT_mult_6_n896) );
  NAND2_X4 MULT_mult_6_U138 ( .A1(MULT_mult_6_n1511), .A2(MULT_mult_6_n1510), 
        .ZN(MULT_mult_6_n1190) );
  NAND2_X2 MULT_mult_6_U137 ( .A1(MULT_mult_6_ab_20__9_), .A2(
        MULT_mult_6_CARRYB_19__9_), .ZN(MULT_mult_6_net81033) );
  NAND2_X4 MULT_mult_6_U136 ( .A1(MULT_mult_6_n391), .A2(MULT_mult_6_n384), 
        .ZN(MULT_mult_6_n390) );
  INV_X8 MULT_mult_6_U135 ( .A(MULT_mult_6_SUMB_12__12_), .ZN(
        MULT_mult_6_net120648) );
  NAND2_X4 MULT_mult_6_U134 ( .A1(MULT_mult_6_ab_16__9_), .A2(
        MULT_mult_6_CARRYB_15__9_), .ZN(MULT_mult_6_n805) );
  NAND3_X4 MULT_mult_6_U133 ( .A1(MULT_mult_6_net81267), .A2(
        MULT_mult_6_net81266), .A3(MULT_mult_6_net81265), .ZN(
        MULT_mult_6_net87619) );
  INV_X8 MULT_mult_6_U132 ( .A(MULT_mult_6_net88878), .ZN(
        MULT_mult_6_SUMB_18__6_) );
  XOR2_X2 MULT_mult_6_U131 ( .A(MULT_mult_6_net88881), .B(
        MULT_mult_6_ab_7__14_), .Z(MULT_mult_6_n46) );
  NAND2_X4 MULT_mult_6_U130 ( .A1(MULT_mult_6_CARRYB_15__5_), .A2(
        MULT_mult_6_ab_16__5_), .ZN(MULT_mult_6_n2071) );
  INV_X4 MULT_mult_6_U129 ( .A(MULT_mult_6_net89168), .ZN(
        MULT_mult_6_net123142) );
  NAND2_X4 MULT_mult_6_U128 ( .A1(MULT_mult_6_n1127), .A2(MULT_mult_6_n1128), 
        .ZN(MULT_mult_6_n1256) );
  NAND2_X4 MULT_mult_6_U127 ( .A1(MULT_mult_6_net85602), .A2(
        MULT_mult_6_net85603), .ZN(MULT_mult_6_SUMB_2__18_) );
  NAND2_X4 MULT_mult_6_U126 ( .A1(MULT_mult_6_CARRYB_9__9_), .A2(
        MULT_mult_6_ab_10__9_), .ZN(MULT_mult_6_n325) );
  NAND2_X4 MULT_mult_6_U125 ( .A1(MULT_mult_6_ab_2__15_), .A2(
        MULT_mult_6_CARRYB_1__15_), .ZN(MULT_mult_6_n1984) );
  INV_X8 MULT_mult_6_U124 ( .A(MULT_mult_6_n194), .ZN(MULT_mult_6_SUMB_10__6_)
         );
  NAND2_X4 MULT_mult_6_U123 ( .A1(MULT_mult_6_CARRYB_11__4_), .A2(
        MULT_mult_6_ab_12__4_), .ZN(MULT_mult_6_n667) );
  AND3_X4 MULT_mult_6_U122 ( .A1(MULT_mult_6_n2007), .A2(MULT_mult_6_n2008), 
        .A3(MULT_mult_6_n2009), .ZN(MULT_mult_6_n45) );
  INV_X8 MULT_mult_6_U121 ( .A(MULT_mult_6_n452), .ZN(
        MULT_mult_6_CARRYB_1__13_) );
  INV_X4 MULT_mult_6_U120 ( .A(MULT_mult_6_net70458), .ZN(MULT_mult_6_n491) );
  AND2_X2 MULT_mult_6_U119 ( .A1(MULT_mult_6_ab_0__28_), .A2(
        MULT_mult_6_ab_1__27_), .ZN(MULT_mult_6_n44) );
  AND2_X2 MULT_mult_6_U118 ( .A1(MULT_mult_6_ab_0__9_), .A2(
        MULT_mult_6_ab_1__8_), .ZN(MULT_mult_6_n43) );
  NAND2_X4 MULT_mult_6_U117 ( .A1(MULT_mult_6_ab_4__8_), .A2(
        MULT_mult_6_CARRYB_3__8_), .ZN(MULT_mult_6_n1944) );
  NAND2_X2 MULT_mult_6_U116 ( .A1(MULT_mult_6_ab_5__7_), .A2(
        MULT_mult_6_CARRYB_4__7_), .ZN(MULT_mult_6_n143) );
  AND2_X2 MULT_mult_6_U115 ( .A1(MULT_mult_6_ab_0__30_), .A2(
        MULT_mult_6_ab_1__29_), .ZN(MULT_mult_6_n42) );
  NOR2_X1 MULT_mult_6_U114 ( .A1(MULT_mult_6_net77898), .A2(
        MULT_mult_6_net70447), .ZN(MULT_mult_6_ab_24__5_) );
  INV_X2 MULT_mult_6_U113 ( .A(MULT_mult_6_ab_24__5_), .ZN(MULT_mult_6_n2195)
         );
  INV_X8 MULT_mult_6_U112 ( .A(MULT_mult_6_n406), .ZN(MULT_mult_6_n420) );
  NOR2_X1 MULT_mult_6_U111 ( .A1(MULT_mult_6_net77914), .A2(
        MULT_mult_6_net70451), .ZN(MULT_mult_6_ab_22__7_) );
  AND2_X2 MULT_mult_6_U110 ( .A1(MULT_mult_6_ab_0__2_), .A2(
        MULT_mult_6_ab_1__1_), .ZN(MULT_mult_6_n41) );
  XOR2_X2 MULT_mult_6_U109 ( .A(MULT_mult_6_ab_1__1_), .B(MULT_mult_6_ab_0__2_), .Z(MULT_mult_6_n40) );
  NAND2_X4 MULT_mult_6_U108 ( .A1(MULT_mult_6_ab_5__22_), .A2(
        MULT_mult_6_CARRYB_4__22_), .ZN(MULT_mult_6_net80794) );
  INV_X4 MULT_mult_6_U107 ( .A(MULT_mult_6_net92311), .ZN(
        MULT_mult_6_ab_28__2_) );
  NOR2_X2 MULT_mult_6_U106 ( .A1(MULT_mult_6_net81673), .A2(
        MULT_mult_6_net77892), .ZN(MULT_mult_6_n870) );
  AND2_X2 MULT_mult_6_U104 ( .A1(MULT_mult_6_ab_1__24_), .A2(
        MULT_mult_6_ab_0__25_), .ZN(MULT_mult_6_n39) );
  NOR2_X4 MULT_mult_6_U103 ( .A1(MULT_mult_6_net88344), .A2(
        MULT_mult_6_net77964), .ZN(MULT_mult_6_n817) );
  XNOR2_X2 MULT_mult_6_U102 ( .A(MULT_mult_6_SUMB_11__14_), .B(
        MULT_mult_6_n1753), .ZN(MULT_mult_6_n38) );
  XNOR2_X2 MULT_mult_6_U101 ( .A(MULT_mult_6_n2112), .B(
        MULT_mult_6_SUMB_5__18_), .ZN(MULT_mult_6_n37) );
  NAND3_X2 MULT_mult_6_U100 ( .A1(MULT_mult_6_n1796), .A2(MULT_mult_6_n1797), 
        .A3(MULT_mult_6_n1798), .ZN(MULT_mult_6_n36) );
  CLKBUF_X2 MULT_mult_6_U99 ( .A(MULT_mult_6_CARRYB_13__1_), .Z(
        MULT_mult_6_n35) );
  NAND2_X1 MULT_mult_6_U98 ( .A1(MULT_mult_6_ab_9__19_), .A2(
        MULT_mult_6_SUMB_8__20_), .ZN(MULT_mult_6_n2290) );
  INV_X4 MULT_mult_6_U97 ( .A(MULT_mult_6_n33), .ZN(MULT_mult_6_n34) );
  INV_X2 MULT_mult_6_U96 ( .A(MULT_mult_6_SUMB_2__23_), .ZN(MULT_mult_6_n33)
         );
  XNOR2_X2 MULT_mult_6_U95 ( .A(MULT_mult_6_SUMB_7__20_), .B(
        MULT_mult_6_net86231), .ZN(MULT_mult_6_n32) );
  INV_X8 MULT_mult_6_U94 ( .A(MULT_mult_6_n1196), .ZN(MULT_mult_6_n1197) );
  OR2_X4 MULT_mult_6_U93 ( .A1(MULT_mult_6_net70467), .A2(
        MULT_mult_6_net123000), .ZN(MULT_mult_6_n31) );
  XNOR2_X2 MULT_mult_6_U92 ( .A(MULT_mult_6_CARRYB_13__17_), .B(
        MULT_mult_6_n31), .ZN(MULT_mult_6_n1532) );
  INV_X4 MULT_mult_6_U91 ( .A(MULT_mult_6_ab_4__12_), .ZN(MULT_mult_6_n316) );
  NAND2_X1 MULT_mult_6_U90 ( .A1(MULT_mult_6_net88881), .A2(
        MULT_mult_6_SUMB_6__15_), .ZN(MULT_mult_6_net81367) );
  CLKBUF_X3 MULT_mult_6_U89 ( .A(MULT_mult_6_SUMB_6__15_), .Z(
        MULT_mult_6_net93800) );
  NAND2_X2 MULT_mult_6_U88 ( .A1(MULT_mult_6_net123897), .A2(
        MULT_mult_6_net123898), .ZN(MULT_mult_6_n872) );
  NAND2_X2 MULT_mult_6_U87 ( .A1(MULT_mult_6_n1764), .A2(MULT_mult_6_n371), 
        .ZN(MULT_mult_6_n254) );
  NAND2_X4 MULT_mult_6_U86 ( .A1(MULT_mult_6_n1024), .A2(MULT_mult_6_n1025), 
        .ZN(MULT_mult_6_n2335) );
  NAND2_X2 MULT_mult_6_U85 ( .A1(MULT_mult_6_net124949), .A2(
        MULT_mult_6_SUMB_21__4_), .ZN(MULT_mult_6_n503) );
  NAND2_X2 MULT_mult_6_U84 ( .A1(MULT_mult_6_n248), .A2(MULT_mult_6_n249), 
        .ZN(MULT_mult_6_n251) );
  NAND2_X2 MULT_mult_6_U83 ( .A1(MULT_mult_6_SUMB_2__12_), .A2(
        MULT_mult_6_CARRYB_2__11_), .ZN(MULT_mult_6_n2028) );
  INV_X8 MULT_mult_6_U82 ( .A(MULT_mult_6_net77976), .ZN(MULT_mult_6_n331) );
  NOR2_X4 MULT_mult_6_U81 ( .A1(MULT_mult_6_net70460), .A2(MULT_mult_6_n331), 
        .ZN(MULT_mult_6_net124833) );
  NOR2_X4 MULT_mult_6_U80 ( .A1(MULT_mult_6_net70450), .A2(
        MULT_mult_6_net86101), .ZN(MULT_mult_6_ab_1__8_) );
  INV_X4 MULT_mult_6_U79 ( .A(MULT_mult_6_SUMB_20__4_), .ZN(
        MULT_mult_6_net148233) );
  INV_X4 MULT_mult_6_U78 ( .A(MULT_mult_6_CARRYB_25__2_), .ZN(
        MULT_mult_6_net120359) );
  INV_X4 MULT_mult_6_U77 ( .A(MULT_mult_6_net120359), .ZN(MULT_mult_6_n30) );
  INV_X4 MULT_mult_6_U76 ( .A(MULT_mult_6_n47), .ZN(MULT_mult_6_n29) );
  INV_X2 MULT_mult_6_U75 ( .A(MULT_mult_6_CARRYB_11__6_), .ZN(
        MULT_mult_6_n1192) );
  XNOR2_X2 MULT_mult_6_U74 ( .A(MULT_mult_6_CARRYB_26__0_), .B(
        MULT_mult_6_ab_27__0_), .ZN(MULT_mult_6_n192) );
  INV_X4 MULT_mult_6_U73 ( .A(MULT_mult_6_n940), .ZN(MULT_mult_6_n28) );
  XNOR2_X2 MULT_mult_6_U72 ( .A(MULT_mult_6_n28), .B(MULT_mult_6_ab_26__0_), 
        .ZN(MULT_mult_6_n2026) );
  NAND2_X2 MULT_mult_6_U71 ( .A1(MULT_mult_6_n1973), .A2(MULT_mult_6_n1308), 
        .ZN(MULT_mult_6_n226) );
  INV_X8 MULT_mult_6_U70 ( .A(MULT_mult_6_net70491), .ZN(MULT_mult_6_net77976)
         );
  XNOR2_X2 MULT_mult_6_U69 ( .A(MULT_mult_6_CARRYB_24__0_), .B(
        MULT_mult_6_ab_25__0_), .ZN(MULT_mult_6_n27) );
  XNOR2_X2 MULT_mult_6_U68 ( .A(MULT_mult_6_n27), .B(MULT_mult_6_n597), .ZN(
        multOut[6]) );
  XNOR2_X2 MULT_mult_6_U66 ( .A(MULT_mult_6_n2026), .B(MULT_mult_6_n1134), 
        .ZN(multOut[5]) );
  XNOR2_X2 MULT_mult_6_U64 ( .A(MULT_mult_6_n2171), .B(MULT_mult_6_net122087), 
        .ZN(MULT_mult_6_n25) );
  CLKBUF_X2 MULT_mult_6_U63 ( .A(MULT_mult_6_SUMB_18__3_), .Z(MULT_mult_6_n24)
         );
  XNOR2_X2 MULT_mult_6_U62 ( .A(MULT_mult_6_net93713), .B(MULT_mult_6_net83358), .ZN(MULT_mult_6_n23) );
  XNOR2_X2 MULT_mult_6_U61 ( .A(MULT_mult_6_SUMB_22__1_), .B(
        MULT_mult_6_ab_23__0_), .ZN(MULT_mult_6_n22) );
  XNOR2_X2 MULT_mult_6_U60 ( .A(MULT_mult_6_n22), .B(MULT_mult_6_n963), .ZN(
        multOut[8]) );
  INV_X4 MULT_mult_6_U59 ( .A(MULT_mult_6_n962), .ZN(MULT_mult_6_n963) );
  NAND2_X2 MULT_mult_6_U58 ( .A1(MULT_mult_6_CARRYB_21__0_), .A2(
        MULT_mult_6_SUMB_21__1_), .ZN(MULT_mult_6_n1798) );
  NAND3_X4 MULT_mult_6_U57 ( .A1(MULT_mult_6_n732), .A2(MULT_mult_6_n733), 
        .A3(MULT_mult_6_n734), .ZN(MULT_mult_6_CARRYB_3__5_) );
  INV_X2 MULT_mult_6_U56 ( .A(MULT_mult_6_n36), .ZN(MULT_mult_6_n962) );
  XNOR2_X2 MULT_mult_6_U55 ( .A(MULT_mult_6_SUMB_17__2_), .B(
        MULT_mult_6_ab_18__1_), .ZN(MULT_mult_6_n396) );
  INV_X4 MULT_mult_6_U54 ( .A(MULT_mult_6_SUMB_19__2_), .ZN(MULT_mult_6_n21)
         );
  XNOR2_X2 MULT_mult_6_U53 ( .A(MULT_mult_6_n425), .B(MULT_mult_6_n21), .ZN(
        MULT_mult_6_SUMB_20__1_) );
  NAND2_X2 MULT_mult_6_U52 ( .A1(MULT_mult_6_ab_6__3_), .A2(
        MULT_mult_6_CARRYB_5__3_), .ZN(MULT_mult_6_n1566) );
  NAND2_X2 MULT_mult_6_U51 ( .A1(MULT_mult_6_CARRYB_19__2_), .A2(
        MULT_mult_6_SUMB_19__3_), .ZN(MULT_mult_6_n1916) );
  NAND2_X2 MULT_mult_6_U50 ( .A1(MULT_mult_6_CARRYB_13__4_), .A2(
        MULT_mult_6_SUMB_13__5_), .ZN(MULT_mult_6_n2150) );
  CLKBUF_X2 MULT_mult_6_U49 ( .A(MULT_mult_6_CARRYB_19__2_), .Z(
        MULT_mult_6_n20) );
  NAND3_X2 MULT_mult_6_U48 ( .A1(MULT_mult_6_n1995), .A2(MULT_mult_6_n1996), 
        .A3(MULT_mult_6_n1997), .ZN(MULT_mult_6_n19) );
  XNOR2_X2 MULT_mult_6_U47 ( .A(MULT_mult_6_ab_22__0_), .B(
        MULT_mult_6_CARRYB_21__0_), .ZN(MULT_mult_6_n18) );
  XNOR2_X2 MULT_mult_6_U46 ( .A(MULT_mult_6_n18), .B(MULT_mult_6_n1280), .ZN(
        multOut[9]) );
  XOR2_X2 MULT_mult_6_U45 ( .A(MULT_mult_6_n1808), .B(MULT_mult_6_n16), .Z(
        multOut[13]) );
  NAND2_X2 MULT_mult_6_U44 ( .A1(MULT_mult_6_CARRYB_13__2_), .A2(
        MULT_mult_6_SUMB_13__3_), .ZN(MULT_mult_6_net81781) );
  NAND3_X2 MULT_mult_6_U43 ( .A1(MULT_mult_6_n1969), .A2(MULT_mult_6_n1968), 
        .A3(MULT_mult_6_n1967), .ZN(MULT_mult_6_n17) );
  CLKBUF_X3 MULT_mult_6_U42 ( .A(MULT_mult_6_SUMB_17__1_), .Z(MULT_mult_6_n16)
         );
  XNOR2_X2 MULT_mult_6_U41 ( .A(MULT_mult_6_n360), .B(MULT_mult_6_SUMB_20__1_), 
        .ZN(multOut[10]) );
  INV_X2 MULT_mult_6_U39 ( .A(MULT_mult_6_net89110), .ZN(MULT_mult_6_net148015) );
  NAND2_X2 MULT_mult_6_U38 ( .A1(MULT_mult_6_net82255), .A2(
        MULT_mult_6_SUMB_19__10_), .ZN(MULT_mult_6_net81035) );
  INV_X16 MULT_mult_6_U37 ( .A(n5851), .ZN(MULT_mult_6_net70466) );
  INV_X4 MULT_mult_6_U36 ( .A(MULT_mult_6_net85287), .ZN(MULT_mult_6_n13) );
  NAND2_X4 MULT_mult_6_U34 ( .A1(MULT_mult_6_n14), .A2(MULT_mult_6_n15), .ZN(
        MULT_mult_6_net86792) );
  NAND2_X4 MULT_mult_6_U33 ( .A1(MULT_mult_6_n12), .A2(MULT_mult_6_n13), .ZN(
        MULT_mult_6_n15) );
  NAND2_X2 MULT_mult_6_U32 ( .A1(MULT_mult_6_n476), .A2(MULT_mult_6_net85287), 
        .ZN(MULT_mult_6_n14) );
  NAND2_X4 MULT_mult_6_U31 ( .A1(MULT_mult_6_net148302), .A2(
        MULT_mult_6_net149605), .ZN(MULT_mult_6_n626) );
  INV_X32 MULT_mult_6_U28 ( .A(MULT_mult_6_ab_25__2_), .ZN(MULT_mult_6_n10) );
  XNOR2_X2 MULT_mult_6_U27 ( .A(MULT_mult_6_CARRYB_24__2_), .B(MULT_mult_6_n10), .ZN(MULT_mult_6_n9) );
  CLKBUF_X3 MULT_mult_6_U26 ( .A(MULT_mult_6_net87411), .Z(
        MULT_mult_6_net86385) );
  NAND2_X2 MULT_mult_6_U25 ( .A1(MULT_mult_6_ab_3__22_), .A2(
        MULT_mult_6_CARRYB_2__22_), .ZN(MULT_mult_6_n1068) );
  INV_X8 MULT_mult_6_U24 ( .A(MULT_mult_6_CARRYB_3__16_), .ZN(MULT_mult_6_n654) );
  INV_X4 MULT_mult_6_U23 ( .A(MULT_mult_6_n7), .ZN(MULT_mult_6_n8) );
  INV_X2 MULT_mult_6_U22 ( .A(MULT_mult_6_SUMB_18__6_), .ZN(MULT_mult_6_n7) );
  NAND2_X2 MULT_mult_6_U21 ( .A1(MULT_mult_6_n1323), .A2(
        MULT_mult_6_SUMB_12__14_), .ZN(MULT_mult_6_n87) );
  NAND2_X4 MULT_mult_6_U20 ( .A1(MULT_mult_6_net123303), .A2(
        MULT_mult_6_ab_4__16_), .ZN(MULT_mult_6_net80835) );
  NAND2_X2 MULT_mult_6_U19 ( .A1(MULT_mult_6_CARRYB_24__3_), .A2(
        MULT_mult_6_ab_25__3_), .ZN(MULT_mult_6_net81007) );
  INV_X2 MULT_mult_6_U18 ( .A(MULT_mult_6_CARRYB_24__3_), .ZN(
        MULT_mult_6_net121450) );
  INV_X8 MULT_mult_6_U16 ( .A(MULT_mult_6_CARRYB_8__9_), .ZN(MULT_mult_6_n1172) );
  INV_X2 MULT_mult_6_U14 ( .A(MULT_mult_6_n5), .ZN(MULT_mult_6_n6) );
  INV_X2 MULT_mult_6_U13 ( .A(MULT_mult_6_CARRYB_16__7_), .ZN(MULT_mult_6_n5)
         );
  NAND2_X2 MULT_mult_6_U12 ( .A1(MULT_mult_6_n399), .A2(MULT_mult_6_net86629), 
        .ZN(MULT_mult_6_n1412) );
  NAND2_X1 MULT_mult_6_U11 ( .A1(MULT_mult_6_ab_23__7_), .A2(MULT_mult_6_n949), 
        .ZN(MULT_mult_6_net86413) );
  NAND2_X2 MULT_mult_6_U10 ( .A1(MULT_mult_6_ab_5__17_), .A2(
        MULT_mult_6_SUMB_4__18_), .ZN(MULT_mult_6_n2202) );
  NAND2_X4 MULT_mult_6_U9 ( .A1(MULT_mult_6_n534), .A2(MULT_mult_6_n535), .ZN(
        MULT_mult_6_n4) );
  NAND2_X2 MULT_mult_6_U8 ( .A1(MULT_mult_6_net86024), .A2(
        MULT_mult_6_net86023), .ZN(MULT_mult_6_n3) );
  NAND2_X2 MULT_mult_6_U7 ( .A1(MULT_mult_6_CARRYB_29__1_), .A2(
        MULT_mult_6_net81548), .ZN(MULT_mult_6_n836) );
  NAND2_X2 MULT_mult_6_U6 ( .A1(MULT_mult_6_net123427), .A2(
        MULT_mult_6_ab_26__3_), .ZN(MULT_mult_6_n2116) );
  NAND2_X2 MULT_mult_6_U5 ( .A1(MULT_mult_6_SUMB_13__11_), .A2(
        MULT_mult_6_CARRYB_13__10_), .ZN(MULT_mult_6_net82162) );
  NAND2_X2 MULT_mult_6_U4 ( .A1(MULT_mult_6_net89453), .A2(
        MULT_mult_6_ab_30__0_), .ZN(MULT_mult_6_net80473) );
  INV_X2 MULT_mult_6_U3 ( .A(MULT_mult_6_net85094), .ZN(MULT_mult_6_net148179)
         );
  INV_X4 MULT_mult_6_U2 ( .A(MULT_mult_6_CARRYB_10__12_), .ZN(
        MULT_mult_6_net83629) );
  FA_X1 MULT_mult_6_S2_14_8 ( .A(MULT_mult_6_SUMB_13__9_), .B(
        MULT_mult_6_ab_14__8_), .CI(MULT_mult_6_CARRYB_13__8_), .CO(
        MULT_mult_6_CARRYB_14__8_), .S(MULT_mult_6_SUMB_14__8_) );
  FA_X1 MULT_mult_6_S2_17_6 ( .A(MULT_mult_6_CARRYB_16__6_), .B(
        MULT_mult_6_ab_17__6_), .CI(MULT_mult_6_SUMB_16__7_), .CO(
        MULT_mult_6_CARRYB_17__6_), .S(MULT_mult_6_SUMB_17__6_) );
  FA_X1 MULT_mult_6_S2_22_5 ( .A(MULT_mult_6_CARRYB_21__5_), .B(
        MULT_mult_6_ab_22__5_), .CI(MULT_mult_6_SUMB_21__6_), .CO(
        MULT_mult_6_CARRYB_22__5_), .S(MULT_mult_6_SUMB_22__5_) );
  FA_X1 MULT_mult_6_S2_6_14 ( .A(MULT_mult_6_SUMB_5__15_), .B(
        MULT_mult_6_ab_6__14_), .CI(MULT_mult_6_CARRYB_5__14_), .CO(
        MULT_mult_6_CARRYB_6__14_), .S(MULT_mult_6_SUMB_6__14_) );
  FA_X1 MULT_mult_6_S2_20_3 ( .A(MULT_mult_6_SUMB_19__4_), .B(
        MULT_mult_6_ab_20__3_), .CI(MULT_mult_6_CARRYB_19__3_), .CO(
        MULT_mult_6_CARRYB_20__3_), .S(MULT_mult_6_SUMB_20__3_) );
  FA_X1 MULT_mult_6_S2_2_7 ( .A(MULT_mult_6_ab_2__7_), .B(
        MULT_mult_6_CARRYB_1__7_), .CI(MULT_mult_6_SUMB_1__8_), .CO(
        MULT_mult_6_CARRYB_2__7_), .S(MULT_mult_6_SUMB_2__7_) );
  FA_X1 MULT_mult_6_S2_12_1 ( .A(MULT_mult_6_ab_12__1_), .B(
        MULT_mult_6_CARRYB_11__1_), .CI(MULT_mult_6_SUMB_11__2_), .CO(
        MULT_mult_6_CARRYB_12__1_), .S(MULT_mult_6_SUMB_12__1_) );
  FA_X1 MULT_mult_6_S2_7_4 ( .A(MULT_mult_6_ab_7__4_), .B(
        MULT_mult_6_CARRYB_6__4_), .CI(MULT_mult_6_SUMB_6__5_), .CO(
        MULT_mult_6_CARRYB_7__4_), .S(MULT_mult_6_SUMB_7__4_) );
  FA_X1 MULT_mult_6_S2_8_3 ( .A(MULT_mult_6_ab_8__3_), .B(
        MULT_mult_6_CARRYB_7__3_), .CI(MULT_mult_6_SUMB_7__4_), .CO(
        MULT_mult_6_CARRYB_8__3_), .S(MULT_mult_6_SUMB_8__3_) );
  FA_X1 MULT_mult_6_S2_12_15 ( .A(MULT_mult_6_CARRYB_11__15_), .B(
        MULT_mult_6_ab_12__15_), .CI(MULT_mult_6_SUMB_11__16_), .CO(
        MULT_mult_6_CARRYB_12__15_), .S(MULT_mult_6_SUMB_12__15_) );
  FA_X1 MULT_mult_6_S2_6_21 ( .A(MULT_mult_6_CARRYB_5__21_), .B(
        MULT_mult_6_ab_6__21_), .CI(MULT_mult_6_SUMB_5__22_), .CO(
        MULT_mult_6_CARRYB_6__21_), .S(MULT_mult_6_SUMB_6__21_) );
  FA_X1 MULT_mult_6_S2_2_29 ( .A(MULT_mult_6_ab_2__29_), .B(MULT_mult_6_n42), 
        .CI(MULT_mult_6_n355), .S(MULT_mult_6_SUMB_2__29_) );
  FA_X1 MULT_mult_6_S2_2_27 ( .A(MULT_mult_6_ab_2__27_), .B(MULT_mult_6_n44), 
        .CI(MULT_mult_6_SUMB_1__28_), .CO(MULT_mult_6_CARRYB_2__27_), .S(
        MULT_mult_6_SUMB_2__27_) );
  FA_X1 MULT_mult_6_S2_2_26 ( .A(MULT_mult_6_ab_2__26_), .B(
        MULT_mult_6_CARRYB_1__26_), .CI(MULT_mult_6_SUMB_1__27_), .CO(
        MULT_mult_6_CARRYB_2__26_), .S(MULT_mult_6_SUMB_2__26_) );
  FA_X1 MULT_mult_6_S2_2_9 ( .A(MULT_mult_6_ab_2__9_), .B(
        MULT_mult_6_CARRYB_1__9_), .CI(MULT_mult_6_SUMB_1__10_), .CO(
        MULT_mult_6_CARRYB_2__9_), .S(MULT_mult_6_SUMB_2__9_) );
  FA_X1 MULT_mult_6_S2_2_8 ( .A(MULT_mult_6_ab_2__8_), .B(MULT_mult_6_n43), 
        .CI(MULT_mult_6_SUMB_1__9_), .CO(MULT_mult_6_CARRYB_2__8_), .S(
        MULT_mult_6_SUMB_2__8_) );
  FA_X1 MULT_mult_6_S2_2_2 ( .A(MULT_mult_6_ab_2__2_), .B(
        MULT_mult_6_CARRYB_1__2_), .CI(MULT_mult_6_SUMB_1__3_), .CO(
        MULT_mult_6_CARRYB_2__2_), .S(MULT_mult_6_SUMB_2__2_) );
  FA_X1 MULT_mult_6_S2_2_1 ( .A(MULT_mult_6_ab_2__1_), .B(MULT_mult_6_n41), 
        .CI(MULT_mult_6_SUMB_1__2_), .CO(MULT_mult_6_CARRYB_2__1_), .S(
        MULT_mult_6_SUMB_2__1_) );
  FA_X1 MULT_mult_6_S1_2_0 ( .A(MULT_mult_6_ab_2__0_), .B(
        MULT_mult_6_CARRYB_1__0_), .CI(MULT_mult_6_n40), .CO(
        MULT_mult_6_CARRYB_2__0_), .S(multOut[29]) );
  FA_X1 MULT_mult_6_S2_3_28 ( .A(MULT_mult_6_ab_3__28_), .B(
        MULT_mult_6_CARRYB_2__28_), .CI(MULT_mult_6_SUMB_2__29_), .S(
        MULT_mult_6_SUMB_3__28_) );
  FA_X1 MULT_mult_6_S2_3_3 ( .A(MULT_mult_6_ab_3__3_), .B(
        MULT_mult_6_CARRYB_2__3_), .CI(MULT_mult_6_SUMB_2__4_), .CO(
        MULT_mult_6_CARRYB_3__3_), .S(MULT_mult_6_SUMB_3__3_) );
  FA_X1 MULT_mult_6_S2_3_2 ( .A(MULT_mult_6_CARRYB_2__2_), .B(
        MULT_mult_6_ab_3__2_), .CI(MULT_mult_6_SUMB_2__3_), .CO(
        MULT_mult_6_CARRYB_3__2_), .S(MULT_mult_6_SUMB_3__2_) );
  FA_X1 MULT_mult_6_S2_3_1 ( .A(MULT_mult_6_ab_3__1_), .B(
        MULT_mult_6_CARRYB_2__1_), .CI(MULT_mult_6_SUMB_2__2_), .CO(
        MULT_mult_6_CARRYB_3__1_), .S(MULT_mult_6_SUMB_3__1_) );
  FA_X1 MULT_mult_6_S1_3_0 ( .A(MULT_mult_6_ab_3__0_), .B(
        MULT_mult_6_CARRYB_2__0_), .CI(MULT_mult_6_SUMB_2__1_), .CO(
        MULT_mult_6_CARRYB_3__0_), .S(multOut[28]) );
  FA_X1 MULT_mult_6_S2_4_26 ( .A(MULT_mult_6_ab_4__26_), .B(
        MULT_mult_6_CARRYB_3__26_), .CI(MULT_mult_6_SUMB_3__27_), .CO(
        MULT_mult_6_CARRYB_4__26_), .S(MULT_mult_6_SUMB_4__26_) );
  FA_X1 MULT_mult_6_S2_4_4 ( .A(MULT_mult_6_ab_4__4_), .B(
        MULT_mult_6_CARRYB_3__4_), .CI(MULT_mult_6_SUMB_3__5_), .CO(
        MULT_mult_6_CARRYB_4__4_), .S(MULT_mult_6_SUMB_4__4_) );
  FA_X1 MULT_mult_6_S2_4_3 ( .A(MULT_mult_6_ab_4__3_), .B(
        MULT_mult_6_CARRYB_3__3_), .CI(MULT_mult_6_SUMB_3__4_), .CO(
        MULT_mult_6_CARRYB_4__3_), .S(MULT_mult_6_SUMB_4__3_) );
  FA_X1 MULT_mult_6_S2_4_2 ( .A(MULT_mult_6_CARRYB_3__2_), .B(
        MULT_mult_6_ab_4__2_), .CI(MULT_mult_6_SUMB_3__3_), .CO(
        MULT_mult_6_CARRYB_4__2_), .S(MULT_mult_6_SUMB_4__2_) );
  FA_X1 MULT_mult_6_S1_4_0 ( .A(MULT_mult_6_CARRYB_3__0_), .B(
        MULT_mult_6_ab_4__0_), .CI(MULT_mult_6_SUMB_3__1_), .CO(
        MULT_mult_6_CARRYB_4__0_), .S(multOut[27]) );
  FA_X1 MULT_mult_6_S2_5_24 ( .A(MULT_mult_6_ab_5__24_), .B(
        MULT_mult_6_CARRYB_4__24_), .CI(MULT_mult_6_n1185), .CO(
        MULT_mult_6_CARRYB_5__24_), .S(MULT_mult_6_SUMB_5__24_) );
  FA_X1 MULT_mult_6_S2_5_6 ( .A(MULT_mult_6_CARRYB_4__6_), .B(
        MULT_mult_6_ab_5__6_), .CI(MULT_mult_6_SUMB_4__7_), .CO(
        MULT_mult_6_CARRYB_5__6_), .S(MULT_mult_6_SUMB_5__6_) );
  FA_X1 MULT_mult_6_S2_5_4 ( .A(MULT_mult_6_CARRYB_4__4_), .B(
        MULT_mult_6_ab_5__4_), .CI(MULT_mult_6_SUMB_4__5_), .CO(
        MULT_mult_6_CARRYB_5__4_), .S(MULT_mult_6_SUMB_5__4_) );
  FA_X1 MULT_mult_6_S2_5_3 ( .A(MULT_mult_6_ab_5__3_), .B(
        MULT_mult_6_CARRYB_4__3_), .CI(MULT_mult_6_SUMB_4__4_), .CO(
        MULT_mult_6_CARRYB_5__3_), .S(MULT_mult_6_SUMB_5__3_) );
  FA_X1 MULT_mult_6_S2_5_2 ( .A(MULT_mult_6_CARRYB_4__2_), .B(
        MULT_mult_6_ab_5__2_), .CI(MULT_mult_6_SUMB_4__3_), .CO(
        MULT_mult_6_CARRYB_5__2_), .S(MULT_mult_6_SUMB_5__2_) );
  FA_X1 MULT_mult_6_S1_5_0 ( .A(MULT_mult_6_ab_5__0_), .B(
        MULT_mult_6_CARRYB_4__0_), .CI(MULT_mult_6_SUMB_4__1_), .CO(
        MULT_mult_6_CARRYB_5__0_), .S(multOut[26]) );
  FA_X1 MULT_mult_6_S2_6_22 ( .A(MULT_mult_6_CARRYB_5__22_), .B(
        MULT_mult_6_ab_6__22_), .CI(MULT_mult_6_SUMB_5__23_), .CO(
        MULT_mult_6_CARRYB_6__22_), .S(MULT_mult_6_SUMB_6__22_) );
  FA_X1 MULT_mult_6_S2_6_9 ( .A(MULT_mult_6_CARRYB_5__9_), .B(
        MULT_mult_6_ab_6__9_), .CI(MULT_mult_6_SUMB_5__10_), .CO(
        MULT_mult_6_CARRYB_6__9_), .S(MULT_mult_6_SUMB_6__9_) );
  FA_X1 MULT_mult_6_S2_6_2 ( .A(MULT_mult_6_ab_6__2_), .B(
        MULT_mult_6_CARRYB_5__2_), .CI(MULT_mult_6_SUMB_5__3_), .CO(
        MULT_mult_6_CARRYB_6__2_), .S(MULT_mult_6_SUMB_6__2_) );
  FA_X1 MULT_mult_6_S1_6_0 ( .A(MULT_mult_6_ab_6__0_), .B(
        MULT_mult_6_CARRYB_5__0_), .CI(MULT_mult_6_SUMB_5__1_), .CO(
        MULT_mult_6_CARRYB_6__0_), .S(multOut[25]) );
  FA_X1 MULT_mult_6_S2_7_24 ( .A(MULT_mult_6_ab_7__24_), .B(
        MULT_mult_6_CARRYB_6__24_), .CI(MULT_mult_6_SUMB_6__25_), .S(
        MULT_mult_6_SUMB_7__24_) );
  FA_X1 MULT_mult_6_S2_7_2 ( .A(MULT_mult_6_CARRYB_6__2_), .B(
        MULT_mult_6_ab_7__2_), .CI(MULT_mult_6_SUMB_6__3_), .CO(
        MULT_mult_6_CARRYB_7__2_), .S(MULT_mult_6_SUMB_7__2_) );
  FA_X1 MULT_mult_6_S1_7_0 ( .A(MULT_mult_6_ab_7__0_), .B(
        MULT_mult_6_SUMB_6__1_), .CI(MULT_mult_6_CARRYB_6__0_), .CO(
        MULT_mult_6_CARRYB_7__0_), .S(multOut[24]) );
  FA_X1 MULT_mult_6_S2_8_23 ( .A(MULT_mult_6_ab_8__23_), .B(
        MULT_mult_6_CARRYB_7__23_), .CI(MULT_mult_6_SUMB_7__24_), .S(
        MULT_mult_6_SUMB_8__23_) );
  FA_X1 MULT_mult_6_S2_8_21 ( .A(MULT_mult_6_ab_8__21_), .B(
        MULT_mult_6_CARRYB_7__21_), .CI(MULT_mult_6_SUMB_7__22_), .CO(
        MULT_mult_6_CARRYB_8__21_), .S(MULT_mult_6_SUMB_8__21_) );
  FA_X1 MULT_mult_6_S2_8_5 ( .A(MULT_mult_6_CARRYB_7__5_), .B(
        MULT_mult_6_ab_8__5_), .CI(MULT_mult_6_n2375), .CO(
        MULT_mult_6_CARRYB_8__5_), .S(MULT_mult_6_SUMB_8__5_) );
  FA_X1 MULT_mult_6_S2_8_2 ( .A(MULT_mult_6_CARRYB_7__2_), .B(
        MULT_mult_6_ab_8__2_), .CI(MULT_mult_6_SUMB_7__3_), .CO(
        MULT_mult_6_CARRYB_8__2_), .S(MULT_mult_6_SUMB_8__2_) );
  FA_X1 MULT_mult_6_S1_8_0 ( .A(MULT_mult_6_ab_8__0_), .B(
        MULT_mult_6_CARRYB_7__0_), .CI(MULT_mult_6_SUMB_7__1_), .CO(
        MULT_mult_6_CARRYB_8__0_), .S(multOut[23]) );
  FA_X1 MULT_mult_6_S2_9_1 ( .A(MULT_mult_6_ab_9__1_), .B(
        MULT_mult_6_CARRYB_8__1_), .CI(MULT_mult_6_SUMB_8__2_), .CO(
        MULT_mult_6_CARRYB_9__1_), .S(MULT_mult_6_SUMB_9__1_) );
  FA_X1 MULT_mult_6_S1_9_0 ( .A(MULT_mult_6_ab_9__0_), .B(
        MULT_mult_6_CARRYB_8__0_), .CI(MULT_mult_6_SUMB_8__1_), .CO(
        MULT_mult_6_CARRYB_9__0_), .S(multOut[22]) );
  FA_X1 MULT_mult_6_S2_10_7 ( .A(MULT_mult_6_CARRYB_9__7_), .B(
        MULT_mult_6_ab_10__7_), .CI(MULT_mult_6_SUMB_9__8_), .CO(
        MULT_mult_6_CARRYB_10__7_), .S(MULT_mult_6_SUMB_10__7_) );
  FA_X1 MULT_mult_6_S2_10_5 ( .A(MULT_mult_6_CARRYB_9__5_), .B(
        MULT_mult_6_ab_10__5_), .CI(MULT_mult_6_SUMB_9__6_), .CO(
        MULT_mult_6_CARRYB_10__5_), .S(MULT_mult_6_SUMB_10__5_) );
  FA_X1 MULT_mult_6_S1_10_0 ( .A(MULT_mult_6_ab_10__0_), .B(
        MULT_mult_6_CARRYB_9__0_), .CI(MULT_mult_6_SUMB_9__1_), .CO(
        MULT_mult_6_CARRYB_10__0_), .S(multOut[21]) );
  FA_X1 MULT_mult_6_S2_11_19 ( .A(MULT_mult_6_ab_11__19_), .B(
        MULT_mult_6_CARRYB_10__19_), .CI(MULT_mult_6_SUMB_10__20_), .CO(
        MULT_mult_6_CARRYB_11__19_), .S(MULT_mult_6_SUMB_11__19_) );
  FA_X1 MULT_mult_6_S2_11_6 ( .A(MULT_mult_6_CARRYB_10__6_), .B(
        MULT_mult_6_ab_11__6_), .CI(MULT_mult_6_SUMB_10__7_), .CO(
        MULT_mult_6_CARRYB_11__6_), .S(MULT_mult_6_SUMB_11__6_) );
  FA_X1 MULT_mult_6_S2_12_19 ( .A(MULT_mult_6_ab_12__19_), .B(
        MULT_mult_6_CARRYB_11__19_), .CI(MULT_mult_6_SUMB_11__20_), .S(
        MULT_mult_6_SUMB_12__19_) );
  FA_X1 MULT_mult_6_S2_12_18 ( .A(MULT_mult_6_ab_12__18_), .B(
        MULT_mult_6_CARRYB_11__18_), .CI(MULT_mult_6_SUMB_11__19_), .CO(
        MULT_mult_6_CARRYB_12__18_), .S(MULT_mult_6_SUMB_12__18_) );
  FA_X1 MULT_mult_6_S2_13_18 ( .A(MULT_mult_6_ab_13__18_), .B(
        MULT_mult_6_CARRYB_12__18_), .CI(MULT_mult_6_SUMB_12__19_), .S(
        MULT_mult_6_SUMB_13__18_) );
endmodule

