
module pipeline_processor ( clk, reset, DMEM_BUS_OUT, DMEM_BUS_IN, 
        IMEM_BUS_OUT, IMEM_BUS_IN );
  output [0:66] DMEM_BUS_OUT;
  input [0:31] DMEM_BUS_IN;
  output [0:31] IMEM_BUS_OUT;
  input [0:31] IMEM_BUS_IN;
  input clk, reset;
  wire   EXEC_MEM_OUT_109, EXEC_MEM_OUT_110, EXEC_MEM_OUT_111,
         EXEC_MEM_OUT_112, EXEC_MEM_OUT_113, EXEC_MEM_OUT_114,
         EXEC_MEM_OUT_115, EXEC_MEM_OUT_116, EXEC_MEM_OUT_117,
         EXEC_MEM_OUT_118, EXEC_MEM_OUT_119, EXEC_MEM_OUT_120,
         EXEC_MEM_OUT_121, EXEC_MEM_OUT_122, EXEC_MEM_OUT_123,
         EXEC_MEM_OUT_124, EXEC_MEM_OUT_125, EXEC_MEM_OUT_126,
         EXEC_MEM_OUT_127, EXEC_MEM_OUT_128, EXEC_MEM_OUT_129,
         EXEC_MEM_OUT_130, EXEC_MEM_OUT_131, EXEC_MEM_OUT_132,
         EXEC_MEM_OUT_133, EXEC_MEM_OUT_134, EXEC_MEM_OUT_135,
         EXEC_MEM_OUT_136, EXEC_MEM_OUT_137, EXEC_MEM_OUT_138,
         EXEC_MEM_OUT_141, RegWrite_wb_out, IF_ID_REG_IF_ID_REG_N36,
         IF_ID_REG_IF_ID_REG_N35, IF_ID_REG_IF_ID_REG_N34,
         IF_ID_REG_IF_ID_REG_N33, IF_ID_REG_IF_ID_REG_N32,
         IF_ID_REG_IF_ID_REG_N31, IF_ID_REG_IF_ID_REG_N30,
         IF_ID_REG_IF_ID_REG_N29, IF_ID_REG_IF_ID_REG_N28,
         IF_ID_REG_IF_ID_REG_N27, IF_ID_REG_IF_ID_REG_N26,
         IF_ID_REG_IF_ID_REG_N25, IF_ID_REG_IF_ID_REG_N24,
         IF_ID_REG_IF_ID_REG_N23, IF_ID_REG_IF_ID_REG_N22,
         IF_ID_REG_IF_ID_REG_N21, IF_ID_REG_IF_ID_REG_N20,
         IF_ID_REG_IF_ID_REG_N19, IF_ID_REG_IF_ID_REG_N18,
         IF_ID_REG_IF_ID_REG_N17, IF_ID_REG_IF_ID_REG_N16,
         IF_ID_REG_IF_ID_REG_N15, IF_ID_REG_IF_ID_REG_N14,
         IF_ID_REG_IF_ID_REG_N13, IF_ID_REG_IF_ID_REG_N12,
         IF_ID_REG_IF_ID_REG_N11, IF_ID_REG_IF_ID_REG_N10,
         IF_ID_REG_IF_ID_REG_N9, IF_ID_REG_IF_ID_REG_N8,
         IF_ID_REG_IF_ID_REG_N7, IF_ID_REG_IF_ID_REG_N6,
         IF_ID_REG_IF_ID_REG_N5, IF_ID_REG_IF_ID_REG_N4,
         IF_ID_REG_IF_ID_REG_N3, ID_EX_REG_ID_EX_REG_N206,
         ID_EX_REG_ID_EX_REG_N205, ID_EX_REG_ID_EX_REG_N204,
         ID_EX_REG_ID_EX_REG_N203, ID_EX_REG_ID_EX_REG_N202,
         ID_EX_REG_ID_EX_REG_N201, ID_EX_REG_ID_EX_REG_N200,
         ID_EX_REG_ID_EX_REG_N199, ID_EX_REG_ID_EX_REG_N198,
         ID_EX_REG_ID_EX_REG_N197, ID_EX_REG_ID_EX_REG_N196,
         ID_EX_REG_ID_EX_REG_N195, ID_EX_REG_ID_EX_REG_N194,
         ID_EX_REG_ID_EX_REG_N193, ID_EX_REG_ID_EX_REG_N192,
         ID_EX_REG_ID_EX_REG_N191, ID_EX_REG_ID_EX_REG_N190,
         ID_EX_REG_ID_EX_REG_N189, ID_EX_REG_ID_EX_REG_N188,
         ID_EX_REG_ID_EX_REG_N187, ID_EX_REG_ID_EX_REG_N186,
         ID_EX_REG_ID_EX_REG_N185, ID_EX_REG_ID_EX_REG_N184,
         ID_EX_REG_ID_EX_REG_N183, ID_EX_REG_ID_EX_REG_N182,
         ID_EX_REG_ID_EX_REG_N181, ID_EX_REG_ID_EX_REG_N180,
         ID_EX_REG_ID_EX_REG_N179, ID_EX_REG_ID_EX_REG_N178,
         ID_EX_REG_ID_EX_REG_N177, ID_EX_REG_ID_EX_REG_N176,
         ID_EX_REG_ID_EX_REG_N175, ID_EX_REG_ID_EX_REG_N174,
         ID_EX_REG_ID_EX_REG_N173, ID_EX_REG_ID_EX_REG_N172,
         ID_EX_REG_ID_EX_REG_N171, ID_EX_REG_ID_EX_REG_N170,
         ID_EX_REG_ID_EX_REG_N169, ID_EX_REG_ID_EX_REG_N168,
         ID_EX_REG_ID_EX_REG_N167, ID_EX_REG_ID_EX_REG_N166,
         ID_EX_REG_ID_EX_REG_N165, ID_EX_REG_ID_EX_REG_N164,
         ID_EX_REG_ID_EX_REG_N163, ID_EX_REG_ID_EX_REG_N162,
         ID_EX_REG_ID_EX_REG_N161, ID_EX_REG_ID_EX_REG_N160,
         ID_EX_REG_ID_EX_REG_N159, ID_EX_REG_ID_EX_REG_N158,
         ID_EX_REG_ID_EX_REG_N157, ID_EX_REG_ID_EX_REG_N156,
         ID_EX_REG_ID_EX_REG_N155, ID_EX_REG_ID_EX_REG_N154,
         ID_EX_REG_ID_EX_REG_N153, ID_EX_REG_ID_EX_REG_N152,
         ID_EX_REG_ID_EX_REG_N151, ID_EX_REG_ID_EX_REG_N150,
         ID_EX_REG_ID_EX_REG_N149, ID_EX_REG_ID_EX_REG_N148,
         ID_EX_REG_ID_EX_REG_N147, ID_EX_REG_ID_EX_REG_N146,
         ID_EX_REG_ID_EX_REG_N145, ID_EX_REG_ID_EX_REG_N144,
         ID_EX_REG_ID_EX_REG_N143, ID_EX_REG_ID_EX_REG_N142,
         ID_EX_REG_ID_EX_REG_N141, ID_EX_REG_ID_EX_REG_N140,
         ID_EX_REG_ID_EX_REG_N139, ID_EX_REG_ID_EX_REG_N138,
         ID_EX_REG_ID_EX_REG_N137, ID_EX_REG_ID_EX_REG_N136,
         ID_EX_REG_ID_EX_REG_N135, ID_EX_REG_ID_EX_REG_N134,
         ID_EX_REG_ID_EX_REG_N133, ID_EX_REG_ID_EX_REG_N132,
         ID_EX_REG_ID_EX_REG_N131, ID_EX_REG_ID_EX_REG_N130,
         ID_EX_REG_ID_EX_REG_N129, ID_EX_REG_ID_EX_REG_N128,
         ID_EX_REG_ID_EX_REG_N127, ID_EX_REG_ID_EX_REG_N124,
         ID_EX_REG_ID_EX_REG_N120, ID_EX_REG_ID_EX_REG_N119,
         ID_EX_REG_ID_EX_REG_N117, ID_EX_REG_ID_EX_REG_N116,
         ID_EX_REG_ID_EX_REG_N115, ID_EX_REG_ID_EX_REG_N113,
         ID_EX_REG_ID_EX_REG_N99, ID_EX_REG_ID_EX_REG_N98,
         ID_EX_REG_ID_EX_REG_N96, ID_EX_REG_ID_EX_REG_N95,
         ID_EX_REG_ID_EX_REG_N94, ID_EX_REG_ID_EX_REG_N93,
         ID_EX_REG_ID_EX_REG_N92, ID_EX_REG_ID_EX_REG_N91,
         ID_EX_REG_ID_EX_REG_N90, ID_EX_REG_ID_EX_REG_N89,
         ID_EX_REG_ID_EX_REG_N88, ID_EX_REG_ID_EX_REG_N87,
         ID_EX_REG_ID_EX_REG_N86, ID_EX_REG_ID_EX_REG_N85,
         ID_EX_REG_ID_EX_REG_N84, ID_EX_REG_ID_EX_REG_N83,
         ID_EX_REG_ID_EX_REG_N81, ID_EX_REG_ID_EX_REG_N80,
         ID_EX_REG_ID_EX_REG_N79, ID_EX_REG_ID_EX_REG_N76,
         ID_EX_REG_ID_EX_REG_N68, ID_EX_REG_ID_EX_REG_N67,
         ID_EX_REG_ID_EX_REG_N66, ID_EX_REG_ID_EX_REG_N65,
         ID_EX_REG_ID_EX_REG_N64, ID_EX_REG_ID_EX_REG_N63,
         ID_EX_REG_ID_EX_REG_N62, ID_EX_REG_ID_EX_REG_N61,
         ID_EX_REG_ID_EX_REG_N59, ID_EX_REG_ID_EX_REG_N57,
         ID_EX_REG_ID_EX_REG_N56, ID_EX_REG_ID_EX_REG_N55,
         ID_EX_REG_ID_EX_REG_N54, ID_EX_REG_ID_EX_REG_N53,
         ID_EX_REG_ID_EX_REG_N52, ID_EX_REG_ID_EX_REG_N51,
         ID_EX_REG_ID_EX_REG_N50, ID_EX_REG_ID_EX_REG_N49,
         ID_EX_REG_ID_EX_REG_N48, ID_EX_REG_ID_EX_REG_N47,
         ID_EX_REG_ID_EX_REG_N46, ID_EX_REG_ID_EX_REG_N45,
         ID_EX_REG_ID_EX_REG_N44, ID_EX_REG_ID_EX_REG_N43,
         ID_EX_REG_ID_EX_REG_N42, ID_EX_REG_ID_EX_REG_N41,
         ID_EX_REG_ID_EX_REG_N40, ID_EX_REG_ID_EX_REG_N39,
         ID_EX_REG_ID_EX_REG_N38, ID_EX_REG_ID_EX_REG_N37,
         ID_EX_REG_ID_EX_REG_N36, ID_EX_REG_ID_EX_REG_N35,
         ID_EX_REG_ID_EX_REG_N34, ID_EX_REG_ID_EX_REG_N33,
         ID_EX_REG_ID_EX_REG_N32, ID_EX_REG_ID_EX_REG_N31,
         ID_EX_REG_ID_EX_REG_N30, ID_EX_REG_ID_EX_REG_N29,
         ID_EX_REG_ID_EX_REG_N28, ID_EX_REG_ID_EX_REG_N27,
         ID_EX_REG_ID_EX_REG_N26, ID_EX_REG_ID_EX_REG_N25,
         ID_EX_REG_ID_EX_REG_N24, ID_EX_REG_ID_EX_REG_N23,
         ID_EX_REG_ID_EX_REG_N22, ID_EX_REG_ID_EX_REG_N21,
         ID_EX_REG_ID_EX_REG_N20, ID_EX_REG_ID_EX_REG_N19,
         ID_EX_REG_ID_EX_REG_N18, ID_EX_REG_ID_EX_REG_N17,
         ID_EX_REG_ID_EX_REG_N16, ID_EX_REG_ID_EX_REG_N15,
         ID_EX_REG_ID_EX_REG_N14, EXEC_STAGE_imm16_32_16_,
         EX_MEM_REGISTER_EX_MEM_REG_N118, EX_MEM_REGISTER_EX_MEM_REG_N117,
         EX_MEM_REGISTER_EX_MEM_REG_N116, EX_MEM_REGISTER_EX_MEM_REG_N115,
         EX_MEM_REGISTER_EX_MEM_REG_N114, EX_MEM_REGISTER_EX_MEM_REG_N109,
         EX_MEM_REGISTER_EX_MEM_REG_N108, EX_MEM_REGISTER_EX_MEM_REG_N107,
         EX_MEM_REGISTER_EX_MEM_REG_N106, EX_MEM_REGISTER_EX_MEM_REG_N105,
         EX_MEM_REGISTER_EX_MEM_REG_N104, EX_MEM_REGISTER_EX_MEM_REG_N103,
         EX_MEM_REGISTER_EX_MEM_REG_N102, EX_MEM_REGISTER_EX_MEM_REG_N101,
         EX_MEM_REGISTER_EX_MEM_REG_N100, EX_MEM_REGISTER_EX_MEM_REG_N99,
         EX_MEM_REGISTER_EX_MEM_REG_N98, EX_MEM_REGISTER_EX_MEM_REG_N97,
         EX_MEM_REGISTER_EX_MEM_REG_N96, EX_MEM_REGISTER_EX_MEM_REG_N95,
         EX_MEM_REGISTER_EX_MEM_REG_N94, EX_MEM_REGISTER_EX_MEM_REG_N93,
         EX_MEM_REGISTER_EX_MEM_REG_N92, EX_MEM_REGISTER_EX_MEM_REG_N91,
         EX_MEM_REGISTER_EX_MEM_REG_N90, EX_MEM_REGISTER_EX_MEM_REG_N89,
         EX_MEM_REGISTER_EX_MEM_REG_N88, EX_MEM_REGISTER_EX_MEM_REG_N87,
         EX_MEM_REGISTER_EX_MEM_REG_N86, EX_MEM_REGISTER_EX_MEM_REG_N85,
         EX_MEM_REGISTER_EX_MEM_REG_N84, EX_MEM_REGISTER_EX_MEM_REG_N83,
         EX_MEM_REGISTER_EX_MEM_REG_N81, EX_MEM_REGISTER_EX_MEM_REG_N79,
         EX_MEM_REGISTER_EX_MEM_REG_N78, EX_MEM_REGISTER_EX_MEM_REG_N77,
         EX_MEM_REGISTER_EX_MEM_REG_N76, EX_MEM_REGISTER_EX_MEM_REG_N75,
         EX_MEM_REGISTER_EX_MEM_REG_N74, EX_MEM_REGISTER_EX_MEM_REG_N72,
         EX_MEM_REGISTER_EX_MEM_REG_N71, EX_MEM_REGISTER_EX_MEM_REG_N70,
         EX_MEM_REGISTER_EX_MEM_REG_N69, EX_MEM_REGISTER_EX_MEM_REG_N68,
         EX_MEM_REGISTER_EX_MEM_REG_N67, EX_MEM_REGISTER_EX_MEM_REG_N66,
         EX_MEM_REGISTER_EX_MEM_REG_N65, EX_MEM_REGISTER_EX_MEM_REG_N64,
         EX_MEM_REGISTER_EX_MEM_REG_N63, EX_MEM_REGISTER_EX_MEM_REG_N62,
         EX_MEM_REGISTER_EX_MEM_REG_N61, EX_MEM_REGISTER_EX_MEM_REG_N60,
         EX_MEM_REGISTER_EX_MEM_REG_N59, EX_MEM_REGISTER_EX_MEM_REG_N58,
         EX_MEM_REGISTER_EX_MEM_REG_N57, EX_MEM_REGISTER_EX_MEM_REG_N56,
         EX_MEM_REGISTER_EX_MEM_REG_N55, EX_MEM_REGISTER_EX_MEM_REG_N54,
         EX_MEM_REGISTER_EX_MEM_REG_N53, EX_MEM_REGISTER_EX_MEM_REG_N52,
         EX_MEM_REGISTER_EX_MEM_REG_N51, EX_MEM_REGISTER_EX_MEM_REG_N50,
         EX_MEM_REGISTER_EX_MEM_REG_N49, EX_MEM_REGISTER_EX_MEM_REG_N48,
         EX_MEM_REGISTER_EX_MEM_REG_N47, EX_MEM_REGISTER_EX_MEM_REG_N46,
         EX_MEM_REGISTER_EX_MEM_REG_N45, EX_MEM_REGISTER_EX_MEM_REG_N44,
         EX_MEM_REGISTER_EX_MEM_REG_N43, EX_MEM_REGISTER_EX_MEM_REG_N42,
         EX_MEM_REGISTER_EX_MEM_REG_N41, EX_MEM_REGISTER_EX_MEM_REG_N40,
         EX_MEM_REGISTER_EX_MEM_REG_N39, EX_MEM_REGISTER_EX_MEM_REG_N38,
         EX_MEM_REGISTER_EX_MEM_REG_N37, EX_MEM_REGISTER_EX_MEM_REG_N36,
         EX_MEM_REGISTER_EX_MEM_REG_N35, EX_MEM_REGISTER_EX_MEM_REG_N34,
         EX_MEM_REGISTER_EX_MEM_REG_N33, EX_MEM_REGISTER_EX_MEM_REG_N32,
         EX_MEM_REGISTER_EX_MEM_REG_N31, EX_MEM_REGISTER_EX_MEM_REG_N30,
         EX_MEM_REGISTER_EX_MEM_REG_N29, EX_MEM_REGISTER_EX_MEM_REG_N28,
         EX_MEM_REGISTER_EX_MEM_REG_N27, EX_MEM_REGISTER_EX_MEM_REG_N26,
         EX_MEM_REGISTER_EX_MEM_REG_N25, EX_MEM_REGISTER_EX_MEM_REG_N24,
         EX_MEM_REGISTER_EX_MEM_REG_N23, EX_MEM_REGISTER_EX_MEM_REG_N22,
         EX_MEM_REGISTER_EX_MEM_REG_N21, EX_MEM_REGISTER_EX_MEM_REG_N20,
         EX_MEM_REGISTER_EX_MEM_REG_N19, EX_MEM_REGISTER_EX_MEM_REG_N18,
         EX_MEM_REGISTER_EX_MEM_REG_N17, EX_MEM_REGISTER_EX_MEM_REG_N16,
         EX_MEM_REGISTER_EX_MEM_REG_N15, EX_MEM_REGISTER_EX_MEM_REG_N14,
         EX_MEM_REGISTER_EX_MEM_REG_N13, EX_MEM_REGISTER_EX_MEM_REG_N12,
         EX_MEM_REGISTER_EX_MEM_REG_N11, EX_MEM_REGISTER_EX_MEM_REG_N10,
         EX_MEM_REGISTER_EX_MEM_REG_N9, MEM_WB_REG_MEM_WB_REG_N78,
         MEM_WB_REG_MEM_WB_REG_N77, MEM_WB_REG_MEM_WB_REG_N76,
         MEM_WB_REG_MEM_WB_REG_N75, MEM_WB_REG_MEM_WB_REG_N74,
         MEM_WB_REG_MEM_WB_REG_N9, MEM_WB_REG_MEM_WB_REG_N8,
         MEM_WB_REG_MEM_WB_REG_N7, MEM_WB_REG_MEM_WB_REG_N6,
         REG_FILE_reg_out_31__31_, REG_FILE_reg_out_31__30_,
         REG_FILE_reg_out_31__29_, REG_FILE_reg_out_31__28_,
         REG_FILE_reg_out_31__27_, REG_FILE_reg_out_31__26_,
         REG_FILE_reg_out_31__25_, REG_FILE_reg_out_31__24_,
         REG_FILE_reg_out_31__23_, REG_FILE_reg_out_31__22_,
         REG_FILE_reg_out_31__21_, REG_FILE_reg_out_31__20_,
         REG_FILE_reg_out_31__19_, REG_FILE_reg_out_31__18_,
         REG_FILE_reg_out_31__17_, REG_FILE_reg_out_31__16_,
         REG_FILE_reg_out_31__15_, REG_FILE_reg_out_31__14_,
         REG_FILE_reg_out_31__13_, REG_FILE_reg_out_31__12_,
         REG_FILE_reg_out_31__11_, REG_FILE_reg_out_31__10_,
         REG_FILE_reg_out_31__9_, REG_FILE_reg_out_31__8_,
         REG_FILE_reg_out_31__7_, REG_FILE_reg_out_31__6_,
         REG_FILE_reg_out_31__5_, REG_FILE_reg_out_31__4_,
         REG_FILE_reg_out_31__3_, REG_FILE_reg_out_31__2_,
         REG_FILE_reg_out_31__1_, REG_FILE_reg_out_31__0_,
         REG_FILE_reg_out_30__31_, REG_FILE_reg_out_30__30_,
         REG_FILE_reg_out_30__29_, REG_FILE_reg_out_30__28_,
         REG_FILE_reg_out_30__27_, REG_FILE_reg_out_30__26_,
         REG_FILE_reg_out_30__25_, REG_FILE_reg_out_30__24_,
         REG_FILE_reg_out_30__23_, REG_FILE_reg_out_30__22_,
         REG_FILE_reg_out_30__21_, REG_FILE_reg_out_30__20_,
         REG_FILE_reg_out_30__19_, REG_FILE_reg_out_30__18_,
         REG_FILE_reg_out_30__17_, REG_FILE_reg_out_30__16_,
         REG_FILE_reg_out_30__15_, REG_FILE_reg_out_30__14_,
         REG_FILE_reg_out_30__13_, REG_FILE_reg_out_30__12_,
         REG_FILE_reg_out_30__11_, REG_FILE_reg_out_30__10_,
         REG_FILE_reg_out_30__9_, REG_FILE_reg_out_30__8_,
         REG_FILE_reg_out_30__7_, REG_FILE_reg_out_30__6_,
         REG_FILE_reg_out_30__5_, REG_FILE_reg_out_30__4_,
         REG_FILE_reg_out_30__3_, REG_FILE_reg_out_30__2_,
         REG_FILE_reg_out_30__1_, REG_FILE_reg_out_30__0_,
         REG_FILE_reg_out_28__31_, REG_FILE_reg_out_28__30_,
         REG_FILE_reg_out_28__29_, REG_FILE_reg_out_28__28_,
         REG_FILE_reg_out_28__27_, REG_FILE_reg_out_28__26_,
         REG_FILE_reg_out_28__25_, REG_FILE_reg_out_28__24_,
         REG_FILE_reg_out_28__23_, REG_FILE_reg_out_28__22_,
         REG_FILE_reg_out_28__21_, REG_FILE_reg_out_28__20_,
         REG_FILE_reg_out_28__19_, REG_FILE_reg_out_28__18_,
         REG_FILE_reg_out_28__17_, REG_FILE_reg_out_28__16_,
         REG_FILE_reg_out_28__15_, REG_FILE_reg_out_28__14_,
         REG_FILE_reg_out_28__13_, REG_FILE_reg_out_28__12_,
         REG_FILE_reg_out_28__11_, REG_FILE_reg_out_28__10_,
         REG_FILE_reg_out_28__9_, REG_FILE_reg_out_28__8_,
         REG_FILE_reg_out_28__7_, REG_FILE_reg_out_28__6_,
         REG_FILE_reg_out_28__5_, REG_FILE_reg_out_28__4_,
         REG_FILE_reg_out_28__3_, REG_FILE_reg_out_28__2_,
         REG_FILE_reg_out_28__1_, REG_FILE_reg_out_28__0_,
         REG_FILE_reg_out_27__31_, REG_FILE_reg_out_27__30_,
         REG_FILE_reg_out_27__29_, REG_FILE_reg_out_27__28_,
         REG_FILE_reg_out_27__27_, REG_FILE_reg_out_27__26_,
         REG_FILE_reg_out_27__25_, REG_FILE_reg_out_27__24_,
         REG_FILE_reg_out_27__23_, REG_FILE_reg_out_27__22_,
         REG_FILE_reg_out_27__21_, REG_FILE_reg_out_27__20_,
         REG_FILE_reg_out_27__19_, REG_FILE_reg_out_27__18_,
         REG_FILE_reg_out_27__17_, REG_FILE_reg_out_27__16_,
         REG_FILE_reg_out_27__15_, REG_FILE_reg_out_27__14_,
         REG_FILE_reg_out_27__13_, REG_FILE_reg_out_27__12_,
         REG_FILE_reg_out_27__11_, REG_FILE_reg_out_27__10_,
         REG_FILE_reg_out_27__9_, REG_FILE_reg_out_27__8_,
         REG_FILE_reg_out_27__7_, REG_FILE_reg_out_27__6_,
         REG_FILE_reg_out_27__5_, REG_FILE_reg_out_27__4_,
         REG_FILE_reg_out_27__3_, REG_FILE_reg_out_27__2_,
         REG_FILE_reg_out_27__1_, REG_FILE_reg_out_27__0_,
         REG_FILE_reg_out_26__31_, REG_FILE_reg_out_26__30_,
         REG_FILE_reg_out_26__29_, REG_FILE_reg_out_26__28_,
         REG_FILE_reg_out_26__27_, REG_FILE_reg_out_26__26_,
         REG_FILE_reg_out_26__25_, REG_FILE_reg_out_26__24_,
         REG_FILE_reg_out_26__23_, REG_FILE_reg_out_26__22_,
         REG_FILE_reg_out_26__21_, REG_FILE_reg_out_26__20_,
         REG_FILE_reg_out_26__19_, REG_FILE_reg_out_26__18_,
         REG_FILE_reg_out_26__17_, REG_FILE_reg_out_26__16_,
         REG_FILE_reg_out_26__15_, REG_FILE_reg_out_26__14_,
         REG_FILE_reg_out_26__13_, REG_FILE_reg_out_26__12_,
         REG_FILE_reg_out_26__11_, REG_FILE_reg_out_26__10_,
         REG_FILE_reg_out_26__9_, REG_FILE_reg_out_26__8_,
         REG_FILE_reg_out_26__7_, REG_FILE_reg_out_26__6_,
         REG_FILE_reg_out_26__5_, REG_FILE_reg_out_26__4_,
         REG_FILE_reg_out_26__3_, REG_FILE_reg_out_26__2_,
         REG_FILE_reg_out_26__1_, REG_FILE_reg_out_26__0_,
         REG_FILE_reg_out_24__31_, REG_FILE_reg_out_24__30_,
         REG_FILE_reg_out_24__29_, REG_FILE_reg_out_24__28_,
         REG_FILE_reg_out_24__27_, REG_FILE_reg_out_24__26_,
         REG_FILE_reg_out_24__25_, REG_FILE_reg_out_24__24_,
         REG_FILE_reg_out_24__23_, REG_FILE_reg_out_24__22_,
         REG_FILE_reg_out_24__21_, REG_FILE_reg_out_24__20_,
         REG_FILE_reg_out_24__19_, REG_FILE_reg_out_24__18_,
         REG_FILE_reg_out_24__17_, REG_FILE_reg_out_24__16_,
         REG_FILE_reg_out_24__15_, REG_FILE_reg_out_24__14_,
         REG_FILE_reg_out_24__13_, REG_FILE_reg_out_24__12_,
         REG_FILE_reg_out_24__11_, REG_FILE_reg_out_24__10_,
         REG_FILE_reg_out_24__9_, REG_FILE_reg_out_24__8_,
         REG_FILE_reg_out_24__7_, REG_FILE_reg_out_24__6_,
         REG_FILE_reg_out_24__5_, REG_FILE_reg_out_24__4_,
         REG_FILE_reg_out_24__3_, REG_FILE_reg_out_24__2_,
         REG_FILE_reg_out_24__1_, REG_FILE_reg_out_24__0_,
         REG_FILE_reg_out_23__31_, REG_FILE_reg_out_23__30_,
         REG_FILE_reg_out_23__29_, REG_FILE_reg_out_23__28_,
         REG_FILE_reg_out_23__27_, REG_FILE_reg_out_23__26_,
         REG_FILE_reg_out_23__25_, REG_FILE_reg_out_23__24_,
         REG_FILE_reg_out_23__23_, REG_FILE_reg_out_23__22_,
         REG_FILE_reg_out_23__21_, REG_FILE_reg_out_23__20_,
         REG_FILE_reg_out_23__19_, REG_FILE_reg_out_23__18_,
         REG_FILE_reg_out_23__17_, REG_FILE_reg_out_23__16_,
         REG_FILE_reg_out_23__15_, REG_FILE_reg_out_23__14_,
         REG_FILE_reg_out_23__13_, REG_FILE_reg_out_23__12_,
         REG_FILE_reg_out_23__11_, REG_FILE_reg_out_23__10_,
         REG_FILE_reg_out_23__9_, REG_FILE_reg_out_23__8_,
         REG_FILE_reg_out_23__7_, REG_FILE_reg_out_23__6_,
         REG_FILE_reg_out_23__5_, REG_FILE_reg_out_23__4_,
         REG_FILE_reg_out_23__3_, REG_FILE_reg_out_23__2_,
         REG_FILE_reg_out_23__1_, REG_FILE_reg_out_23__0_,
         REG_FILE_reg_out_20__31_, REG_FILE_reg_out_20__30_,
         REG_FILE_reg_out_20__29_, REG_FILE_reg_out_20__28_,
         REG_FILE_reg_out_20__27_, REG_FILE_reg_out_20__26_,
         REG_FILE_reg_out_20__25_, REG_FILE_reg_out_20__24_,
         REG_FILE_reg_out_20__23_, REG_FILE_reg_out_20__22_,
         REG_FILE_reg_out_20__21_, REG_FILE_reg_out_20__20_,
         REG_FILE_reg_out_20__19_, REG_FILE_reg_out_20__18_,
         REG_FILE_reg_out_20__17_, REG_FILE_reg_out_20__16_,
         REG_FILE_reg_out_20__15_, REG_FILE_reg_out_20__14_,
         REG_FILE_reg_out_20__13_, REG_FILE_reg_out_20__12_,
         REG_FILE_reg_out_20__11_, REG_FILE_reg_out_20__10_,
         REG_FILE_reg_out_20__9_, REG_FILE_reg_out_20__8_,
         REG_FILE_reg_out_20__7_, REG_FILE_reg_out_20__6_,
         REG_FILE_reg_out_20__5_, REG_FILE_reg_out_20__4_,
         REG_FILE_reg_out_20__3_, REG_FILE_reg_out_20__2_,
         REG_FILE_reg_out_20__1_, REG_FILE_reg_out_20__0_,
         REG_FILE_reg_out_19__31_, REG_FILE_reg_out_19__30_,
         REG_FILE_reg_out_19__29_, REG_FILE_reg_out_19__28_,
         REG_FILE_reg_out_19__27_, REG_FILE_reg_out_19__26_,
         REG_FILE_reg_out_19__25_, REG_FILE_reg_out_19__24_,
         REG_FILE_reg_out_19__23_, REG_FILE_reg_out_19__22_,
         REG_FILE_reg_out_19__21_, REG_FILE_reg_out_19__20_,
         REG_FILE_reg_out_19__19_, REG_FILE_reg_out_19__18_,
         REG_FILE_reg_out_19__17_, REG_FILE_reg_out_19__16_,
         REG_FILE_reg_out_19__15_, REG_FILE_reg_out_19__14_,
         REG_FILE_reg_out_19__13_, REG_FILE_reg_out_19__12_,
         REG_FILE_reg_out_19__11_, REG_FILE_reg_out_19__10_,
         REG_FILE_reg_out_19__9_, REG_FILE_reg_out_19__8_,
         REG_FILE_reg_out_19__7_, REG_FILE_reg_out_19__6_,
         REG_FILE_reg_out_19__5_, REG_FILE_reg_out_19__4_,
         REG_FILE_reg_out_19__3_, REG_FILE_reg_out_19__2_,
         REG_FILE_reg_out_19__1_, REG_FILE_reg_out_19__0_,
         REG_FILE_reg_out_16__31_, REG_FILE_reg_out_16__30_,
         REG_FILE_reg_out_16__29_, REG_FILE_reg_out_16__28_,
         REG_FILE_reg_out_16__27_, REG_FILE_reg_out_16__26_,
         REG_FILE_reg_out_16__25_, REG_FILE_reg_out_16__24_,
         REG_FILE_reg_out_16__23_, REG_FILE_reg_out_16__22_,
         REG_FILE_reg_out_16__21_, REG_FILE_reg_out_16__20_,
         REG_FILE_reg_out_16__19_, REG_FILE_reg_out_16__18_,
         REG_FILE_reg_out_16__17_, REG_FILE_reg_out_16__16_,
         REG_FILE_reg_out_16__15_, REG_FILE_reg_out_16__14_,
         REG_FILE_reg_out_16__13_, REG_FILE_reg_out_16__12_,
         REG_FILE_reg_out_16__11_, REG_FILE_reg_out_16__10_,
         REG_FILE_reg_out_16__9_, REG_FILE_reg_out_16__8_,
         REG_FILE_reg_out_16__7_, REG_FILE_reg_out_16__6_,
         REG_FILE_reg_out_16__5_, REG_FILE_reg_out_16__4_,
         REG_FILE_reg_out_16__3_, REG_FILE_reg_out_16__2_,
         REG_FILE_reg_out_16__1_, REG_FILE_reg_out_16__0_,
         REG_FILE_reg_out_15__31_, REG_FILE_reg_out_15__30_,
         REG_FILE_reg_out_15__29_, REG_FILE_reg_out_15__28_,
         REG_FILE_reg_out_15__27_, REG_FILE_reg_out_15__26_,
         REG_FILE_reg_out_15__25_, REG_FILE_reg_out_15__24_,
         REG_FILE_reg_out_15__23_, REG_FILE_reg_out_15__22_,
         REG_FILE_reg_out_15__21_, REG_FILE_reg_out_15__20_,
         REG_FILE_reg_out_15__19_, REG_FILE_reg_out_15__18_,
         REG_FILE_reg_out_15__17_, REG_FILE_reg_out_15__16_,
         REG_FILE_reg_out_15__15_, REG_FILE_reg_out_15__14_,
         REG_FILE_reg_out_15__13_, REG_FILE_reg_out_15__12_,
         REG_FILE_reg_out_15__11_, REG_FILE_reg_out_15__10_,
         REG_FILE_reg_out_15__9_, REG_FILE_reg_out_15__8_,
         REG_FILE_reg_out_15__7_, REG_FILE_reg_out_15__6_,
         REG_FILE_reg_out_15__5_, REG_FILE_reg_out_15__4_,
         REG_FILE_reg_out_15__3_, REG_FILE_reg_out_15__2_,
         REG_FILE_reg_out_15__1_, REG_FILE_reg_out_15__0_,
         REG_FILE_reg_out_14__31_, REG_FILE_reg_out_14__30_,
         REG_FILE_reg_out_14__29_, REG_FILE_reg_out_14__28_,
         REG_FILE_reg_out_14__27_, REG_FILE_reg_out_14__26_,
         REG_FILE_reg_out_14__25_, REG_FILE_reg_out_14__24_,
         REG_FILE_reg_out_14__23_, REG_FILE_reg_out_14__22_,
         REG_FILE_reg_out_14__21_, REG_FILE_reg_out_14__20_,
         REG_FILE_reg_out_14__19_, REG_FILE_reg_out_14__18_,
         REG_FILE_reg_out_14__17_, REG_FILE_reg_out_14__16_,
         REG_FILE_reg_out_14__15_, REG_FILE_reg_out_14__14_,
         REG_FILE_reg_out_14__13_, REG_FILE_reg_out_14__12_,
         REG_FILE_reg_out_14__11_, REG_FILE_reg_out_14__10_,
         REG_FILE_reg_out_14__9_, REG_FILE_reg_out_14__8_,
         REG_FILE_reg_out_14__7_, REG_FILE_reg_out_14__6_,
         REG_FILE_reg_out_14__5_, REG_FILE_reg_out_14__4_,
         REG_FILE_reg_out_14__3_, REG_FILE_reg_out_14__2_,
         REG_FILE_reg_out_14__1_, REG_FILE_reg_out_14__0_,
         REG_FILE_reg_out_12__31_, REG_FILE_reg_out_12__30_,
         REG_FILE_reg_out_12__29_, REG_FILE_reg_out_12__28_,
         REG_FILE_reg_out_12__27_, REG_FILE_reg_out_12__26_,
         REG_FILE_reg_out_12__25_, REG_FILE_reg_out_12__24_,
         REG_FILE_reg_out_12__23_, REG_FILE_reg_out_12__22_,
         REG_FILE_reg_out_12__21_, REG_FILE_reg_out_12__20_,
         REG_FILE_reg_out_12__19_, REG_FILE_reg_out_12__18_,
         REG_FILE_reg_out_12__17_, REG_FILE_reg_out_12__16_,
         REG_FILE_reg_out_12__15_, REG_FILE_reg_out_12__14_,
         REG_FILE_reg_out_12__13_, REG_FILE_reg_out_12__12_,
         REG_FILE_reg_out_12__11_, REG_FILE_reg_out_12__10_,
         REG_FILE_reg_out_12__9_, REG_FILE_reg_out_12__8_,
         REG_FILE_reg_out_12__7_, REG_FILE_reg_out_12__6_,
         REG_FILE_reg_out_12__5_, REG_FILE_reg_out_12__4_,
         REG_FILE_reg_out_12__3_, REG_FILE_reg_out_12__2_,
         REG_FILE_reg_out_12__1_, REG_FILE_reg_out_12__0_,
         REG_FILE_reg_out_11__31_, REG_FILE_reg_out_11__30_,
         REG_FILE_reg_out_11__29_, REG_FILE_reg_out_11__28_,
         REG_FILE_reg_out_11__27_, REG_FILE_reg_out_11__26_,
         REG_FILE_reg_out_11__25_, REG_FILE_reg_out_11__24_,
         REG_FILE_reg_out_11__23_, REG_FILE_reg_out_11__22_,
         REG_FILE_reg_out_11__21_, REG_FILE_reg_out_11__20_,
         REG_FILE_reg_out_11__19_, REG_FILE_reg_out_11__18_,
         REG_FILE_reg_out_11__17_, REG_FILE_reg_out_11__16_,
         REG_FILE_reg_out_11__15_, REG_FILE_reg_out_11__14_,
         REG_FILE_reg_out_11__13_, REG_FILE_reg_out_11__12_,
         REG_FILE_reg_out_11__11_, REG_FILE_reg_out_11__10_,
         REG_FILE_reg_out_11__9_, REG_FILE_reg_out_11__8_,
         REG_FILE_reg_out_11__7_, REG_FILE_reg_out_11__6_,
         REG_FILE_reg_out_11__5_, REG_FILE_reg_out_11__4_,
         REG_FILE_reg_out_11__3_, REG_FILE_reg_out_11__2_,
         REG_FILE_reg_out_11__1_, REG_FILE_reg_out_11__0_,
         REG_FILE_reg_out_10__31_, REG_FILE_reg_out_10__30_,
         REG_FILE_reg_out_10__29_, REG_FILE_reg_out_10__28_,
         REG_FILE_reg_out_10__27_, REG_FILE_reg_out_10__26_,
         REG_FILE_reg_out_10__25_, REG_FILE_reg_out_10__24_,
         REG_FILE_reg_out_10__23_, REG_FILE_reg_out_10__22_,
         REG_FILE_reg_out_10__21_, REG_FILE_reg_out_10__20_,
         REG_FILE_reg_out_10__19_, REG_FILE_reg_out_10__18_,
         REG_FILE_reg_out_10__17_, REG_FILE_reg_out_10__16_,
         REG_FILE_reg_out_10__15_, REG_FILE_reg_out_10__14_,
         REG_FILE_reg_out_10__13_, REG_FILE_reg_out_10__12_,
         REG_FILE_reg_out_10__11_, REG_FILE_reg_out_10__10_,
         REG_FILE_reg_out_10__9_, REG_FILE_reg_out_10__8_,
         REG_FILE_reg_out_10__7_, REG_FILE_reg_out_10__6_,
         REG_FILE_reg_out_10__5_, REG_FILE_reg_out_10__4_,
         REG_FILE_reg_out_10__3_, REG_FILE_reg_out_10__2_,
         REG_FILE_reg_out_10__1_, REG_FILE_reg_out_10__0_,
         REG_FILE_reg_out_8__31_, REG_FILE_reg_out_8__30_,
         REG_FILE_reg_out_8__29_, REG_FILE_reg_out_8__28_,
         REG_FILE_reg_out_8__27_, REG_FILE_reg_out_8__26_,
         REG_FILE_reg_out_8__25_, REG_FILE_reg_out_8__24_,
         REG_FILE_reg_out_8__23_, REG_FILE_reg_out_8__22_,
         REG_FILE_reg_out_8__21_, REG_FILE_reg_out_8__20_,
         REG_FILE_reg_out_8__19_, REG_FILE_reg_out_8__18_,
         REG_FILE_reg_out_8__17_, REG_FILE_reg_out_8__16_,
         REG_FILE_reg_out_8__15_, REG_FILE_reg_out_8__14_,
         REG_FILE_reg_out_8__13_, REG_FILE_reg_out_8__12_,
         REG_FILE_reg_out_8__11_, REG_FILE_reg_out_8__10_,
         REG_FILE_reg_out_8__9_, REG_FILE_reg_out_8__8_,
         REG_FILE_reg_out_8__7_, REG_FILE_reg_out_8__6_,
         REG_FILE_reg_out_8__5_, REG_FILE_reg_out_8__4_,
         REG_FILE_reg_out_8__3_, REG_FILE_reg_out_8__2_,
         REG_FILE_reg_out_8__1_, REG_FILE_reg_out_8__0_,
         REG_FILE_reg_out_7__31_, REG_FILE_reg_out_7__30_,
         REG_FILE_reg_out_7__29_, REG_FILE_reg_out_7__28_,
         REG_FILE_reg_out_7__27_, REG_FILE_reg_out_7__26_,
         REG_FILE_reg_out_7__25_, REG_FILE_reg_out_7__24_,
         REG_FILE_reg_out_7__23_, REG_FILE_reg_out_7__22_,
         REG_FILE_reg_out_7__21_, REG_FILE_reg_out_7__20_,
         REG_FILE_reg_out_7__19_, REG_FILE_reg_out_7__18_,
         REG_FILE_reg_out_7__17_, REG_FILE_reg_out_7__16_,
         REG_FILE_reg_out_7__15_, REG_FILE_reg_out_7__14_,
         REG_FILE_reg_out_7__13_, REG_FILE_reg_out_7__12_,
         REG_FILE_reg_out_7__11_, REG_FILE_reg_out_7__10_,
         REG_FILE_reg_out_7__9_, REG_FILE_reg_out_7__8_,
         REG_FILE_reg_out_7__7_, REG_FILE_reg_out_7__6_,
         REG_FILE_reg_out_7__5_, REG_FILE_reg_out_7__4_,
         REG_FILE_reg_out_7__3_, REG_FILE_reg_out_7__2_,
         REG_FILE_reg_out_7__1_, REG_FILE_reg_out_7__0_,
         REG_FILE_reg_out_6__31_, REG_FILE_reg_out_6__30_,
         REG_FILE_reg_out_6__29_, REG_FILE_reg_out_6__28_,
         REG_FILE_reg_out_6__27_, REG_FILE_reg_out_6__26_,
         REG_FILE_reg_out_6__25_, REG_FILE_reg_out_6__24_,
         REG_FILE_reg_out_6__23_, REG_FILE_reg_out_6__22_,
         REG_FILE_reg_out_6__21_, REG_FILE_reg_out_6__20_,
         REG_FILE_reg_out_6__19_, REG_FILE_reg_out_6__18_,
         REG_FILE_reg_out_6__17_, REG_FILE_reg_out_6__16_,
         REG_FILE_reg_out_6__15_, REG_FILE_reg_out_6__14_,
         REG_FILE_reg_out_6__13_, REG_FILE_reg_out_6__12_,
         REG_FILE_reg_out_6__11_, REG_FILE_reg_out_6__10_,
         REG_FILE_reg_out_6__9_, REG_FILE_reg_out_6__8_,
         REG_FILE_reg_out_6__7_, REG_FILE_reg_out_6__6_,
         REG_FILE_reg_out_6__5_, REG_FILE_reg_out_6__4_,
         REG_FILE_reg_out_6__3_, REG_FILE_reg_out_6__2_,
         REG_FILE_reg_out_6__1_, REG_FILE_reg_out_6__0_,
         REG_FILE_reg_out_4__31_, REG_FILE_reg_out_4__30_,
         REG_FILE_reg_out_4__29_, REG_FILE_reg_out_4__28_,
         REG_FILE_reg_out_4__27_, REG_FILE_reg_out_4__26_,
         REG_FILE_reg_out_4__25_, REG_FILE_reg_out_4__24_,
         REG_FILE_reg_out_4__23_, REG_FILE_reg_out_4__22_,
         REG_FILE_reg_out_4__21_, REG_FILE_reg_out_4__20_,
         REG_FILE_reg_out_4__19_, REG_FILE_reg_out_4__18_,
         REG_FILE_reg_out_4__17_, REG_FILE_reg_out_4__16_,
         REG_FILE_reg_out_4__15_, REG_FILE_reg_out_4__14_,
         REG_FILE_reg_out_4__13_, REG_FILE_reg_out_4__12_,
         REG_FILE_reg_out_4__11_, REG_FILE_reg_out_4__10_,
         REG_FILE_reg_out_4__9_, REG_FILE_reg_out_4__8_,
         REG_FILE_reg_out_4__7_, REG_FILE_reg_out_4__6_,
         REG_FILE_reg_out_4__5_, REG_FILE_reg_out_4__4_,
         REG_FILE_reg_out_4__3_, REG_FILE_reg_out_4__2_,
         REG_FILE_reg_out_4__1_, REG_FILE_reg_out_4__0_,
         REG_FILE_reg_out_3__31_, REG_FILE_reg_out_3__30_,
         REG_FILE_reg_out_3__29_, REG_FILE_reg_out_3__28_,
         REG_FILE_reg_out_3__27_, REG_FILE_reg_out_3__26_,
         REG_FILE_reg_out_3__25_, REG_FILE_reg_out_3__24_,
         REG_FILE_reg_out_3__23_, REG_FILE_reg_out_3__22_,
         REG_FILE_reg_out_3__21_, REG_FILE_reg_out_3__20_,
         REG_FILE_reg_out_3__19_, REG_FILE_reg_out_3__18_,
         REG_FILE_reg_out_3__17_, REG_FILE_reg_out_3__16_,
         REG_FILE_reg_out_3__15_, REG_FILE_reg_out_3__14_,
         REG_FILE_reg_out_3__13_, REG_FILE_reg_out_3__12_,
         REG_FILE_reg_out_3__11_, REG_FILE_reg_out_3__10_,
         REG_FILE_reg_out_3__9_, REG_FILE_reg_out_3__8_,
         REG_FILE_reg_out_3__7_, REG_FILE_reg_out_3__6_,
         REG_FILE_reg_out_3__5_, REG_FILE_reg_out_3__4_,
         REG_FILE_reg_out_3__3_, REG_FILE_reg_out_3__2_,
         REG_FILE_reg_out_3__1_, REG_FILE_reg_out_3__0_,
         REG_FILE_reg_out_2__31_, REG_FILE_reg_out_2__30_,
         REG_FILE_reg_out_2__29_, REG_FILE_reg_out_2__28_,
         REG_FILE_reg_out_2__27_, REG_FILE_reg_out_2__26_,
         REG_FILE_reg_out_2__25_, REG_FILE_reg_out_2__24_,
         REG_FILE_reg_out_2__23_, REG_FILE_reg_out_2__22_,
         REG_FILE_reg_out_2__21_, REG_FILE_reg_out_2__20_,
         REG_FILE_reg_out_2__19_, REG_FILE_reg_out_2__18_,
         REG_FILE_reg_out_2__17_, REG_FILE_reg_out_2__16_,
         REG_FILE_reg_out_2__15_, REG_FILE_reg_out_2__14_,
         REG_FILE_reg_out_2__13_, REG_FILE_reg_out_2__12_,
         REG_FILE_reg_out_2__11_, REG_FILE_reg_out_2__10_,
         REG_FILE_reg_out_2__9_, REG_FILE_reg_out_2__8_,
         REG_FILE_reg_out_2__7_, REG_FILE_reg_out_2__6_,
         REG_FILE_reg_out_2__5_, REG_FILE_reg_out_2__4_,
         REG_FILE_reg_out_2__3_, REG_FILE_reg_out_2__2_,
         REG_FILE_reg_out_2__1_, REG_FILE_reg_out_2__0_,
         REG_FILE_reg_out_0__31_, REG_FILE_reg_out_0__30_,
         REG_FILE_reg_out_0__29_, REG_FILE_reg_out_0__28_,
         REG_FILE_reg_out_0__27_, REG_FILE_reg_out_0__26_,
         REG_FILE_reg_out_0__25_, REG_FILE_reg_out_0__24_,
         REG_FILE_reg_out_0__23_, REG_FILE_reg_out_0__22_,
         REG_FILE_reg_out_0__21_, REG_FILE_reg_out_0__20_,
         REG_FILE_reg_out_0__19_, REG_FILE_reg_out_0__18_,
         REG_FILE_reg_out_0__17_, REG_FILE_reg_out_0__16_,
         REG_FILE_reg_out_0__15_, REG_FILE_reg_out_0__14_,
         REG_FILE_reg_out_0__13_, REG_FILE_reg_out_0__12_,
         REG_FILE_reg_out_0__11_, REG_FILE_reg_out_0__10_,
         REG_FILE_reg_out_0__9_, REG_FILE_reg_out_0__8_,
         REG_FILE_reg_out_0__7_, REG_FILE_reg_out_0__6_,
         REG_FILE_reg_out_0__5_, REG_FILE_reg_out_0__4_,
         REG_FILE_reg_out_0__3_, REG_FILE_reg_out_0__2_,
         REG_FILE_reg_out_0__1_, REG_FILE_reg_out_0__0_,
         IF_STAGE_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         n1541, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1598, n1601, n1602, n1604, n1605, n1609, n1629, n1630,
         n1631, n1632, n1633, n1634, n1641, n1652, n1654, n1656, n1659, n1660,
         n1996, n2008, n2012, n3077, n3078, n3080, n3084, n3087, n3090, n3092,
         n3093, n3096, n3098, n3099, n3101, n3103, n3105, n3107, n3110, n3112,
         n3114, n3126, n3128, n3131, n3133, n3135, n3146, n3148, n3150, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3378, n3385,
         n3386, n3387, n3388, n3390, n3391, n3392, n3393, n3394, n3397, n3399,
         n3402, n3403, n3405, n3407, n3408, n3409, n3410, n3412, n3413, n3414,
         n3415, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3595, n3596, n3597, n3598, n3599, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3638, n3639, n3640, n3641, n3642, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3681, n3682, n3683, n3684, n3685, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3721, n3722, n3723, n3725, n3726, n3727, n3728, n3729, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3934, n3935, n3936, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4064, n4065, n4066, n4067, n4068, n4069,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4096, n4098, n4099, n4100, n4102, n4103, n4104, n4105,
         n4106, n4108, n4110, n4111, n4112, n4113, n4114, n4115, n4117, n4118,
         n4119, n4120, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4133, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4155, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4178, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4200, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4223, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4837, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n5398, n5399, n5400, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5665,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7346,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300;
  wire   [0:37] IF_ID_OUT;
  wire   [0:9] offset_26_id;
  wire   [32:202] ID_EXEC_OUT;
  wire   [0:31] nextPC_ex_out;
  wire   [0:4] destReg_ex_out;
  wire   [0:1] DSize_ex_out;
  wire   [101:106] EXEC_MEM_IN;
  wire   [37:106] MEM_WB_OUT;
  wire   [0:4] destReg_wb_out;
  wire   [16:31] ID_STAGE_imm16_aluA;
  wire   [6:15] EXEC_STAGE_imm26_32;
  wire   [16:31] WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf;

  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_32_ ( .D(IF_ID_REG_IF_ID_REG_N34), .CK(
        clk), .RN(n7787), .Q(IF_ID_OUT[32]), .QN(n6865) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_34_ ( .D(IF_ID_REG_IF_ID_REG_N32), .CK(
        clk), .RN(n7785), .Q(IF_ID_OUT[34]), .QN(n6347) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_59_ ( .D(IF_ID_REG_IF_ID_REG_N7), .CK(
        clk), .RN(n7776), .Q(ID_STAGE_imm16_aluA[27]), .QN(n6898) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_60_ ( .D(IF_ID_REG_IF_ID_REG_N6), .CK(
        clk), .RN(n7791), .Q(ID_STAGE_imm16_aluA[28]), .QN(n6862) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_62_ ( .D(IF_ID_REG_IF_ID_REG_N4), .CK(
        clk), .RN(n7777), .Q(ID_STAGE_imm16_aluA[30]), .QN(n6011) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_33_ ( .D(IF_ID_REG_IF_ID_REG_N33), .CK(
        clk), .RN(n7784), .Q(IF_ID_OUT[33]), .QN(n6343) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_35_ ( .D(IF_ID_REG_IF_ID_REG_N31), .CK(
        clk), .RN(n7778), .Q(IF_ID_OUT[35]), .QN(n6881) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_38_ ( .D(IF_ID_REG_IF_ID_REG_N28), .CK(
        clk), .RN(n7787), .Q(offset_26_id[0]), .QN(n6886) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_39_ ( .D(IF_ID_REG_IF_ID_REG_N27), .CK(
        clk), .RN(n7783), .Q(offset_26_id[1]), .QN(n6016) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_40_ ( .D(IF_ID_REG_IF_ID_REG_N26), .CK(
        clk), .RN(n7779), .Q(offset_26_id[2]), .QN(n5857) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_41_ ( .D(IF_ID_REG_IF_ID_REG_N25), .CK(
        clk), .RN(n7788), .Q(offset_26_id[3]), .QN(n6868) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_42_ ( .D(IF_ID_REG_IF_ID_REG_N24), .CK(
        clk), .RN(n7779), .Q(offset_26_id[4]), .QN(n6348) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_43_ ( .D(IF_ID_REG_IF_ID_REG_N23), .CK(
        clk), .RN(n7789), .Q(offset_26_id[5]), .QN(n6014) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_44_ ( .D(IF_ID_REG_IF_ID_REG_N22), .CK(
        clk), .RN(n7778), .Q(offset_26_id[6]), .QN(n6351) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_46_ ( .D(IF_ID_REG_IF_ID_REG_N20), .CK(
        clk), .RN(n7788), .Q(offset_26_id[8]), .QN(n5856) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_47_ ( .D(IF_ID_REG_IF_ID_REG_N19), .CK(
        clk), .RN(n7788), .Q(offset_26_id[9]), .QN(n5861) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_48_ ( .D(IF_ID_REG_IF_ID_REG_N18), .CK(
        clk), .RN(n7785), .Q(ID_STAGE_imm16_aluA[16]), .QN(n6891) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_49_ ( .D(IF_ID_REG_IF_ID_REG_N17), .CK(
        clk), .RN(n7790), .Q(ID_STAGE_imm16_aluA[17]), .QN(n6992) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_51_ ( .D(IF_ID_REG_IF_ID_REG_N15), .CK(
        clk), .RN(n7776), .Q(ID_STAGE_imm16_aluA[19]), .QN(n6022) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_52_ ( .D(IF_ID_REG_IF_ID_REG_N14), .CK(
        clk), .RN(n7784), .Q(ID_STAGE_imm16_aluA[20]), .QN(n6353) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_53_ ( .D(IF_ID_REG_IF_ID_REG_N13), .CK(
        clk), .RN(n7791), .QN(n6899) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_56_ ( .D(IF_ID_REG_IF_ID_REG_N10), .CK(
        clk), .RN(n7780), .Q(ID_STAGE_imm16_aluA[24]), .QN(n7216) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_77_ ( .D(DMEM_BUS_IN[8]), .CK(clk), 
        .RN(n7788), .QN(n6996) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_72_ ( .D(DMEM_BUS_IN[3]), .CK(clk), 
        .RN(n7788), .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[19]), .QN(n6991)
         );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_70_ ( .D(DMEM_BUS_IN[1]), .CK(clk), 
        .RN(n7788), .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[17]), .QN(n6997)
         );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_69_ ( .D(DMEM_BUS_IN[0]), .CK(clk), 
        .RN(n7788), .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[16]), .QN(n6352)
         );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__31_), .QN(n6276) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_95_ ( .D(n1586), .CK(clk), .RN(n7792), 
        .Q(ID_EXEC_OUT[95]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_82_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N100), .CK(clk), .RN(n7793), .Q(
        DMEM_BUS_OUT[13]), .QN(n6043) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_50_ ( .D(DMEM_BUS_OUT[13]), .CK(clk), 
        .RN(n7788), .Q(MEM_WB_OUT[50]), .QN(n6820) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_81_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N101), .CK(clk), .RN(n7788), .Q(
        DMEM_BUS_OUT[12]), .QN(n6024) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_49_ ( .D(DMEM_BUS_OUT[12]), .CK(clk), 
        .RN(n7788), .Q(MEM_WB_OUT[49]), .QN(n6821) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_80_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N102), .CK(clk), .RN(n7776), .Q(
        DMEM_BUS_OUT[11]), .QN(n6019) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_48_ ( .D(DMEM_BUS_OUT[11]), .CK(clk), 
        .RN(n7790), .Q(MEM_WB_OUT[48]), .QN(n6822) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_79_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N103), .CK(clk), .RN(n7791), .Q(
        DMEM_BUS_OUT[10]), .QN(n5923) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_47_ ( .D(DMEM_BUS_OUT[10]), .CK(clk), 
        .RN(n7780), .Q(MEM_WB_OUT[47]), .QN(n6823) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_78_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N104), .CK(clk), .RN(n7789), .Q(
        DMEM_BUS_OUT[9]), .QN(n5953) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_46_ ( .D(DMEM_BUS_OUT[9]), .CK(clk), 
        .RN(n7793), .Q(MEM_WB_OUT[46]), .QN(n6824) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_83_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N99), .CK(clk), .RN(n7777), .Q(
        DMEM_BUS_OUT[14]), .QN(n6017) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_51_ ( .D(DMEM_BUS_OUT[14]), .CK(clk), 
        .RN(n7793), .Q(MEM_WB_OUT[51]), .QN(n6819) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_100_ ( .D(n10293), .CK(clk), .RN(
        n7782), .Q(DMEM_BUS_OUT[31]), .QN(n6018) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_68_ ( .D(DMEM_BUS_OUT[31]), .CK(clk), 
        .RN(n7788), .Q(MEM_WB_OUT[68]), .QN(n6813) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_97_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N85), .CK(clk), .RN(n7792), .Q(
        DMEM_BUS_OUT[28]), .QN(n5919) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_65_ ( .D(DMEM_BUS_OUT[28]), .CK(clk), 
        .RN(n7792), .Q(MEM_WB_OUT[65]), .QN(n6321) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_76_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N106), .CK(clk), .RN(n7792), .Q(
        DMEM_BUS_OUT[7]), .QN(n5920) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_44_ ( .D(DMEM_BUS_OUT[7]), .CK(clk), 
        .RN(n7792), .Q(MEM_WB_OUT[44]), .QN(n6825) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_77_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N105), .CK(clk), .RN(n7792), .Q(
        DMEM_BUS_OUT[8]), .QN(n5922) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_45_ ( .D(DMEM_BUS_OUT[8]), .CK(clk), 
        .RN(n7792), .QN(n7033) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_75_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N107), .CK(clk), .RN(n7792), .Q(
        DMEM_BUS_OUT[6]), .QN(n5921) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_43_ ( .D(DMEM_BUS_OUT[6]), .CK(clk), 
        .RN(n7792), .Q(MEM_WB_OUT[43]), .QN(n6814) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_74_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N108), .CK(clk), .RN(n7792), .Q(
        DMEM_BUS_OUT[5]), .QN(n5914) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_42_ ( .D(DMEM_BUS_OUT[5]), .CK(clk), 
        .RN(n7792), .Q(MEM_WB_OUT[42]), .QN(n6815) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_89_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N93), .CK(clk), .RN(n7792), .Q(
        DMEM_BUS_OUT[20]), .QN(n6025) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_57_ ( .D(DMEM_BUS_OUT[20]), .CK(clk), 
        .RN(n7792), .Q(MEM_WB_OUT[57]), .QN(n6808) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_84_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N98), .CK(clk), .RN(n7792), .Q(
        DMEM_BUS_OUT[15]), .QN(n6042) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_52_ ( .D(DMEM_BUS_OUT[15]), .CK(clk), 
        .RN(n7793), .Q(MEM_WB_OUT[52]), .QN(n6818) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_91_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N91), .CK(clk), .RN(n7793), .Q(
        DMEM_BUS_OUT[22]), .QN(n5917) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_59_ ( .D(DMEM_BUS_OUT[22]), .CK(clk), 
        .RN(n7793), .Q(MEM_WB_OUT[59]), .QN(n6318) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_90_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N92), .CK(clk), .RN(n7793), .Q(
        DMEM_BUS_OUT[21]), .QN(n5918) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_58_ ( .D(DMEM_BUS_OUT[21]), .CK(clk), 
        .RN(n7793), .Q(MEM_WB_OUT[58]), .QN(n6319) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_86_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N96), .CK(clk), .RN(n7793), .Q(
        DMEM_BUS_OUT[17]), .QN(n6033) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_54_ ( .D(DMEM_BUS_OUT[17]), .CK(clk), 
        .RN(n7793), .Q(MEM_WB_OUT[54]), .QN(n6810) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_72_ ( .D(n10294), .CK(clk), .RN(
        n7793), .Q(DMEM_BUS_OUT[3]), .QN(n5952) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_40_ ( .D(DMEM_BUS_OUT[3]), .CK(clk), 
        .RN(n7793), .Q(MEM_WB_OUT[40]), .QN(n6826) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_71_ ( .D(n10295), .CK(clk), .RN(
        n7793), .Q(DMEM_BUS_OUT[2]), .QN(n5926) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_39_ ( .D(DMEM_BUS_OUT[2]), .CK(clk), 
        .RN(n7793), .Q(MEM_WB_OUT[39]), .QN(n6827) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_70_ ( .D(n10297), .CK(clk), .RN(
        n7793), .Q(DMEM_BUS_OUT[1]), .QN(n5948) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_38_ ( .D(DMEM_BUS_OUT[1]), .CK(clk), 
        .RN(n7793), .QN(n7034) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_73_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N109), .CK(clk), .RN(n7793), .Q(
        DMEM_BUS_OUT[4]), .QN(n5925) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_41_ ( .D(DMEM_BUS_OUT[4]), .CK(clk), 
        .RN(n7793), .Q(MEM_WB_OUT[41]), .QN(n6816) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_87_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N95), .CK(clk), .RN(n7789), .Q(
        DMEM_BUS_OUT[18]), .QN(n6032) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_55_ ( .D(DMEM_BUS_OUT[18]), .CK(clk), 
        .RN(n7785), .Q(MEM_WB_OUT[55]), .QN(n6809) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_69_ ( .D(n10298), .CK(clk), .RN(
        n7788), .Q(DMEM_BUS_OUT[0]), .QN(n5888) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_37_ ( .D(DMEM_BUS_OUT[0]), .CK(clk), 
        .RN(n7785), .Q(MEM_WB_OUT[37]), .QN(n6817) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_85_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N97), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[16]), .QN(n6030) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_53_ ( .D(DMEM_BUS_OUT[16]), .CK(clk), 
        .RN(n7783), .Q(MEM_WB_OUT[53]), .QN(n6811) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_99_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N83), .CK(clk), .RN(n7778), .Q(
        DMEM_BUS_OUT[30]), .QN(n5889) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_67_ ( .D(DMEM_BUS_OUT[30]), .CK(clk), 
        .RN(n7776), .Q(MEM_WB_OUT[67]), .QN(n6266) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_98_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N84), .CK(clk), .RN(n7786), .Q(
        DMEM_BUS_OUT[29]), .QN(n5885) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_66_ ( .D(DMEM_BUS_OUT[29]), .CK(clk), 
        .RN(n7787), .Q(MEM_WB_OUT[66]), .QN(n6320) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_93_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N89), .CK(clk), .RN(n7792), .Q(
        DMEM_BUS_OUT[24]), .QN(n5887) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_61_ ( .D(DMEM_BUS_OUT[24]), .CK(clk), 
        .RN(n7784), .Q(MEM_WB_OUT[61]), .QN(n6325) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_92_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N90), .CK(clk), .RN(n7781), .Q(
        DMEM_BUS_OUT[23]), .QN(n5886) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_60_ ( .D(DMEM_BUS_OUT[23]), .CK(clk), 
        .RN(n7777), .Q(MEM_WB_OUT[60]), .QN(n6330) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_147_ ( .D(ID_EX_REG_ID_EX_REG_N59), .CK(
        clk), .RN(n7776), .Q(ID_EXEC_OUT[147]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_143_ ( .D(ID_EX_REG_ID_EX_REG_N63), .CK(
        clk), .RN(n7794), .Q(EXEC_MEM_IN[101]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_149_ ( .D(ID_EX_REG_ID_EX_REG_N57), .CK(
        clk), .RN(n7794), .Q(EXEC_MEM_IN[103]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_150_ ( .D(ID_EX_REG_ID_EX_REG_N56), .CK(
        clk), .RN(n7794), .Q(EXEC_MEM_IN[104]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_151_ ( .D(ID_EX_REG_ID_EX_REG_N55), .CK(
        clk), .RN(n7787), .Q(EXEC_MEM_IN[105]), .QN(n5869) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_191_ ( .D(ID_EX_REG_ID_EX_REG_N15), .CK(
        clk), .RN(n7794), .QN(n7280) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_135_ ( .D(n1598), .CK(clk), .RN(n7794), 
        .QN(n7301) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_109_ ( .D(n1598), .CK(clk), .RN(n7794), 
        .QN(n6849) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_153_ ( .D(ID_EX_REG_ID_EX_REG_N53), .CK(
        clk), .RN(n7794), .Q(ID_EXEC_OUT[153]), .QN(n6481) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_148_ ( .D(n6010), .CK(clk), .RN(n7794), 
        .QN(n6461) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_98_ ( .D(n1609), .CK(clk), .RN(n7794), 
        .Q(EXEC_STAGE_imm26_32[8]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_124_ ( .D(n1609), .CK(clk), .RN(n7792), 
        .QN(n7294) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_102_ ( .D(n1605), .CK(clk), .RN(n7792), 
        .Q(EXEC_STAGE_imm26_32[12]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_128_ ( .D(n1605), .CK(clk), .RN(n7792), 
        .QN(n7291) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_103_ ( .D(n1604), .CK(clk), .RN(n7792), 
        .Q(EXEC_STAGE_imm26_32[13]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_129_ ( .D(n1604), .CK(clk), .RN(n7791), 
        .QN(n7299) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_105_ ( .D(n1602), .CK(clk), .RN(n7791), 
        .Q(EXEC_STAGE_imm26_32[15]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_131_ ( .D(n1602), .CK(clk), .RN(n7791), 
        .QN(n7296) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_106_ ( .D(n1601), .CK(clk), .RN(n7791), 
        .QN(n7304) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_132_ ( .D(n1601), .CK(clk), .RN(n7791), 
        .QN(n7295) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_101_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N81), .CK(clk), .RN(n7791), .Q(
        MEM_WB_REG_MEM_WB_REG_N9) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_103_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N79), .CK(clk), .RN(n7791), .Q(
        MEM_WB_REG_MEM_WB_REG_N8), .QN(n6908) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_102_ ( .D(MEM_WB_REG_MEM_WB_REG_N8), 
        .CK(clk), .RN(n7791), .Q(RegWrite_wb_out) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_104_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N78), .CK(clk), .RN(n7791), .Q(
        MEM_WB_REG_MEM_WB_REG_N7) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_116_ ( .D(ID_EX_REG_ID_EX_REG_N90), .CK(
        clk), .RN(n7791), .QN(n6851) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_197_ ( .D(ID_EX_REG_ID_EX_REG_N90), .CK(
        clk), .RN(n7791), .Q(ID_EXEC_OUT[197]), .QN(n7330) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_117_ ( .D(ID_EX_REG_ID_EX_REG_N89), .CK(
        clk), .RN(n7791), .QN(n6854) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_118_ ( .D(ID_EX_REG_ID_EX_REG_N88), .CK(
        clk), .RN(n7791), .QN(n6859) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_138_ ( .D(ID_EX_REG_ID_EX_REG_N68), .CK(
        clk), .RN(n7790), .Q(destReg_ex_out[0]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_139_ ( .D(ID_EX_REG_ID_EX_REG_N67), .CK(
        clk), .RN(n7790), .Q(destReg_ex_out[1]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_140_ ( .D(ID_EX_REG_ID_EX_REG_N66), .CK(
        clk), .RN(n7790), .Q(destReg_ex_out[2]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_141_ ( .D(ID_EX_REG_ID_EX_REG_N65), .CK(
        clk), .RN(n7790), .Q(destReg_ex_out[3]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_142_ ( .D(ID_EX_REG_ID_EX_REG_N64), .CK(
        clk), .RN(n7790), .Q(destReg_ex_out[4]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_36_ ( .D(MEM_WB_REG_MEM_WB_REG_N74), 
        .CK(clk), .RN(n7790), .Q(destReg_wb_out[4]), .QN(n7334) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_119_ ( .D(ID_EX_REG_ID_EX_REG_N87), .CK(
        clk), .RN(n7790), .QN(n6857) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_200_ ( .D(ID_EX_REG_ID_EX_REG_N87), .CK(
        clk), .RN(n7790), .Q(ID_EXEC_OUT[200]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_152_ ( .D(ID_EX_REG_ID_EX_REG_N54), .CK(
        clk), .RN(n7788), .Q(EXEC_MEM_IN[106]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_106_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N76), .CK(clk), .RN(n7777), .Q(
        MEM_WB_REG_MEM_WB_REG_N6) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_104_ ( .D(MEM_WB_REG_MEM_WB_REG_N6), 
        .CK(clk), .RN(n7785), .QN(n6913) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_154_ ( .D(ID_EX_REG_ID_EX_REG_N52), .CK(
        clk), .RN(n7793), .Q(DSize_ex_out[0]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_107_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N75), .CK(clk), .RN(n7781), .Q(
        DMEM_BUS_OUT[65]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_155_ ( .D(ID_EX_REG_ID_EX_REG_N51), .CK(
        clk), .RN(n7782), .Q(DSize_ex_out[1]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_108_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N74), .CK(clk), .RN(n7783), .Q(
        DMEM_BUS_OUT[66]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6448) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__12_), .QN(n6263) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__12_), .QN(n6560) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__12_), .QN(n6749) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6458) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__12_), .QN(n5988) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__12_), .QN(n6622) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__12_), .QN(n7177) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__12_), .QN(n6180) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__12_), .QN(n6790) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6079) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__12_), .QN(n5989) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__12_), .QN(n6789) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__12_), .QN(n5969) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6447) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__12_), .QN(n6262) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__12_), .QN(n6232) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5942) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6391) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__12_), .QN(n6601) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6126) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__12_), .QN(n6692) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6107) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6058) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__12_), .QN(n6240) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__12_), .QN(n6748) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__12_), .QN(n6181) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6080) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__12_), .QN(n5907) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__12_), .QN(n6788) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__12_), .QN(n5970) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__12_), .QN(n6241) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_76_ ( .D(ID_EX_REG_ID_EX_REG_N130), .CK(
        clk), .RN(n7791), .Q(ID_EXEC_OUT[76]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6405) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__4_), .QN(n6258) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__4_), .QN(n6526) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__4_), .QN(n6713) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6115) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__4_), .QN(n6197) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__4_), .QN(n6203) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__4_), .QN(n6272) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__4_), .QN(n6155) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__4_), .QN(n6297) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5929) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__4_), .QN(n5975) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__4_), .QN(n6289) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__4_), .QN(n5959) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6097) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__4_), .QN(n6253) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__4_), .QN(n6542) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6367) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6051) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__4_), .QN(n6193) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6464) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__4_), .QN(n6249) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6090) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6402) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__4_), .QN(n6635) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__4_), .QN(n6705) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__4_), .QN(n6487) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6047) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__4_), .QN(n6534) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__4_), .QN(n6281) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__4_), .QN(n6147) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__4_), .QN(n6627) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_68_ ( .D(ID_EX_REG_ID_EX_REG_N138), .CK(
        clk), .RN(n7786), .Q(ID_EXEC_OUT[68]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6974) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__10_), .QN(n6265) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__10_), .QN(n6559) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__10_), .QN(n6747) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6460) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__10_), .QN(n5992) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__10_), .QN(n6621) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__10_), .QN(n7176) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__10_), .QN(n6183) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__10_), .QN(n6787) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6082) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__10_), .QN(n5993) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__10_), .QN(n6786) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__10_), .QN(n5971) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6449) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__10_), .QN(n6264) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__10_), .QN(n6236) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5943) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6395) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__10_), .QN(n5991) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6127) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__10_), .QN(n6693) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6108) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6059) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__10_), .QN(n6242) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__10_), .QN(n6746) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__10_), .QN(n6184) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6396) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__10_), .QN(n5994) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__10_), .QN(n6785) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__10_), .QN(n5972) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__10_), .QN(n6243) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_74_ ( .D(ID_EX_REG_ID_EX_REG_N132), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[74]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6946) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__2_), .QN(n6001) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__2_), .QN(n6524) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__2_), .QN(n6711) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6113) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__2_), .QN(n5981) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__2_), .QN(n6201) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__2_), .QN(n6270) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__2_), .QN(n6153) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__2_), .QN(n6295) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5894) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__2_), .QN(n5904) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__2_), .QN(n6287) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__2_), .QN(n5957) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6095) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__2_), .QN(n5998) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__2_), .QN(n6540) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6365) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6049) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__2_), .QN(n5974) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6462) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__2_), .QN(n6247) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6088) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6400) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__2_), .QN(n6633) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__2_), .QN(n6703) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__2_), .QN(n6485) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6358) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__2_), .QN(n6532) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__2_), .QN(n6279) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__2_), .QN(n6145) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__2_), .QN(n6625) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_66_ ( .D(ID_EX_REG_ID_EX_REG_N140), .CK(
        clk), .RN(n7790), .Q(ID_EXEC_OUT[66]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6112) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__8_), .QN(n6698) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__8_), .QN(n6558) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__8_), .QN(n6745) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5883) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__8_), .QN(n5995) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__8_), .QN(n6620) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__8_), .QN(n6744) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__8_), .QN(n6518) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__8_), .QN(n6784) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6084) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__8_), .QN(n6607) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__8_), .QN(n7207) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__8_), .QN(n7011) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6978) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__8_), .QN(n7134) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__8_), .QN(n6606) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6398) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5878) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__8_), .QN(n6238) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6133) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__8_), .QN(n7133) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6977) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6111) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__8_), .QN(n6696) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__8_), .QN(n6743) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__8_), .QN(n6519) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5879) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__8_), .QN(n6239) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__8_), .QN(n7206) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__8_), .QN(n7012) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__8_), .QN(n6697) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_72_ ( .D(ID_EX_REG_ID_EX_REG_N134), .CK(
        clk), .RN(n7784), .Q(ID_EXEC_OUT[72]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6949) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__6_), .QN(n6260) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__6_), .QN(n6528) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__6_), .QN(n6715) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6117) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__6_), .QN(n6198) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__6_), .QN(n6205) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__6_), .QN(n6274) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__6_), .QN(n6157) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__6_), .QN(n6299) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5931) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__6_), .QN(n5977) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__6_), .QN(n6291) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__6_), .QN(n5961) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6099) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__6_), .QN(n6255) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__6_), .QN(n6544) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6369) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6053) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__6_), .QN(n6195) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6466) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__6_), .QN(n6251) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6092) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6404) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__6_), .QN(n6637) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__6_), .QN(n6707) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__6_), .QN(n6489) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6361) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__6_), .QN(n6536) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__6_), .QN(n6283) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__6_), .QN(n6149) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__6_), .QN(n6629) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_70_ ( .D(ID_EX_REG_ID_EX_REG_N136), .CK(
        clk), .RN(n7780), .Q(ID_EXEC_OUT[70]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6948) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__5_), .QN(n6259) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__5_), .QN(n6527) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__5_), .QN(n6714) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6116) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__5_), .QN(n5983) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__5_), .QN(n6204) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__5_), .QN(n6273) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__5_), .QN(n6156) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__5_), .QN(n6298) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5930) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__5_), .QN(n5976) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__5_), .QN(n6290) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__5_), .QN(n5960) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6098) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__5_), .QN(n6254) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__5_), .QN(n6543) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6368) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6052) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__5_), .QN(n6194) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6465) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__5_), .QN(n6250) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6091) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6403) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__5_), .QN(n6636) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__5_), .QN(n6706) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__5_), .QN(n6488) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6360) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__5_), .QN(n6535) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__5_), .QN(n6282) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__5_), .QN(n6148) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__5_), .QN(n6628) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_69_ ( .D(ID_EX_REG_ID_EX_REG_N137), .CK(
        clk), .RN(n7776), .Q(ID_EXEC_OUT[69]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6973) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__11_), .QN(n7129) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__11_), .QN(n7047) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__11_), .QN(n7175) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6459) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__11_), .QN(n5990) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__11_), .QN(n7098) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__11_), .QN(n7174) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__11_), .QN(n7031) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__11_), .QN(n7205) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6393) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__11_), .QN(n6234) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__11_), .QN(n7204) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__11_), .QN(n6173) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6972) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__11_), .QN(n7128) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__11_), .QN(n6602) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6081) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6392) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__11_), .QN(n6233) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6986) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__11_), .QN(n7127) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6971) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6922) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__11_), .QN(n7089) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__11_), .QN(n6742) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__11_), .QN(n6182) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6394) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__11_), .QN(n6235) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__11_), .QN(n7203) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__11_), .QN(n7009) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__11_), .QN(n7090) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_75_ ( .D(ID_EX_REG_ID_EX_REG_N131), .CK(
        clk), .RN(n7779), .Q(ID_EXEC_OUT[75]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6947) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__3_), .QN(n6002) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__3_), .QN(n6525) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__3_), .QN(n6712) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6114) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__3_), .QN(n5982) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__3_), .QN(n6202) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__3_), .QN(n6271) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__3_), .QN(n6154) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__3_), .QN(n6296) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5928) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__3_), .QN(n5905) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__3_), .QN(n6288) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__3_), .QN(n5958) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6096) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__3_), .QN(n5999) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__3_), .QN(n6541) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6366) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6050) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__3_), .QN(n5901) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6463) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__3_), .QN(n6248) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6089) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6401) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__3_), .QN(n6634) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__3_), .QN(n6704) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__3_), .QN(n6486) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6359) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__3_), .QN(n6533) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__3_), .QN(n6280) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__3_), .QN(n6146) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__3_), .QN(n6626) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_67_ ( .D(ID_EX_REG_ID_EX_REG_N139), .CK(
        clk), .RN(n7777), .Q(ID_EXEC_OUT[67]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6110) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__9_), .QN(n7132) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__9_), .QN(n7046) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__9_), .QN(n7173) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6980) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__9_), .QN(n7074) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__9_), .QN(n7097) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__9_), .QN(n7172) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__9_), .QN(n7032) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__9_), .QN(n7202) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6083) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__9_), .QN(n6604) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__9_), .QN(n7201) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__9_), .QN(n6502) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6976) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__9_), .QN(n7131) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__9_), .QN(n6603) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6397) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5876) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__9_), .QN(n6237) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6132) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__9_), .QN(n7130) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6975) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6109) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__9_), .QN(n6694) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__9_), .QN(n6741) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__9_), .QN(n6517) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5877) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__9_), .QN(n6605) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__9_), .QN(n7200) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__9_), .QN(n7010) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__9_), .QN(n6695) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_73_ ( .D(ID_EX_REG_ID_EX_REG_N133), .CK(
        clk), .RN(n7781), .Q(ID_EXEC_OUT[73]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6102) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__1_), .QN(n6000) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__1_), .QN(n6523) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__1_), .QN(n6710) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5880) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__1_), .QN(n5980) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__1_), .QN(n6200) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__1_), .QN(n6269) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__1_), .QN(n6152) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__1_), .QN(n6294) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5927) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__1_), .QN(n5903) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__1_), .QN(n6286) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__1_), .QN(n5956) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6094) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__1_), .QN(n5997) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__1_), .QN(n6539) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6364) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6048) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__1_), .QN(n5900) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6128) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__1_), .QN(n6246) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6087) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6399) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__1_), .QN(n6632) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__1_), .QN(n6702) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__1_), .QN(n6484) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5891) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__1_), .QN(n6531) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__1_), .QN(n6278) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__1_), .QN(n6144) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__1_), .QN(n6624) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_65_ ( .D(ID_EX_REG_ID_EX_REG_N141), .CK(
        clk), .RN(n7781), .Q(ID_EXEC_OUT[65]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6101) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__0_), .QN(n6257) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__0_), .QN(n6522) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__0_), .QN(n6709) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5897) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__0_), .QN(n5979) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__0_), .QN(n6199) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__0_), .QN(n6268) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__0_), .QN(n6151) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__0_), .QN(n6293) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5893) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__0_), .QN(n5902) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__0_), .QN(n6285) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__0_), .QN(n5955) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5945) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__0_), .QN(n5996) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__0_), .QN(n6538) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6363) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5892) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__0_), .QN(n5973) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5954) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__0_), .QN(n6245) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6086) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5944) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__0_), .QN(n6631) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__0_), .QN(n6701) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__0_), .QN(n6483) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5890) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__0_), .QN(n6530) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__0_), .QN(n6277) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__0_), .QN(n6143) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__0_), .QN(n6623) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_64_ ( .D(ID_EX_REG_ID_EX_REG_N142), .CK(
        clk), .RN(n7781), .Q(ID_EXEC_OUT[64]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6950) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__7_), .QN(n6261) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__7_), .QN(n6529) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__7_), .QN(n6716) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5881) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__7_), .QN(n5984) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__7_), .QN(n6206) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__7_), .QN(n6275) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__7_), .QN(n6158) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__7_), .QN(n6300) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5932) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__7_), .QN(n5978) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__7_), .QN(n6292) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__7_), .QN(n5962) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6100) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__7_), .QN(n6256) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__7_), .QN(n6545) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6370) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5870) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__7_), .QN(n6196) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6129) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__7_), .QN(n6252) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6093) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6085) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__7_), .QN(n6638) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__7_), .QN(n6708) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__7_), .QN(n6490) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6362) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__7_), .QN(n6537) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__7_), .QN(n6284) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__7_), .QN(n6150) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__7_), .QN(n6630) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_71_ ( .D(ID_EX_REG_ID_EX_REG_N135), .CK(
        clk), .RN(n7781), .Q(ID_EXEC_OUT[71]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6407) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__31_), .QN(n6642) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__31_), .QN(n6557) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__31_), .QN(n6740) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6118) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__31_), .QN(n5985) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__31_), .QN(n6619) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__31_), .QN(n6503) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__31_), .QN(n6783) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6372) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__31_), .QN(n6207) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__31_), .QN(n7199) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__31_), .QN(n7002) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6952) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__31_), .QN(n6641) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__31_), .QN(n6561) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6371) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6060) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__31_), .QN(n5906) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6468) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__31_), .QN(n7099) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6951) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6406) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__31_), .QN(n6639) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__31_), .QN(n6739) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__31_), .QN(n6504) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6061) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__31_), .QN(n6208) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__31_), .QN(n7198) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__31_), .QN(n7003) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__31_), .QN(n6640) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6955) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__30_), .QN(n7102) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__30_), .QN(n7045) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__30_), .QN(n7171) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5898) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__30_), .QN(n7048) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__30_), .QN(n7096) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__30_), .QN(n7170) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__30_), .QN(n7013) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__30_), .QN(n7197) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6374) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__30_), .QN(n6563) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__30_), .QN(n7196) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__30_), .QN(n6491) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6954) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__30_), .QN(n7101) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__30_), .QN(n6562) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6373) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6062) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__30_), .QN(n6209) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6130) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__30_), .QN(n7100) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6953) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6408) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__30_), .QN(n6643) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__30_), .QN(n6738) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__30_), .QN(n6505) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6375) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__30_), .QN(n6564) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__30_), .QN(n7195) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__30_), .QN(n7004) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__30_), .QN(n6644) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_190_ ( .D(ID_EX_REG_ID_EX_REG_N16), .CK(
        clk), .RN(n7781), .QN(n6834) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6958) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__29_), .QN(n7105) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__29_), .QN(n7044) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__29_), .QN(n7169) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5899) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__29_), .QN(n6567) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__29_), .QN(n7095) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__29_), .QN(n7168) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__29_), .QN(n7014) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__29_), .QN(n7194) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6378) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__29_), .QN(n6568) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__29_), .QN(n7193) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__29_), .QN(n6492) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6957) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__29_), .QN(n7104) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__29_), .QN(n6565) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6377) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6376) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__29_), .QN(n6566) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6123) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__29_), .QN(n7103) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6956) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6919) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__29_), .QN(n7075) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__29_), .QN(n6737) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__29_), .QN(n6506) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5871) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__29_), .QN(n6569) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__29_), .QN(n7192) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__29_), .QN(n7005) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__29_), .QN(n7076) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_93_ ( .D(ID_EX_REG_ID_EX_REG_N113), .CK(
        clk), .RN(n7781), .Q(ID_EXEC_OUT[93]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6961) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__28_), .QN(n7108) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__28_), .QN(n7043) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__28_), .QN(n7167) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5882) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__28_), .QN(n6572) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__28_), .QN(n7094) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__28_), .QN(n7166) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__28_), .QN(n7015) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__28_), .QN(n7191) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5934) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__28_), .QN(n6573) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__28_), .QN(n7190) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__28_), .QN(n6493) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6960) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__28_), .QN(n7107) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__28_), .QN(n6570) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6379) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5872) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__28_), .QN(n6571) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6124) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__28_), .QN(n7106) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6959) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6920) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__28_), .QN(n7077) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__28_), .QN(n6736) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__28_), .QN(n6507) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5873) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__28_), .QN(n6574) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__28_), .QN(n7189) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__28_), .QN(n7006) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__28_), .QN(n7078) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_188_ ( .D(ID_EX_REG_ID_EX_REG_N18), .CK(
        clk), .RN(n7781), .QN(n6836) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6415) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__24_), .QN(n7117) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__24_), .QN(n7042) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__24_), .QN(n7165) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6119) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__24_), .QN(n7053) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__24_), .QN(n7093) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__24_), .QN(n7164) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__24_), .QN(n7021) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__24_), .QN(n7188) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6066) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__24_), .QN(n6584) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__24_), .QN(n7187) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__24_), .QN(n6496) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6414) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__24_), .QN(n7116) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__24_), .QN(n6583) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6382) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6065) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__24_), .QN(n6213) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6469) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__24_), .QN(n7115) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6964) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6413) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__24_), .QN(n6650) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__24_), .QN(n6735) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__24_), .QN(n6509) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6067) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__24_), .QN(n6585) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__24_), .QN(n7186) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__24_), .QN(n7007) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__24_), .QN(n6651) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_184_ ( .D(ID_EX_REG_ID_EX_REG_N22), .CK(
        clk), .RN(n7781), .QN(n6840) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6970) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__15_), .QN(n7126) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__15_), .QN(n7041) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__15_), .QN(n7163) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6456) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__15_), .QN(n6596) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__15_), .QN(n7092) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__15_), .QN(n7162) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__15_), .QN(n7030) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__15_), .QN(n7185) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6388) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__15_), .QN(n6597) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__15_), .QN(n7184) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__15_), .QN(n6172) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6969) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__15_), .QN(n7125) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__15_), .QN(n6594) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6073) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6387) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__15_), .QN(n6595) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6984) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__15_), .QN(n7124) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6968) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6921) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__15_), .QN(n7085) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__15_), .QN(n6734) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__15_), .QN(n6175) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6389) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__15_), .QN(n6598) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__15_), .QN(n7183) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__15_), .QN(n7008) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__15_), .QN(n7086) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_79_ ( .D(ID_EX_REG_ID_EX_REG_N127), .CK(
        clk), .RN(n7781), .Q(ID_EXEC_OUT[79]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6443) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__14_), .QN(n6686) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__14_), .QN(n7040) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__14_), .QN(n7161) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6457) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__14_), .QN(n6600) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__14_), .QN(n6618) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__14_), .QN(n7160) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__14_), .QN(n6176) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__14_), .QN(n6782) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6074) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__14_), .QN(n6226) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__14_), .QN(n6781) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__14_), .QN(n5965) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6442) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__14_), .QN(n6685) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__14_), .QN(n6225) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5940) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6390) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__14_), .QN(n6599) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6985) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__14_), .QN(n6684) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6105) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6057) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__14_), .QN(n7087) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__14_), .QN(n6733) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__14_), .QN(n6177) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6075) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__14_), .QN(n6227) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__14_), .QN(n6780) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__14_), .QN(n5966) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__14_), .QN(n7088) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_78_ ( .D(ID_EX_REG_ID_EX_REG_N128), .CK(
        clk), .RN(n7781), .Q(ID_EXEC_OUT[78]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6446) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__13_), .QN(n6691) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__13_), .QN(n7039) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__13_), .QN(n7159) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6979) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__13_), .QN(n7073) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__13_), .QN(n6617) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__13_), .QN(n7158) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__13_), .QN(n6178) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__13_), .QN(n6779) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6077) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__13_), .QN(n6230) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__13_), .QN(n6778) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__13_), .QN(n5967) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6445) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__13_), .QN(n6690) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__13_), .QN(n6228) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5941) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6076) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__13_), .QN(n6229) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6475) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__13_), .QN(n6687) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6106) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6444) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__13_), .QN(n6688) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__13_), .QN(n6732) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__13_), .QN(n6179) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6078) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__13_), .QN(n6231) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__13_), .QN(n6777) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__13_), .QN(n5968) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__13_), .QN(n6689) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_77_ ( .D(ID_EX_REG_ID_EX_REG_N129), .CK(
        clk), .RN(n7781), .Q(ID_EXEC_OUT[77]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6965) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__23_), .QN(n6656) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__23_), .QN(n6556) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__23_), .QN(n6731) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6453) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__23_), .QN(n6214) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__23_), .QN(n6616) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__23_), .QN(n7157) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__23_), .QN(n6510) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__23_), .QN(n6776) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6068) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__23_), .QN(n6215) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__23_), .QN(n6775) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__23_), .QN(n6162) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6417) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__23_), .QN(n6655) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__23_), .QN(n7054) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6927) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6383) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__23_), .QN(n7055) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6982) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__23_), .QN(n6652) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6416) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6055) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__23_), .QN(n6653) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__23_), .QN(n7156) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__23_), .QN(n7022) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6384) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__23_), .QN(n7056) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__23_), .QN(n6774) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__23_), .QN(n6497) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__23_), .QN(n6654) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_87_ ( .D(ID_EX_REG_ID_EX_REG_N119), .CK(
        clk), .RN(n7781), .Q(ID_EXEC_OUT[87]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6421) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__22_), .QN(n6661) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__22_), .QN(n6555) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__22_), .QN(n6730) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6120) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__22_), .QN(n6216) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__22_), .QN(n6615) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__22_), .QN(n7155) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__22_), .QN(n6511) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__22_), .QN(n6773) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6069) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__22_), .QN(n6217) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__22_), .QN(n6772) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__22_), .QN(n6163) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6420) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__22_), .QN(n6660) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__22_), .QN(n7057) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6929) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6928) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__22_), .QN(n7058) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6470) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__22_), .QN(n6657) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6419) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6418) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__22_), .QN(n6658) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__22_), .QN(n7154) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__22_), .QN(n7023) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6930) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__22_), .QN(n7059) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__22_), .QN(n6771) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__22_), .QN(n6498) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__22_), .QN(n6659) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_86_ ( .D(ID_EX_REG_ID_EX_REG_N120), .CK(
        clk), .RN(n7781), .Q(ID_EXEC_OUT[86]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6425) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__21_), .QN(n6666) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__21_), .QN(n6554) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__21_), .QN(n6729) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6121) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__21_), .QN(n6218) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__21_), .QN(n6614) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__21_), .QN(n7153) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__21_), .QN(n6512) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__21_), .QN(n6770) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6070) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__21_), .QN(n6219) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__21_), .QN(n6769) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__21_), .QN(n6164) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6424) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__21_), .QN(n6665) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__21_), .QN(n7060) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6932) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6931) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__21_), .QN(n7061) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6471) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__21_), .QN(n6662) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6423) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6422) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__21_), .QN(n6663) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__21_), .QN(n7152) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__21_), .QN(n7024) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6933) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__21_), .QN(n7062) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__21_), .QN(n6768) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__21_), .QN(n6499) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__21_), .QN(n6664) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_181_ ( .D(ID_EX_REG_ID_EX_REG_N25), .CK(
        clk), .RN(n7781), .QN(n6843) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6429) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__20_), .QN(n6671) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__20_), .QN(n6553) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__20_), .QN(n6728) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5950) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__20_), .QN(n6220) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__20_), .QN(n6613) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__20_), .QN(n7151) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__20_), .QN(n6513) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__20_), .QN(n6767) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5936) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__20_), .QN(n6221) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__20_), .QN(n6766) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__20_), .QN(n6165) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6428) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__20_), .QN(n6670) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__20_), .QN(n7063) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6935) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6934) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__20_), .QN(n7064) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6472) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__20_), .QN(n6667) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6427) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6426) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__20_), .QN(n6668) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__20_), .QN(n7150) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__20_), .QN(n7025) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6936) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__20_), .QN(n7065) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__20_), .QN(n6765) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__20_), .QN(n6500) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__20_), .QN(n6669) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_180_ ( .D(ID_EX_REG_ID_EX_REG_N26), .CK(
        clk), .RN(n7780), .QN(n7270) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6435) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__18_), .QN(n6677) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__18_), .QN(n6552) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__18_), .QN(n6727) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5951) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__18_), .QN(n6223) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__18_), .QN(n6612) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__18_), .QN(n7149) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__18_), .QN(n6515) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__18_), .QN(n6764) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5939) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__18_), .QN(n6224) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__18_), .QN(n6763) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__18_), .QN(n6168) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6434) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__18_), .QN(n6676) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__18_), .QN(n7066) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6938) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6937) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__18_), .QN(n7067) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6473) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__18_), .QN(n6673) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6433) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6432) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__18_), .QN(n6674) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__18_), .QN(n7148) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__18_), .QN(n7027) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6939) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__18_), .QN(n7068) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__18_), .QN(n6762) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__18_), .QN(n6501) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__18_), .QN(n6675) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_82_ ( .D(ID_EX_REG_ID_EX_REG_N124), .CK(
        clk), .RN(n7780), .Q(ID_EXEC_OUT[82]) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6439) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__17_), .QN(n6680) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__17_), .QN(n6551) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__17_), .QN(n6726) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6122) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__17_), .QN(n6591) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__17_), .QN(n6611) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__17_), .QN(n7147) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__17_), .QN(n6516) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__17_), .QN(n6761) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6071) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__17_), .QN(n5986) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__17_), .QN(n6760) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__17_), .QN(n6169) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6438) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__17_), .QN(n6679) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__17_), .QN(n7069) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6941) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6940) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__17_), .QN(n6590) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6474) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__17_), .QN(n6678) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6437) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6436) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__17_), .QN(n7122) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__17_), .QN(n7146) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__17_), .QN(n7028) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6942) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__17_), .QN(n7070) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__17_), .QN(n6759) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__17_), .QN(n6170) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__17_), .QN(n7123) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_177_ ( .D(ID_EX_REG_ID_EX_REG_N29), .CK(
        clk), .RN(n7780), .QN(n7273) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6441) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__16_), .QN(n6683) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__16_), .QN(n6550) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__16_), .QN(n6725) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6455) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__16_), .QN(n6593) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__16_), .QN(n6610) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__16_), .QN(n7145) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__16_), .QN(n6174) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__16_), .QN(n6758) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6072) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__16_), .QN(n5987) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__16_), .QN(n6757) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__16_), .QN(n5964) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6440) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__16_), .QN(n6682) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__16_), .QN(n7071) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6944) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6943) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__16_), .QN(n6592) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6983) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__16_), .QN(n6681) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6104) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6056) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__16_), .QN(n7083) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__16_), .QN(n7144) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__16_), .QN(n7029) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6945) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__16_), .QN(n7072) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__16_), .QN(n6756) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__16_), .QN(n6171) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__16_), .QN(n7084) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_176_ ( .D(ID_EX_REG_ID_EX_REG_N30), .CK(
        clk), .RN(n7780), .QN(n7274) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_156_ ( .D(ID_EX_REG_ID_EX_REG_N50), .CK(
        clk), .RN(n7780), .Q(ID_EXEC_OUT[156]), .QN(n6863) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_120_ ( .D(ID_EX_REG_ID_EX_REG_N86), .CK(
        clk), .RN(n7780), .QN(n6856) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_201_ ( .D(ID_EX_REG_ID_EX_REG_N86), .CK(
        clk), .RN(n7780), .Q(ID_EXEC_OUT[201]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_160_ ( .D(ID_EX_REG_ID_EX_REG_N46), .CK(
        clk), .RN(n7780), .Q(ID_EXEC_OUT[160]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_161_ ( .D(ID_EX_REG_ID_EX_REG_N45), .CK(
        clk), .RN(n7780), .Q(ID_EXEC_OUT[161]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_162_ ( .D(ID_EX_REG_ID_EX_REG_N44), .CK(
        clk), .RN(n7780), .Q(ID_EXEC_OUT[162]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_163_ ( .D(ID_EX_REG_ID_EX_REG_N43), .CK(
        clk), .RN(n7780), .Q(ID_EXEC_OUT[163]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_164_ ( .D(ID_EX_REG_ID_EX_REG_N42), .CK(
        clk), .RN(n7780), .Q(ID_EXEC_OUT[164]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_165_ ( .D(ID_EX_REG_ID_EX_REG_N41), .CK(
        clk), .RN(n7780), .Q(ID_EXEC_OUT[165]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_166_ ( .D(ID_EX_REG_ID_EX_REG_N40), .CK(
        clk), .RN(n7780), .Q(ID_EXEC_OUT[166]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_121_ ( .D(ID_EX_REG_ID_EX_REG_N85), .CK(
        clk), .RN(n7779), .QN(n6858) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_202_ ( .D(ID_EX_REG_ID_EX_REG_N85), .CK(
        clk), .RN(n7779), .Q(ID_EXEC_OUT[202]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_167_ ( .D(ID_EX_REG_ID_EX_REG_N39), .CK(
        clk), .RN(n7779), .Q(ID_EXEC_OUT[167]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_168_ ( .D(ID_EX_REG_ID_EX_REG_N38), .CK(
        clk), .RN(n7779), .Q(ID_EXEC_OUT[168]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_169_ ( .D(ID_EX_REG_ID_EX_REG_N37), .CK(
        clk), .RN(n7779), .Q(ID_EXEC_OUT[169]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_170_ ( .D(ID_EX_REG_ID_EX_REG_N36), .CK(
        clk), .RN(n7779), .Q(ID_EXEC_OUT[170]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_171_ ( .D(ID_EX_REG_ID_EX_REG_N35), .CK(
        clk), .RN(n7779), .QN(n7279) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_172_ ( .D(ID_EX_REG_ID_EX_REG_N34), .CK(
        clk), .RN(n7779), .QN(n7278) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_173_ ( .D(ID_EX_REG_ID_EX_REG_N33), .CK(
        clk), .RN(n7779), .QN(n7277) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_174_ ( .D(ID_EX_REG_ID_EX_REG_N32), .CK(
        clk), .RN(n7779), .QN(n7276) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_175_ ( .D(ID_EX_REG_ID_EX_REG_N31), .CK(
        clk), .RN(n7779), .QN(n7275) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_178_ ( .D(ID_EX_REG_ID_EX_REG_N28), .CK(
        clk), .RN(n7779), .QN(n7272) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_182_ ( .D(ID_EX_REG_ID_EX_REG_N24), .CK(
        clk), .RN(n7779), .QN(n6842) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_183_ ( .D(ID_EX_REG_ID_EX_REG_N23), .CK(
        clk), .RN(n7779), .QN(n6841) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_189_ ( .D(ID_EX_REG_ID_EX_REG_N17), .CK(
        clk), .RN(n7779), .QN(n6835) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_145_ ( .D(ID_EX_REG_ID_EX_REG_N61), .CK(
        clk), .RN(n7779), .Q(ID_EXEC_OUT[145]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_144_ ( .D(ID_EX_REG_ID_EX_REG_N62), .CK(
        clk), .RN(n7779), .Q(EXEC_MEM_IN[102]), .QN(n6031) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_112_ ( .D(ID_EX_REG_ID_EX_REG_N94), .CK(
        clk), .RN(n7778), .QN(n6847) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_193_ ( .D(ID_EX_REG_ID_EX_REG_N94), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[193]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_113_ ( .D(ID_EX_REG_ID_EX_REG_N93), .CK(
        clk), .RN(n7778), .QN(n6855) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_194_ ( .D(ID_EX_REG_ID_EX_REG_N93), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[194]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_32_ ( .D(ID_EX_REG_ID_EX_REG_N174), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[32]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_33_ ( .D(ID_EX_REG_ID_EX_REG_N173), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[33]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_34_ ( .D(ID_EX_REG_ID_EX_REG_N172), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[34]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_35_ ( .D(ID_EX_REG_ID_EX_REG_N171), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[35]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_36_ ( .D(ID_EX_REG_ID_EX_REG_N170), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[36]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_37_ ( .D(ID_EX_REG_ID_EX_REG_N169), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[37]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_38_ ( .D(ID_EX_REG_ID_EX_REG_N168), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[38]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_39_ ( .D(ID_EX_REG_ID_EX_REG_N167), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[39]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_40_ ( .D(ID_EX_REG_ID_EX_REG_N166), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[40]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_41_ ( .D(ID_EX_REG_ID_EX_REG_N165), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[41]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_42_ ( .D(ID_EX_REG_ID_EX_REG_N164), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[42]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_43_ ( .D(ID_EX_REG_ID_EX_REG_N163), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[43]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_44_ ( .D(ID_EX_REG_ID_EX_REG_N162), .CK(
        clk), .RN(n7777), .Q(ID_EXEC_OUT[44]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_45_ ( .D(ID_EX_REG_ID_EX_REG_N161), .CK(
        clk), .RN(n7777), .Q(ID_EXEC_OUT[45]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_46_ ( .D(ID_EX_REG_ID_EX_REG_N160), .CK(
        clk), .RN(n7777), .Q(ID_EXEC_OUT[46]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_47_ ( .D(ID_EX_REG_ID_EX_REG_N159), .CK(
        clk), .RN(n7777), .Q(ID_EXEC_OUT[47]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_50_ ( .D(ID_EX_REG_ID_EX_REG_N156), .CK(
        clk), .RN(n7777), .Q(ID_EXEC_OUT[50]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_54_ ( .D(ID_EX_REG_ID_EX_REG_N152), .CK(
        clk), .RN(n7777), .Q(ID_EXEC_OUT[54]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_55_ ( .D(ID_EX_REG_ID_EX_REG_N151), .CK(
        clk), .RN(n7777), .Q(ID_EXEC_OUT[55]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_61_ ( .D(ID_EX_REG_ID_EX_REG_N145), .CK(
        clk), .RN(n7777), .Q(ID_EXEC_OUT[61]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_107_ ( .D(ID_EX_REG_ID_EX_REG_N99), .CK(
        clk), .RN(n7777), .QN(n6845) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_133_ ( .D(ID_EX_REG_ID_EX_REG_N99), .CK(
        clk), .RN(n7777), .QN(n7298) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_108_ ( .D(ID_EX_REG_ID_EX_REG_N98), .CK(
        clk), .RN(n7777), .QN(n6850) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_134_ ( .D(ID_EX_REG_ID_EX_REG_N98), .CK(
        clk), .RN(n7777), .QN(n7303) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_60_ ( .D(ID_EX_REG_ID_EX_REG_N146), .CK(
        clk), .RN(n7777), .Q(ID_EXEC_OUT[60]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_92_ ( .D(n1584), .CK(clk), .RN(n7777), 
        .Q(ID_EXEC_OUT[92]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_110_ ( .D(ID_EX_REG_ID_EX_REG_N96), .CK(
        clk), .RN(n7777), .QN(n6848) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_136_ ( .D(ID_EX_REG_ID_EX_REG_N96), .CK(
        clk), .RN(n7777), .QN(n7300) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_62_ ( .D(ID_EX_REG_ID_EX_REG_N144), .CK(
        clk), .RN(n7793), .Q(ID_EXEC_OUT[62]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_94_ ( .D(n1585), .CK(clk), .RN(n7777), 
        .Q(ID_EXEC_OUT[94]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_111_ ( .D(ID_EX_REG_ID_EX_REG_N95), .CK(
        clk), .RN(n7789), .QN(n6846) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_137_ ( .D(ID_EX_REG_ID_EX_REG_N95), .CK(
        clk), .RN(n7784), .QN(n7302) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_63_ ( .D(ID_EX_REG_ID_EX_REG_N143), .CK(
        clk), .RN(n7781), .Q(ID_EXEC_OUT[63]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_122_ ( .D(ID_EX_REG_ID_EX_REG_N84), .CK(
        clk), .RN(n7788), .Q(EXEC_STAGE_imm16_32_16_), .QN(n6833) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_96_ ( .D(ID_EX_REG_ID_EX_REG_N84), .CK(
        clk), .RN(n7785), .Q(EXEC_STAGE_imm26_32[6]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_48_ ( .D(ID_EX_REG_ID_EX_REG_N158), .CK(
        clk), .RN(n7792), .Q(ID_EXEC_OUT[48]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_80_ ( .D(n1578), .CK(clk), .RN(n7780), 
        .Q(ID_EXEC_OUT[80]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_114_ ( .D(ID_EX_REG_ID_EX_REG_N92), .CK(
        clk), .RN(n7789), .QN(n6853) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_195_ ( .D(ID_EX_REG_ID_EX_REG_N92), .CK(
        clk), .RN(n7786), .Q(ID_EXEC_OUT[195]), .QN(n7332) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_123_ ( .D(ID_EX_REG_ID_EX_REG_N83), .CK(
        clk), .RN(n7786), .QN(n7289) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_97_ ( .D(ID_EX_REG_ID_EX_REG_N83), .CK(
        clk), .RN(n7787), .Q(EXEC_STAGE_imm26_32[7]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_49_ ( .D(ID_EX_REG_ID_EX_REG_N157), .CK(
        clk), .RN(n7791), .Q(ID_EXEC_OUT[49]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_81_ ( .D(n1579), .CK(clk), .RN(n7790), 
        .Q(ID_EXEC_OUT[81]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_125_ ( .D(ID_EX_REG_ID_EX_REG_N81), .CK(
        clk), .RN(n7782), .QN(n7293) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_99_ ( .D(ID_EX_REG_ID_EX_REG_N81), .CK(
        clk), .RN(n7783), .Q(EXEC_STAGE_imm26_32[9]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_126_ ( .D(ID_EX_REG_ID_EX_REG_N80), .CK(
        clk), .RN(n7776), .QN(n7292) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_100_ ( .D(ID_EX_REG_ID_EX_REG_N80), .CK(
        clk), .RN(n7776), .Q(EXEC_STAGE_imm26_32[10]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_52_ ( .D(ID_EX_REG_ID_EX_REG_N154), .CK(
        clk), .RN(n7776), .Q(ID_EXEC_OUT[52]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_84_ ( .D(n1581), .CK(clk), .RN(n7776), 
        .Q(ID_EXEC_OUT[84]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_127_ ( .D(ID_EX_REG_ID_EX_REG_N79), .CK(
        clk), .RN(n7776), .QN(n7290) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_101_ ( .D(ID_EX_REG_ID_EX_REG_N79), .CK(
        clk), .RN(n7776), .Q(EXEC_STAGE_imm26_32[11]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_53_ ( .D(ID_EX_REG_ID_EX_REG_N153), .CK(
        clk), .RN(n7776), .Q(ID_EXEC_OUT[53]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_85_ ( .D(n1582), .CK(clk), .RN(n7776), 
        .Q(ID_EXEC_OUT[85]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_130_ ( .D(ID_EX_REG_ID_EX_REG_N76), .CK(
        clk), .RN(n7776), .QN(n7297) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_104_ ( .D(ID_EX_REG_ID_EX_REG_N76), .CK(
        clk), .RN(n7776), .Q(EXEC_STAGE_imm26_32[14]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_56_ ( .D(ID_EX_REG_ID_EX_REG_N150), .CK(
        clk), .RN(n7776), .Q(ID_EXEC_OUT[56]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_88_ ( .D(n1583), .CK(clk), .RN(n7776), 
        .QN(n7227) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_115_ ( .D(ID_EX_REG_ID_EX_REG_N91), .CK(
        clk), .RN(n7776), .QN(n6852) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_196_ ( .D(ID_EX_REG_ID_EX_REG_N91), .CK(
        clk), .RN(n7776), .Q(ID_EXEC_OUT[196]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_105_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N77), .CK(clk), .RN(n7776), .Q(
        DMEM_BUS_OUT[64]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_140_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N42), .CK(clk), .RN(n7776), .QN(n7283) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[31]), .QN(n6477) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_31_ ( .D(ID_EX_REG_ID_EX_REG_N175), .CK(
        clk), .RN(n7775), .Q(nextPC_ex_out[31]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_139_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N43), .CK(clk), .RN(n7775), .QN(n7282) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[30]), .QN(n6476) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_30_ ( .D(ID_EX_REG_ID_EX_REG_N176), .CK(
        clk), .RN(n7775), .Q(nextPC_ex_out[30]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_138_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N44), .CK(clk), .RN(n7775), .Q(
        EXEC_MEM_OUT_138) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[29]), .QN(n6882) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_29_ ( .D(ID_EX_REG_ID_EX_REG_N177), .CK(
        clk), .RN(n7775), .Q(nextPC_ex_out[29]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_28_ ( .D(ID_EX_REG_ID_EX_REG_N178), .CK(
        clk), .RN(n7775), .Q(nextPC_ex_out[28]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_137_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N45), .CK(clk), .RN(n7775), .Q(
        EXEC_MEM_OUT_137) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[28]), .QN(n6890) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_96_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N86), .CK(clk), .RN(n7775), .Q(
        DMEM_BUS_OUT[27]), .QN(n5912) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_64_ ( .D(DMEM_BUS_OUT[27]), .CK(clk), 
        .RN(n7775), .Q(MEM_WB_OUT[64]), .QN(n6324) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5947) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__27_), .QN(n6647) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__27_), .QN(n6549) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__27_), .QN(n6724) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5949) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__27_), .QN(n6576) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__27_), .QN(n6609) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__27_), .QN(n7143) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__27_), .QN(n6508) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__27_), .QN(n6755) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5874) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__27_), .QN(n6210) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__27_), .QN(n6754) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__27_), .QN(n6159) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5946) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__27_), .QN(n6646) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__27_), .QN(n7049) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6923) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5935) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__27_), .QN(n6575) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6131) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__27_), .QN(n6645) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6409) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6962) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__27_), .QN(n7109) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__27_), .QN(n7142) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__27_), .QN(n7016) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6924) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__27_), .QN(n7050) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__27_), .QN(n6753) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__27_), .QN(n6494) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__27_), .QN(n7110) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_187_ ( .D(ID_EX_REG_ID_EX_REG_N19), .CK(
        clk), .RN(n7775), .QN(n6837) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_91_ ( .D(ID_EX_REG_ID_EX_REG_N115), .CK(
        clk), .RN(n7775), .Q(ID_EXEC_OUT[91]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_59_ ( .D(ID_EX_REG_ID_EX_REG_N147), .CK(
        clk), .RN(n7777), .Q(ID_EXEC_OUT[59]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_136_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N46), .CK(clk), .RN(n7792), .Q(
        EXEC_MEM_OUT_136) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[27]), .QN(n6905) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_27_ ( .D(ID_EX_REG_ID_EX_REG_N179), .CK(
        clk), .RN(n7778), .Q(nextPC_ex_out[27]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_95_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N87), .CK(clk), .RN(n7783), .Q(
        DMEM_BUS_OUT[26]), .QN(n5924) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_63_ ( .D(DMEM_BUS_OUT[26]), .CK(clk), 
        .RN(n7778), .Q(MEM_WB_OUT[63]), .QN(n6322) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6411) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__26_), .QN(n6649) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__26_), .QN(n6548) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__26_), .QN(n6723) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6451) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__26_), .QN(n6578) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__26_), .QN(n6608) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__26_), .QN(n6722) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__26_), .QN(n7017) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__26_), .QN(n6752) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5875) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__26_), .QN(n6211) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__26_), .QN(n7182) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__26_), .QN(n6160) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5896) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__26_), .QN(n7111) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__26_), .QN(n7051) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6926) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6925) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__26_), .QN(n6577) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6981) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__26_), .QN(n6648) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6410) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5933) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__26_), .QN(n7079) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__26_), .QN(n7141) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__26_), .QN(n7018) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6063) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__26_), .QN(n7052) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__26_), .QN(n6751) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__26_), .QN(n6495) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__26_), .QN(n7080) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_186_ ( .D(ID_EX_REG_ID_EX_REG_N20), .CK(
        clk), .RN(n7781), .QN(n6838) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_90_ ( .D(ID_EX_REG_ID_EX_REG_N116), .CK(
        clk), .RN(n7784), .Q(ID_EXEC_OUT[90]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_58_ ( .D(ID_EX_REG_ID_EX_REG_N148), .CK(
        clk), .RN(n7787), .Q(ID_EXEC_OUT[58]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_135_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N47), .CK(clk), .RN(n7787), .Q(
        EXEC_MEM_OUT_135) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_26_ ( .D(ID_EX_REG_ID_EX_REG_N180), .CK(
        clk), .RN(n7787), .Q(nextPC_ex_out[26]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_94_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N88), .CK(clk), .RN(n7787), .Q(
        DMEM_BUS_OUT[25]), .QN(n5916) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_62_ ( .D(DMEM_BUS_OUT[25]), .CK(clk), 
        .RN(n7787), .Q(MEM_WB_OUT[62]), .QN(n6323) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6412) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__25_), .QN(n7114) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__25_), .QN(n6547) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__25_), .QN(n6721) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6452) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__25_), .QN(n6581) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__25_), .QN(n6244) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__25_), .QN(n6720) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__25_), .QN(n7019) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__25_), .QN(n7181) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5895) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__25_), .QN(n6212) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__25_), .QN(n7180) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__25_), .QN(n5963) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6103) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__25_), .QN(n7113) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__25_), .QN(n6579) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6381) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6380) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__25_), .QN(n6580) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6125) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__25_), .QN(n7112) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6963) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6054) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__25_), .QN(n7081) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__25_), .QN(n7140) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__25_), .QN(n7020) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6064) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__25_), .QN(n6582) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__25_), .QN(n7179) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__25_), .QN(n6161) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__25_), .QN(n7082) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_185_ ( .D(ID_EX_REG_ID_EX_REG_N21), .CK(
        clk), .RN(n7787), .QN(n6839) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_89_ ( .D(ID_EX_REG_ID_EX_REG_N117), .CK(
        clk), .RN(n7787), .Q(ID_EXEC_OUT[89]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_57_ ( .D(ID_EX_REG_ID_EX_REG_N149), .CK(
        clk), .RN(n7787), .Q(ID_EXEC_OUT[57]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_134_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N48), .CK(clk), .RN(n7787), .Q(
        EXEC_MEM_OUT_134) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[25]), .QN(n6915) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_25_ ( .D(ID_EX_REG_ID_EX_REG_N181), .CK(
        clk), .RN(n7787), .Q(nextPC_ex_out[25]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_133_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N49), .CK(clk), .RN(n7787), .Q(
        EXEC_MEM_OUT_133) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[24]), .QN(n6885) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_24_ ( .D(ID_EX_REG_ID_EX_REG_N182), .CK(
        clk), .RN(n7787), .Q(nextPC_ex_out[24]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_132_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N50), .CK(clk), .RN(n7787), .Q(
        EXEC_MEM_OUT_132) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[23]), .QN(n6910) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_23_ ( .D(ID_EX_REG_ID_EX_REG_N183), .CK(
        clk), .RN(n7787), .Q(nextPC_ex_out[23]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_22_ ( .D(n1550), .CK(clk), .RN(n7786), 
        .Q(IF_ID_OUT[22]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_22_ ( .D(ID_EX_REG_ID_EX_REG_N184), .CK(
        clk), .RN(n7786), .Q(nextPC_ex_out[22]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_131_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N51), .CK(clk), .RN(n7786), .Q(
        EXEC_MEM_OUT_131) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_21_ ( .D(n1551), .CK(clk), .RN(n7786), 
        .Q(IF_ID_OUT[21]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_21_ ( .D(ID_EX_REG_ID_EX_REG_N185), .CK(
        clk), .RN(n7786), .Q(nextPC_ex_out[21]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_130_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N52), .CK(clk), .RN(n7786), .Q(
        EXEC_MEM_OUT_130) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[21]), .QN(n6914) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_20_ ( .D(ID_EX_REG_ID_EX_REG_N186), .CK(
        clk), .RN(n7786), .Q(nextPC_ex_out[20]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_129_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N53), .CK(clk), .RN(n7786), .Q(
        EXEC_MEM_OUT_129) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[20]), .QN(n6884) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_88_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N94), .CK(clk), .RN(n7786), .Q(
        DMEM_BUS_OUT[19]), .QN(n6026) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_56_ ( .D(DMEM_BUS_OUT[19]), .CK(clk), 
        .RN(n7786), .Q(MEM_WB_OUT[56]), .QN(n6812) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6431) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__19_), .QN(n7121) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__19_), .QN(n6546) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__19_), .QN(n6719) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6454) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__19_), .QN(n6588) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__19_), .QN(n7091) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__19_), .QN(n6718) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__19_), .QN(n6514) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_2__19_), .QN(n6302) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5937) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_28__19_), .QN(n6222) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__19_), .QN(n6750) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__19_), .QN(n6166) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6430) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__19_), .QN(n6672) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__19_), .QN(n6586) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6386) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6385) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__19_), .QN(n6587) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6987) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__19_), .QN(n7118) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6967) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n6966) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__19_), .QN(n7119) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__19_), .QN(n6717) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__19_), .QN(n7026) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n5938) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__19_), .QN(n6589) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__19_), .QN(n7178) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__19_), .QN(n6167) );
  DFF_X1 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__19_), .QN(n7120) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_179_ ( .D(ID_EX_REG_ID_EX_REG_N27), .CK(
        clk), .RN(n7786), .QN(n7271) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_83_ ( .D(n1580), .CK(clk), .RN(n7786), 
        .Q(ID_EXEC_OUT[83]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_51_ ( .D(ID_EX_REG_ID_EX_REG_N155), .CK(
        clk), .RN(n7786), .Q(ID_EXEC_OUT[51]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_128_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N54), .CK(clk), .RN(n7786), .Q(
        EXEC_MEM_OUT_128) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[19]), .QN(n6909) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_19_ ( .D(ID_EX_REG_ID_EX_REG_N187), .CK(
        clk), .RN(n7786), .Q(nextPC_ex_out[19]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_18_ ( .D(ID_EX_REG_ID_EX_REG_N188), .CK(
        clk), .RN(n7785), .Q(nextPC_ex_out[18]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_127_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N55), .CK(clk), .RN(n7785), .Q(
        EXEC_MEM_OUT_127) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[18]), .QN(n6877) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_17_ ( .D(ID_EX_REG_ID_EX_REG_N189), .CK(
        clk), .RN(n7785), .Q(nextPC_ex_out[17]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_126_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N56), .CK(clk), .RN(n7785), .Q(
        EXEC_MEM_OUT_126) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[17]), .QN(n6041) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_16_ ( .D(ID_EX_REG_ID_EX_REG_N190), .CK(
        clk), .RN(n7785), .Q(nextPC_ex_out[16]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_125_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N57), .CK(clk), .RN(n7785), .Q(
        EXEC_MEM_OUT_125) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[16]), .QN(n6021) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_15_ ( .D(ID_EX_REG_ID_EX_REG_N191), .CK(
        clk), .RN(n7785), .QN(n7215) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_124_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N58), .CK(clk), .RN(n7785), .Q(
        EXEC_MEM_OUT_124) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[15]), .QN(n6039) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_14_ ( .D(ID_EX_REG_ID_EX_REG_N192), .CK(
        clk), .RN(n7785), .Q(nextPC_ex_out[14]), .QN(n7136) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_123_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N59), .CK(clk), .RN(n7785), .Q(
        EXEC_MEM_OUT_123) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[14]), .QN(n5909) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_13_ ( .D(ID_EX_REG_ID_EX_REG_N193), .CK(
        clk), .RN(n7785), .Q(nextPC_ex_out[13]), .QN(n7137) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_122_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N60), .CK(clk), .RN(n7784), .Q(
        EXEC_MEM_OUT_122) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[13]), .QN(n6040) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_12_ ( .D(ID_EX_REG_ID_EX_REG_N194), .CK(
        clk), .RN(n7784), .QN(n7211) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_121_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N61), .CK(clk), .RN(n7784), .Q(
        EXEC_MEM_OUT_121) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[12]), .QN(n6020) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_11_ ( .D(ID_EX_REG_ID_EX_REG_N195), .CK(
        clk), .RN(n7784), .Q(nextPC_ex_out[11]), .QN(n7221) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_120_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N62), .CK(clk), .RN(n7784), .Q(
        EXEC_MEM_OUT_120) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[11]), .QN(n6038) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_10_ ( .D(ID_EX_REG_ID_EX_REG_N196), .CK(
        clk), .RN(n7784), .Q(nextPC_ex_out[10]), .QN(n6801) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_119_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N63), .CK(clk), .RN(n7784), .Q(
        EXEC_MEM_OUT_119) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_9_ ( .D(ID_EX_REG_ID_EX_REG_N197), .CK(
        clk), .RN(n7784), .Q(nextPC_ex_out[9]), .QN(n6802) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_118_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N64), .CK(clk), .RN(n7784), .Q(
        EXEC_MEM_OUT_118) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[9]), .QN(n6907) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_8_ ( .D(ID_EX_REG_ID_EX_REG_N198), .CK(
        clk), .RN(n7784), .Q(nextPC_ex_out[8]), .QN(n7222) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_117_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N65), .CK(clk), .RN(n7784), .Q(
        EXEC_MEM_OUT_117) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[8]), .QN(n6888) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_7_ ( .D(ID_EX_REG_ID_EX_REG_N199), .CK(
        clk), .RN(n7778), .Q(nextPC_ex_out[7]), .QN(n6803) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_116_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N66), .CK(clk), .RN(n7786), .Q(
        EXEC_MEM_OUT_116) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[7]), .QN(n6902) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_6_ ( .D(ID_EX_REG_ID_EX_REG_N200), .CK(
        clk), .RN(n7793), .Q(nextPC_ex_out[6]), .QN(n6699) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_115_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N67), .CK(clk), .RN(n7783), .Q(
        EXEC_MEM_OUT_115) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[6]), .QN(n6015) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_5_ ( .D(ID_EX_REG_ID_EX_REG_N201), .CK(
        clk), .RN(n7784), .QN(n7212) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_114_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N68), .CK(clk), .RN(n7788), .Q(
        EXEC_MEM_OUT_114) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[5]), .QN(n6906) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_4_ ( .D(ID_EX_REG_ID_EX_REG_N202), .CK(
        clk), .RN(n7785), .Q(nextPC_ex_out[4]), .QN(n7220) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_113_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N69), .CK(clk), .RN(n7782), .Q(
        EXEC_MEM_OUT_113) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[4]), .QN(n6887) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_3_ ( .D(ID_EX_REG_ID_EX_REG_N203), .CK(
        clk), .RN(n7790), .Q(nextPC_ex_out[3]), .QN(n7217) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_112_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N70), .CK(clk), .RN(n7791), .Q(
        EXEC_MEM_OUT_112) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[3]), .QN(n6901) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_2_ ( .D(ID_EX_REG_ID_EX_REG_N204), .CK(
        clk), .RN(n7779), .Q(nextPC_ex_out[2]), .QN(n7219) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_111_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N71), .CK(clk), .RN(n7783), .Q(
        EXEC_MEM_OUT_111) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[2]), .QN(n6894) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_1_ ( .D(ID_EX_REG_ID_EX_REG_N205), .CK(
        clk), .RN(n7783), .Q(nextPC_ex_out[1]), .QN(n7218) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_110_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N72), .CK(clk), .RN(n7783), .Q(
        EXEC_MEM_OUT_110) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[1]), .QN(n6995) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_0_ ( .D(ID_EX_REG_ID_EX_REG_N206), .CK(
        clk), .RN(n7783), .Q(nextPC_ex_out[0]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_109_ ( .D(n10296), .CK(clk), .RN(
        n7783), .Q(EXEC_MEM_OUT_109) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[0]), .QN(n7135) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_173_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N9), .CK(clk), .RN(n7783), .Q(
        DMEM_BUS_OUT[63]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_142_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N40), .CK(clk), .RN(n7783), .Q(
        DMEM_BUS_OUT[32]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_143_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N39), .CK(clk), .RN(n7783), .Q(
        DMEM_BUS_OUT[33]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_144_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N38), .CK(clk), .RN(n7783), .Q(
        DMEM_BUS_OUT[34]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_145_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N37), .CK(clk), .RN(n7783), .Q(
        DMEM_BUS_OUT[35]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_146_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N36), .CK(clk), .RN(n7783), .Q(
        DMEM_BUS_OUT[36]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_147_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N35), .CK(clk), .RN(n7783), .Q(
        DMEM_BUS_OUT[37]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_148_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N34), .CK(clk), .RN(n7783), .Q(
        DMEM_BUS_OUT[38]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_149_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N33), .CK(clk), .RN(n7783), .Q(
        DMEM_BUS_OUT[39]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_150_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N32), .CK(clk), .RN(n7783), .Q(
        DMEM_BUS_OUT[40]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_151_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N31), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[41]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_152_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N30), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[42]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_153_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N29), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[43]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_154_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N28), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[44]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_155_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N27), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[45]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_156_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N26), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[46]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_157_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N25), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[47]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_158_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N24), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[48]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_159_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N23), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[49]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_160_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N22), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[50]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_161_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N21), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[51]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_162_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N20), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[52]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_163_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N19), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[53]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_164_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N18), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[54]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_165_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N17), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[55]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_166_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N16), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[56]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_167_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N15), .CK(clk), .RN(n7782), .Q(
        DMEM_BUS_OUT[57]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_168_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N14), .CK(clk), .RN(n7781), .Q(
        DMEM_BUS_OUT[58]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_169_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N13), .CK(clk), .RN(n7781), .Q(
        DMEM_BUS_OUT[59]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_170_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N12), .CK(clk), .RN(n7781), .Q(
        DMEM_BUS_OUT[60]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_171_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N11), .CK(clk), .RN(n7784), .Q(
        DMEM_BUS_OUT[61]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_172_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N10), .CK(clk), .RN(n7775), .Q(
        DMEM_BUS_OUT[62]) );
  OAI22_X2 U3 ( .A1(n7761), .A2(n6950), .B1(n7760), .B2(n7758), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U4 ( .A1(n7761), .A2(n6949), .B1(n7760), .B2(n5868), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5 ( .A1(n7761), .A2(n6948), .B1(n7760), .B2(n7756), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6 ( .A1(n7761), .A2(n6405), .B1(n7760), .B2(n5867), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7 ( .A1(n7761), .A2(n6947), .B1(n7760), .B2(n7754), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U10 ( .A1(n7761), .A2(n6946), .B1(n7760), .B2(n5866), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U21 ( .A1(n7761), .A2(n6102), .B1(n7760), .B2(n7752), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U32 ( .A1(n7761), .A2(n6101), .B1(n7760), .B2(n7750), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U37 ( .A1(n7757), .A2(n7747), .B1(n7745), .B2(n6261), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U38 ( .A1(n5868), .A2(n7747), .B1(n7745), .B2(n6260), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U39 ( .A1(n7755), .A2(n7747), .B1(n7746), .B2(n6259), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U40 ( .A1(n5867), .A2(n7747), .B1(n7745), .B2(n6258), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U41 ( .A1(n7753), .A2(n7747), .B1(n7746), .B2(n6002), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U44 ( .A1(n5866), .A2(n7747), .B1(n7745), .B2(n6001), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U55 ( .A1(n7751), .A2(n7747), .B1(n7745), .B2(n6000), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U66 ( .A1(n7749), .A2(n3078), .B1(n7746), .B2(n6257), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U71 ( .A1(n7757), .A2(n7743), .B1(n7742), .B2(n6529), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U72 ( .A1(n5868), .A2(n7744), .B1(n7742), .B2(n6528), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U73 ( .A1(n7755), .A2(n7743), .B1(n7742), .B2(n6527), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U74 ( .A1(n5867), .A2(n7744), .B1(n7742), .B2(n6526), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U75 ( .A1(n7753), .A2(n7743), .B1(n7742), .B2(n6525), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U78 ( .A1(n5866), .A2(n7744), .B1(n7742), .B2(n6524), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U89 ( .A1(n7751), .A2(n7743), .B1(n7742), .B2(n6523), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U100 ( .A1(n7749), .A2(n7744), .B1(n7742), .B2(n6522), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U105 ( .A1(n7757), .A2(n7740), .B1(n7738), .B2(n6716), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U106 ( .A1(n5868), .A2(n7739), .B1(n7738), .B2(n6715), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U107 ( .A1(n7755), .A2(n7740), .B1(n7738), .B2(n6714), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U108 ( .A1(n5867), .A2(n7739), .B1(n7738), .B2(n6713), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U109 ( .A1(n7753), .A2(n7740), .B1(n7738), .B2(n6712), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U112 ( .A1(n5866), .A2(n7739), .B1(n7738), .B2(n6711), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U123 ( .A1(n7751), .A2(n7740), .B1(n7738), .B2(n6710), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U134 ( .A1(n7749), .A2(n7739), .B1(n7738), .B2(n6709), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U139 ( .A1(n7757), .A2(n7735), .B1(n7734), .B2(n5881), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U140 ( .A1(n5868), .A2(n7736), .B1(n7734), .B2(n6117), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U141 ( .A1(n7755), .A2(n7735), .B1(n7734), .B2(n6116), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U142 ( .A1(n5867), .A2(n7736), .B1(n7734), .B2(n6115), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U143 ( .A1(n7753), .A2(n7735), .B1(n7734), .B2(n6114), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U146 ( .A1(n5866), .A2(n7736), .B1(n7734), .B2(n6113), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U157 ( .A1(n7751), .A2(n7735), .B1(n7734), .B2(n5880), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U168 ( .A1(n7749), .A2(n7736), .B1(n7734), .B2(n5897), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U173 ( .A1(n7757), .A2(n3090), .B1(n7730), .B2(n5984), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U174 ( .A1(n5868), .A2(n7732), .B1(n7730), .B2(n6198), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U175 ( .A1(n7755), .A2(n3090), .B1(n7730), .B2(n5983), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U176 ( .A1(n5867), .A2(n7732), .B1(n7730), .B2(n6197), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U177 ( .A1(n7753), .A2(n3090), .B1(n7730), .B2(n5982), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U180 ( .A1(n5866), .A2(n7732), .B1(n7730), .B2(n5981), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U191 ( .A1(n7751), .A2(n3090), .B1(n7730), .B2(n5980), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U202 ( .A1(n7749), .A2(n7732), .B1(n7730), .B2(n5979), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U208 ( .A1(n7757), .A2(n7727), .B1(n7726), .B2(n6206), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U209 ( .A1(n5868), .A2(n7727), .B1(n7725), .B2(n6205), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U210 ( .A1(n7755), .A2(n7727), .B1(n7726), .B2(n6204), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U211 ( .A1(n5867), .A2(n7727), .B1(n7725), .B2(n6203), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U212 ( .A1(n7753), .A2(n7727), .B1(n7726), .B2(n6202), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U215 ( .A1(n5866), .A2(n7727), .B1(n7725), .B2(n6201), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U226 ( .A1(n7751), .A2(n7727), .B1(n7725), .B2(n6200), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U237 ( .A1(n7749), .A2(n7727), .B1(n7725), .B2(n6199), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U242 ( .A1(n7757), .A2(n7723), .B1(n7720), .B2(n6275), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U243 ( .A1(n5868), .A2(n7722), .B1(n7721), .B2(n6274), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U244 ( .A1(n7755), .A2(n7723), .B1(n7720), .B2(n6273), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U245 ( .A1(n5867), .A2(n7722), .B1(n7721), .B2(n6272), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U246 ( .A1(n7753), .A2(n7723), .B1(n7720), .B2(n6271), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U249 ( .A1(n5866), .A2(n7722), .B1(n7721), .B2(n6270), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U260 ( .A1(n7751), .A2(n7723), .B1(n7720), .B2(n6269), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U271 ( .A1(n7749), .A2(n7722), .B1(n7721), .B2(n6268), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U273 ( .A1(n3098), .A2(n3084), .ZN(n3096) );
  OAI22_X2 U276 ( .A1(n7757), .A2(n3099), .B1(n7717), .B2(n6158), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U277 ( .A1(n5868), .A2(n7718), .B1(n7716), .B2(n6157), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U278 ( .A1(n7755), .A2(n3099), .B1(n7717), .B2(n6156), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U279 ( .A1(n5867), .A2(n3099), .B1(n7716), .B2(n6155), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U280 ( .A1(n7753), .A2(n3099), .B1(n7717), .B2(n6154), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U283 ( .A1(n5866), .A2(n3099), .B1(n7716), .B2(n6153), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U294 ( .A1(n7751), .A2(n3099), .B1(n7717), .B2(n6152), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U305 ( .A1(n7749), .A2(n3099), .B1(n7716), .B2(n6151), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U307 ( .A1(n3098), .A2(n3087), .ZN(n3099) );
  OAI22_X2 U310 ( .A1(n7757), .A2(n7714), .B1(n7713), .B2(n6300), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U311 ( .A1(n5868), .A2(n7714), .B1(n7712), .B2(n6299), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U312 ( .A1(n7755), .A2(n7714), .B1(n7713), .B2(n6298), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U313 ( .A1(n5867), .A2(n7714), .B1(n7712), .B2(n6297), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U314 ( .A1(n7753), .A2(n7714), .B1(n7713), .B2(n6296), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U317 ( .A1(n5866), .A2(n7714), .B1(n7712), .B2(n6295), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U328 ( .A1(n7751), .A2(n7714), .B1(n7712), .B2(n6294), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U339 ( .A1(n7749), .A2(n7714), .B1(n7712), .B2(n6293), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U344 ( .A1(n7758), .A2(n7710), .B1(n7708), .B2(n5932), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U345 ( .A1(n5868), .A2(n7710), .B1(n7708), .B2(n5931), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U346 ( .A1(n7756), .A2(n7710), .B1(n7709), .B2(n5930), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U347 ( .A1(n5867), .A2(n7710), .B1(n7708), .B2(n5929), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U348 ( .A1(n7754), .A2(n3103), .B1(n7709), .B2(n5928), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U351 ( .A1(n5866), .A2(n7710), .B1(n7708), .B2(n5894), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U362 ( .A1(n7752), .A2(n7710), .B1(n7708), .B2(n5927), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U373 ( .A1(n7750), .A2(n7710), .B1(n7709), .B2(n5893), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U375 ( .A1(n3098), .A2(n3077), .ZN(n3103) );
  OAI22_X2 U378 ( .A1(n7758), .A2(n7706), .B1(n7704), .B2(n5978), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U379 ( .A1(n5868), .A2(n7706), .B1(n7704), .B2(n5977), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U380 ( .A1(n7756), .A2(n7706), .B1(n7705), .B2(n5976), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U381 ( .A1(n5867), .A2(n7706), .B1(n7704), .B2(n5975), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U382 ( .A1(n7754), .A2(n7706), .B1(n7705), .B2(n5905), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U385 ( .A1(n5866), .A2(n7706), .B1(n7704), .B2(n5904), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U396 ( .A1(n7752), .A2(n3105), .B1(n7705), .B2(n5903), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U407 ( .A1(n7750), .A2(n7706), .B1(n7704), .B2(n5902), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U409 ( .A1(n3098), .A2(n3080), .ZN(n3105) );
  OAI22_X2 U413 ( .A1(n7758), .A2(n3107), .B1(n7701), .B2(n6292), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U414 ( .A1(n5868), .A2(n7702), .B1(n7700), .B2(n6291), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U415 ( .A1(n7756), .A2(n3107), .B1(n7701), .B2(n6290), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U416 ( .A1(n5867), .A2(n3107), .B1(n7700), .B2(n6289), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U417 ( .A1(n7754), .A2(n3107), .B1(n7701), .B2(n6288), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U420 ( .A1(n5866), .A2(n3107), .B1(n7700), .B2(n6287), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U431 ( .A1(n7752), .A2(n3107), .B1(n7701), .B2(n6286), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U442 ( .A1(n7750), .A2(n3107), .B1(n7700), .B2(n6285), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U447 ( .A1(n7758), .A2(n3110), .B1(n7697), .B2(n5962), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U448 ( .A1(n5868), .A2(n7698), .B1(n7696), .B2(n5961), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U449 ( .A1(n7756), .A2(n3110), .B1(n7697), .B2(n5960), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U450 ( .A1(n5867), .A2(n3110), .B1(n7696), .B2(n5959), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U451 ( .A1(n7754), .A2(n3110), .B1(n7697), .B2(n5958), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U454 ( .A1(n5866), .A2(n3110), .B1(n7696), .B2(n5957), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U465 ( .A1(n7752), .A2(n3110), .B1(n7697), .B2(n5956), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U476 ( .A1(n7750), .A2(n3110), .B1(n7696), .B2(n5955), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U481 ( .A1(n7758), .A2(n7694), .B1(n7692), .B2(n6100), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U482 ( .A1(n5868), .A2(n7694), .B1(n7692), .B2(n6099), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U483 ( .A1(n7756), .A2(n7694), .B1(n7693), .B2(n6098), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U484 ( .A1(n5867), .A2(n7694), .B1(n7692), .B2(n6097), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U485 ( .A1(n7754), .A2(n7694), .B1(n7693), .B2(n6096), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U488 ( .A1(n5866), .A2(n7694), .B1(n7692), .B2(n6095), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U499 ( .A1(n7752), .A2(n7694), .B1(n7693), .B2(n6094), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U510 ( .A1(n7750), .A2(n7694), .B1(n7692), .B2(n5945), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U515 ( .A1(n7758), .A2(n7690), .B1(n7688), .B2(n6256), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U516 ( .A1(n5868), .A2(n7690), .B1(n7688), .B2(n6255), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U517 ( .A1(n7756), .A2(n7690), .B1(n7689), .B2(n6254), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U518 ( .A1(n5867), .A2(n7690), .B1(n7688), .B2(n6253), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U519 ( .A1(n7754), .A2(n7690), .B1(n7689), .B2(n5999), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U522 ( .A1(n5866), .A2(n7690), .B1(n7688), .B2(n5998), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U533 ( .A1(n7752), .A2(n7690), .B1(n7688), .B2(n5997), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U544 ( .A1(n7750), .A2(n7690), .B1(n7689), .B2(n5996), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U550 ( .A1(n7758), .A2(n7686), .B1(n7685), .B2(n6545), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U551 ( .A1(n5868), .A2(n7687), .B1(n7685), .B2(n6544), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U552 ( .A1(n7756), .A2(n7686), .B1(n7685), .B2(n6543), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U553 ( .A1(n5867), .A2(n7687), .B1(n7685), .B2(n6542), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U554 ( .A1(n7754), .A2(n7686), .B1(n7685), .B2(n6541), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U557 ( .A1(n5866), .A2(n7687), .B1(n7685), .B2(n6540), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U568 ( .A1(n7752), .A2(n7686), .B1(n7685), .B2(n6539), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U579 ( .A1(n7750), .A2(n7687), .B1(n7685), .B2(n6538), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U584 ( .A1(n7758), .A2(n7682), .B1(n7681), .B2(n6370), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U585 ( .A1(n5868), .A2(n7683), .B1(n7681), .B2(n6369), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U586 ( .A1(n7756), .A2(n7682), .B1(n7681), .B2(n6368), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U587 ( .A1(n5867), .A2(n7683), .B1(n7681), .B2(n6367), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U588 ( .A1(n7754), .A2(n7682), .B1(n7681), .B2(n6366), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U591 ( .A1(n5866), .A2(n7683), .B1(n7681), .B2(n6365), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U602 ( .A1(n7752), .A2(n7682), .B1(n7681), .B2(n6364), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U613 ( .A1(n7750), .A2(n7683), .B1(n7681), .B2(n6363), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U618 ( .A1(n7758), .A2(n7678), .B1(n7677), .B2(n5870), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U619 ( .A1(n5868), .A2(n7679), .B1(n7677), .B2(n6053), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U620 ( .A1(n7756), .A2(n7678), .B1(n7677), .B2(n6052), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U621 ( .A1(n5867), .A2(n7679), .B1(n7677), .B2(n6051), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U622 ( .A1(n7754), .A2(n7678), .B1(n7677), .B2(n6050), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U625 ( .A1(n5866), .A2(n7679), .B1(n7677), .B2(n6049), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U636 ( .A1(n7752), .A2(n7678), .B1(n7677), .B2(n6048), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U647 ( .A1(n7750), .A2(n7679), .B1(n7677), .B2(n5892), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U652 ( .A1(n7758), .A2(n7674), .B1(n7673), .B2(n6196), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U653 ( .A1(n5868), .A2(n7675), .B1(n7673), .B2(n6195), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U654 ( .A1(n7756), .A2(n7674), .B1(n7673), .B2(n6194), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U655 ( .A1(n5867), .A2(n7675), .B1(n7673), .B2(n6193), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U656 ( .A1(n7754), .A2(n7674), .B1(n7673), .B2(n5901), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U659 ( .A1(n5866), .A2(n7675), .B1(n7673), .B2(n5974), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U670 ( .A1(n7752), .A2(n7674), .B1(n7673), .B2(n5900), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U681 ( .A1(n7750), .A2(n7675), .B1(n7673), .B2(n5973), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U687 ( .A1(n7758), .A2(n7670), .B1(n7669), .B2(n6129), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U688 ( .A1(n5868), .A2(n7670), .B1(n7669), .B2(n6466), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U689 ( .A1(n7756), .A2(n7670), .B1(n7669), .B2(n6465), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U690 ( .A1(n5867), .A2(n7670), .B1(n7669), .B2(n6464), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U691 ( .A1(n7754), .A2(n7670), .B1(n7668), .B2(n6463), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U694 ( .A1(n5866), .A2(n7670), .B1(n7669), .B2(n6462), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U705 ( .A1(n7752), .A2(n7670), .B1(n7668), .B2(n6128), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U716 ( .A1(n7750), .A2(n7670), .B1(n7669), .B2(n5954), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U721 ( .A1(n7757), .A2(n3128), .B1(n7665), .B2(n6252), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U722 ( .A1(n5868), .A2(n7666), .B1(n7664), .B2(n6251), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U723 ( .A1(n7755), .A2(n3128), .B1(n7665), .B2(n6250), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U724 ( .A1(n5867), .A2(n3128), .B1(n7664), .B2(n6249), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U725 ( .A1(n7753), .A2(n3128), .B1(n7665), .B2(n6248), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U728 ( .A1(n5866), .A2(n3128), .B1(n7664), .B2(n6247), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U739 ( .A1(n7751), .A2(n3128), .B1(n7665), .B2(n6246), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U750 ( .A1(n7749), .A2(n3128), .B1(n7664), .B2(n6245), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U755 ( .A1(n7757), .A2(n3131), .B1(n7661), .B2(n6093), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U756 ( .A1(n5868), .A2(n7662), .B1(n7660), .B2(n6092), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U757 ( .A1(n7755), .A2(n3131), .B1(n7661), .B2(n6091), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U758 ( .A1(n5867), .A2(n3131), .B1(n7660), .B2(n6090), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U759 ( .A1(n7753), .A2(n3131), .B1(n7661), .B2(n6089), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U762 ( .A1(n5866), .A2(n3131), .B1(n7660), .B2(n6088), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U773 ( .A1(n7751), .A2(n3131), .B1(n7661), .B2(n6087), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U784 ( .A1(n7749), .A2(n3131), .B1(n7660), .B2(n6086), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U789 ( .A1(n7757), .A2(n7658), .B1(n7657), .B2(n6085), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U790 ( .A1(n5868), .A2(n7658), .B1(n7657), .B2(n6404), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U791 ( .A1(n7755), .A2(n7658), .B1(n7657), .B2(n6403), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U792 ( .A1(n5867), .A2(n7658), .B1(n7657), .B2(n6402), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U793 ( .A1(n7753), .A2(n7658), .B1(n7656), .B2(n6401), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U796 ( .A1(n5866), .A2(n7658), .B1(n7657), .B2(n6400), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U807 ( .A1(n7751), .A2(n7658), .B1(n7656), .B2(n6399), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U818 ( .A1(n7749), .A2(n7658), .B1(n7657), .B2(n5944), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U823 ( .A1(n7757), .A2(n7654), .B1(n7653), .B2(n6638), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U824 ( .A1(n5868), .A2(n7654), .B1(n7653), .B2(n6637), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U825 ( .A1(n7755), .A2(n7654), .B1(n7653), .B2(n6636), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U826 ( .A1(n5867), .A2(n7654), .B1(n7653), .B2(n6635), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U827 ( .A1(n7753), .A2(n7654), .B1(n7652), .B2(n6634), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U830 ( .A1(n5866), .A2(n7654), .B1(n7653), .B2(n6633), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U841 ( .A1(n7751), .A2(n7654), .B1(n7652), .B2(n6632), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U852 ( .A1(n7749), .A2(n7654), .B1(n7653), .B2(n6631), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U858 ( .A1(n7757), .A2(n7650), .B1(n7649), .B2(n6708), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U859 ( .A1(n5868), .A2(n7651), .B1(n7649), .B2(n6707), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U860 ( .A1(n7755), .A2(n7650), .B1(n7649), .B2(n6706), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U861 ( .A1(n5867), .A2(n7651), .B1(n7649), .B2(n6705), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U862 ( .A1(n7753), .A2(n7650), .B1(n7649), .B2(n6704), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U865 ( .A1(n5866), .A2(n7651), .B1(n7649), .B2(n6703), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U876 ( .A1(n7751), .A2(n7650), .B1(n7649), .B2(n6702), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U887 ( .A1(n7749), .A2(n7651), .B1(n7649), .B2(n6701), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U892 ( .A1(n7757), .A2(n7646), .B1(n7645), .B2(n6490), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U893 ( .A1(n5868), .A2(n7647), .B1(n7645), .B2(n6489), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U894 ( .A1(n7755), .A2(n7646), .B1(n7645), .B2(n6488), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U895 ( .A1(n5867), .A2(n7647), .B1(n7645), .B2(n6487), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U896 ( .A1(n7753), .A2(n7646), .B1(n7645), .B2(n6486), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U899 ( .A1(n5866), .A2(n7647), .B1(n7645), .B2(n6485), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U910 ( .A1(n7751), .A2(n7646), .B1(n7645), .B2(n6484), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U921 ( .A1(n7749), .A2(n7647), .B1(n7645), .B2(n6483), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U926 ( .A1(n7757), .A2(n7642), .B1(n7641), .B2(n6362), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U927 ( .A1(n5868), .A2(n7643), .B1(n7641), .B2(n6361), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U928 ( .A1(n7755), .A2(n7642), .B1(n7641), .B2(n6360), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U929 ( .A1(n5867), .A2(n7643), .B1(n7641), .B2(n6047), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U930 ( .A1(n7753), .A2(n7642), .B1(n7641), .B2(n6359), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U933 ( .A1(n5866), .A2(n7643), .B1(n7641), .B2(n6358), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U944 ( .A1(n7751), .A2(n7642), .B1(n7641), .B2(n5891), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U955 ( .A1(n7749), .A2(n7643), .B1(n7641), .B2(n5890), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U961 ( .A1(n7757), .A2(n7638), .B1(n7637), .B2(n6537), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U962 ( .A1(n5868), .A2(n7639), .B1(n7637), .B2(n6536), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U963 ( .A1(n7755), .A2(n7638), .B1(n7637), .B2(n6535), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U964 ( .A1(n5867), .A2(n7639), .B1(n7637), .B2(n6534), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U965 ( .A1(n7753), .A2(n7638), .B1(n7637), .B2(n6533), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U968 ( .A1(n5866), .A2(n7639), .B1(n7637), .B2(n6532), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U979 ( .A1(n7751), .A2(n7638), .B1(n7637), .B2(n6531), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U990 ( .A1(n7749), .A2(n7639), .B1(n7637), .B2(n6530), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  AND2_X2 U994 ( .A1(n7321), .A2(RegWrite_wb_out), .ZN(n3092) );
  OAI22_X2 U997 ( .A1(n7757), .A2(n3146), .B1(n7633), .B2(n6284), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U998 ( .A1(n5868), .A2(n7634), .B1(n7632), .B2(n6283), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U999 ( .A1(n7755), .A2(n3146), .B1(n7633), .B2(n6282), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1000 ( .A1(n5867), .A2(n3146), .B1(n7632), .B2(n6281), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1001 ( .A1(n7753), .A2(n3146), .B1(n7633), .B2(n6280), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1004 ( .A1(n5866), .A2(n3146), .B1(n7632), .B2(n6279), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1015 ( .A1(n7751), .A2(n3146), .B1(n7633), .B2(n6278), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1026 ( .A1(n7749), .A2(n3146), .B1(n7632), .B2(n6277), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  AND2_X2 U1029 ( .A1(n7310), .A2(n7335), .ZN(n3084) );
  OAI22_X2 U1032 ( .A1(n7757), .A2(n3148), .B1(n7629), .B2(n6150), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1033 ( .A1(n5868), .A2(n7630), .B1(n7628), .B2(n6149), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1034 ( .A1(n7755), .A2(n3148), .B1(n7629), .B2(n6148), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1035 ( .A1(n5867), .A2(n3148), .B1(n7628), .B2(n6147), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1036 ( .A1(n7753), .A2(n3148), .B1(n7629), .B2(n6146), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1039 ( .A1(n5866), .A2(n3148), .B1(n7628), .B2(n6145), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1050 ( .A1(n7751), .A2(n3148), .B1(n7629), .B2(n6144), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1061 ( .A1(n7749), .A2(n3148), .B1(n7628), .B2(n6143), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  AND2_X2 U1065 ( .A1(n7310), .A2(n7334), .ZN(n3087) );
  OAI22_X2 U1070 ( .A1(n7757), .A2(n7626), .B1(n7625), .B2(n6630), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1072 ( .A1(n5868), .A2(n7626), .B1(n7625), .B2(n6629), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1074 ( .A1(n7755), .A2(n7626), .B1(n7625), .B2(n6628), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1076 ( .A1(n5867), .A2(n7626), .B1(n7625), .B2(n6627), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1078 ( .A1(n7753), .A2(n7626), .B1(n7624), .B2(n6626), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1084 ( .A1(n5866), .A2(n7626), .B1(n7625), .B2(n6625), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1106 ( .A1(n7751), .A2(n7626), .B1(n7624), .B2(n6624), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1128 ( .A1(n7749), .A2(n7626), .B1(n7625), .B2(n6623), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI221_X2 U1135 ( .B1(n7622), .B2(n6907), .C1(n7619), .C2(n3170), .A(n3171), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1136 ( .A1(EXEC_MEM_OUT_118), .A2(n1541), .ZN(n3171) );
  OAI221_X2 U1137 ( .B1(n7621), .B2(n6888), .C1(n3169), .C2(n3172), .A(n3173), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1138 ( .A1(EXEC_MEM_OUT_117), .A2(n1541), .ZN(n3173) );
  OAI221_X2 U1139 ( .B1(n7621), .B2(n6902), .C1(n3169), .C2(n3174), .A(n3175), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1140 ( .A1(EXEC_MEM_OUT_116), .A2(n1541), .ZN(n3175) );
  OAI221_X2 U1141 ( .B1(n7621), .B2(n6015), .C1(n3169), .C2(n3176), .A(n3177), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1142 ( .A1(EXEC_MEM_OUT_115), .A2(n1541), .ZN(n3177) );
  OAI221_X2 U1143 ( .B1(n7621), .B2(n6906), .C1(n3169), .C2(n3178), .A(n3179), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1144 ( .A1(EXEC_MEM_OUT_114), .A2(n1541), .ZN(n3179) );
  OAI221_X2 U1145 ( .B1(n7621), .B2(n6887), .C1(n3169), .C2(n3180), .A(n3181), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1146 ( .A1(EXEC_MEM_OUT_113), .A2(n1541), .ZN(n3181) );
  OAI221_X2 U1147 ( .B1(n7621), .B2(n6901), .C1(n3169), .C2(n3182), .A(n3183), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1148 ( .A1(EXEC_MEM_OUT_112), .A2(n1541), .ZN(n3183) );
  OAI22_X2 U1149 ( .A1(n3184), .A2(n7283), .B1(n3185), .B2(n6477), .ZN(
        IF_STAGE_PC_REG_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1150 ( .A1(n3184), .A2(n7282), .B1(n3185), .B2(n6476), .ZN(
        IF_STAGE_PC_REG_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  AND2_X2 U1151 ( .A1(n3169), .A2(n7621), .ZN(n3185) );
  OAI221_X2 U1152 ( .B1(n7621), .B2(n6894), .C1(n7619), .C2(n3186), .A(n3187), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1153 ( .A1(EXEC_MEM_OUT_111), .A2(n1541), .ZN(n3187) );
  OAI221_X2 U1154 ( .B1(n7621), .B2(n6882), .C1(n3169), .C2(n3188), .A(n3189), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1155 ( .A1(EXEC_MEM_OUT_138), .A2(n1541), .ZN(n3189) );
  OAI221_X2 U1156 ( .B1(n7621), .B2(n6890), .C1(n3169), .C2(n3190), .A(n3191), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1157 ( .A1(EXEC_MEM_OUT_137), .A2(n1541), .ZN(n3191) );
  OAI221_X2 U1158 ( .B1(n7621), .B2(n6905), .C1(n3169), .C2(n3192), .A(n3193), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1159 ( .A1(EXEC_MEM_OUT_136), .A2(n1541), .ZN(n3193) );
  OAI221_X2 U1160 ( .B1(n7622), .B2(n2012), .C1(n7619), .C2(n3194), .A(n3195), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1161 ( .A1(EXEC_MEM_OUT_135), .A2(n1541), .ZN(n3195) );
  OAI221_X2 U1162 ( .B1(n7622), .B2(n6915), .C1(n7619), .C2(n3196), .A(n3197), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1163 ( .A1(EXEC_MEM_OUT_134), .A2(n1541), .ZN(n3197) );
  OAI221_X2 U1164 ( .B1(n7622), .B2(n6885), .C1(n7619), .C2(n3198), .A(n3199), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1165 ( .A1(EXEC_MEM_OUT_133), .A2(n1541), .ZN(n3199) );
  OAI221_X2 U1166 ( .B1(n7622), .B2(n6910), .C1(n7619), .C2(n3200), .A(n3201), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1167 ( .A1(EXEC_MEM_OUT_132), .A2(n1541), .ZN(n3201) );
  OAI221_X2 U1168 ( .B1(n7622), .B2(n2008), .C1(n7619), .C2(n3202), .A(n3203), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1169 ( .A1(EXEC_MEM_OUT_131), .A2(n1541), .ZN(n3203) );
  OAI221_X2 U1170 ( .B1(n7622), .B2(n6914), .C1(n7619), .C2(n3204), .A(n3205), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1171 ( .A1(EXEC_MEM_OUT_130), .A2(n1541), .ZN(n3205) );
  OAI221_X2 U1172 ( .B1(n7622), .B2(n6884), .C1(n7619), .C2(n3206), .A(n3207), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1173 ( .A1(EXEC_MEM_OUT_129), .A2(n1541), .ZN(n3207) );
  OAI221_X2 U1174 ( .B1(n7622), .B2(n6995), .C1(n7619), .C2(n3208), .A(n3209), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1175 ( .A1(EXEC_MEM_OUT_110), .A2(n1541), .ZN(n3209) );
  OAI221_X2 U1176 ( .B1(n7622), .B2(n6909), .C1(n7619), .C2(n3210), .A(n3211), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1177 ( .A1(EXEC_MEM_OUT_128), .A2(n1541), .ZN(n3211) );
  OAI221_X2 U1178 ( .B1(n7622), .B2(n6877), .C1(n7619), .C2(n3212), .A(n3213), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1179 ( .A1(EXEC_MEM_OUT_127), .A2(n1541), .ZN(n3213) );
  OAI221_X2 U1180 ( .B1(n7621), .B2(n6041), .C1(n7619), .C2(n3214), .A(n3215), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1181 ( .A1(EXEC_MEM_OUT_126), .A2(n1541), .ZN(n3215) );
  OAI221_X2 U1182 ( .B1(n7621), .B2(n6021), .C1(n7619), .C2(n3216), .A(n3217), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1183 ( .A1(EXEC_MEM_OUT_125), .A2(n1541), .ZN(n3217) );
  OAI221_X2 U1184 ( .B1(n7621), .B2(n6039), .C1(n7619), .C2(n3218), .A(n3219), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1185 ( .A1(EXEC_MEM_OUT_124), .A2(n1541), .ZN(n3219) );
  OAI221_X2 U1186 ( .B1(n7621), .B2(n5909), .C1(n7619), .C2(n3220), .A(n3221), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1187 ( .A1(EXEC_MEM_OUT_123), .A2(n1541), .ZN(n3221) );
  OAI221_X2 U1188 ( .B1(n7621), .B2(n6040), .C1(n7619), .C2(n3222), .A(n3223), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1189 ( .A1(EXEC_MEM_OUT_122), .A2(n1541), .ZN(n3223) );
  OAI221_X2 U1190 ( .B1(n7621), .B2(n6020), .C1(n7619), .C2(n3224), .A(n3225), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1191 ( .A1(EXEC_MEM_OUT_121), .A2(n1541), .ZN(n3225) );
  OAI221_X2 U1192 ( .B1(n7621), .B2(n6038), .C1(n7619), .C2(n3226), .A(n3227), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1193 ( .A1(EXEC_MEM_OUT_120), .A2(n1541), .ZN(n3227) );
  OAI221_X2 U1194 ( .B1(n7621), .B2(n1996), .C1(n7619), .C2(n3228), .A(n3229), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI221_X2 U1196 ( .B1(n7621), .B2(n7135), .C1(n3169), .C2(n3230), .A(n3231), 
        .ZN(IF_STAGE_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1197 ( .A1(EXEC_MEM_OUT_109), .A2(n1541), .ZN(n3231) );
  NAND2_X2 U1199 ( .A1(n7796), .A2(n7774), .ZN(n3169) );
  AND2_X2 U1201 ( .A1(IMEM_BUS_IN[25]), .A2(n7617), .ZN(IF_ID_REG_IF_ID_REG_N9) );
  AND2_X2 U1202 ( .A1(IMEM_BUS_IN[26]), .A2(n7617), .ZN(IF_ID_REG_IF_ID_REG_N8) );
  AND2_X2 U1203 ( .A1(IMEM_BUS_IN[27]), .A2(n7617), .ZN(IF_ID_REG_IF_ID_REG_N7) );
  NAND2_X2 U1204 ( .A1(n3233), .A2(n7616), .ZN(n3230) );
  XOR2_X2 U1205 ( .A(n7135), .B(n3234), .Z(n3233) );
  NAND2_X2 U1206 ( .A1(n3235), .A2(IMEM_BUS_OUT[1]), .ZN(n3234) );
  NAND2_X2 U1207 ( .A1(n3236), .A2(n7616), .ZN(n3208) );
  XOR2_X2 U1208 ( .A(IMEM_BUS_OUT[1]), .B(n3235), .Z(n3236) );
  NAND2_X2 U1210 ( .A1(n3238), .A2(n7616), .ZN(n3186) );
  XOR2_X2 U1211 ( .A(n6894), .B(n3237), .Z(n3238) );
  NAND2_X2 U1213 ( .A1(n3240), .A2(n7616), .ZN(n3182) );
  XOR2_X2 U1214 ( .A(n6901), .B(n3241), .Z(n3240) );
  NAND2_X2 U1215 ( .A1(n3239), .A2(IMEM_BUS_OUT[4]), .ZN(n3241) );
  NAND2_X2 U1216 ( .A1(n3242), .A2(n7616), .ZN(n3180) );
  XOR2_X2 U1217 ( .A(IMEM_BUS_OUT[4]), .B(n3239), .Z(n3242) );
  NAND2_X2 U1219 ( .A1(n3244), .A2(n7616), .ZN(n3178) );
  XOR2_X2 U1220 ( .A(IMEM_BUS_OUT[5]), .B(n3245), .Z(n3244) );
  NAND2_X2 U1222 ( .A1(n3246), .A2(n7616), .ZN(n3176) );
  XOR2_X2 U1223 ( .A(n6015), .B(n3243), .Z(n3246) );
  AND2_X2 U1225 ( .A1(IMEM_BUS_IN[28]), .A2(n7617), .ZN(IF_ID_REG_IF_ID_REG_N6) );
  NAND2_X2 U1226 ( .A1(n3248), .A2(n7616), .ZN(n3174) );
  XOR2_X2 U1227 ( .A(n6902), .B(n3249), .Z(n3248) );
  NAND2_X2 U1228 ( .A1(n3247), .A2(IMEM_BUS_OUT[8]), .ZN(n3249) );
  NAND2_X2 U1229 ( .A1(n3250), .A2(n7616), .ZN(n3172) );
  XOR2_X2 U1230 ( .A(IMEM_BUS_OUT[8]), .B(n3247), .Z(n3250) );
  NAND2_X2 U1232 ( .A1(n3252), .A2(n7616), .ZN(n3170) );
  XOR2_X2 U1233 ( .A(IMEM_BUS_OUT[9]), .B(n3253), .Z(n3252) );
  NAND2_X2 U1235 ( .A1(n3254), .A2(n7616), .ZN(n3228) );
  XOR2_X2 U1236 ( .A(n1996), .B(n3251), .Z(n3254) );
  NAND2_X2 U1238 ( .A1(n3256), .A2(n7616), .ZN(n3226) );
  XOR2_X2 U1239 ( .A(n6038), .B(n3257), .Z(n3256) );
  NAND2_X2 U1240 ( .A1(IMEM_BUS_OUT[12]), .A2(n3255), .ZN(n3257) );
  NAND2_X2 U1241 ( .A1(n3258), .A2(n7616), .ZN(n3224) );
  XOR2_X2 U1242 ( .A(IMEM_BUS_OUT[12]), .B(n3255), .Z(n3258) );
  NAND2_X2 U1244 ( .A1(n3260), .A2(n7616), .ZN(n3222) );
  XOR2_X2 U1245 ( .A(IMEM_BUS_OUT[13]), .B(n3261), .Z(n3260) );
  NAND2_X2 U1247 ( .A1(n3262), .A2(n7616), .ZN(n3220) );
  XOR2_X2 U1248 ( .A(n5909), .B(n3259), .Z(n3262) );
  NAND2_X2 U1250 ( .A1(n3264), .A2(n7616), .ZN(n3218) );
  XOR2_X2 U1251 ( .A(n6039), .B(n3265), .Z(n3264) );
  NAND2_X2 U1252 ( .A1(IMEM_BUS_OUT[16]), .A2(n3263), .ZN(n3265) );
  NAND2_X2 U1253 ( .A1(n3266), .A2(n7616), .ZN(n3216) );
  XOR2_X2 U1254 ( .A(IMEM_BUS_OUT[16]), .B(n3263), .Z(n3266) );
  AND2_X2 U1256 ( .A1(IMEM_BUS_IN[29]), .A2(n7617), .ZN(IF_ID_REG_IF_ID_REG_N5) );
  NAND2_X2 U1257 ( .A1(n3268), .A2(n7616), .ZN(n3214) );
  XOR2_X2 U1258 ( .A(IMEM_BUS_OUT[17]), .B(n3269), .Z(n3268) );
  NAND2_X2 U1260 ( .A1(n3270), .A2(n7616), .ZN(n3212) );
  XOR2_X2 U1261 ( .A(n6877), .B(n3267), .Z(n3270) );
  NAND2_X2 U1263 ( .A1(n3272), .A2(n7616), .ZN(n3210) );
  XOR2_X2 U1264 ( .A(n6909), .B(n3273), .Z(n3272) );
  NAND2_X2 U1265 ( .A1(IMEM_BUS_OUT[20]), .A2(n3271), .ZN(n3273) );
  NAND2_X2 U1266 ( .A1(n3274), .A2(n7616), .ZN(n3206) );
  XOR2_X2 U1267 ( .A(IMEM_BUS_OUT[20]), .B(n3271), .Z(n3274) );
  NAND2_X2 U1269 ( .A1(n3276), .A2(n7617), .ZN(n3204) );
  XOR2_X2 U1270 ( .A(IMEM_BUS_OUT[21]), .B(n3277), .Z(n3276) );
  NAND2_X2 U1272 ( .A1(n3278), .A2(n7617), .ZN(n3202) );
  XOR2_X2 U1273 ( .A(n2008), .B(n3275), .Z(n3278) );
  NAND2_X2 U1275 ( .A1(n3280), .A2(n7617), .ZN(n3200) );
  XOR2_X2 U1276 ( .A(n6910), .B(n3281), .Z(n3280) );
  NAND2_X2 U1277 ( .A1(IMEM_BUS_OUT[24]), .A2(n3279), .ZN(n3281) );
  NAND2_X2 U1278 ( .A1(n3282), .A2(n7617), .ZN(n3198) );
  XOR2_X2 U1279 ( .A(IMEM_BUS_OUT[24]), .B(n3279), .Z(n3282) );
  NAND2_X2 U1281 ( .A1(n3284), .A2(n7617), .ZN(n3196) );
  XOR2_X2 U1282 ( .A(IMEM_BUS_OUT[25]), .B(n3285), .Z(n3284) );
  NAND2_X2 U1284 ( .A1(n3286), .A2(n7617), .ZN(n3194) );
  XOR2_X2 U1285 ( .A(n2012), .B(n3283), .Z(n3286) );
  AND2_X2 U1287 ( .A1(IMEM_BUS_IN[30]), .A2(n7617), .ZN(IF_ID_REG_IF_ID_REG_N4) );
  NAND2_X2 U1288 ( .A1(n3287), .A2(n7617), .ZN(n3192) );
  XOR2_X2 U1289 ( .A(n6905), .B(n3288), .Z(n3287) );
  NAND2_X2 U1290 ( .A1(IMEM_BUS_OUT[29]), .A2(IMEM_BUS_OUT[28]), .ZN(n3288) );
  NAND2_X2 U1291 ( .A1(n3289), .A2(n7617), .ZN(n3190) );
  XOR2_X2 U1292 ( .A(IMEM_BUS_OUT[29]), .B(IMEM_BUS_OUT[28]), .Z(n3289) );
  NAND2_X2 U1293 ( .A1(n7616), .A2(n6882), .ZN(n3188) );
  AND2_X2 U1297 ( .A1(n7617), .A2(IMEM_BUS_IN[1]), .ZN(IF_ID_REG_IF_ID_REG_N33) );
  AND2_X2 U1299 ( .A1(n7617), .A2(IMEM_BUS_IN[3]), .ZN(IF_ID_REG_IF_ID_REG_N31) );
  AND2_X2 U1300 ( .A1(n7617), .A2(IMEM_BUS_IN[4]), .ZN(IF_ID_REG_IF_ID_REG_N30) );
  AND2_X2 U1301 ( .A1(IMEM_BUS_IN[31]), .A2(n7617), .ZN(IF_ID_REG_IF_ID_REG_N3) );
  AND2_X2 U1303 ( .A1(n7617), .A2(IMEM_BUS_IN[6]), .ZN(IF_ID_REG_IF_ID_REG_N28) );
  AND2_X2 U1304 ( .A1(n7617), .A2(IMEM_BUS_IN[7]), .ZN(IF_ID_REG_IF_ID_REG_N27) );
  AND2_X2 U1305 ( .A1(n7617), .A2(IMEM_BUS_IN[8]), .ZN(IF_ID_REG_IF_ID_REG_N26) );
  AND2_X2 U1306 ( .A1(n7617), .A2(IMEM_BUS_IN[9]), .ZN(IF_ID_REG_IF_ID_REG_N25) );
  AND2_X2 U1307 ( .A1(n7617), .A2(IMEM_BUS_IN[10]), .ZN(
        IF_ID_REG_IF_ID_REG_N24) );
  AND2_X2 U1308 ( .A1(n7617), .A2(IMEM_BUS_IN[11]), .ZN(
        IF_ID_REG_IF_ID_REG_N23) );
  AND2_X2 U1309 ( .A1(n7617), .A2(IMEM_BUS_IN[12]), .ZN(
        IF_ID_REG_IF_ID_REG_N22) );
  AND2_X2 U1310 ( .A1(n7617), .A2(IMEM_BUS_IN[13]), .ZN(
        IF_ID_REG_IF_ID_REG_N21) );
  AND2_X2 U1311 ( .A1(n7617), .A2(IMEM_BUS_IN[14]), .ZN(
        IF_ID_REG_IF_ID_REG_N20) );
  AND2_X2 U1312 ( .A1(n7617), .A2(IMEM_BUS_IN[15]), .ZN(
        IF_ID_REG_IF_ID_REG_N19) );
  AND2_X2 U1313 ( .A1(IMEM_BUS_IN[16]), .A2(n7617), .ZN(
        IF_ID_REG_IF_ID_REG_N18) );
  AND2_X2 U1314 ( .A1(IMEM_BUS_IN[17]), .A2(n7617), .ZN(
        IF_ID_REG_IF_ID_REG_N17) );
  AND2_X2 U1315 ( .A1(IMEM_BUS_IN[18]), .A2(n7617), .ZN(
        IF_ID_REG_IF_ID_REG_N16) );
  AND2_X2 U1316 ( .A1(IMEM_BUS_IN[19]), .A2(n7617), .ZN(
        IF_ID_REG_IF_ID_REG_N15) );
  AND2_X2 U1317 ( .A1(IMEM_BUS_IN[20]), .A2(n7617), .ZN(
        IF_ID_REG_IF_ID_REG_N14) );
  AND2_X2 U1318 ( .A1(IMEM_BUS_IN[21]), .A2(n7617), .ZN(
        IF_ID_REG_IF_ID_REG_N13) );
  AND2_X2 U1319 ( .A1(IMEM_BUS_IN[22]), .A2(n7617), .ZN(
        IF_ID_REG_IF_ID_REG_N12) );
  AND2_X2 U1320 ( .A1(IMEM_BUS_IN[23]), .A2(n7617), .ZN(
        IF_ID_REG_IF_ID_REG_N11) );
  AND2_X2 U1321 ( .A1(IMEM_BUS_IN[24]), .A2(n7617), .ZN(
        IF_ID_REG_IF_ID_REG_N10) );
  NAND4_X2 U1323 ( .A1(IMEM_BUS_IN[4]), .A2(n3294), .A3(n1574), .A4(n1575), 
        .ZN(n3293) );
  XNOR2_X2 U1325 ( .A(n5848), .B(IMEM_BUS_IN[8]), .ZN(n3298) );
  XNOR2_X2 U1326 ( .A(n3300), .B(IMEM_BUS_IN[6]), .ZN(n3297) );
  XNOR2_X2 U1327 ( .A(n3301), .B(IMEM_BUS_IN[7]), .ZN(n3296) );
  XNOR2_X2 U1332 ( .A(n5848), .B(IMEM_BUS_IN[13]), .ZN(n3310) );
  XNOR2_X2 U1333 ( .A(n3300), .B(IMEM_BUS_IN[11]), .ZN(n3309) );
  XNOR2_X2 U1334 ( .A(n3301), .B(IMEM_BUS_IN[12]), .ZN(n3308) );
  OAI211_X2 U1335 ( .C1(n3311), .C2(n1573), .A(n3312), .B(n3313), .ZN(n3307)
         );
  NAND4_X2 U1338 ( .A1(IMEM_BUS_IN[2]), .A2(IMEM_BUS_IN[0]), .A3(n3294), .A4(
        n3314), .ZN(n3303) );
  NAND2_X2 U1339 ( .A1(IMEM_BUS_IN[4]), .A2(n1576), .ZN(n3314) );
  AND4_X2 U1340 ( .A1(n1576), .A2(n1575), .A3(n1574), .A4(n3294), .ZN(n3311)
         );
  AOI221_X2 U1346 ( .B1(n5850), .B2(offset_26_id[5]), .C1(n1591), .C2(
        ID_STAGE_imm16_aluA[16]), .A(n3316), .ZN(n3300) );
  AOI221_X2 U1348 ( .B1(n5850), .B2(offset_26_id[6]), .C1(n1591), .C2(
        ID_STAGE_imm16_aluA[17]), .A(n3316), .ZN(n3301) );
  AOI221_X2 U1350 ( .B1(n5850), .B2(offset_26_id[7]), .C1(n1591), .C2(
        ID_STAGE_imm16_aluA[18]), .A(n3316), .ZN(n3299) );
  AOI221_X2 U1352 ( .B1(n5850), .B2(offset_26_id[8]), .C1(n1591), .C2(
        ID_STAGE_imm16_aluA[19]), .A(n3316), .ZN(n3306) );
  NAND2_X2 U1358 ( .A1(n3318), .A2(n7305), .ZN(n3317) );
  NOR4_X2 U1359 ( .A1(n3318), .A2(n3319), .A3(n3320), .A4(n3321), .ZN(
        ID_EX_REG_ID_EX_REG_N57) );
  AND2_X2 U1361 ( .A1(n3316), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N63) );
  AND2_X2 U1363 ( .A1(n3323), .A2(n3324), .ZN(n3318) );
  AND2_X2 U1364 ( .A1(n7305), .A2(n3292), .ZN(ID_EX_REG_ID_EX_REG_N56) );
  AND2_X2 U1367 ( .A1(n7305), .A2(n3319), .ZN(ID_EX_REG_ID_EX_REG_N55) );
  NOR4_X2 U1369 ( .A1(IF_ID_OUT[35]), .A2(EXEC_MEM_OUT_141), .A3(n6865), .A4(
        n1592), .ZN(ID_EX_REG_ID_EX_REG_N54) );
  NOR4_X2 U1370 ( .A1(n3327), .A2(n3328), .A3(n1592), .A4(n6011), .ZN(
        ID_EX_REG_ID_EX_REG_N53) );
  NAND4_X2 U1371 ( .A1(n3329), .A2(n3330), .A3(IF_ID_OUT[37]), .A4(n6012), 
        .ZN(n3327) );
  XOR2_X2 U1372 ( .A(ID_STAGE_imm16_aluA[28]), .B(ID_STAGE_imm16_aluA[27]), 
        .Z(n3330) );
  NOR4_X2 U1373 ( .A1(EXEC_MEM_OUT_141), .A2(n6346), .A3(n3326), .A4(n6864), 
        .ZN(ID_EX_REG_ID_EX_REG_N52) );
  NOR4_X2 U1375 ( .A1(EXEC_MEM_OUT_141), .A2(n3331), .A3(n6346), .A4(n6865), 
        .ZN(ID_EX_REG_ID_EX_REG_N51) );
  NOR4_X2 U1378 ( .A1(n3333), .A2(n3334), .A3(n3335), .A4(n3336), .ZN(n3332)
         );
  NOR4_X2 U1381 ( .A1(n3333), .A2(n3338), .A3(n3339), .A4(n3340), .ZN(n3337)
         );
  OR4_X2 U1384 ( .A1(n3343), .A2(n3344), .A3(n3345), .A4(n3346), .ZN(n3333) );
  AOI221_X2 U1386 ( .B1(n3350), .B2(n1589), .C1(n1660), .C2(n1654), .A(n3343), 
        .ZN(n3349) );
  OAI22_X2 U1391 ( .A1(n3357), .A2(n3353), .B1(n3358), .B2(n3359), .ZN(n3335)
         );
  NAND2_X2 U1392 ( .A1(ID_STAGE_imm16_aluA[30]), .A2(n1594), .ZN(n3359) );
  NOR4_X2 U1394 ( .A1(n3361), .A2(n3356), .A3(n3336), .A4(n3340), .ZN(n3360)
         );
  NAND2_X2 U1395 ( .A1(IF_ID_OUT[37]), .A2(n6864), .ZN(n3362) );
  OAI221_X2 U1396 ( .B1(n3364), .B2(n3357), .C1(n6864), .C2(n3351), .A(n3365), 
        .ZN(n3336) );
  OR3_X2 U1397 ( .A1(n3366), .A2(ID_STAGE_imm16_aluA[30]), .A3(n3358), .ZN(
        n3365) );
  OR4_X2 U1398 ( .A1(n3339), .A2(n3334), .A3(n3367), .A4(n3345), .ZN(n3356) );
  NAND2_X2 U1401 ( .A1(IF_ID_OUT[36]), .A2(n6346), .ZN(n3353) );
  OR3_X2 U1403 ( .A1(n3363), .A2(n3364), .A3(n6343), .ZN(n3371) );
  NAND2_X2 U1409 ( .A1(ID_STAGE_imm16_aluA[30]), .A2(n3375), .ZN(n3374) );
  OAI211_X2 U1411 ( .C1(ID_STAGE_imm16_aluA[28]), .C2(n3355), .A(n3376), .B(
        n1577), .ZN(n3361) );
  OAI22_X2 U1412 ( .A1(n3364), .A2(n3368), .B1(ID_STAGE_imm16_aluA[31]), .B2(
        n3370), .ZN(n3344) );
  AND3_X2 U1416 ( .A1(n1591), .A2(n6898), .A3(ID_STAGE_imm16_aluA[26]), .ZN(
        n3373) );
  AND2_X2 U1445 ( .A1(IF_ID_OUT[0]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N206)
         );
  AND2_X2 U1446 ( .A1(IF_ID_OUT[1]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N205)
         );
  AND2_X2 U1447 ( .A1(IF_ID_OUT[2]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N204)
         );
  AND2_X2 U1448 ( .A1(IF_ID_OUT[3]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N203)
         );
  AND2_X2 U1449 ( .A1(IF_ID_OUT[4]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N202)
         );
  AND2_X2 U1450 ( .A1(IF_ID_OUT[5]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N201)
         );
  AND2_X2 U1451 ( .A1(IF_ID_OUT[6]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N200)
         );
  AND2_X2 U1453 ( .A1(IF_ID_OUT[7]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N199)
         );
  AND2_X2 U1454 ( .A1(IF_ID_OUT[8]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N198)
         );
  AND2_X2 U1455 ( .A1(IF_ID_OUT[9]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N197)
         );
  AND2_X2 U1456 ( .A1(IF_ID_OUT[10]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N196) );
  AND2_X2 U1457 ( .A1(IF_ID_OUT[11]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N195) );
  AND2_X2 U1458 ( .A1(IF_ID_OUT[12]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N194) );
  AND2_X2 U1459 ( .A1(IF_ID_OUT[13]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N193) );
  AND2_X2 U1460 ( .A1(IF_ID_OUT[14]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N192) );
  AND2_X2 U1461 ( .A1(IF_ID_OUT[15]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N191) );
  AND2_X2 U1462 ( .A1(IF_ID_OUT[16]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N190) );
  AND2_X2 U1464 ( .A1(IF_ID_OUT[17]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N189) );
  AND2_X2 U1465 ( .A1(IF_ID_OUT[18]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N188) );
  AND2_X2 U1466 ( .A1(IF_ID_OUT[19]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N187) );
  AND2_X2 U1467 ( .A1(IF_ID_OUT[20]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N186) );
  AND2_X2 U1468 ( .A1(IF_ID_OUT[21]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N185) );
  AND2_X2 U1469 ( .A1(IF_ID_OUT[22]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N184) );
  AND2_X2 U1470 ( .A1(IF_ID_OUT[23]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N183) );
  AND2_X2 U1471 ( .A1(IF_ID_OUT[24]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N182) );
  AND2_X2 U1472 ( .A1(IF_ID_OUT[25]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N181) );
  AND2_X2 U1473 ( .A1(IF_ID_OUT[26]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N180) );
  AND2_X2 U1475 ( .A1(IF_ID_OUT[27]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N179) );
  AND2_X2 U1476 ( .A1(IF_ID_OUT[28]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N178) );
  AND2_X2 U1477 ( .A1(IF_ID_OUT[29]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N177) );
  AND2_X2 U1478 ( .A1(IF_ID_OUT[30]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N176) );
  AND2_X2 U1479 ( .A1(IF_ID_OUT[31]), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N175) );
  NAND4_X2 U1480 ( .A1(n3385), .A2(n3386), .A3(n3387), .A4(n3388), .ZN(
        ID_EX_REG_ID_EX_REG_N174) );
  AOI221_X2 U1483 ( .B1(n7606), .B2(REG_FILE_reg_out_3__0_), .C1(n7599), .C2(
        REG_FILE_reg_out_7__0_), .A(n3397), .ZN(n3394) );
  OAI22_X2 U1484 ( .A1(n5897), .A2(n7592), .B1(n5954), .B2(n7588), .ZN(n3397)
         );
  AOI22_X2 U1485 ( .A1(n7573), .A2(REG_FILE_reg_out_2__0_), .B1(n7566), .B2(
        REG_FILE_reg_out_6__0_), .ZN(n3393) );
  AOI22_X2 U1486 ( .A1(n7769), .A2(REG_FILE_reg_out_0__0_), .B1(n7576), .B2(
        REG_FILE_reg_out_4__0_), .ZN(n3392) );
  OAI221_X2 U1488 ( .B1(n6143), .B2(n7570), .C1(n6483), .C2(n7564), .A(n3407), 
        .ZN(n3403) );
  AOI22_X2 U1489 ( .A1(n7763), .A2(REG_FILE_reg_out_8__0_), .B1(n7576), .B2(
        REG_FILE_reg_out_12__0_), .ZN(n3407) );
  OAI221_X2 U1490 ( .B1(n6101), .B2(n7587), .C1(n5890), .C2(n7597), .A(n3408), 
        .ZN(n3402) );
  AOI22_X2 U1491 ( .A1(n7607), .A2(REG_FILE_reg_out_11__0_), .B1(n7600), .B2(
        REG_FILE_reg_out_15__0_), .ZN(n3408) );
  OAI221_X2 U1493 ( .B1(n5955), .B2(n7571), .C1(n6151), .C2(n7564), .A(n3412), 
        .ZN(n3410) );
  AOI22_X2 U1494 ( .A1(n7769), .A2(REG_FILE_reg_out_24__0_), .B1(n7576), .B2(
        REG_FILE_reg_out_28__0_), .ZN(n3412) );
  OAI221_X2 U1495 ( .B1(n5945), .B2(n7587), .C1(n5893), .C2(n7595), .A(n3413), 
        .ZN(n3409) );
  AOI22_X2 U1496 ( .A1(n7606), .A2(REG_FILE_reg_out_27__0_), .B1(n7600), .B2(
        REG_FILE_reg_out_31__0_), .ZN(n3413) );
  OAI221_X2 U1498 ( .B1(n6086), .B2(n7570), .C1(n6363), .C2(n7564), .A(n3417), 
        .ZN(n3415) );
  AOI22_X2 U1499 ( .A1(n7769), .A2(REG_FILE_reg_out_16__0_), .B1(n7576), .B2(
        REG_FILE_reg_out_20__0_), .ZN(n3417) );
  OAI221_X2 U1500 ( .B1(n5944), .B2(n7587), .C1(n5892), .C2(n7595), .A(n3418), 
        .ZN(n3414) );
  AOI22_X2 U1501 ( .A1(n7608), .A2(REG_FILE_reg_out_19__0_), .B1(n7600), .B2(
        REG_FILE_reg_out_23__0_), .ZN(n3418) );
  NAND4_X2 U1502 ( .A1(n3419), .A2(n3420), .A3(n3421), .A4(n3422), .ZN(
        ID_EX_REG_ID_EX_REG_N173) );
  AOI221_X2 U1505 ( .B1(n7611), .B2(REG_FILE_reg_out_3__1_), .C1(n7604), .C2(
        REG_FILE_reg_out_7__1_), .A(n3427), .ZN(n3426) );
  OAI22_X2 U1506 ( .A1(n5880), .A2(n7593), .B1(n6128), .B2(n7588), .ZN(n3427)
         );
  AOI22_X2 U1507 ( .A1(n7573), .A2(REG_FILE_reg_out_2__1_), .B1(n7566), .B2(
        REG_FILE_reg_out_6__1_), .ZN(n3425) );
  AOI22_X2 U1508 ( .A1(n7770), .A2(REG_FILE_reg_out_0__1_), .B1(n7576), .B2(
        REG_FILE_reg_out_4__1_), .ZN(n3424) );
  OAI221_X2 U1510 ( .B1(n6144), .B2(n7571), .C1(n6484), .C2(n7564), .A(n3431), 
        .ZN(n3430) );
  AOI22_X2 U1511 ( .A1(n7763), .A2(REG_FILE_reg_out_8__1_), .B1(n7576), .B2(
        REG_FILE_reg_out_12__1_), .ZN(n3431) );
  OAI221_X2 U1512 ( .B1(n6102), .B2(n7587), .C1(n5891), .C2(n7597), .A(n3432), 
        .ZN(n3429) );
  AOI22_X2 U1513 ( .A1(n7606), .A2(REG_FILE_reg_out_11__1_), .B1(n7600), .B2(
        REG_FILE_reg_out_15__1_), .ZN(n3432) );
  OAI221_X2 U1515 ( .B1(n5956), .B2(n7570), .C1(n6152), .C2(n7564), .A(n3435), 
        .ZN(n3434) );
  AOI22_X2 U1516 ( .A1(n7770), .A2(REG_FILE_reg_out_24__1_), .B1(n7576), .B2(
        REG_FILE_reg_out_28__1_), .ZN(n3435) );
  OAI221_X2 U1517 ( .B1(n6094), .B2(n7587), .C1(n5927), .C2(n7597), .A(n3436), 
        .ZN(n3433) );
  AOI22_X2 U1518 ( .A1(n7607), .A2(REG_FILE_reg_out_27__1_), .B1(n7600), .B2(
        REG_FILE_reg_out_31__1_), .ZN(n3436) );
  OAI221_X2 U1520 ( .B1(n6087), .B2(n7571), .C1(n6364), .C2(n7564), .A(n3439), 
        .ZN(n3438) );
  AOI22_X2 U1521 ( .A1(n7770), .A2(REG_FILE_reg_out_16__1_), .B1(n7578), .B2(
        REG_FILE_reg_out_20__1_), .ZN(n3439) );
  OAI221_X2 U1522 ( .B1(n6399), .B2(n7587), .C1(n6048), .C2(n7597), .A(n3440), 
        .ZN(n3437) );
  AOI22_X2 U1523 ( .A1(n7608), .A2(REG_FILE_reg_out_19__1_), .B1(n7600), .B2(
        REG_FILE_reg_out_23__1_), .ZN(n3440) );
  NAND4_X2 U1524 ( .A1(n3441), .A2(n3442), .A3(n3443), .A4(n3444), .ZN(
        ID_EX_REG_ID_EX_REG_N172) );
  AOI221_X2 U1527 ( .B1(n7610), .B2(REG_FILE_reg_out_3__2_), .C1(n7604), .C2(
        REG_FILE_reg_out_7__2_), .A(n3449), .ZN(n3448) );
  OAI22_X2 U1528 ( .A1(n6113), .A2(n7598), .B1(n6462), .B2(n7588), .ZN(n3449)
         );
  AOI22_X2 U1529 ( .A1(n7573), .A2(REG_FILE_reg_out_2__2_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__2_), .ZN(n3447) );
  AOI22_X2 U1530 ( .A1(n7770), .A2(REG_FILE_reg_out_0__2_), .B1(n7578), .B2(
        REG_FILE_reg_out_4__2_), .ZN(n3446) );
  OAI221_X2 U1532 ( .B1(n6145), .B2(n7570), .C1(n6485), .C2(n7564), .A(n3452), 
        .ZN(n3451) );
  AOI22_X2 U1533 ( .A1(n7770), .A2(REG_FILE_reg_out_8__2_), .B1(n7577), .B2(
        REG_FILE_reg_out_12__2_), .ZN(n3452) );
  OAI221_X2 U1534 ( .B1(n6946), .B2(n7585), .C1(n6358), .C2(n7596), .A(n3453), 
        .ZN(n3450) );
  AOI22_X2 U1535 ( .A1(n7607), .A2(REG_FILE_reg_out_11__2_), .B1(n7600), .B2(
        REG_FILE_reg_out_15__2_), .ZN(n3453) );
  OAI221_X2 U1537 ( .B1(n5957), .B2(n7571), .C1(n6153), .C2(n7564), .A(n3456), 
        .ZN(n3455) );
  AOI22_X2 U1538 ( .A1(n7770), .A2(REG_FILE_reg_out_24__2_), .B1(n7578), .B2(
        REG_FILE_reg_out_28__2_), .ZN(n3456) );
  OAI221_X2 U1539 ( .B1(n6095), .B2(n7585), .C1(n5894), .C2(n7596), .A(n3457), 
        .ZN(n3454) );
  AOI22_X2 U1540 ( .A1(n7607), .A2(REG_FILE_reg_out_27__2_), .B1(n7601), .B2(
        REG_FILE_reg_out_31__2_), .ZN(n3457) );
  OAI221_X2 U1542 ( .B1(n6088), .B2(n7571), .C1(n6365), .C2(n7564), .A(n3460), 
        .ZN(n3459) );
  AOI22_X2 U1543 ( .A1(n7770), .A2(REG_FILE_reg_out_16__2_), .B1(n7577), .B2(
        REG_FILE_reg_out_20__2_), .ZN(n3460) );
  OAI221_X2 U1544 ( .B1(n6400), .B2(n7586), .C1(n6049), .C2(n7595), .A(n3461), 
        .ZN(n3458) );
  AOI22_X2 U1545 ( .A1(n7607), .A2(REG_FILE_reg_out_19__2_), .B1(n7600), .B2(
        REG_FILE_reg_out_23__2_), .ZN(n3461) );
  NAND4_X2 U1546 ( .A1(n3462), .A2(n3463), .A3(n3464), .A4(n3465), .ZN(
        ID_EX_REG_ID_EX_REG_N171) );
  AOI221_X2 U1549 ( .B1(n7611), .B2(REG_FILE_reg_out_3__3_), .C1(n7604), .C2(
        REG_FILE_reg_out_7__3_), .A(n3470), .ZN(n3469) );
  OAI22_X2 U1550 ( .A1(n6114), .A2(n7598), .B1(n6463), .B2(n7588), .ZN(n3470)
         );
  AOI22_X2 U1551 ( .A1(n7573), .A2(REG_FILE_reg_out_2__3_), .B1(n7566), .B2(
        REG_FILE_reg_out_6__3_), .ZN(n3468) );
  AOI22_X2 U1552 ( .A1(n7770), .A2(REG_FILE_reg_out_0__3_), .B1(n7577), .B2(
        REG_FILE_reg_out_4__3_), .ZN(n3467) );
  OAI221_X2 U1554 ( .B1(n6146), .B2(n7571), .C1(n6486), .C2(n7564), .A(n3474), 
        .ZN(n3473) );
  AOI22_X2 U1555 ( .A1(n7770), .A2(REG_FILE_reg_out_8__3_), .B1(n7578), .B2(
        REG_FILE_reg_out_12__3_), .ZN(n3474) );
  OAI221_X2 U1556 ( .B1(n6947), .B2(n7586), .C1(n6359), .C2(n7595), .A(n3475), 
        .ZN(n3472) );
  AOI22_X2 U1557 ( .A1(n7607), .A2(REG_FILE_reg_out_11__3_), .B1(n7600), .B2(
        REG_FILE_reg_out_15__3_), .ZN(n3475) );
  OAI221_X2 U1559 ( .B1(n5958), .B2(n7571), .C1(n6154), .C2(n7563), .A(n3478), 
        .ZN(n3477) );
  AOI22_X2 U1560 ( .A1(n7770), .A2(REG_FILE_reg_out_24__3_), .B1(n7577), .B2(
        REG_FILE_reg_out_28__3_), .ZN(n3478) );
  OAI221_X2 U1561 ( .B1(n6096), .B2(n7585), .C1(n5928), .C2(n7594), .A(n3479), 
        .ZN(n3476) );
  AOI22_X2 U1562 ( .A1(n7607), .A2(REG_FILE_reg_out_27__3_), .B1(n7601), .B2(
        REG_FILE_reg_out_31__3_), .ZN(n3479) );
  OAI221_X2 U1564 ( .B1(n6089), .B2(n7571), .C1(n6366), .C2(n7563), .A(n3482), 
        .ZN(n3481) );
  AOI22_X2 U1565 ( .A1(n7770), .A2(REG_FILE_reg_out_16__3_), .B1(n7578), .B2(
        REG_FILE_reg_out_20__3_), .ZN(n3482) );
  OAI221_X2 U1566 ( .B1(n6401), .B2(n7585), .C1(n6050), .C2(n7594), .A(n3483), 
        .ZN(n3480) );
  AOI22_X2 U1567 ( .A1(n7608), .A2(REG_FILE_reg_out_19__3_), .B1(n7600), .B2(
        REG_FILE_reg_out_23__3_), .ZN(n3483) );
  NAND4_X2 U1568 ( .A1(n3484), .A2(n3485), .A3(n3486), .A4(n3487), .ZN(
        ID_EX_REG_ID_EX_REG_N170) );
  AOI221_X2 U1571 ( .B1(n7610), .B2(REG_FILE_reg_out_3__4_), .C1(n7604), .C2(
        REG_FILE_reg_out_7__4_), .A(n3492), .ZN(n3491) );
  OAI22_X2 U1572 ( .A1(n6115), .A2(n7598), .B1(n6464), .B2(n7588), .ZN(n3492)
         );
  AOI22_X2 U1573 ( .A1(n7573), .A2(REG_FILE_reg_out_2__4_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__4_), .ZN(n3490) );
  AOI22_X2 U1574 ( .A1(n7770), .A2(REG_FILE_reg_out_0__4_), .B1(n7578), .B2(
        REG_FILE_reg_out_4__4_), .ZN(n3489) );
  OAI221_X2 U1576 ( .B1(n6147), .B2(n7571), .C1(n6487), .C2(n7564), .A(n3495), 
        .ZN(n3494) );
  AOI22_X2 U1577 ( .A1(n7770), .A2(REG_FILE_reg_out_8__4_), .B1(n7577), .B2(
        REG_FILE_reg_out_12__4_), .ZN(n3495) );
  OAI221_X2 U1578 ( .B1(n6405), .B2(n7583), .C1(n6047), .C2(n7594), .A(n3496), 
        .ZN(n3493) );
  AOI22_X2 U1579 ( .A1(n7607), .A2(REG_FILE_reg_out_11__4_), .B1(n7601), .B2(
        REG_FILE_reg_out_15__4_), .ZN(n3496) );
  OAI221_X2 U1581 ( .B1(n5959), .B2(n7571), .C1(n6155), .C2(n7564), .A(n3499), 
        .ZN(n3498) );
  AOI22_X2 U1582 ( .A1(n7769), .A2(REG_FILE_reg_out_24__4_), .B1(n7576), .B2(
        REG_FILE_reg_out_28__4_), .ZN(n3499) );
  OAI221_X2 U1583 ( .B1(n6097), .B2(n7583), .C1(n5929), .C2(n7595), .A(n3500), 
        .ZN(n3497) );
  AOI22_X2 U1584 ( .A1(n7607), .A2(REG_FILE_reg_out_27__4_), .B1(n7601), .B2(
        REG_FILE_reg_out_31__4_), .ZN(n3500) );
  OAI221_X2 U1586 ( .B1(n6090), .B2(n7571), .C1(n6367), .C2(n7564), .A(n3503), 
        .ZN(n3502) );
  AOI22_X2 U1587 ( .A1(n7769), .A2(REG_FILE_reg_out_16__4_), .B1(n7576), .B2(
        REG_FILE_reg_out_20__4_), .ZN(n3503) );
  OAI221_X2 U1588 ( .B1(n6402), .B2(n7584), .C1(n6051), .C2(n7593), .A(n3504), 
        .ZN(n3501) );
  AOI22_X2 U1589 ( .A1(n7607), .A2(REG_FILE_reg_out_19__4_), .B1(n7601), .B2(
        REG_FILE_reg_out_23__4_), .ZN(n3504) );
  NAND4_X2 U1591 ( .A1(n3505), .A2(n3506), .A3(n3507), .A4(n3508), .ZN(
        ID_EX_REG_ID_EX_REG_N169) );
  AOI221_X2 U1594 ( .B1(n7611), .B2(REG_FILE_reg_out_3__5_), .C1(n7604), .C2(
        REG_FILE_reg_out_7__5_), .A(n3513), .ZN(n3512) );
  OAI22_X2 U1595 ( .A1(n6116), .A2(n7598), .B1(n6465), .B2(n7588), .ZN(n3513)
         );
  AOI22_X2 U1596 ( .A1(n7573), .A2(REG_FILE_reg_out_2__5_), .B1(n7566), .B2(
        REG_FILE_reg_out_6__5_), .ZN(n3511) );
  AOI22_X2 U1597 ( .A1(n7769), .A2(REG_FILE_reg_out_0__5_), .B1(n7576), .B2(
        REG_FILE_reg_out_4__5_), .ZN(n3510) );
  OAI221_X2 U1599 ( .B1(n6148), .B2(n7571), .C1(n6488), .C2(n7564), .A(n3517), 
        .ZN(n3516) );
  AOI22_X2 U1600 ( .A1(n7769), .A2(REG_FILE_reg_out_8__5_), .B1(n7576), .B2(
        REG_FILE_reg_out_12__5_), .ZN(n3517) );
  OAI221_X2 U1601 ( .B1(n6948), .B2(n7584), .C1(n6360), .C2(n7593), .A(n3518), 
        .ZN(n3515) );
  AOI22_X2 U1602 ( .A1(n7607), .A2(REG_FILE_reg_out_11__5_), .B1(n7601), .B2(
        REG_FILE_reg_out_15__5_), .ZN(n3518) );
  OAI221_X2 U1604 ( .B1(n5960), .B2(n7571), .C1(n6156), .C2(n7563), .A(n3521), 
        .ZN(n3520) );
  AOI22_X2 U1605 ( .A1(n7769), .A2(REG_FILE_reg_out_24__5_), .B1(n7576), .B2(
        REG_FILE_reg_out_28__5_), .ZN(n3521) );
  OAI221_X2 U1606 ( .B1(n6098), .B2(n7584), .C1(n5930), .C2(n7592), .A(n3522), 
        .ZN(n3519) );
  AOI22_X2 U1607 ( .A1(n7607), .A2(REG_FILE_reg_out_27__5_), .B1(n7601), .B2(
        REG_FILE_reg_out_31__5_), .ZN(n3522) );
  OAI221_X2 U1609 ( .B1(n6091), .B2(n7571), .C1(n6368), .C2(n7563), .A(n3525), 
        .ZN(n3524) );
  AOI22_X2 U1610 ( .A1(n7769), .A2(REG_FILE_reg_out_16__5_), .B1(n7576), .B2(
        REG_FILE_reg_out_20__5_), .ZN(n3525) );
  OAI221_X2 U1611 ( .B1(n6403), .B2(n7584), .C1(n6052), .C2(n7592), .A(n3526), 
        .ZN(n3523) );
  AOI22_X2 U1612 ( .A1(n7607), .A2(REG_FILE_reg_out_19__5_), .B1(n7601), .B2(
        REG_FILE_reg_out_23__5_), .ZN(n3526) );
  NAND4_X2 U1613 ( .A1(n3527), .A2(n3528), .A3(n3529), .A4(n3530), .ZN(
        ID_EX_REG_ID_EX_REG_N168) );
  AOI221_X2 U1616 ( .B1(n7610), .B2(REG_FILE_reg_out_3__6_), .C1(n7604), .C2(
        REG_FILE_reg_out_7__6_), .A(n3535), .ZN(n3534) );
  OAI22_X2 U1617 ( .A1(n6117), .A2(n7593), .B1(n6466), .B2(n7588), .ZN(n3535)
         );
  AOI22_X2 U1618 ( .A1(n7573), .A2(REG_FILE_reg_out_2__6_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__6_), .ZN(n3533) );
  AOI22_X2 U1619 ( .A1(n7769), .A2(REG_FILE_reg_out_0__6_), .B1(n7576), .B2(
        REG_FILE_reg_out_4__6_), .ZN(n3532) );
  OAI221_X2 U1621 ( .B1(n6149), .B2(n7571), .C1(n6489), .C2(n7564), .A(n3538), 
        .ZN(n3537) );
  AOI22_X2 U1622 ( .A1(n7769), .A2(REG_FILE_reg_out_8__6_), .B1(n7576), .B2(
        REG_FILE_reg_out_12__6_), .ZN(n3538) );
  OAI221_X2 U1623 ( .B1(n6949), .B2(n7586), .C1(n6361), .C2(n7595), .A(n3539), 
        .ZN(n3536) );
  AOI22_X2 U1624 ( .A1(n7607), .A2(REG_FILE_reg_out_11__6_), .B1(n7603), .B2(
        REG_FILE_reg_out_15__6_), .ZN(n3539) );
  OAI221_X2 U1626 ( .B1(n5961), .B2(n7570), .C1(n6157), .C2(n7563), .A(n3542), 
        .ZN(n3541) );
  AOI22_X2 U1627 ( .A1(n7769), .A2(REG_FILE_reg_out_24__6_), .B1(n7576), .B2(
        REG_FILE_reg_out_28__6_), .ZN(n3542) );
  OAI221_X2 U1628 ( .B1(n6099), .B2(n7584), .C1(n5931), .C2(n7592), .A(n3543), 
        .ZN(n3540) );
  AOI22_X2 U1629 ( .A1(n7607), .A2(REG_FILE_reg_out_27__6_), .B1(n7601), .B2(
        REG_FILE_reg_out_31__6_), .ZN(n3543) );
  OAI221_X2 U1631 ( .B1(n6092), .B2(n7570), .C1(n6369), .C2(n7563), .A(n3546), 
        .ZN(n3545) );
  AOI22_X2 U1632 ( .A1(n7769), .A2(REG_FILE_reg_out_16__6_), .B1(n7576), .B2(
        REG_FILE_reg_out_20__6_), .ZN(n3546) );
  OAI221_X2 U1633 ( .B1(n6404), .B2(n7584), .C1(n6053), .C2(n7592), .A(n3547), 
        .ZN(n3544) );
  AOI22_X2 U1634 ( .A1(n7607), .A2(REG_FILE_reg_out_19__6_), .B1(n7601), .B2(
        REG_FILE_reg_out_23__6_), .ZN(n3547) );
  NAND4_X2 U1635 ( .A1(n3548), .A2(n3549), .A3(n3550), .A4(n3551), .ZN(
        ID_EX_REG_ID_EX_REG_N167) );
  AOI221_X2 U1638 ( .B1(n7608), .B2(REG_FILE_reg_out_3__7_), .C1(n7605), .C2(
        REG_FILE_reg_out_7__7_), .A(n3556), .ZN(n3555) );
  OAI22_X2 U1639 ( .A1(n5881), .A2(n7598), .B1(n6129), .B2(n7588), .ZN(n3556)
         );
  AOI22_X2 U1640 ( .A1(n7573), .A2(REG_FILE_reg_out_2__7_), .B1(n7565), .B2(
        REG_FILE_reg_out_6__7_), .ZN(n3554) );
  AOI22_X2 U1641 ( .A1(n7769), .A2(REG_FILE_reg_out_0__7_), .B1(n7576), .B2(
        REG_FILE_reg_out_4__7_), .ZN(n3553) );
  OAI221_X2 U1643 ( .B1(n6150), .B2(n7570), .C1(n6490), .C2(n7563), .A(n3560), 
        .ZN(n3559) );
  AOI22_X2 U1644 ( .A1(n7768), .A2(REG_FILE_reg_out_8__7_), .B1(n7581), .B2(
        REG_FILE_reg_out_12__7_), .ZN(n3560) );
  OAI221_X2 U1645 ( .B1(n6950), .B2(n7584), .C1(n6362), .C2(n7592), .A(n3561), 
        .ZN(n3558) );
  AOI22_X2 U1646 ( .A1(n7608), .A2(REG_FILE_reg_out_11__7_), .B1(n7603), .B2(
        REG_FILE_reg_out_15__7_), .ZN(n3561) );
  OAI221_X2 U1648 ( .B1(n5962), .B2(n7570), .C1(n6158), .C2(n7563), .A(n3564), 
        .ZN(n3563) );
  AOI22_X2 U1649 ( .A1(n7765), .A2(REG_FILE_reg_out_24__7_), .B1(n7582), .B2(
        REG_FILE_reg_out_28__7_), .ZN(n3564) );
  OAI221_X2 U1650 ( .B1(n6100), .B2(n7584), .C1(n5932), .C2(n7592), .A(n3565), 
        .ZN(n3562) );
  AOI22_X2 U1651 ( .A1(n7607), .A2(REG_FILE_reg_out_27__7_), .B1(n7603), .B2(
        REG_FILE_reg_out_31__7_), .ZN(n3565) );
  OAI221_X2 U1653 ( .B1(n6093), .B2(n7570), .C1(n6370), .C2(n7563), .A(n3568), 
        .ZN(n3567) );
  AOI22_X2 U1654 ( .A1(n7767), .A2(REG_FILE_reg_out_16__7_), .B1(n7579), .B2(
        REG_FILE_reg_out_20__7_), .ZN(n3568) );
  OAI221_X2 U1655 ( .B1(n6085), .B2(n7584), .C1(n5870), .C2(n7592), .A(n3569), 
        .ZN(n3566) );
  AOI22_X2 U1656 ( .A1(n7607), .A2(REG_FILE_reg_out_19__7_), .B1(n7602), .B2(
        REG_FILE_reg_out_23__7_), .ZN(n3569) );
  AOI221_X2 U1660 ( .B1(n7610), .B2(REG_FILE_reg_out_3__8_), .C1(n7600), .C2(
        REG_FILE_reg_out_7__8_), .A(n3578), .ZN(n3577) );
  OAI22_X2 U1661 ( .A1(n5883), .A2(n7596), .B1(n6133), .B2(n7588), .ZN(n3578)
         );
  AOI22_X2 U1662 ( .A1(n7573), .A2(REG_FILE_reg_out_2__8_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__8_), .ZN(n3576) );
  AOI22_X2 U1663 ( .A1(n7768), .A2(REG_FILE_reg_out_0__8_), .B1(n7581), .B2(
        REG_FILE_reg_out_4__8_), .ZN(n3575) );
  OAI221_X2 U1665 ( .B1(n7012), .B2(n7570), .C1(n6519), .C2(n7563), .A(n3581), 
        .ZN(n3580) );
  AOI22_X2 U1666 ( .A1(n7766), .A2(REG_FILE_reg_out_8__8_), .B1(n7581), .B2(
        REG_FILE_reg_out_12__8_), .ZN(n3581) );
  OAI221_X2 U1667 ( .B1(n6112), .B2(n7584), .C1(n5879), .C2(n7592), .A(n3582), 
        .ZN(n3579) );
  AOI22_X2 U1668 ( .A1(n7608), .A2(REG_FILE_reg_out_11__8_), .B1(n7602), .B2(
        REG_FILE_reg_out_15__8_), .ZN(n3582) );
  OAI221_X2 U1670 ( .B1(n7011), .B2(n7570), .C1(n6518), .C2(n7563), .A(n3585), 
        .ZN(n3584) );
  AOI22_X2 U1671 ( .A1(n7766), .A2(REG_FILE_reg_out_24__8_), .B1(n7581), .B2(
        REG_FILE_reg_out_28__8_), .ZN(n3585) );
  OAI221_X2 U1672 ( .B1(n6978), .B2(n7584), .C1(n6084), .C2(n7592), .A(n3586), 
        .ZN(n3583) );
  AOI22_X2 U1673 ( .A1(n7608), .A2(REG_FILE_reg_out_27__8_), .B1(n7603), .B2(
        REG_FILE_reg_out_31__8_), .ZN(n3586) );
  OAI221_X2 U1675 ( .B1(n6977), .B2(n7570), .C1(n6398), .C2(n7563), .A(n3589), 
        .ZN(n3588) );
  AOI22_X2 U1676 ( .A1(n7768), .A2(REG_FILE_reg_out_16__8_), .B1(n7582), .B2(
        REG_FILE_reg_out_20__8_), .ZN(n3589) );
  OAI221_X2 U1677 ( .B1(n6111), .B2(n7584), .C1(n5878), .C2(n7592), .A(n3590), 
        .ZN(n3587) );
  AOI22_X2 U1678 ( .A1(n7608), .A2(REG_FILE_reg_out_19__8_), .B1(n7603), .B2(
        REG_FILE_reg_out_23__8_), .ZN(n3590) );
  AOI221_X2 U1682 ( .B1(n7611), .B2(REG_FILE_reg_out_3__9_), .C1(n7602), .C2(
        REG_FILE_reg_out_7__9_), .A(n3599), .ZN(n3598) );
  OAI22_X2 U1683 ( .A1(n6980), .A2(n7596), .B1(n6132), .B2(n7588), .ZN(n3599)
         );
  AOI22_X2 U1684 ( .A1(n7573), .A2(REG_FILE_reg_out_2__9_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__9_), .ZN(n3597) );
  AOI22_X2 U1685 ( .A1(n7765), .A2(REG_FILE_reg_out_0__9_), .B1(n7579), .B2(
        REG_FILE_reg_out_4__9_), .ZN(n3596) );
  OAI221_X2 U1687 ( .B1(n7010), .B2(n7570), .C1(n6517), .C2(n7563), .A(n3603), 
        .ZN(n3602) );
  AOI22_X2 U1688 ( .A1(n7766), .A2(REG_FILE_reg_out_8__9_), .B1(n7582), .B2(
        REG_FILE_reg_out_12__9_), .ZN(n3603) );
  OAI221_X2 U1689 ( .B1(n6110), .B2(n7584), .C1(n5877), .C2(n7593), .A(n3604), 
        .ZN(n3601) );
  AOI22_X2 U1690 ( .A1(n7608), .A2(REG_FILE_reg_out_11__9_), .B1(n7602), .B2(
        REG_FILE_reg_out_15__9_), .ZN(n3604) );
  OAI221_X2 U1692 ( .B1(n6502), .B2(n7570), .C1(n7032), .C2(n7563), .A(n3607), 
        .ZN(n3606) );
  AOI22_X2 U1693 ( .A1(n7765), .A2(REG_FILE_reg_out_24__9_), .B1(n7582), .B2(
        REG_FILE_reg_out_28__9_), .ZN(n3607) );
  OAI221_X2 U1694 ( .B1(n6976), .B2(n7584), .C1(n6083), .C2(n7593), .A(n3608), 
        .ZN(n3605) );
  AOI22_X2 U1695 ( .A1(n7608), .A2(REG_FILE_reg_out_27__9_), .B1(n7603), .B2(
        REG_FILE_reg_out_31__9_), .ZN(n3608) );
  OAI221_X2 U1697 ( .B1(n6975), .B2(n7570), .C1(n6397), .C2(n7563), .A(n3611), 
        .ZN(n3610) );
  AOI22_X2 U1698 ( .A1(n7767), .A2(REG_FILE_reg_out_16__9_), .B1(n7581), .B2(
        REG_FILE_reg_out_20__9_), .ZN(n3611) );
  OAI221_X2 U1699 ( .B1(n6109), .B2(n7584), .C1(n5876), .C2(n7593), .A(n3612), 
        .ZN(n3609) );
  AOI22_X2 U1700 ( .A1(n7608), .A2(REG_FILE_reg_out_19__9_), .B1(n7603), .B2(
        REG_FILE_reg_out_23__9_), .ZN(n3612) );
  AOI221_X2 U1704 ( .B1(n7608), .B2(REG_FILE_reg_out_3__10_), .C1(n7600), .C2(
        REG_FILE_reg_out_7__10_), .A(n3621), .ZN(n3620) );
  OAI22_X2 U1705 ( .A1(n6460), .A2(n7596), .B1(n6127), .B2(n7588), .ZN(n3621)
         );
  AOI22_X2 U1706 ( .A1(n7573), .A2(REG_FILE_reg_out_2__10_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__10_), .ZN(n3619) );
  AOI22_X2 U1707 ( .A1(n7768), .A2(REG_FILE_reg_out_0__10_), .B1(n7582), .B2(
        REG_FILE_reg_out_4__10_), .ZN(n3618) );
  OAI221_X2 U1709 ( .B1(n5972), .B2(n7569), .C1(n6184), .C2(n7562), .A(n3624), 
        .ZN(n3623) );
  AOI22_X2 U1710 ( .A1(n7768), .A2(REG_FILE_reg_out_8__10_), .B1(n7582), .B2(
        REG_FILE_reg_out_12__10_), .ZN(n3624) );
  OAI221_X2 U1711 ( .B1(n6974), .B2(n7584), .C1(n6396), .C2(n7593), .A(n3625), 
        .ZN(n3622) );
  AOI22_X2 U1712 ( .A1(n7608), .A2(REG_FILE_reg_out_11__10_), .B1(n7602), .B2(
        REG_FILE_reg_out_15__10_), .ZN(n3625) );
  OAI221_X2 U1714 ( .B1(n5971), .B2(n7569), .C1(n6183), .C2(n7562), .A(n3628), 
        .ZN(n3627) );
  AOI22_X2 U1715 ( .A1(n7768), .A2(REG_FILE_reg_out_24__10_), .B1(n7582), .B2(
        REG_FILE_reg_out_28__10_), .ZN(n3628) );
  OAI221_X2 U1716 ( .B1(n6449), .B2(n7587), .C1(n6082), .C2(n7593), .A(n3629), 
        .ZN(n3626) );
  AOI22_X2 U1717 ( .A1(n7608), .A2(REG_FILE_reg_out_27__10_), .B1(n7602), .B2(
        REG_FILE_reg_out_31__10_), .ZN(n3629) );
  OAI221_X2 U1719 ( .B1(n6108), .B2(n7568), .C1(n5943), .C2(n7562), .A(n3632), 
        .ZN(n3631) );
  AOI22_X2 U1720 ( .A1(n7768), .A2(REG_FILE_reg_out_16__10_), .B1(n7582), .B2(
        REG_FILE_reg_out_20__10_), .ZN(n3632) );
  OAI221_X2 U1721 ( .B1(n6059), .B2(n7584), .C1(n6395), .C2(n7593), .A(n3633), 
        .ZN(n3630) );
  AOI22_X2 U1722 ( .A1(n7609), .A2(REG_FILE_reg_out_19__10_), .B1(n7602), .B2(
        REG_FILE_reg_out_23__10_), .ZN(n3633) );
  AOI221_X2 U1726 ( .B1(n7608), .B2(REG_FILE_reg_out_3__11_), .C1(n7602), .C2(
        REG_FILE_reg_out_7__11_), .A(n3642), .ZN(n3641) );
  OAI22_X2 U1727 ( .A1(n6459), .A2(n7596), .B1(n6986), .B2(n7588), .ZN(n3642)
         );
  AOI22_X2 U1728 ( .A1(n7573), .A2(REG_FILE_reg_out_2__11_), .B1(n7566), .B2(
        REG_FILE_reg_out_6__11_), .ZN(n3640) );
  AOI22_X2 U1729 ( .A1(n7768), .A2(REG_FILE_reg_out_0__11_), .B1(n7582), .B2(
        REG_FILE_reg_out_4__11_), .ZN(n3639) );
  OAI221_X2 U1731 ( .B1(n7009), .B2(n7568), .C1(n6182), .C2(n7562), .A(n3646), 
        .ZN(n3645) );
  AOI22_X2 U1732 ( .A1(n7768), .A2(REG_FILE_reg_out_8__11_), .B1(n7582), .B2(
        REG_FILE_reg_out_12__11_), .ZN(n3646) );
  OAI221_X2 U1733 ( .B1(n6973), .B2(n7584), .C1(n6394), .C2(n7593), .A(n3647), 
        .ZN(n3644) );
  AOI22_X2 U1734 ( .A1(n7609), .A2(REG_FILE_reg_out_11__11_), .B1(n7602), .B2(
        REG_FILE_reg_out_15__11_), .ZN(n3647) );
  OAI221_X2 U1736 ( .B1(n6173), .B2(n7568), .C1(n7031), .C2(n7562), .A(n3650), 
        .ZN(n3649) );
  AOI22_X2 U1737 ( .A1(n7768), .A2(REG_FILE_reg_out_24__11_), .B1(n7582), .B2(
        REG_FILE_reg_out_28__11_), .ZN(n3650) );
  OAI221_X2 U1738 ( .B1(n6972), .B2(n7584), .C1(n6393), .C2(n7593), .A(n3651), 
        .ZN(n3648) );
  AOI22_X2 U1739 ( .A1(n7609), .A2(REG_FILE_reg_out_27__11_), .B1(n7602), .B2(
        REG_FILE_reg_out_31__11_), .ZN(n3651) );
  OAI221_X2 U1741 ( .B1(n6971), .B2(n7568), .C1(n6081), .C2(n7562), .A(n3654), 
        .ZN(n3653) );
  AOI22_X2 U1742 ( .A1(n7768), .A2(REG_FILE_reg_out_16__11_), .B1(n7582), .B2(
        REG_FILE_reg_out_20__11_), .ZN(n3654) );
  OAI221_X2 U1743 ( .B1(n6922), .B2(n7584), .C1(n6392), .C2(n7593), .A(n3655), 
        .ZN(n3652) );
  AOI22_X2 U1744 ( .A1(n7609), .A2(REG_FILE_reg_out_19__11_), .B1(n7602), .B2(
        REG_FILE_reg_out_23__11_), .ZN(n3655) );
  AOI221_X2 U1748 ( .B1(n7606), .B2(REG_FILE_reg_out_3__12_), .C1(n7599), .C2(
        REG_FILE_reg_out_7__12_), .A(n3664), .ZN(n3663) );
  OAI22_X2 U1749 ( .A1(n6458), .A2(n7596), .B1(n6126), .B2(n7588), .ZN(n3664)
         );
  AOI22_X2 U1750 ( .A1(n7573), .A2(REG_FILE_reg_out_2__12_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__12_), .ZN(n3662) );
  AOI22_X2 U1751 ( .A1(n7768), .A2(REG_FILE_reg_out_0__12_), .B1(n7582), .B2(
        REG_FILE_reg_out_4__12_), .ZN(n3661) );
  OAI221_X2 U1753 ( .B1(n5970), .B2(n7569), .C1(n6181), .C2(n7562), .A(n3667), 
        .ZN(n3666) );
  AOI22_X2 U1754 ( .A1(n7768), .A2(REG_FILE_reg_out_8__12_), .B1(n7582), .B2(
        REG_FILE_reg_out_12__12_), .ZN(n3667) );
  OAI221_X2 U1755 ( .B1(n6448), .B2(n7583), .C1(n6080), .C2(n7595), .A(n3668), 
        .ZN(n3665) );
  AOI22_X2 U1756 ( .A1(n7609), .A2(REG_FILE_reg_out_11__12_), .B1(n7602), .B2(
        REG_FILE_reg_out_15__12_), .ZN(n3668) );
  OAI221_X2 U1758 ( .B1(n5969), .B2(n7569), .C1(n6180), .C2(n7562), .A(n3671), 
        .ZN(n3670) );
  AOI22_X2 U1759 ( .A1(n7768), .A2(REG_FILE_reg_out_24__12_), .B1(n7582), .B2(
        REG_FILE_reg_out_28__12_), .ZN(n3671) );
  OAI221_X2 U1760 ( .B1(n6447), .B2(n7583), .C1(n6079), .C2(n7594), .A(n3672), 
        .ZN(n3669) );
  AOI22_X2 U1761 ( .A1(n7609), .A2(REG_FILE_reg_out_27__12_), .B1(n7602), .B2(
        REG_FILE_reg_out_31__12_), .ZN(n3672) );
  OAI221_X2 U1763 ( .B1(n6107), .B2(n7569), .C1(n5942), .C2(n7562), .A(n3675), 
        .ZN(n3674) );
  AOI22_X2 U1764 ( .A1(n7767), .A2(REG_FILE_reg_out_16__12_), .B1(n7581), .B2(
        REG_FILE_reg_out_20__12_), .ZN(n3675) );
  OAI221_X2 U1765 ( .B1(n6058), .B2(n7583), .C1(n6391), .C2(n7594), .A(n3676), 
        .ZN(n3673) );
  AOI22_X2 U1766 ( .A1(n7609), .A2(REG_FILE_reg_out_19__12_), .B1(n7603), .B2(
        REG_FILE_reg_out_23__12_), .ZN(n3676) );
  AOI221_X2 U1770 ( .B1(n7606), .B2(REG_FILE_reg_out_3__13_), .C1(n7599), .C2(
        REG_FILE_reg_out_7__13_), .A(n3685), .ZN(n3684) );
  OAI22_X2 U1771 ( .A1(n6979), .A2(n7596), .B1(n6475), .B2(n7588), .ZN(n3685)
         );
  AOI22_X2 U1772 ( .A1(n7573), .A2(REG_FILE_reg_out_2__13_), .B1(n7565), .B2(
        REG_FILE_reg_out_6__13_), .ZN(n3683) );
  AOI22_X2 U1773 ( .A1(n7767), .A2(REG_FILE_reg_out_0__13_), .B1(n7581), .B2(
        REG_FILE_reg_out_4__13_), .ZN(n3682) );
  OAI221_X2 U1775 ( .B1(n5968), .B2(n7568), .C1(n6179), .C2(n7562), .A(n3689), 
        .ZN(n3688) );
  AOI22_X2 U1776 ( .A1(n7767), .A2(REG_FILE_reg_out_8__13_), .B1(n7581), .B2(
        REG_FILE_reg_out_12__13_), .ZN(n3689) );
  OAI221_X2 U1777 ( .B1(n6446), .B2(n7583), .C1(n6078), .C2(n7594), .A(n3690), 
        .ZN(n3687) );
  AOI22_X2 U1778 ( .A1(n7609), .A2(REG_FILE_reg_out_11__13_), .B1(n7603), .B2(
        REG_FILE_reg_out_15__13_), .ZN(n3690) );
  OAI221_X2 U1780 ( .B1(n5967), .B2(n7568), .C1(n6178), .C2(n7562), .A(n3693), 
        .ZN(n3692) );
  AOI22_X2 U1781 ( .A1(n7767), .A2(REG_FILE_reg_out_24__13_), .B1(n7581), .B2(
        REG_FILE_reg_out_28__13_), .ZN(n3693) );
  OAI221_X2 U1782 ( .B1(n6445), .B2(n7583), .C1(n6077), .C2(n7594), .A(n3694), 
        .ZN(n3691) );
  AOI22_X2 U1783 ( .A1(n7609), .A2(REG_FILE_reg_out_27__13_), .B1(n7603), .B2(
        REG_FILE_reg_out_31__13_), .ZN(n3694) );
  OAI221_X2 U1785 ( .B1(n6106), .B2(n7569), .C1(n5941), .C2(n7562), .A(n3697), 
        .ZN(n3696) );
  AOI22_X2 U1786 ( .A1(n7767), .A2(REG_FILE_reg_out_16__13_), .B1(n7581), .B2(
        REG_FILE_reg_out_20__13_), .ZN(n3697) );
  OAI221_X2 U1787 ( .B1(n6444), .B2(n7583), .C1(n6076), .C2(n7595), .A(n3698), 
        .ZN(n3695) );
  AOI22_X2 U1788 ( .A1(n7609), .A2(REG_FILE_reg_out_19__13_), .B1(n7603), .B2(
        REG_FILE_reg_out_23__13_), .ZN(n3698) );
  AOI221_X2 U1792 ( .B1(n7606), .B2(REG_FILE_reg_out_3__14_), .C1(n7599), .C2(
        REG_FILE_reg_out_7__14_), .A(n3707), .ZN(n3706) );
  OAI22_X2 U1793 ( .A1(n6457), .A2(n7596), .B1(n6985), .B2(n7588), .ZN(n3707)
         );
  AOI22_X2 U1794 ( .A1(n7573), .A2(REG_FILE_reg_out_2__14_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__14_), .ZN(n3705) );
  AOI22_X2 U1795 ( .A1(n7767), .A2(REG_FILE_reg_out_0__14_), .B1(n7581), .B2(
        REG_FILE_reg_out_4__14_), .ZN(n3704) );
  OAI221_X2 U1797 ( .B1(n5966), .B2(n7569), .C1(n6177), .C2(n7561), .A(n3710), 
        .ZN(n3709) );
  AOI22_X2 U1798 ( .A1(n7767), .A2(REG_FILE_reg_out_8__14_), .B1(n7581), .B2(
        REG_FILE_reg_out_12__14_), .ZN(n3710) );
  OAI221_X2 U1799 ( .B1(n6443), .B2(n7583), .C1(n6075), .C2(n7594), .A(n3711), 
        .ZN(n3708) );
  AOI22_X2 U1800 ( .A1(n7609), .A2(REG_FILE_reg_out_11__14_), .B1(n7603), .B2(
        REG_FILE_reg_out_15__14_), .ZN(n3711) );
  OAI221_X2 U1802 ( .B1(n5965), .B2(n7569), .C1(n6176), .C2(n7562), .A(n3714), 
        .ZN(n3713) );
  AOI22_X2 U1803 ( .A1(n7767), .A2(REG_FILE_reg_out_24__14_), .B1(n7581), .B2(
        REG_FILE_reg_out_28__14_), .ZN(n3714) );
  OAI221_X2 U1804 ( .B1(n6442), .B2(n7583), .C1(n6074), .C2(n7595), .A(n3715), 
        .ZN(n3712) );
  AOI22_X2 U1805 ( .A1(n7609), .A2(REG_FILE_reg_out_27__14_), .B1(n7603), .B2(
        REG_FILE_reg_out_31__14_), .ZN(n3715) );
  OAI221_X2 U1807 ( .B1(n6105), .B2(n7569), .C1(n5940), .C2(n7561), .A(n3718), 
        .ZN(n3717) );
  AOI22_X2 U1808 ( .A1(n7767), .A2(REG_FILE_reg_out_16__14_), .B1(n7581), .B2(
        REG_FILE_reg_out_20__14_), .ZN(n3718) );
  OAI221_X2 U1809 ( .B1(n6057), .B2(n7583), .C1(n6390), .C2(n7595), .A(n3719), 
        .ZN(n3716) );
  AOI22_X2 U1810 ( .A1(n7609), .A2(REG_FILE_reg_out_19__14_), .B1(n7603), .B2(
        REG_FILE_reg_out_23__14_), .ZN(n3719) );
  AOI221_X2 U1815 ( .B1(n7606), .B2(REG_FILE_reg_out_3__15_), .C1(n7599), .C2(
        REG_FILE_reg_out_7__15_), .A(n3729), .ZN(n3728) );
  OAI22_X2 U1816 ( .A1(n6456), .A2(n7598), .B1(n6984), .B2(n7589), .ZN(n3729)
         );
  AOI22_X2 U1817 ( .A1(n7573), .A2(REG_FILE_reg_out_2__15_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__15_), .ZN(n3727) );
  AOI22_X2 U1818 ( .A1(n7767), .A2(REG_FILE_reg_out_0__15_), .B1(n7581), .B2(
        REG_FILE_reg_out_4__15_), .ZN(n3726) );
  OAI221_X2 U1820 ( .B1(n7008), .B2(n7569), .C1(n6175), .C2(n7562), .A(n3733), 
        .ZN(n3732) );
  AOI22_X2 U1821 ( .A1(n7767), .A2(REG_FILE_reg_out_8__15_), .B1(n7581), .B2(
        REG_FILE_reg_out_12__15_), .ZN(n3733) );
  OAI221_X2 U1822 ( .B1(n6970), .B2(n7585), .C1(n6389), .C2(n7594), .A(n3734), 
        .ZN(n3731) );
  AOI22_X2 U1823 ( .A1(n7609), .A2(REG_FILE_reg_out_11__15_), .B1(n7603), .B2(
        REG_FILE_reg_out_15__15_), .ZN(n3734) );
  OAI221_X2 U1825 ( .B1(n6172), .B2(n7569), .C1(n7030), .C2(n7561), .A(n3737), 
        .ZN(n3736) );
  AOI22_X2 U1826 ( .A1(n7766), .A2(REG_FILE_reg_out_24__15_), .B1(n7580), .B2(
        REG_FILE_reg_out_28__15_), .ZN(n3737) );
  OAI221_X2 U1827 ( .B1(n6969), .B2(n7585), .C1(n6388), .C2(n7594), .A(n3738), 
        .ZN(n3735) );
  AOI22_X2 U1828 ( .A1(n7609), .A2(REG_FILE_reg_out_27__15_), .B1(n7603), .B2(
        REG_FILE_reg_out_31__15_), .ZN(n3738) );
  OAI221_X2 U1830 ( .B1(n6968), .B2(n7569), .C1(n6073), .C2(n7562), .A(n3741), 
        .ZN(n3740) );
  AOI22_X2 U1831 ( .A1(n7766), .A2(REG_FILE_reg_out_16__15_), .B1(n7580), .B2(
        REG_FILE_reg_out_20__15_), .ZN(n3741) );
  OAI221_X2 U1832 ( .B1(n6921), .B2(n7585), .C1(n6387), .C2(n7594), .A(n3742), 
        .ZN(n3739) );
  AOI22_X2 U1833 ( .A1(n7609), .A2(REG_FILE_reg_out_19__15_), .B1(n7603), .B2(
        REG_FILE_reg_out_23__15_), .ZN(n3742) );
  AOI221_X2 U1837 ( .B1(n7606), .B2(REG_FILE_reg_out_3__16_), .C1(n7601), .C2(
        REG_FILE_reg_out_7__16_), .A(n3752), .ZN(n3751) );
  OAI22_X2 U1838 ( .A1(n6455), .A2(n7598), .B1(n6983), .B2(n7589), .ZN(n3752)
         );
  AOI22_X2 U1839 ( .A1(n7573), .A2(REG_FILE_reg_out_2__16_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__16_), .ZN(n3750) );
  AOI22_X2 U1840 ( .A1(n7766), .A2(REG_FILE_reg_out_0__16_), .B1(n7580), .B2(
        REG_FILE_reg_out_4__16_), .ZN(n3749) );
  OAI221_X2 U1842 ( .B1(n6171), .B2(n7569), .C1(n7029), .C2(n7561), .A(n3755), 
        .ZN(n3754) );
  AOI22_X2 U1843 ( .A1(n7766), .A2(REG_FILE_reg_out_8__16_), .B1(n7580), .B2(
        REG_FILE_reg_out_12__16_), .ZN(n3755) );
  OAI221_X2 U1844 ( .B1(n6441), .B2(n7585), .C1(n6945), .C2(n7594), .A(n3756), 
        .ZN(n3753) );
  AOI22_X2 U1845 ( .A1(n7609), .A2(REG_FILE_reg_out_11__16_), .B1(n7604), .B2(
        REG_FILE_reg_out_15__16_), .ZN(n3756) );
  OAI221_X2 U1847 ( .B1(n5964), .B2(n7569), .C1(n6174), .C2(n7561), .A(n3759), 
        .ZN(n3758) );
  AOI22_X2 U1848 ( .A1(n7766), .A2(REG_FILE_reg_out_24__16_), .B1(n7580), .B2(
        REG_FILE_reg_out_28__16_), .ZN(n3759) );
  OAI221_X2 U1849 ( .B1(n6440), .B2(n7585), .C1(n6072), .C2(n7594), .A(n3760), 
        .ZN(n3757) );
  AOI22_X2 U1850 ( .A1(n7609), .A2(REG_FILE_reg_out_27__16_), .B1(n7600), .B2(
        REG_FILE_reg_out_31__16_), .ZN(n3760) );
  OAI221_X2 U1852 ( .B1(n6104), .B2(n7569), .C1(n6944), .C2(n7561), .A(n3763), 
        .ZN(n3762) );
  AOI22_X2 U1853 ( .A1(n7766), .A2(REG_FILE_reg_out_16__16_), .B1(n7580), .B2(
        REG_FILE_reg_out_20__16_), .ZN(n3763) );
  OAI221_X2 U1854 ( .B1(n6056), .B2(n7585), .C1(n6943), .C2(n7594), .A(n3764), 
        .ZN(n3761) );
  AOI22_X2 U1855 ( .A1(n7610), .A2(REG_FILE_reg_out_19__16_), .B1(n7602), .B2(
        REG_FILE_reg_out_23__16_), .ZN(n3764) );
  AOI221_X2 U1859 ( .B1(n7606), .B2(REG_FILE_reg_out_3__17_), .C1(n7599), .C2(
        REG_FILE_reg_out_7__17_), .A(n3773), .ZN(n3772) );
  OAI22_X2 U1860 ( .A1(n6122), .A2(n7598), .B1(n6474), .B2(n7589), .ZN(n3773)
         );
  AOI22_X2 U1861 ( .A1(n7573), .A2(REG_FILE_reg_out_2__17_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__17_), .ZN(n3771) );
  AOI22_X2 U1862 ( .A1(n7766), .A2(REG_FILE_reg_out_0__17_), .B1(n7580), .B2(
        REG_FILE_reg_out_4__17_), .ZN(n3770) );
  OAI221_X2 U1864 ( .B1(n6170), .B2(n7569), .C1(n7028), .C2(n7562), .A(n3776), 
        .ZN(n3775) );
  AOI22_X2 U1865 ( .A1(n7766), .A2(REG_FILE_reg_out_8__17_), .B1(n7580), .B2(
        REG_FILE_reg_out_12__17_), .ZN(n3776) );
  OAI221_X2 U1866 ( .B1(n6439), .B2(n7585), .C1(n6942), .C2(n7594), .A(n3777), 
        .ZN(n3774) );
  AOI22_X2 U1867 ( .A1(n7610), .A2(REG_FILE_reg_out_11__17_), .B1(n7604), .B2(
        REG_FILE_reg_out_15__17_), .ZN(n3777) );
  OAI221_X2 U1869 ( .B1(n6169), .B2(n7568), .C1(n6516), .C2(n7561), .A(n3780), 
        .ZN(n3779) );
  AOI22_X2 U1870 ( .A1(n7766), .A2(REG_FILE_reg_out_24__17_), .B1(n7580), .B2(
        REG_FILE_reg_out_28__17_), .ZN(n3780) );
  OAI221_X2 U1871 ( .B1(n6438), .B2(n7585), .C1(n6071), .C2(n7594), .A(n3781), 
        .ZN(n3778) );
  AOI22_X2 U1872 ( .A1(n7610), .A2(REG_FILE_reg_out_27__17_), .B1(n7604), .B2(
        REG_FILE_reg_out_31__17_), .ZN(n3781) );
  OAI221_X2 U1874 ( .B1(n6437), .B2(n7568), .C1(n6941), .C2(n7561), .A(n3784), 
        .ZN(n3783) );
  AOI22_X2 U1875 ( .A1(n7766), .A2(REG_FILE_reg_out_16__17_), .B1(n7580), .B2(
        REG_FILE_reg_out_20__17_), .ZN(n3784) );
  OAI221_X2 U1876 ( .B1(n6436), .B2(n7585), .C1(n6940), .C2(n7594), .A(n3785), 
        .ZN(n3782) );
  AOI22_X2 U1877 ( .A1(n7610), .A2(REG_FILE_reg_out_19__17_), .B1(n7600), .B2(
        REG_FILE_reg_out_23__17_), .ZN(n3785) );
  AOI221_X2 U1881 ( .B1(n7606), .B2(REG_FILE_reg_out_3__18_), .C1(n7599), .C2(
        REG_FILE_reg_out_7__18_), .A(n3794), .ZN(n3793) );
  OAI22_X2 U1882 ( .A1(n5951), .A2(n7598), .B1(n6473), .B2(n7589), .ZN(n3794)
         );
  AOI22_X2 U1883 ( .A1(n7573), .A2(REG_FILE_reg_out_2__18_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__18_), .ZN(n3792) );
  AOI22_X2 U1884 ( .A1(n7766), .A2(REG_FILE_reg_out_0__18_), .B1(n7580), .B2(
        REG_FILE_reg_out_4__18_), .ZN(n3791) );
  OAI221_X2 U1886 ( .B1(n6501), .B2(n7568), .C1(n7027), .C2(n7561), .A(n3797), 
        .ZN(n3796) );
  AOI22_X2 U1887 ( .A1(n7765), .A2(REG_FILE_reg_out_8__18_), .B1(n7580), .B2(
        REG_FILE_reg_out_12__18_), .ZN(n3797) );
  OAI221_X2 U1888 ( .B1(n6435), .B2(n7586), .C1(n6939), .C2(n7595), .A(n3798), 
        .ZN(n3795) );
  AOI22_X2 U1889 ( .A1(n7610), .A2(REG_FILE_reg_out_11__18_), .B1(n7600), .B2(
        REG_FILE_reg_out_15__18_), .ZN(n3798) );
  OAI221_X2 U1891 ( .B1(n6168), .B2(n7568), .C1(n6515), .C2(n7561), .A(n3801), 
        .ZN(n3800) );
  AOI22_X2 U1892 ( .A1(n7765), .A2(REG_FILE_reg_out_24__18_), .B1(n7580), .B2(
        REG_FILE_reg_out_28__18_), .ZN(n3801) );
  OAI221_X2 U1893 ( .B1(n6434), .B2(n7586), .C1(n5939), .C2(n7595), .A(n3802), 
        .ZN(n3799) );
  AOI22_X2 U1894 ( .A1(n7610), .A2(REG_FILE_reg_out_27__18_), .B1(n7602), .B2(
        REG_FILE_reg_out_31__18_), .ZN(n3802) );
  OAI221_X2 U1896 ( .B1(n6433), .B2(n7568), .C1(n6938), .C2(n7561), .A(n3805), 
        .ZN(n3804) );
  AOI22_X2 U1897 ( .A1(n7765), .A2(REG_FILE_reg_out_16__18_), .B1(n7580), .B2(
        REG_FILE_reg_out_20__18_), .ZN(n3805) );
  OAI221_X2 U1898 ( .B1(n6432), .B2(n7586), .C1(n6937), .C2(n7595), .A(n3806), 
        .ZN(n3803) );
  AOI22_X2 U1899 ( .A1(n7610), .A2(REG_FILE_reg_out_19__18_), .B1(n7602), .B2(
        REG_FILE_reg_out_23__18_), .ZN(n3806) );
  AOI221_X2 U1903 ( .B1(n7606), .B2(REG_FILE_reg_out_3__19_), .C1(n7599), .C2(
        REG_FILE_reg_out_7__19_), .A(n3815), .ZN(n3814) );
  OAI22_X2 U1904 ( .A1(n6454), .A2(n7598), .B1(n6987), .B2(n7589), .ZN(n3815)
         );
  AOI22_X2 U1905 ( .A1(n7573), .A2(REG_FILE_reg_out_2__19_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__19_), .ZN(n3813) );
  AOI22_X2 U1906 ( .A1(n7765), .A2(REG_FILE_reg_out_0__19_), .B1(n7580), .B2(
        REG_FILE_reg_out_4__19_), .ZN(n3812) );
  OAI221_X2 U1908 ( .B1(n6167), .B2(n7568), .C1(n7026), .C2(n7561), .A(n3818), 
        .ZN(n3817) );
  AOI22_X2 U1909 ( .A1(n7765), .A2(REG_FILE_reg_out_8__19_), .B1(n7580), .B2(
        REG_FILE_reg_out_12__19_), .ZN(n3818) );
  OAI221_X2 U1910 ( .B1(n6431), .B2(n7586), .C1(n5938), .C2(n7595), .A(n3819), 
        .ZN(n3816) );
  AOI22_X2 U1911 ( .A1(n7610), .A2(REG_FILE_reg_out_11__19_), .B1(n7604), .B2(
        REG_FILE_reg_out_15__19_), .ZN(n3819) );
  OAI221_X2 U1913 ( .B1(n6166), .B2(n7568), .C1(n6514), .C2(n7561), .A(n3822), 
        .ZN(n3821) );
  AOI22_X2 U1914 ( .A1(n7765), .A2(REG_FILE_reg_out_24__19_), .B1(n7580), .B2(
        REG_FILE_reg_out_28__19_), .ZN(n3822) );
  OAI221_X2 U1915 ( .B1(n6430), .B2(n7586), .C1(n5937), .C2(n7595), .A(n3823), 
        .ZN(n3820) );
  AOI22_X2 U1916 ( .A1(n7610), .A2(REG_FILE_reg_out_27__19_), .B1(n7604), .B2(
        REG_FILE_reg_out_31__19_), .ZN(n3823) );
  OAI221_X2 U1918 ( .B1(n6967), .B2(n7568), .C1(n6386), .C2(n7561), .A(n3826), 
        .ZN(n3825) );
  AOI22_X2 U1919 ( .A1(n7765), .A2(REG_FILE_reg_out_16__19_), .B1(n7580), .B2(
        REG_FILE_reg_out_20__19_), .ZN(n3826) );
  OAI221_X2 U1920 ( .B1(n6966), .B2(n7586), .C1(n6385), .C2(n7595), .A(n3827), 
        .ZN(n3824) );
  AOI22_X2 U1921 ( .A1(n7610), .A2(REG_FILE_reg_out_19__19_), .B1(n7604), .B2(
        REG_FILE_reg_out_23__19_), .ZN(n3827) );
  AOI221_X2 U1925 ( .B1(n7606), .B2(REG_FILE_reg_out_3__20_), .C1(n7599), .C2(
        REG_FILE_reg_out_7__20_), .A(n3836), .ZN(n3835) );
  OAI22_X2 U1926 ( .A1(n5950), .A2(n7598), .B1(n6472), .B2(n7589), .ZN(n3836)
         );
  AOI22_X2 U1927 ( .A1(n7573), .A2(REG_FILE_reg_out_2__20_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__20_), .ZN(n3834) );
  AOI22_X2 U1928 ( .A1(n7765), .A2(REG_FILE_reg_out_0__20_), .B1(n7580), .B2(
        REG_FILE_reg_out_4__20_), .ZN(n3833) );
  OAI221_X2 U1930 ( .B1(n6500), .B2(n7568), .C1(n7025), .C2(n7561), .A(n3839), 
        .ZN(n3838) );
  AOI22_X2 U1931 ( .A1(n7765), .A2(REG_FILE_reg_out_8__20_), .B1(n7580), .B2(
        REG_FILE_reg_out_12__20_), .ZN(n3839) );
  OAI221_X2 U1932 ( .B1(n6429), .B2(n7586), .C1(n6936), .C2(n7595), .A(n3840), 
        .ZN(n3837) );
  AOI22_X2 U1933 ( .A1(n7611), .A2(REG_FILE_reg_out_11__20_), .B1(n7604), .B2(
        REG_FILE_reg_out_15__20_), .ZN(n3840) );
  OAI221_X2 U1935 ( .B1(n6165), .B2(n7568), .C1(n6513), .C2(n7561), .A(n3843), 
        .ZN(n3842) );
  AOI22_X2 U1936 ( .A1(n7765), .A2(REG_FILE_reg_out_24__20_), .B1(n7580), .B2(
        REG_FILE_reg_out_28__20_), .ZN(n3843) );
  OAI221_X2 U1937 ( .B1(n6428), .B2(n7586), .C1(n5936), .C2(n7595), .A(n3844), 
        .ZN(n3841) );
  AOI22_X2 U1938 ( .A1(n7611), .A2(REG_FILE_reg_out_27__20_), .B1(n7604), .B2(
        REG_FILE_reg_out_31__20_), .ZN(n3844) );
  OAI221_X2 U1940 ( .B1(n6427), .B2(n7568), .C1(n6935), .C2(n7561), .A(n3847), 
        .ZN(n3846) );
  AOI22_X2 U1941 ( .A1(n7765), .A2(REG_FILE_reg_out_16__20_), .B1(n7580), .B2(
        REG_FILE_reg_out_20__20_), .ZN(n3847) );
  OAI221_X2 U1942 ( .B1(n6426), .B2(n7586), .C1(n6934), .C2(n7596), .A(n3848), 
        .ZN(n3845) );
  AOI22_X2 U1943 ( .A1(n7611), .A2(REG_FILE_reg_out_19__20_), .B1(n7604), .B2(
        REG_FILE_reg_out_23__20_), .ZN(n3848) );
  AOI221_X2 U1947 ( .B1(n7606), .B2(REG_FILE_reg_out_3__21_), .C1(n7599), .C2(
        REG_FILE_reg_out_7__21_), .A(n3857), .ZN(n3856) );
  OAI22_X2 U1948 ( .A1(n6121), .A2(n7598), .B1(n6471), .B2(n7589), .ZN(n3857)
         );
  AOI22_X2 U1949 ( .A1(n7573), .A2(REG_FILE_reg_out_2__21_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__21_), .ZN(n3855) );
  AOI22_X2 U1950 ( .A1(n7765), .A2(REG_FILE_reg_out_0__21_), .B1(n7579), .B2(
        REG_FILE_reg_out_4__21_), .ZN(n3854) );
  OAI221_X2 U1952 ( .B1(n6499), .B2(n7570), .C1(n7024), .C2(n7560), .A(n3860), 
        .ZN(n3859) );
  AOI22_X2 U1953 ( .A1(n7765), .A2(REG_FILE_reg_out_8__21_), .B1(n7579), .B2(
        REG_FILE_reg_out_12__21_), .ZN(n3860) );
  OAI221_X2 U1954 ( .B1(n6425), .B2(n7586), .C1(n6933), .C2(n7596), .A(n3861), 
        .ZN(n3858) );
  AOI22_X2 U1955 ( .A1(n7611), .A2(REG_FILE_reg_out_11__21_), .B1(n7604), .B2(
        REG_FILE_reg_out_15__21_), .ZN(n3861) );
  OAI221_X2 U1957 ( .B1(n6164), .B2(n7569), .C1(n6512), .C2(n7560), .A(n3864), 
        .ZN(n3863) );
  AOI22_X2 U1958 ( .A1(n7765), .A2(REG_FILE_reg_out_24__21_), .B1(n7579), .B2(
        REG_FILE_reg_out_28__21_), .ZN(n3864) );
  OAI221_X2 U1959 ( .B1(n6424), .B2(n7585), .C1(n6070), .C2(n7596), .A(n3865), 
        .ZN(n3862) );
  AOI22_X2 U1960 ( .A1(n7611), .A2(REG_FILE_reg_out_27__21_), .B1(n7604), .B2(
        REG_FILE_reg_out_31__21_), .ZN(n3865) );
  OAI221_X2 U1962 ( .B1(n6423), .B2(n7571), .C1(n6932), .C2(n7559), .A(n3868), 
        .ZN(n3867) );
  AOI22_X2 U1963 ( .A1(n7765), .A2(REG_FILE_reg_out_16__21_), .B1(n7579), .B2(
        REG_FILE_reg_out_20__21_), .ZN(n3868) );
  OAI221_X2 U1964 ( .B1(n6422), .B2(n7585), .C1(n6931), .C2(n7596), .A(n3869), 
        .ZN(n3866) );
  AOI22_X2 U1965 ( .A1(n7611), .A2(REG_FILE_reg_out_19__21_), .B1(n7604), .B2(
        REG_FILE_reg_out_23__21_), .ZN(n3869) );
  AOI221_X2 U1969 ( .B1(n7606), .B2(REG_FILE_reg_out_3__22_), .C1(n7605), .C2(
        REG_FILE_reg_out_7__22_), .A(n3878), .ZN(n3877) );
  OAI22_X2 U1970 ( .A1(n6120), .A2(n7598), .B1(n6470), .B2(n7589), .ZN(n3878)
         );
  AOI22_X2 U1971 ( .A1(n7573), .A2(REG_FILE_reg_out_2__22_), .B1(n7565), .B2(
        REG_FILE_reg_out_6__22_), .ZN(n3876) );
  AOI22_X2 U1972 ( .A1(n7765), .A2(REG_FILE_reg_out_0__22_), .B1(n7579), .B2(
        REG_FILE_reg_out_4__22_), .ZN(n3875) );
  OAI221_X2 U1974 ( .B1(n6498), .B2(n7569), .C1(n7023), .C2(n7559), .A(n3881), 
        .ZN(n3880) );
  AOI22_X2 U1975 ( .A1(n7765), .A2(REG_FILE_reg_out_8__22_), .B1(n7579), .B2(
        REG_FILE_reg_out_12__22_), .ZN(n3881) );
  OAI221_X2 U1976 ( .B1(n6421), .B2(n7585), .C1(n6930), .C2(n7596), .A(n3882), 
        .ZN(n3879) );
  AOI22_X2 U1977 ( .A1(n7611), .A2(REG_FILE_reg_out_11__22_), .B1(n7605), .B2(
        REG_FILE_reg_out_15__22_), .ZN(n3882) );
  OAI221_X2 U1979 ( .B1(n6163), .B2(n7568), .C1(n6511), .C2(n7559), .A(n3885), 
        .ZN(n3884) );
  AOI22_X2 U1980 ( .A1(n7765), .A2(REG_FILE_reg_out_24__22_), .B1(n7579), .B2(
        REG_FILE_reg_out_28__22_), .ZN(n3885) );
  OAI221_X2 U1981 ( .B1(n6420), .B2(n7586), .C1(n6069), .C2(n7596), .A(n3886), 
        .ZN(n3883) );
  AOI22_X2 U1982 ( .A1(n7611), .A2(REG_FILE_reg_out_27__22_), .B1(n7605), .B2(
        REG_FILE_reg_out_31__22_), .ZN(n3886) );
  OAI221_X2 U1984 ( .B1(n6419), .B2(n7570), .C1(n6929), .C2(n7560), .A(n3889), 
        .ZN(n3888) );
  AOI22_X2 U1985 ( .A1(n7765), .A2(REG_FILE_reg_out_16__22_), .B1(n7579), .B2(
        REG_FILE_reg_out_20__22_), .ZN(n3889) );
  OAI221_X2 U1986 ( .B1(n6418), .B2(n7586), .C1(n6928), .C2(n7596), .A(n3890), 
        .ZN(n3887) );
  AOI22_X2 U1987 ( .A1(n7611), .A2(REG_FILE_reg_out_19__22_), .B1(n7605), .B2(
        REG_FILE_reg_out_23__22_), .ZN(n3890) );
  AOI221_X2 U1991 ( .B1(n7606), .B2(REG_FILE_reg_out_3__23_), .C1(n7601), .C2(
        REG_FILE_reg_out_7__23_), .A(n3899), .ZN(n3898) );
  OAI22_X2 U1992 ( .A1(n6453), .A2(n7598), .B1(n6982), .B2(n7589), .ZN(n3899)
         );
  AOI22_X2 U1993 ( .A1(n7573), .A2(REG_FILE_reg_out_2__23_), .B1(n7565), .B2(
        REG_FILE_reg_out_6__23_), .ZN(n3897) );
  AOI22_X2 U1994 ( .A1(n7765), .A2(REG_FILE_reg_out_0__23_), .B1(n7579), .B2(
        REG_FILE_reg_out_4__23_), .ZN(n3896) );
  OAI221_X2 U1996 ( .B1(n6497), .B2(n7571), .C1(n7022), .C2(n7559), .A(n3902), 
        .ZN(n3901) );
  AOI22_X2 U1997 ( .A1(n7765), .A2(REG_FILE_reg_out_8__23_), .B1(n7579), .B2(
        REG_FILE_reg_out_12__23_), .ZN(n3902) );
  OAI221_X2 U1998 ( .B1(n6965), .B2(n7586), .C1(n6384), .C2(n7596), .A(n3903), 
        .ZN(n3900) );
  AOI22_X2 U1999 ( .A1(n7610), .A2(REG_FILE_reg_out_11__23_), .B1(n7605), .B2(
        REG_FILE_reg_out_15__23_), .ZN(n3903) );
  OAI221_X2 U2001 ( .B1(n6162), .B2(n7571), .C1(n6510), .C2(n7560), .A(n3906), 
        .ZN(n3905) );
  AOI22_X2 U2002 ( .A1(n7765), .A2(REG_FILE_reg_out_24__23_), .B1(n7579), .B2(
        REG_FILE_reg_out_28__23_), .ZN(n3906) );
  OAI221_X2 U2003 ( .B1(n6417), .B2(n7585), .C1(n6068), .C2(n7596), .A(n3907), 
        .ZN(n3904) );
  AOI22_X2 U2004 ( .A1(n7611), .A2(REG_FILE_reg_out_27__23_), .B1(n7605), .B2(
        REG_FILE_reg_out_31__23_), .ZN(n3907) );
  OAI221_X2 U2006 ( .B1(n6416), .B2(n7571), .C1(n6927), .C2(n7559), .A(n3910), 
        .ZN(n3909) );
  AOI22_X2 U2007 ( .A1(n7763), .A2(REG_FILE_reg_out_16__23_), .B1(n7579), .B2(
        REG_FILE_reg_out_20__23_), .ZN(n3910) );
  OAI221_X2 U2008 ( .B1(n6055), .B2(n7587), .C1(n6383), .C2(n7597), .A(n3911), 
        .ZN(n3908) );
  AOI22_X2 U2009 ( .A1(n7610), .A2(REG_FILE_reg_out_19__23_), .B1(n7605), .B2(
        REG_FILE_reg_out_23__23_), .ZN(n3911) );
  AOI221_X2 U2013 ( .B1(n7606), .B2(REG_FILE_reg_out_3__24_), .C1(n7601), .C2(
        REG_FILE_reg_out_7__24_), .A(n3920), .ZN(n3919) );
  OAI22_X2 U2014 ( .A1(n6119), .A2(n7598), .B1(n6469), .B2(n7589), .ZN(n3920)
         );
  AOI22_X2 U2015 ( .A1(n7573), .A2(REG_FILE_reg_out_2__24_), .B1(n7565), .B2(
        REG_FILE_reg_out_6__24_), .ZN(n3918) );
  AOI22_X2 U2016 ( .A1(n7763), .A2(REG_FILE_reg_out_0__24_), .B1(n7579), .B2(
        REG_FILE_reg_out_4__24_), .ZN(n3917) );
  OAI221_X2 U2018 ( .B1(n7007), .B2(n7570), .C1(n6509), .C2(n7560), .A(n3923), 
        .ZN(n3922) );
  AOI22_X2 U2019 ( .A1(n7763), .A2(REG_FILE_reg_out_8__24_), .B1(n7582), .B2(
        REG_FILE_reg_out_12__24_), .ZN(n3923) );
  OAI221_X2 U2020 ( .B1(n6415), .B2(n7587), .C1(n6067), .C2(n7597), .A(n3924), 
        .ZN(n3921) );
  AOI22_X2 U2021 ( .A1(n7611), .A2(REG_FILE_reg_out_11__24_), .B1(n7605), .B2(
        REG_FILE_reg_out_15__24_), .ZN(n3924) );
  OAI221_X2 U2023 ( .B1(n6496), .B2(n7570), .C1(n7021), .C2(n7559), .A(n3927), 
        .ZN(n3926) );
  AOI22_X2 U2024 ( .A1(n7763), .A2(REG_FILE_reg_out_24__24_), .B1(n7582), .B2(
        REG_FILE_reg_out_28__24_), .ZN(n3927) );
  OAI221_X2 U2025 ( .B1(n6414), .B2(n7587), .C1(n6066), .C2(n7597), .A(n3928), 
        .ZN(n3925) );
  AOI22_X2 U2026 ( .A1(n7610), .A2(REG_FILE_reg_out_27__24_), .B1(n7605), .B2(
        REG_FILE_reg_out_31__24_), .ZN(n3928) );
  OAI221_X2 U2028 ( .B1(n6964), .B2(n7568), .C1(n6382), .C2(n7560), .A(n3931), 
        .ZN(n3930) );
  AOI22_X2 U2029 ( .A1(n7763), .A2(REG_FILE_reg_out_16__24_), .B1(n7582), .B2(
        REG_FILE_reg_out_20__24_), .ZN(n3931) );
  OAI221_X2 U2030 ( .B1(n6413), .B2(n7587), .C1(n6065), .C2(n7597), .A(n3932), 
        .ZN(n3929) );
  AOI22_X2 U2031 ( .A1(n7610), .A2(REG_FILE_reg_out_19__24_), .B1(n7605), .B2(
        REG_FILE_reg_out_23__24_), .ZN(n3932) );
  AOI221_X2 U2036 ( .B1(n7606), .B2(REG_FILE_reg_out_3__25_), .C1(n7600), .C2(
        REG_FILE_reg_out_7__25_), .A(n3942), .ZN(n3941) );
  OAI22_X2 U2037 ( .A1(n6452), .A2(n7598), .B1(n6125), .B2(n7589), .ZN(n3942)
         );
  AOI22_X2 U2038 ( .A1(n7573), .A2(REG_FILE_reg_out_2__25_), .B1(n7565), .B2(
        REG_FILE_reg_out_6__25_), .ZN(n3940) );
  AOI22_X2 U2039 ( .A1(n7763), .A2(REG_FILE_reg_out_0__25_), .B1(n7577), .B2(
        REG_FILE_reg_out_4__25_), .ZN(n3939) );
  OAI221_X2 U2041 ( .B1(n6161), .B2(n7568), .C1(n7020), .C2(n7560), .A(n3945), 
        .ZN(n3944) );
  AOI22_X2 U2042 ( .A1(n7763), .A2(REG_FILE_reg_out_8__25_), .B1(n7581), .B2(
        REG_FILE_reg_out_12__25_), .ZN(n3945) );
  OAI221_X2 U2043 ( .B1(n6412), .B2(n7587), .C1(n6064), .C2(n7597), .A(n3946), 
        .ZN(n3943) );
  AOI22_X2 U2044 ( .A1(n7608), .A2(REG_FILE_reg_out_11__25_), .B1(n7600), .B2(
        REG_FILE_reg_out_15__25_), .ZN(n3946) );
  OAI221_X2 U2046 ( .B1(n5963), .B2(n7571), .C1(n7019), .C2(n7560), .A(n3949), 
        .ZN(n3948) );
  AOI22_X2 U2047 ( .A1(n7763), .A2(REG_FILE_reg_out_24__25_), .B1(n7581), .B2(
        REG_FILE_reg_out_28__25_), .ZN(n3949) );
  OAI221_X2 U2048 ( .B1(n6103), .B2(n7587), .C1(n5895), .C2(n7597), .A(n3950), 
        .ZN(n3947) );
  AOI22_X2 U2049 ( .A1(n7611), .A2(REG_FILE_reg_out_27__25_), .B1(n7605), .B2(
        REG_FILE_reg_out_31__25_), .ZN(n3950) );
  OAI221_X2 U2051 ( .B1(n6963), .B2(n7568), .C1(n6381), .C2(n7560), .A(n3953), 
        .ZN(n3952) );
  AOI22_X2 U2052 ( .A1(n7763), .A2(REG_FILE_reg_out_16__25_), .B1(n7579), .B2(
        REG_FILE_reg_out_20__25_), .ZN(n3953) );
  OAI221_X2 U2053 ( .B1(n6054), .B2(n7587), .C1(n6380), .C2(n7597), .A(n3954), 
        .ZN(n3951) );
  AOI22_X2 U2054 ( .A1(n7611), .A2(REG_FILE_reg_out_19__25_), .B1(n7605), .B2(
        REG_FILE_reg_out_23__25_), .ZN(n3954) );
  AOI221_X2 U2058 ( .B1(n7606), .B2(REG_FILE_reg_out_3__26_), .C1(n7600), .C2(
        REG_FILE_reg_out_7__26_), .A(n3963), .ZN(n3962) );
  OAI22_X2 U2059 ( .A1(n6451), .A2(n7598), .B1(n6981), .B2(n7589), .ZN(n3963)
         );
  AOI22_X2 U2060 ( .A1(n7573), .A2(REG_FILE_reg_out_2__26_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__26_), .ZN(n3961) );
  AOI22_X2 U2061 ( .A1(n7763), .A2(REG_FILE_reg_out_0__26_), .B1(n7578), .B2(
        REG_FILE_reg_out_4__26_), .ZN(n3960) );
  OAI221_X2 U2063 ( .B1(n6495), .B2(n7571), .C1(n7018), .C2(n7560), .A(n3966), 
        .ZN(n3965) );
  AOI22_X2 U2064 ( .A1(n7763), .A2(REG_FILE_reg_out_8__26_), .B1(n7579), .B2(
        REG_FILE_reg_out_12__26_), .ZN(n3966) );
  OAI221_X2 U2065 ( .B1(n6411), .B2(n7587), .C1(n6063), .C2(n7597), .A(n3967), 
        .ZN(n3964) );
  AOI22_X2 U2066 ( .A1(n7611), .A2(REG_FILE_reg_out_11__26_), .B1(n7604), .B2(
        REG_FILE_reg_out_15__26_), .ZN(n3967) );
  OAI221_X2 U2068 ( .B1(n6160), .B2(n7570), .C1(n7017), .C2(n7560), .A(n3970), 
        .ZN(n3969) );
  AOI22_X2 U2069 ( .A1(n7763), .A2(REG_FILE_reg_out_24__26_), .B1(n7578), .B2(
        REG_FILE_reg_out_28__26_), .ZN(n3970) );
  OAI221_X2 U2070 ( .B1(n5896), .B2(n7587), .C1(n5875), .C2(n7597), .A(n3971), 
        .ZN(n3968) );
  AOI22_X2 U2071 ( .A1(n7611), .A2(REG_FILE_reg_out_27__26_), .B1(n7604), .B2(
        REG_FILE_reg_out_31__26_), .ZN(n3971) );
  OAI221_X2 U2073 ( .B1(n6410), .B2(n7571), .C1(n6926), .C2(n7560), .A(n3974), 
        .ZN(n3973) );
  AOI22_X2 U2074 ( .A1(n7764), .A2(REG_FILE_reg_out_16__26_), .B1(n7578), .B2(
        REG_FILE_reg_out_20__26_), .ZN(n3974) );
  OAI221_X2 U2075 ( .B1(n5933), .B2(n7587), .C1(n6925), .C2(n7597), .A(n3975), 
        .ZN(n3972) );
  AOI22_X2 U2076 ( .A1(n7611), .A2(REG_FILE_reg_out_19__26_), .B1(n7604), .B2(
        REG_FILE_reg_out_23__26_), .ZN(n3975) );
  AOI221_X2 U2080 ( .B1(n7606), .B2(REG_FILE_reg_out_3__27_), .C1(n7601), .C2(
        REG_FILE_reg_out_7__27_), .A(n3984), .ZN(n3983) );
  OAI22_X2 U2081 ( .A1(n5949), .A2(n7591), .B1(n6131), .B2(n7589), .ZN(n3984)
         );
  AOI22_X2 U2082 ( .A1(n7573), .A2(REG_FILE_reg_out_2__27_), .B1(n7566), .B2(
        REG_FILE_reg_out_6__27_), .ZN(n3982) );
  AOI22_X2 U2083 ( .A1(n7770), .A2(REG_FILE_reg_out_0__27_), .B1(n7578), .B2(
        REG_FILE_reg_out_4__27_), .ZN(n3981) );
  OAI221_X2 U2085 ( .B1(n6494), .B2(n7570), .C1(n7016), .C2(n7560), .A(n3987), 
        .ZN(n3986) );
  AOI22_X2 U2086 ( .A1(n7764), .A2(REG_FILE_reg_out_8__27_), .B1(n7578), .B2(
        REG_FILE_reg_out_12__27_), .ZN(n3987) );
  OAI221_X2 U2087 ( .B1(n5947), .B2(n7587), .C1(n6924), .C2(n7597), .A(n3988), 
        .ZN(n3985) );
  AOI22_X2 U2088 ( .A1(n7610), .A2(REG_FILE_reg_out_11__27_), .B1(n7600), .B2(
        REG_FILE_reg_out_15__27_), .ZN(n3988) );
  OAI221_X2 U2090 ( .B1(n6159), .B2(n7568), .C1(n6508), .C2(n7560), .A(n3991), 
        .ZN(n3990) );
  AOI22_X2 U2091 ( .A1(n7763), .A2(REG_FILE_reg_out_24__27_), .B1(n7578), .B2(
        REG_FILE_reg_out_28__27_), .ZN(n3991) );
  OAI221_X2 U2092 ( .B1(n5946), .B2(n7587), .C1(n5874), .C2(n7596), .A(n3992), 
        .ZN(n3989) );
  AOI22_X2 U2093 ( .A1(n7610), .A2(REG_FILE_reg_out_27__27_), .B1(n7604), .B2(
        REG_FILE_reg_out_31__27_), .ZN(n3992) );
  OAI221_X2 U2095 ( .B1(n6409), .B2(n7570), .C1(n6923), .C2(n7560), .A(n3995), 
        .ZN(n3994) );
  AOI22_X2 U2096 ( .A1(n7764), .A2(REG_FILE_reg_out_16__27_), .B1(n7578), .B2(
        REG_FILE_reg_out_20__27_), .ZN(n3995) );
  OAI221_X2 U2097 ( .B1(n6962), .B2(n7587), .C1(n5935), .C2(n7597), .A(n3996), 
        .ZN(n3993) );
  AOI22_X2 U2098 ( .A1(n7609), .A2(REG_FILE_reg_out_19__27_), .B1(n7602), .B2(
        REG_FILE_reg_out_23__27_), .ZN(n3996) );
  AOI221_X2 U2102 ( .B1(n7606), .B2(REG_FILE_reg_out_3__28_), .C1(n7601), .C2(
        REG_FILE_reg_out_7__28_), .A(n4005), .ZN(n4004) );
  OAI22_X2 U2103 ( .A1(n5882), .A2(n7591), .B1(n6124), .B2(n7589), .ZN(n4005)
         );
  AOI22_X2 U2104 ( .A1(n7573), .A2(REG_FILE_reg_out_2__28_), .B1(n7565), .B2(
        REG_FILE_reg_out_6__28_), .ZN(n4003) );
  AOI22_X2 U2105 ( .A1(n7763), .A2(REG_FILE_reg_out_0__28_), .B1(n7578), .B2(
        REG_FILE_reg_out_4__28_), .ZN(n4002) );
  OAI221_X2 U2107 ( .B1(n7006), .B2(n7568), .C1(n6507), .C2(n7560), .A(n4008), 
        .ZN(n4007) );
  AOI22_X2 U2108 ( .A1(n7764), .A2(REG_FILE_reg_out_8__28_), .B1(n7578), .B2(
        REG_FILE_reg_out_12__28_), .ZN(n4008) );
  OAI221_X2 U2109 ( .B1(n6961), .B2(n7587), .C1(n5873), .C2(n7597), .A(n4009), 
        .ZN(n4006) );
  AOI22_X2 U2110 ( .A1(n7609), .A2(REG_FILE_reg_out_11__28_), .B1(n7603), .B2(
        REG_FILE_reg_out_15__28_), .ZN(n4009) );
  OAI221_X2 U2112 ( .B1(n6493), .B2(n7569), .C1(n7015), .C2(n7559), .A(n4012), 
        .ZN(n4011) );
  AOI22_X2 U2113 ( .A1(n7764), .A2(REG_FILE_reg_out_24__28_), .B1(n7578), .B2(
        REG_FILE_reg_out_28__28_), .ZN(n4012) );
  OAI221_X2 U2114 ( .B1(n6960), .B2(n7587), .C1(n5934), .C2(n7594), .A(n4013), 
        .ZN(n4010) );
  AOI22_X2 U2115 ( .A1(n7609), .A2(REG_FILE_reg_out_27__28_), .B1(n7603), .B2(
        REG_FILE_reg_out_31__28_), .ZN(n4013) );
  OAI221_X2 U2117 ( .B1(n6959), .B2(n7569), .C1(n6379), .C2(n7559), .A(n4016), 
        .ZN(n4015) );
  AOI22_X2 U2118 ( .A1(n7764), .A2(REG_FILE_reg_out_16__28_), .B1(n7578), .B2(
        REG_FILE_reg_out_20__28_), .ZN(n4016) );
  OAI221_X2 U2119 ( .B1(n6920), .B2(n7587), .C1(n5872), .C2(n7597), .A(n4017), 
        .ZN(n4014) );
  AOI22_X2 U2120 ( .A1(n7609), .A2(REG_FILE_reg_out_19__28_), .B1(n7602), .B2(
        REG_FILE_reg_out_23__28_), .ZN(n4017) );
  AOI221_X2 U2124 ( .B1(n7606), .B2(REG_FILE_reg_out_3__29_), .C1(n7601), .C2(
        REG_FILE_reg_out_7__29_), .A(n4026), .ZN(n4025) );
  OAI22_X2 U2125 ( .A1(n5899), .A2(n7591), .B1(n6123), .B2(n7589), .ZN(n4026)
         );
  AOI22_X2 U2126 ( .A1(n7573), .A2(REG_FILE_reg_out_2__29_), .B1(n7565), .B2(
        REG_FILE_reg_out_6__29_), .ZN(n4024) );
  AOI22_X2 U2127 ( .A1(n7767), .A2(REG_FILE_reg_out_0__29_), .B1(n7578), .B2(
        REG_FILE_reg_out_4__29_), .ZN(n4023) );
  OAI221_X2 U2129 ( .B1(n7005), .B2(n7569), .C1(n6506), .C2(n7559), .A(n4029), 
        .ZN(n4028) );
  AOI22_X2 U2130 ( .A1(n7764), .A2(REG_FILE_reg_out_8__29_), .B1(n7577), .B2(
        REG_FILE_reg_out_12__29_), .ZN(n4029) );
  OAI221_X2 U2131 ( .B1(n6958), .B2(n7587), .C1(n5871), .C2(n7594), .A(n4030), 
        .ZN(n4027) );
  AOI22_X2 U2132 ( .A1(n7609), .A2(REG_FILE_reg_out_11__29_), .B1(n7602), .B2(
        REG_FILE_reg_out_15__29_), .ZN(n4030) );
  OAI221_X2 U2134 ( .B1(n6492), .B2(n7571), .C1(n7014), .C2(n7559), .A(n4033), 
        .ZN(n4032) );
  AOI22_X2 U2135 ( .A1(n7764), .A2(REG_FILE_reg_out_24__29_), .B1(n7577), .B2(
        REG_FILE_reg_out_28__29_), .ZN(n4033) );
  OAI221_X2 U2136 ( .B1(n6957), .B2(n7587), .C1(n6378), .C2(n7597), .A(n4034), 
        .ZN(n4031) );
  AOI22_X2 U2137 ( .A1(n7608), .A2(REG_FILE_reg_out_27__29_), .B1(n7603), .B2(
        REG_FILE_reg_out_31__29_), .ZN(n4034) );
  OAI221_X2 U2139 ( .B1(n6956), .B2(n7569), .C1(n6377), .C2(n7559), .A(n4037), 
        .ZN(n4036) );
  AOI22_X2 U2140 ( .A1(n7764), .A2(REG_FILE_reg_out_16__29_), .B1(n7577), .B2(
        REG_FILE_reg_out_20__29_), .ZN(n4037) );
  OAI221_X2 U2141 ( .B1(n6919), .B2(n7587), .C1(n6376), .C2(n7597), .A(n4038), 
        .ZN(n4035) );
  AOI22_X2 U2142 ( .A1(n7608), .A2(REG_FILE_reg_out_19__29_), .B1(n7602), .B2(
        REG_FILE_reg_out_23__29_), .ZN(n4038) );
  AOI221_X2 U2146 ( .B1(n7606), .B2(REG_FILE_reg_out_3__30_), .C1(n7601), .C2(
        REG_FILE_reg_out_7__30_), .A(n4047), .ZN(n4046) );
  OAI22_X2 U2147 ( .A1(n5898), .A2(n7591), .B1(n6130), .B2(n7589), .ZN(n4047)
         );
  AOI22_X2 U2148 ( .A1(n7573), .A2(REG_FILE_reg_out_2__30_), .B1(n6009), .B2(
        REG_FILE_reg_out_6__30_), .ZN(n4045) );
  AOI22_X2 U2149 ( .A1(n7764), .A2(REG_FILE_reg_out_0__30_), .B1(n7577), .B2(
        REG_FILE_reg_out_4__30_), .ZN(n4044) );
  OAI221_X2 U2151 ( .B1(n7004), .B2(n7571), .C1(n6505), .C2(n7559), .A(n4050), 
        .ZN(n4049) );
  AOI22_X2 U2152 ( .A1(n7764), .A2(REG_FILE_reg_out_8__30_), .B1(n7577), .B2(
        REG_FILE_reg_out_12__30_), .ZN(n4050) );
  OAI221_X2 U2153 ( .B1(n6955), .B2(n7587), .C1(n6375), .C2(n7597), .A(n4051), 
        .ZN(n4048) );
  AOI22_X2 U2154 ( .A1(n7607), .A2(REG_FILE_reg_out_11__30_), .B1(n7601), .B2(
        REG_FILE_reg_out_15__30_), .ZN(n4051) );
  OAI221_X2 U2156 ( .B1(n6491), .B2(n7570), .C1(n7013), .C2(n7559), .A(n4054), 
        .ZN(n4053) );
  AOI22_X2 U2157 ( .A1(n7764), .A2(REG_FILE_reg_out_24__30_), .B1(n7577), .B2(
        REG_FILE_reg_out_28__30_), .ZN(n4054) );
  OAI221_X2 U2158 ( .B1(n6954), .B2(n7587), .C1(n6374), .C2(n7597), .A(n4055), 
        .ZN(n4052) );
  AOI22_X2 U2159 ( .A1(n7608), .A2(REG_FILE_reg_out_27__30_), .B1(n7603), .B2(
        REG_FILE_reg_out_31__30_), .ZN(n4055) );
  OAI221_X2 U2161 ( .B1(n6953), .B2(n7569), .C1(n6373), .C2(n7559), .A(n4058), 
        .ZN(n4057) );
  AOI22_X2 U2162 ( .A1(n7764), .A2(REG_FILE_reg_out_16__30_), .B1(n7577), .B2(
        REG_FILE_reg_out_20__30_), .ZN(n4058) );
  OAI221_X2 U2163 ( .B1(n6408), .B2(n7587), .C1(n6062), .C2(n7597), .A(n4059), 
        .ZN(n4056) );
  AOI22_X2 U2164 ( .A1(n7607), .A2(REG_FILE_reg_out_19__30_), .B1(n7601), .B2(
        REG_FILE_reg_out_23__30_), .ZN(n4059) );
  AOI221_X2 U2168 ( .B1(n7606), .B2(REG_FILE_reg_out_3__31_), .C1(n7601), .C2(
        REG_FILE_reg_out_7__31_), .A(n4068), .ZN(n4067) );
  OAI22_X2 U2169 ( .A1(n6118), .A2(n7596), .B1(n6468), .B2(n7588), .ZN(n4068)
         );
  AOI22_X2 U2170 ( .A1(n7573), .A2(REG_FILE_reg_out_2__31_), .B1(n7566), .B2(
        REG_FILE_reg_out_6__31_), .ZN(n4066) );
  AOI22_X2 U2171 ( .A1(n7764), .A2(REG_FILE_reg_out_0__31_), .B1(n7577), .B2(
        REG_FILE_reg_out_4__31_), .ZN(n4065) );
  AND3_X2 U2172 ( .A1(n7774), .A2(n6016), .A3(n4069), .ZN(n3390) );
  OAI221_X2 U2177 ( .B1(n7003), .B2(n7570), .C1(n6504), .C2(n7559), .A(n4073), 
        .ZN(n4072) );
  AOI22_X2 U2178 ( .A1(n7764), .A2(REG_FILE_reg_out_8__31_), .B1(n7577), .B2(
        REG_FILE_reg_out_12__31_), .ZN(n4073) );
  OAI221_X2 U2179 ( .B1(n6407), .B2(n7587), .C1(n6061), .C2(n7597), .A(n4074), 
        .ZN(n4071) );
  AOI22_X2 U2180 ( .A1(n7607), .A2(REG_FILE_reg_out_11__31_), .B1(n7600), .B2(
        REG_FILE_reg_out_15__31_), .ZN(n4074) );
  OAI221_X2 U2183 ( .B1(n7002), .B2(n7569), .C1(n6503), .C2(n7559), .A(n4078), 
        .ZN(n4076) );
  AOI22_X2 U2184 ( .A1(n7764), .A2(REG_FILE_reg_out_24__31_), .B1(n7577), .B2(
        REG_FILE_reg_out_28__31_), .ZN(n4078) );
  OAI221_X2 U2185 ( .B1(n6952), .B2(n7587), .C1(n6372), .C2(n7597), .A(n4079), 
        .ZN(n4075) );
  AOI22_X2 U2186 ( .A1(n7606), .A2(REG_FILE_reg_out_27__31_), .B1(n7600), .B2(
        REG_FILE_reg_out_31__31_), .ZN(n4079) );
  XOR2_X2 U2196 ( .A(n7321), .B(n5857), .Z(n4082) );
  OAI221_X2 U2197 ( .B1(n6951), .B2(n7569), .C1(n6371), .C2(n7559), .A(n4088), 
        .ZN(n4081) );
  AOI22_X2 U2198 ( .A1(n7764), .A2(REG_FILE_reg_out_16__31_), .B1(n7577), .B2(
        REG_FILE_reg_out_20__31_), .ZN(n4088) );
  NAND2_X2 U2201 ( .A1(n4091), .A2(n5857), .ZN(n3405) );
  OAI221_X2 U2203 ( .B1(n6406), .B2(n7584), .C1(n6060), .C2(n7592), .A(n4092), 
        .ZN(n4080) );
  AOI22_X2 U2204 ( .A1(n7609), .A2(REG_FILE_reg_out_19__31_), .B1(n7602), .B2(
        REG_FILE_reg_out_23__31_), .ZN(n4092) );
  NAND2_X2 U2209 ( .A1(n4094), .A2(n5857), .ZN(n3399) );
  AOI221_X2 U2215 ( .B1(n7485), .B2(REG_FILE_reg_out_11__0_), .C1(n7500), .C2(
        REG_FILE_reg_out_15__0_), .A(n4108), .ZN(n4106) );
  OAI22_X2 U2216 ( .A1(n5890), .A2(n7545), .B1(n6101), .B2(n7536), .ZN(n4108)
         );
  AOI221_X2 U2217 ( .B1(n7501), .B2(REG_FILE_reg_out_10__0_), .C1(n7516), .C2(
        REG_FILE_reg_out_14__0_), .A(n4111), .ZN(n4105) );
  OAI22_X2 U2218 ( .A1(n6530), .A2(n7527), .B1(n6257), .B2(n7521), .ZN(n4111)
         );
  AOI221_X2 U2220 ( .B1(n7485), .B2(REG_FILE_reg_out_27__0_), .C1(n7500), .C2(
        REG_FILE_reg_out_31__0_), .A(n4117), .ZN(n4115) );
  OAI22_X2 U2221 ( .A1(n5893), .A2(n7545), .B1(n5945), .B2(n7542), .ZN(n4117)
         );
  AOI221_X2 U2222 ( .B1(n7501), .B2(REG_FILE_reg_out_26__0_), .C1(n7516), .C2(
        REG_FILE_reg_out_30__0_), .A(n4118), .ZN(n4114) );
  OAI22_X2 U2223 ( .A1(n5902), .A2(n7527), .B1(n5996), .B2(n7525), .ZN(n4118)
         );
  AOI221_X2 U2225 ( .B1(n7485), .B2(REG_FILE_reg_out_3__0_), .C1(n7498), .C2(
        REG_FILE_reg_out_7__0_), .A(n4122), .ZN(n4120) );
  OAI22_X2 U2226 ( .A1(n5897), .A2(n7545), .B1(n5954), .B2(n7537), .ZN(n4122)
         );
  AOI221_X2 U2227 ( .B1(n7501), .B2(REG_FILE_reg_out_2__0_), .C1(n7516), .C2(
        REG_FILE_reg_out_6__0_), .A(n4123), .ZN(n4119) );
  OAI22_X2 U2228 ( .A1(n5979), .A2(n7527), .B1(n6623), .B2(n7523), .ZN(n4123)
         );
  NOR4_X2 U2229 ( .A1(n4124), .A2(n4125), .A3(n4126), .A4(n4127), .ZN(n4098)
         );
  OAI22_X2 U2230 ( .A1(n5973), .A2(n7533), .B1(n6631), .B2(n7523), .ZN(n4127)
         );
  OAI22_X2 U2231 ( .A1(n6363), .A2(n4128), .B1(n6086), .B2(n7508), .ZN(n4126)
         );
  OAI22_X2 U2232 ( .A1(n5892), .A2(n7546), .B1(n5944), .B2(n7543), .ZN(n4125)
         );
  OAI22_X2 U2233 ( .A1(n6538), .A2(n4130), .B1(n6245), .B2(n7492), .ZN(n4124)
         );
  AOI221_X2 U2238 ( .B1(n7485), .B2(REG_FILE_reg_out_11__1_), .C1(n7500), .C2(
        REG_FILE_reg_out_15__1_), .A(n4140), .ZN(n4139) );
  OAI22_X2 U2239 ( .A1(n5891), .A2(n7545), .B1(n6102), .B2(n7536), .ZN(n4140)
         );
  AOI221_X2 U2240 ( .B1(n7501), .B2(REG_FILE_reg_out_10__1_), .C1(n7516), .C2(
        REG_FILE_reg_out_14__1_), .A(n4141), .ZN(n4138) );
  OAI22_X2 U2241 ( .A1(n6531), .A2(n7527), .B1(n6000), .B2(n7524), .ZN(n4141)
         );
  AOI221_X2 U2243 ( .B1(n7485), .B2(REG_FILE_reg_out_27__1_), .C1(n7500), .C2(
        REG_FILE_reg_out_31__1_), .A(n4144), .ZN(n4143) );
  OAI22_X2 U2244 ( .A1(n5927), .A2(n7545), .B1(n6094), .B2(n7541), .ZN(n4144)
         );
  AOI221_X2 U2245 ( .B1(n7501), .B2(REG_FILE_reg_out_26__1_), .C1(n7516), .C2(
        REG_FILE_reg_out_30__1_), .A(n4145), .ZN(n4142) );
  OAI22_X2 U2246 ( .A1(n5903), .A2(n7527), .B1(n5997), .B2(n7525), .ZN(n4145)
         );
  AOI221_X2 U2248 ( .B1(n7485), .B2(REG_FILE_reg_out_3__1_), .C1(n7500), .C2(
        REG_FILE_reg_out_7__1_), .A(n4148), .ZN(n4147) );
  OAI22_X2 U2249 ( .A1(n5880), .A2(n7545), .B1(n6128), .B2(n7544), .ZN(n4148)
         );
  AOI221_X2 U2250 ( .B1(n7501), .B2(REG_FILE_reg_out_2__1_), .C1(n7514), .C2(
        REG_FILE_reg_out_6__1_), .A(n4149), .ZN(n4146) );
  OAI22_X2 U2251 ( .A1(n5980), .A2(n7527), .B1(n6624), .B2(n7523), .ZN(n4149)
         );
  NOR4_X2 U2252 ( .A1(n4150), .A2(n4151), .A3(n4152), .A4(n4153), .ZN(n4133)
         );
  OAI22_X2 U2253 ( .A1(n5900), .A2(n7531), .B1(n6632), .B2(n7524), .ZN(n4153)
         );
  OAI22_X2 U2254 ( .A1(n6364), .A2(n4128), .B1(n6087), .B2(n7508), .ZN(n4152)
         );
  OAI22_X2 U2255 ( .A1(n6048), .A2(n7548), .B1(n6399), .B2(n7537), .ZN(n4151)
         );
  OAI22_X2 U2256 ( .A1(n6539), .A2(n4130), .B1(n6246), .B2(n7492), .ZN(n4150)
         );
  AOI221_X2 U2261 ( .B1(n7485), .B2(REG_FILE_reg_out_11__2_), .C1(n7500), .C2(
        REG_FILE_reg_out_15__2_), .A(n4163), .ZN(n4162) );
  OAI22_X2 U2262 ( .A1(n6358), .A2(n7552), .B1(n6946), .B2(n7536), .ZN(n4163)
         );
  AOI221_X2 U2263 ( .B1(n7501), .B2(REG_FILE_reg_out_10__2_), .C1(n7516), .C2(
        REG_FILE_reg_out_14__2_), .A(n4164), .ZN(n4161) );
  OAI22_X2 U2264 ( .A1(n6532), .A2(n7534), .B1(n6001), .B2(n7525), .ZN(n4164)
         );
  AOI221_X2 U2266 ( .B1(n7485), .B2(REG_FILE_reg_out_27__2_), .C1(n7500), .C2(
        REG_FILE_reg_out_31__2_), .A(n4167), .ZN(n4166) );
  OAI22_X2 U2267 ( .A1(n5894), .A2(n7552), .B1(n6095), .B2(n7537), .ZN(n4167)
         );
  AOI221_X2 U2268 ( .B1(n7501), .B2(REG_FILE_reg_out_26__2_), .C1(n7516), .C2(
        REG_FILE_reg_out_30__2_), .A(n4168), .ZN(n4165) );
  OAI22_X2 U2269 ( .A1(n5904), .A2(n7534), .B1(n5998), .B2(n7525), .ZN(n4168)
         );
  AOI221_X2 U2271 ( .B1(n7490), .B2(REG_FILE_reg_out_3__2_), .C1(n7494), .C2(
        REG_FILE_reg_out_7__2_), .A(n4171), .ZN(n4170) );
  OAI22_X2 U2272 ( .A1(n6113), .A2(n7546), .B1(n6462), .B2(n7536), .ZN(n4171)
         );
  AOI221_X2 U2273 ( .B1(n7506), .B2(REG_FILE_reg_out_2__2_), .C1(n7510), .C2(
        REG_FILE_reg_out_6__2_), .A(n4172), .ZN(n4169) );
  OAI22_X2 U2274 ( .A1(n5981), .A2(n7534), .B1(n6625), .B2(n7523), .ZN(n4172)
         );
  NOR4_X2 U2275 ( .A1(n4173), .A2(n4174), .A3(n4175), .A4(n4176), .ZN(n4155)
         );
  OAI22_X2 U2276 ( .A1(n5974), .A2(n7531), .B1(n6633), .B2(n7525), .ZN(n4176)
         );
  OAI22_X2 U2277 ( .A1(n6365), .A2(n4128), .B1(n6088), .B2(n7508), .ZN(n4175)
         );
  OAI22_X2 U2278 ( .A1(n6049), .A2(n7548), .B1(n6400), .B2(n7536), .ZN(n4174)
         );
  OAI22_X2 U2279 ( .A1(n6540), .A2(n4130), .B1(n6247), .B2(n7492), .ZN(n4173)
         );
  AOI221_X2 U2287 ( .B1(n7493), .B2(REG_FILE_reg_out_11__3_), .C1(n7494), .C2(
        REG_FILE_reg_out_15__3_), .A(n4185), .ZN(n4184) );
  OAI22_X2 U2288 ( .A1(n6359), .A2(n7552), .B1(n6947), .B2(n7536), .ZN(n4185)
         );
  AOI221_X2 U2289 ( .B1(n7509), .B2(REG_FILE_reg_out_10__3_), .C1(n7510), .C2(
        REG_FILE_reg_out_14__3_), .A(n4186), .ZN(n4183) );
  OAI22_X2 U2290 ( .A1(n6533), .A2(n7534), .B1(n6002), .B2(n7525), .ZN(n4186)
         );
  AOI221_X2 U2292 ( .B1(n7493), .B2(REG_FILE_reg_out_27__3_), .C1(n7494), .C2(
        REG_FILE_reg_out_31__3_), .A(n4189), .ZN(n4188) );
  OAI22_X2 U2293 ( .A1(n5928), .A2(n7545), .B1(n6096), .B2(n7536), .ZN(n4189)
         );
  AOI221_X2 U2294 ( .B1(n7509), .B2(REG_FILE_reg_out_26__3_), .C1(n7510), .C2(
        REG_FILE_reg_out_30__3_), .A(n4190), .ZN(n4187) );
  OAI22_X2 U2295 ( .A1(n5905), .A2(n7534), .B1(n5999), .B2(n7524), .ZN(n4190)
         );
  AOI221_X2 U2297 ( .B1(n7493), .B2(REG_FILE_reg_out_3__3_), .C1(n7494), .C2(
        REG_FILE_reg_out_7__3_), .A(n4193), .ZN(n4192) );
  OAI22_X2 U2298 ( .A1(n6114), .A2(n7546), .B1(n6463), .B2(n7536), .ZN(n4193)
         );
  AOI221_X2 U2299 ( .B1(n7509), .B2(REG_FILE_reg_out_2__3_), .C1(n7510), .C2(
        REG_FILE_reg_out_6__3_), .A(n4194), .ZN(n4191) );
  OAI22_X2 U2300 ( .A1(n5982), .A2(n7534), .B1(n6626), .B2(n7523), .ZN(n4194)
         );
  NOR4_X2 U2301 ( .A1(n4195), .A2(n4196), .A3(n4197), .A4(n4198), .ZN(n4178)
         );
  OAI22_X2 U2302 ( .A1(n5901), .A2(n7528), .B1(n6634), .B2(n7523), .ZN(n4198)
         );
  OAI22_X2 U2303 ( .A1(n6366), .A2(n4128), .B1(n6089), .B2(n7508), .ZN(n4197)
         );
  OAI22_X2 U2304 ( .A1(n6050), .A2(n7547), .B1(n6401), .B2(n4110), .ZN(n4196)
         );
  OAI22_X2 U2305 ( .A1(n6541), .A2(n4130), .B1(n6248), .B2(n7492), .ZN(n4195)
         );
  AOI221_X2 U2310 ( .B1(n7493), .B2(REG_FILE_reg_out_11__4_), .C1(n7494), .C2(
        REG_FILE_reg_out_15__4_), .A(n4208), .ZN(n4207) );
  OAI22_X2 U2311 ( .A1(n6047), .A2(n7552), .B1(n6405), .B2(n7536), .ZN(n4208)
         );
  AOI221_X2 U2312 ( .B1(n7509), .B2(REG_FILE_reg_out_10__4_), .C1(n7510), .C2(
        REG_FILE_reg_out_14__4_), .A(n4209), .ZN(n4206) );
  OAI22_X2 U2313 ( .A1(n6534), .A2(n7534), .B1(n6258), .B2(n7521), .ZN(n4209)
         );
  AOI221_X2 U2315 ( .B1(n7493), .B2(REG_FILE_reg_out_27__4_), .C1(n7494), .C2(
        REG_FILE_reg_out_31__4_), .A(n4212), .ZN(n4211) );
  OAI22_X2 U2316 ( .A1(n5929), .A2(n7552), .B1(n6097), .B2(n7537), .ZN(n4212)
         );
  AOI221_X2 U2317 ( .B1(n7509), .B2(REG_FILE_reg_out_26__4_), .C1(n7510), .C2(
        REG_FILE_reg_out_30__4_), .A(n4213), .ZN(n4210) );
  OAI22_X2 U2318 ( .A1(n5975), .A2(n7534), .B1(n6253), .B2(n7521), .ZN(n4213)
         );
  AOI221_X2 U2320 ( .B1(n7490), .B2(REG_FILE_reg_out_3__4_), .C1(n7494), .C2(
        REG_FILE_reg_out_7__4_), .A(n4216), .ZN(n4215) );
  OAI22_X2 U2321 ( .A1(n6115), .A2(n7552), .B1(n6464), .B2(n7544), .ZN(n4216)
         );
  AOI221_X2 U2322 ( .B1(n7509), .B2(REG_FILE_reg_out_2__4_), .C1(n7510), .C2(
        REG_FILE_reg_out_6__4_), .A(n4217), .ZN(n4214) );
  OAI22_X2 U2323 ( .A1(n6197), .A2(n7534), .B1(n6627), .B2(n7521), .ZN(n4217)
         );
  NOR4_X2 U2324 ( .A1(n4218), .A2(n4219), .A3(n4220), .A4(n4221), .ZN(n4200)
         );
  OAI22_X2 U2325 ( .A1(n6193), .A2(n7534), .B1(n6635), .B2(n7521), .ZN(n4221)
         );
  OAI22_X2 U2326 ( .A1(n6367), .A2(n4128), .B1(n6090), .B2(n7508), .ZN(n4220)
         );
  OAI22_X2 U2327 ( .A1(n6051), .A2(n7552), .B1(n6402), .B2(n7544), .ZN(n4219)
         );
  OAI22_X2 U2328 ( .A1(n6542), .A2(n4130), .B1(n6249), .B2(n7492), .ZN(n4218)
         );
  AOI221_X2 U2333 ( .B1(n7493), .B2(REG_FILE_reg_out_11__5_), .C1(n7494), .C2(
        REG_FILE_reg_out_15__5_), .A(n4230), .ZN(n4229) );
  OAI22_X2 U2334 ( .A1(n6360), .A2(n7552), .B1(n6948), .B2(n7544), .ZN(n4230)
         );
  AOI221_X2 U2335 ( .B1(n7509), .B2(REG_FILE_reg_out_10__5_), .C1(n7510), .C2(
        REG_FILE_reg_out_14__5_), .A(n4231), .ZN(n4228) );
  OAI22_X2 U2336 ( .A1(n6535), .A2(n7534), .B1(n6259), .B2(n7521), .ZN(n4231)
         );
  AOI221_X2 U2338 ( .B1(n7493), .B2(REG_FILE_reg_out_27__5_), .C1(n7494), .C2(
        REG_FILE_reg_out_31__5_), .A(n4234), .ZN(n4233) );
  OAI22_X2 U2339 ( .A1(n5930), .A2(n7552), .B1(n6098), .B2(n7544), .ZN(n4234)
         );
  AOI221_X2 U2340 ( .B1(n7509), .B2(REG_FILE_reg_out_26__5_), .C1(n7510), .C2(
        REG_FILE_reg_out_30__5_), .A(n4235), .ZN(n4232) );
  OAI22_X2 U2341 ( .A1(n5976), .A2(n7534), .B1(n6254), .B2(n7521), .ZN(n4235)
         );
  AOI221_X2 U2343 ( .B1(n7493), .B2(REG_FILE_reg_out_3__5_), .C1(n7494), .C2(
        REG_FILE_reg_out_7__5_), .A(n4238), .ZN(n4237) );
  OAI22_X2 U2344 ( .A1(n6116), .A2(n7552), .B1(n6465), .B2(n7544), .ZN(n4238)
         );
  AOI221_X2 U2345 ( .B1(n7506), .B2(REG_FILE_reg_out_2__5_), .C1(n7510), .C2(
        REG_FILE_reg_out_6__5_), .A(n4239), .ZN(n4236) );
  OAI22_X2 U2346 ( .A1(n5983), .A2(n7534), .B1(n6628), .B2(n7521), .ZN(n4239)
         );
  NOR4_X2 U2347 ( .A1(n4240), .A2(n4241), .A3(n4242), .A4(n4243), .ZN(n4223)
         );
  OAI22_X2 U2348 ( .A1(n6194), .A2(n7534), .B1(n6636), .B2(n7521), .ZN(n4243)
         );
  OAI22_X2 U2349 ( .A1(n6368), .A2(n4128), .B1(n6091), .B2(n7508), .ZN(n4242)
         );
  OAI22_X2 U2350 ( .A1(n6052), .A2(n7552), .B1(n6403), .B2(n7544), .ZN(n4241)
         );
  OAI22_X2 U2351 ( .A1(n6543), .A2(n4130), .B1(n6250), .B2(n7492), .ZN(n4240)
         );
  AOI221_X2 U2356 ( .B1(n7489), .B2(REG_FILE_reg_out_11__6_), .C1(n7495), .C2(
        REG_FILE_reg_out_15__6_), .A(n4253), .ZN(n4252) );
  OAI22_X2 U2357 ( .A1(n6361), .A2(n7552), .B1(n6949), .B2(n7544), .ZN(n4253)
         );
  AOI221_X2 U2358 ( .B1(n7505), .B2(REG_FILE_reg_out_10__6_), .C1(n7513), .C2(
        REG_FILE_reg_out_14__6_), .A(n4254), .ZN(n4251) );
  OAI22_X2 U2359 ( .A1(n6536), .A2(n7534), .B1(n6260), .B2(n7521), .ZN(n4254)
         );
  AOI221_X2 U2361 ( .B1(n7490), .B2(REG_FILE_reg_out_27__6_), .C1(n7498), .C2(
        REG_FILE_reg_out_31__6_), .A(n4257), .ZN(n4256) );
  OAI22_X2 U2362 ( .A1(n5931), .A2(n7552), .B1(n6099), .B2(n7544), .ZN(n4257)
         );
  AOI221_X2 U2363 ( .B1(n7506), .B2(REG_FILE_reg_out_26__6_), .C1(n7514), .C2(
        REG_FILE_reg_out_30__6_), .A(n4258), .ZN(n4255) );
  OAI22_X2 U2364 ( .A1(n5977), .A2(n7534), .B1(n6255), .B2(n7521), .ZN(n4258)
         );
  AOI221_X2 U2366 ( .B1(n7490), .B2(REG_FILE_reg_out_3__6_), .C1(n7498), .C2(
        REG_FILE_reg_out_7__6_), .A(n4261), .ZN(n4260) );
  OAI22_X2 U2367 ( .A1(n6117), .A2(n7552), .B1(n6466), .B2(n7544), .ZN(n4261)
         );
  AOI221_X2 U2368 ( .B1(n7506), .B2(REG_FILE_reg_out_2__6_), .C1(n7514), .C2(
        REG_FILE_reg_out_6__6_), .A(n4262), .ZN(n4259) );
  OAI22_X2 U2369 ( .A1(n6198), .A2(n7534), .B1(n6629), .B2(n7521), .ZN(n4262)
         );
  OAI22_X2 U2371 ( .A1(n6195), .A2(n7534), .B1(n6637), .B2(n7521), .ZN(n4266)
         );
  OAI22_X2 U2372 ( .A1(n6369), .A2(n7515), .B1(n6092), .B2(n7508), .ZN(n4265)
         );
  OAI22_X2 U2373 ( .A1(n6053), .A2(n7552), .B1(n6404), .B2(n7544), .ZN(n4264)
         );
  OAI22_X2 U2374 ( .A1(n6544), .A2(n7499), .B1(n6251), .B2(n7492), .ZN(n4263)
         );
  AOI221_X2 U2379 ( .B1(n7490), .B2(REG_FILE_reg_out_11__7_), .C1(n7498), .C2(
        REG_FILE_reg_out_15__7_), .A(n4275), .ZN(n4274) );
  OAI22_X2 U2380 ( .A1(n6362), .A2(n7552), .B1(n6950), .B2(n7544), .ZN(n4275)
         );
  AOI221_X2 U2381 ( .B1(n7506), .B2(REG_FILE_reg_out_10__7_), .C1(n7514), .C2(
        REG_FILE_reg_out_14__7_), .A(n4276), .ZN(n4273) );
  OAI22_X2 U2382 ( .A1(n6537), .A2(n7534), .B1(n6261), .B2(n7521), .ZN(n4276)
         );
  AOI221_X2 U2384 ( .B1(n7490), .B2(REG_FILE_reg_out_27__7_), .C1(n7498), .C2(
        REG_FILE_reg_out_31__7_), .A(n4279), .ZN(n4278) );
  OAI22_X2 U2385 ( .A1(n5932), .A2(n7548), .B1(n6100), .B2(n7539), .ZN(n4279)
         );
  AOI221_X2 U2386 ( .B1(n7506), .B2(REG_FILE_reg_out_26__7_), .C1(n7514), .C2(
        REG_FILE_reg_out_30__7_), .A(n4280), .ZN(n4277) );
  OAI22_X2 U2387 ( .A1(n5978), .A2(n7533), .B1(n6256), .B2(n7521), .ZN(n4280)
         );
  AOI221_X2 U2389 ( .B1(n7490), .B2(REG_FILE_reg_out_3__7_), .C1(n7498), .C2(
        REG_FILE_reg_out_7__7_), .A(n4283), .ZN(n4282) );
  OAI22_X2 U2390 ( .A1(n5881), .A2(n7547), .B1(n6129), .B2(n7539), .ZN(n4283)
         );
  AOI221_X2 U2391 ( .B1(n7506), .B2(REG_FILE_reg_out_2__7_), .C1(n7514), .C2(
        REG_FILE_reg_out_6__7_), .A(n4284), .ZN(n4281) );
  OAI22_X2 U2392 ( .A1(n5984), .A2(n7533), .B1(n6630), .B2(n7521), .ZN(n4284)
         );
  OAI22_X2 U2394 ( .A1(n6196), .A2(n7533), .B1(n6638), .B2(n7521), .ZN(n4288)
         );
  OAI22_X2 U2395 ( .A1(n6370), .A2(n7515), .B1(n6093), .B2(n7508), .ZN(n4287)
         );
  OAI22_X2 U2396 ( .A1(n5870), .A2(n7547), .B1(n6085), .B2(n7544), .ZN(n4286)
         );
  OAI22_X2 U2397 ( .A1(n6545), .A2(n7499), .B1(n6252), .B2(n7492), .ZN(n4285)
         );
  AOI221_X2 U2402 ( .B1(n7490), .B2(REG_FILE_reg_out_11__8_), .C1(n7498), .C2(
        REG_FILE_reg_out_15__8_), .A(n4298), .ZN(n4297) );
  OAI22_X2 U2403 ( .A1(n5879), .A2(n7550), .B1(n6112), .B2(n7539), .ZN(n4298)
         );
  AOI221_X2 U2404 ( .B1(n7506), .B2(REG_FILE_reg_out_10__8_), .C1(n7514), .C2(
        REG_FILE_reg_out_14__8_), .A(n4299), .ZN(n4296) );
  OAI22_X2 U2405 ( .A1(n6239), .A2(n7533), .B1(n6698), .B2(n7521), .ZN(n4299)
         );
  AOI221_X2 U2407 ( .B1(n7490), .B2(REG_FILE_reg_out_27__8_), .C1(n7498), .C2(
        REG_FILE_reg_out_31__8_), .A(n4302), .ZN(n4301) );
  OAI22_X2 U2408 ( .A1(n6084), .A2(n7548), .B1(n6978), .B2(n7539), .ZN(n4302)
         );
  AOI221_X2 U2409 ( .B1(n7506), .B2(REG_FILE_reg_out_26__8_), .C1(n7514), .C2(
        REG_FILE_reg_out_30__8_), .A(n4303), .ZN(n4300) );
  OAI22_X2 U2410 ( .A1(n6607), .A2(n7533), .B1(n7134), .B2(n7521), .ZN(n4303)
         );
  AOI221_X2 U2412 ( .B1(n7490), .B2(REG_FILE_reg_out_3__8_), .C1(n7498), .C2(
        REG_FILE_reg_out_7__8_), .A(n4306), .ZN(n4305) );
  OAI22_X2 U2413 ( .A1(n5883), .A2(n7549), .B1(n6133), .B2(n7539), .ZN(n4306)
         );
  AOI221_X2 U2414 ( .B1(n7506), .B2(REG_FILE_reg_out_2__8_), .C1(n7514), .C2(
        REG_FILE_reg_out_6__8_), .A(n4307), .ZN(n4304) );
  OAI22_X2 U2415 ( .A1(n5995), .A2(n7533), .B1(n6697), .B2(n7522), .ZN(n4307)
         );
  OAI22_X2 U2417 ( .A1(n6238), .A2(n7533), .B1(n6696), .B2(n7522), .ZN(n4311)
         );
  OAI22_X2 U2418 ( .A1(n6398), .A2(n4128), .B1(n6977), .B2(n7508), .ZN(n4310)
         );
  OAI22_X2 U2419 ( .A1(n5878), .A2(n7548), .B1(n6111), .B2(n7539), .ZN(n4309)
         );
  OAI22_X2 U2420 ( .A1(n6606), .A2(n4130), .B1(n7133), .B2(n7492), .ZN(n4308)
         );
  AOI221_X2 U2425 ( .B1(n7490), .B2(REG_FILE_reg_out_11__9_), .C1(n7498), .C2(
        REG_FILE_reg_out_15__9_), .A(n4320), .ZN(n4319) );
  OAI22_X2 U2426 ( .A1(n5877), .A2(n7551), .B1(n6110), .B2(n7539), .ZN(n4320)
         );
  AOI221_X2 U2427 ( .B1(n7506), .B2(REG_FILE_reg_out_10__9_), .C1(n7514), .C2(
        REG_FILE_reg_out_14__9_), .A(n4321), .ZN(n4318) );
  OAI22_X2 U2428 ( .A1(n6605), .A2(n7533), .B1(n7132), .B2(n7522), .ZN(n4321)
         );
  AOI221_X2 U2430 ( .B1(n7490), .B2(REG_FILE_reg_out_27__9_), .C1(n7498), .C2(
        REG_FILE_reg_out_31__9_), .A(n4324), .ZN(n4323) );
  OAI22_X2 U2431 ( .A1(n6083), .A2(n7548), .B1(n6976), .B2(n7539), .ZN(n4324)
         );
  AOI221_X2 U2432 ( .B1(n7506), .B2(REG_FILE_reg_out_26__9_), .C1(n7514), .C2(
        REG_FILE_reg_out_30__9_), .A(n4325), .ZN(n4322) );
  OAI22_X2 U2433 ( .A1(n6604), .A2(n7533), .B1(n7131), .B2(n7522), .ZN(n4325)
         );
  AOI221_X2 U2435 ( .B1(n7490), .B2(REG_FILE_reg_out_3__9_), .C1(n7498), .C2(
        REG_FILE_reg_out_7__9_), .A(n4328), .ZN(n4327) );
  OAI22_X2 U2436 ( .A1(n6980), .A2(n7548), .B1(n6132), .B2(n7539), .ZN(n4328)
         );
  AOI221_X2 U2437 ( .B1(n7506), .B2(REG_FILE_reg_out_2__9_), .C1(n7514), .C2(
        REG_FILE_reg_out_6__9_), .A(n4329), .ZN(n4326) );
  OAI22_X2 U2438 ( .A1(n7074), .A2(n7533), .B1(n6695), .B2(n7522), .ZN(n4329)
         );
  OAI22_X2 U2440 ( .A1(n6237), .A2(n7533), .B1(n6694), .B2(n7522), .ZN(n4333)
         );
  OAI22_X2 U2441 ( .A1(n6397), .A2(n4128), .B1(n6975), .B2(n7508), .ZN(n4332)
         );
  OAI22_X2 U2442 ( .A1(n5876), .A2(n7549), .B1(n6109), .B2(n7543), .ZN(n4331)
         );
  OAI22_X2 U2443 ( .A1(n6603), .A2(n4130), .B1(n7130), .B2(n7492), .ZN(n4330)
         );
  AOI221_X2 U2448 ( .B1(n7489), .B2(REG_FILE_reg_out_11__10_), .C1(n7497), 
        .C2(REG_FILE_reg_out_15__10_), .A(n4343), .ZN(n4342) );
  OAI22_X2 U2449 ( .A1(n6396), .A2(n7551), .B1(n6974), .B2(n7543), .ZN(n4343)
         );
  AOI221_X2 U2450 ( .B1(n7505), .B2(REG_FILE_reg_out_10__10_), .C1(n7511), 
        .C2(REG_FILE_reg_out_14__10_), .A(n4344), .ZN(n4341) );
  OAI22_X2 U2451 ( .A1(n5994), .A2(n7532), .B1(n6265), .B2(n7522), .ZN(n4344)
         );
  AOI221_X2 U2453 ( .B1(n7489), .B2(REG_FILE_reg_out_27__10_), .C1(n7497), 
        .C2(REG_FILE_reg_out_31__10_), .A(n4347), .ZN(n4346) );
  OAI22_X2 U2454 ( .A1(n6082), .A2(n7551), .B1(n6449), .B2(n7543), .ZN(n4347)
         );
  AOI221_X2 U2455 ( .B1(n7505), .B2(REG_FILE_reg_out_26__10_), .C1(n7511), 
        .C2(REG_FILE_reg_out_30__10_), .A(n4348), .ZN(n4345) );
  OAI22_X2 U2456 ( .A1(n5993), .A2(n7532), .B1(n6264), .B2(n7522), .ZN(n4348)
         );
  AOI221_X2 U2458 ( .B1(n7489), .B2(REG_FILE_reg_out_3__10_), .C1(n7497), .C2(
        REG_FILE_reg_out_7__10_), .A(n4351), .ZN(n4350) );
  OAI22_X2 U2459 ( .A1(n6460), .A2(n7551), .B1(n6127), .B2(n7543), .ZN(n4351)
         );
  AOI221_X2 U2460 ( .B1(n7505), .B2(REG_FILE_reg_out_2__10_), .C1(n7511), .C2(
        REG_FILE_reg_out_6__10_), .A(n4352), .ZN(n4349) );
  OAI22_X2 U2461 ( .A1(n5992), .A2(n7531), .B1(n6243), .B2(n7522), .ZN(n4352)
         );
  OAI22_X2 U2463 ( .A1(n5991), .A2(n7532), .B1(n6242), .B2(n7522), .ZN(n4356)
         );
  OAI22_X2 U2464 ( .A1(n5943), .A2(n4128), .B1(n6108), .B2(n7508), .ZN(n4355)
         );
  OAI22_X2 U2465 ( .A1(n6395), .A2(n7551), .B1(n6059), .B2(n7543), .ZN(n4354)
         );
  OAI22_X2 U2466 ( .A1(n6236), .A2(n4130), .B1(n6693), .B2(n7492), .ZN(n4353)
         );
  AOI221_X2 U2471 ( .B1(n7489), .B2(REG_FILE_reg_out_11__11_), .C1(n7497), 
        .C2(REG_FILE_reg_out_15__11_), .A(n4365), .ZN(n4364) );
  OAI22_X2 U2472 ( .A1(n6394), .A2(n7551), .B1(n6973), .B2(n7543), .ZN(n4365)
         );
  AOI221_X2 U2473 ( .B1(n7505), .B2(REG_FILE_reg_out_10__11_), .C1(n7511), 
        .C2(REG_FILE_reg_out_14__11_), .A(n4366), .ZN(n4363) );
  OAI22_X2 U2474 ( .A1(n6235), .A2(n7532), .B1(n7129), .B2(n7522), .ZN(n4366)
         );
  AOI221_X2 U2476 ( .B1(n7489), .B2(REG_FILE_reg_out_27__11_), .C1(n7497), 
        .C2(REG_FILE_reg_out_31__11_), .A(n4369), .ZN(n4368) );
  OAI22_X2 U2477 ( .A1(n6393), .A2(n7551), .B1(n6972), .B2(n7543), .ZN(n4369)
         );
  AOI221_X2 U2478 ( .B1(n7505), .B2(REG_FILE_reg_out_26__11_), .C1(n7511), 
        .C2(REG_FILE_reg_out_30__11_), .A(n4370), .ZN(n4367) );
  OAI22_X2 U2479 ( .A1(n6234), .A2(n7532), .B1(n7128), .B2(n7522), .ZN(n4370)
         );
  AOI221_X2 U2481 ( .B1(n7489), .B2(REG_FILE_reg_out_3__11_), .C1(n7497), .C2(
        REG_FILE_reg_out_7__11_), .A(n4373), .ZN(n4372) );
  OAI22_X2 U2482 ( .A1(n6459), .A2(n7551), .B1(n6986), .B2(n7543), .ZN(n4373)
         );
  AOI221_X2 U2483 ( .B1(n7505), .B2(REG_FILE_reg_out_2__11_), .C1(n7511), .C2(
        REG_FILE_reg_out_6__11_), .A(n4374), .ZN(n4371) );
  OAI22_X2 U2484 ( .A1(n5990), .A2(n7532), .B1(n7090), .B2(n7522), .ZN(n4374)
         );
  OAI22_X2 U2486 ( .A1(n6233), .A2(n7531), .B1(n7089), .B2(n7522), .ZN(n4378)
         );
  OAI22_X2 U2487 ( .A1(n6081), .A2(n4128), .B1(n6971), .B2(n7508), .ZN(n4377)
         );
  OAI22_X2 U2488 ( .A1(n6392), .A2(n7551), .B1(n6922), .B2(n7543), .ZN(n4376)
         );
  OAI22_X2 U2489 ( .A1(n6602), .A2(n4130), .B1(n7127), .B2(n7492), .ZN(n4375)
         );
  AOI221_X2 U2494 ( .B1(n7489), .B2(REG_FILE_reg_out_11__12_), .C1(n7497), 
        .C2(REG_FILE_reg_out_15__12_), .A(n4388), .ZN(n4387) );
  OAI22_X2 U2495 ( .A1(n6080), .A2(n7551), .B1(n6448), .B2(n7543), .ZN(n4388)
         );
  AOI221_X2 U2496 ( .B1(n7505), .B2(REG_FILE_reg_out_10__12_), .C1(n7511), 
        .C2(REG_FILE_reg_out_14__12_), .A(n4389), .ZN(n4386) );
  OAI22_X2 U2497 ( .A1(n5907), .A2(n7532), .B1(n6263), .B2(n7522), .ZN(n4389)
         );
  AOI221_X2 U2499 ( .B1(n7489), .B2(REG_FILE_reg_out_27__12_), .C1(n7497), 
        .C2(REG_FILE_reg_out_31__12_), .A(n4392), .ZN(n4391) );
  OAI22_X2 U2500 ( .A1(n6079), .A2(n7551), .B1(n6447), .B2(n7543), .ZN(n4392)
         );
  AOI221_X2 U2501 ( .B1(n7505), .B2(REG_FILE_reg_out_26__12_), .C1(n7511), 
        .C2(REG_FILE_reg_out_30__12_), .A(n4393), .ZN(n4390) );
  OAI22_X2 U2502 ( .A1(n5989), .A2(n7531), .B1(n6262), .B2(n7522), .ZN(n4393)
         );
  AOI221_X2 U2504 ( .B1(n7489), .B2(REG_FILE_reg_out_3__12_), .C1(n7497), .C2(
        REG_FILE_reg_out_7__12_), .A(n4396), .ZN(n4395) );
  OAI22_X2 U2505 ( .A1(n6458), .A2(n7551), .B1(n6126), .B2(n7543), .ZN(n4396)
         );
  AOI221_X2 U2506 ( .B1(n7505), .B2(REG_FILE_reg_out_2__12_), .C1(n7511), .C2(
        REG_FILE_reg_out_6__12_), .A(n4397), .ZN(n4394) );
  OAI22_X2 U2507 ( .A1(n5988), .A2(n7531), .B1(n6241), .B2(n7522), .ZN(n4397)
         );
  OAI22_X2 U2509 ( .A1(n6601), .A2(n7532), .B1(n6240), .B2(n7522), .ZN(n4401)
         );
  OAI22_X2 U2510 ( .A1(n5942), .A2(n7515), .B1(n6107), .B2(n7507), .ZN(n4400)
         );
  OAI22_X2 U2511 ( .A1(n6391), .A2(n7550), .B1(n6058), .B2(n7543), .ZN(n4399)
         );
  OAI22_X2 U2512 ( .A1(n6232), .A2(n7499), .B1(n6692), .B2(n7491), .ZN(n4398)
         );
  AOI221_X2 U2518 ( .B1(n7489), .B2(REG_FILE_reg_out_11__13_), .C1(n7497), 
        .C2(REG_FILE_reg_out_15__13_), .A(n4410), .ZN(n4409) );
  OAI22_X2 U2519 ( .A1(n6078), .A2(n7550), .B1(n6446), .B2(n7543), .ZN(n4410)
         );
  AOI221_X2 U2520 ( .B1(n7505), .B2(REG_FILE_reg_out_10__13_), .C1(n7511), 
        .C2(REG_FILE_reg_out_14__13_), .A(n4411), .ZN(n4408) );
  OAI22_X2 U2521 ( .A1(n6231), .A2(n7532), .B1(n6691), .B2(n7525), .ZN(n4411)
         );
  AOI221_X2 U2523 ( .B1(n7489), .B2(REG_FILE_reg_out_27__13_), .C1(n7497), 
        .C2(REG_FILE_reg_out_31__13_), .A(n4414), .ZN(n4413) );
  OAI22_X2 U2524 ( .A1(n6077), .A2(n7550), .B1(n6445), .B2(n7543), .ZN(n4414)
         );
  AOI221_X2 U2525 ( .B1(n7505), .B2(REG_FILE_reg_out_26__13_), .C1(n7511), 
        .C2(REG_FILE_reg_out_30__13_), .A(n4415), .ZN(n4412) );
  OAI22_X2 U2526 ( .A1(n6230), .A2(n7532), .B1(n6690), .B2(n7525), .ZN(n4415)
         );
  AOI221_X2 U2528 ( .B1(n7488), .B2(REG_FILE_reg_out_3__13_), .C1(n7494), .C2(
        REG_FILE_reg_out_7__13_), .A(n4418), .ZN(n4417) );
  OAI22_X2 U2529 ( .A1(n6979), .A2(n7550), .B1(n6475), .B2(n7543), .ZN(n4418)
         );
  AOI221_X2 U2530 ( .B1(n7504), .B2(REG_FILE_reg_out_2__13_), .C1(n7510), .C2(
        REG_FILE_reg_out_6__13_), .A(n4419), .ZN(n4416) );
  OAI22_X2 U2531 ( .A1(n7073), .A2(n7532), .B1(n6689), .B2(n7525), .ZN(n4419)
         );
  OAI22_X2 U2533 ( .A1(n6229), .A2(n7532), .B1(n6688), .B2(n7525), .ZN(n4423)
         );
  OAI22_X2 U2534 ( .A1(n5941), .A2(n7515), .B1(n6106), .B2(n7507), .ZN(n4422)
         );
  OAI22_X2 U2535 ( .A1(n6076), .A2(n7550), .B1(n6444), .B2(n7543), .ZN(n4421)
         );
  OAI22_X2 U2536 ( .A1(n6228), .A2(n7499), .B1(n6687), .B2(n7491), .ZN(n4420)
         );
  AOI221_X2 U2541 ( .B1(n7488), .B2(REG_FILE_reg_out_11__14_), .C1(n7494), 
        .C2(REG_FILE_reg_out_15__14_), .A(n4433), .ZN(n4432) );
  OAI22_X2 U2542 ( .A1(n6075), .A2(n7550), .B1(n6443), .B2(n7543), .ZN(n4433)
         );
  AOI221_X2 U2543 ( .B1(n7504), .B2(REG_FILE_reg_out_10__14_), .C1(n7510), 
        .C2(REG_FILE_reg_out_14__14_), .A(n4434), .ZN(n4431) );
  OAI22_X2 U2544 ( .A1(n6227), .A2(n7532), .B1(n6686), .B2(n7525), .ZN(n4434)
         );
  AOI221_X2 U2546 ( .B1(n7488), .B2(REG_FILE_reg_out_27__14_), .C1(n7494), 
        .C2(REG_FILE_reg_out_31__14_), .A(n4437), .ZN(n4436) );
  OAI22_X2 U2547 ( .A1(n6074), .A2(n7550), .B1(n6442), .B2(n7543), .ZN(n4437)
         );
  AOI221_X2 U2548 ( .B1(n7504), .B2(REG_FILE_reg_out_26__14_), .C1(n7510), 
        .C2(REG_FILE_reg_out_30__14_), .A(n4438), .ZN(n4435) );
  OAI22_X2 U2549 ( .A1(n6226), .A2(n7532), .B1(n6685), .B2(n7525), .ZN(n4438)
         );
  AOI221_X2 U2551 ( .B1(n7488), .B2(REG_FILE_reg_out_3__14_), .C1(n7494), .C2(
        REG_FILE_reg_out_7__14_), .A(n4441), .ZN(n4440) );
  OAI22_X2 U2552 ( .A1(n6457), .A2(n7550), .B1(n6985), .B2(n7543), .ZN(n4441)
         );
  AOI221_X2 U2553 ( .B1(n7504), .B2(REG_FILE_reg_out_2__14_), .C1(n7510), .C2(
        REG_FILE_reg_out_6__14_), .A(n4442), .ZN(n4439) );
  OAI22_X2 U2554 ( .A1(n6600), .A2(n7532), .B1(n7088), .B2(n7521), .ZN(n4442)
         );
  OAI22_X2 U2556 ( .A1(n6599), .A2(n7532), .B1(n7087), .B2(n7521), .ZN(n4446)
         );
  OAI22_X2 U2557 ( .A1(n5940), .A2(n7515), .B1(n6105), .B2(n7507), .ZN(n4445)
         );
  OAI22_X2 U2558 ( .A1(n6390), .A2(n7550), .B1(n6057), .B2(n7543), .ZN(n4444)
         );
  OAI22_X2 U2559 ( .A1(n6225), .A2(n7499), .B1(n6684), .B2(n7491), .ZN(n4443)
         );
  AOI221_X2 U2566 ( .B1(n7488), .B2(REG_FILE_reg_out_11__15_), .C1(n7494), 
        .C2(REG_FILE_reg_out_15__15_), .A(n4458), .ZN(n4457) );
  OAI22_X2 U2567 ( .A1(n6389), .A2(n7550), .B1(n6970), .B2(n7543), .ZN(n4458)
         );
  AOI221_X2 U2568 ( .B1(n7504), .B2(REG_FILE_reg_out_10__15_), .C1(n7510), 
        .C2(REG_FILE_reg_out_14__15_), .A(n4459), .ZN(n4456) );
  OAI22_X2 U2569 ( .A1(n6598), .A2(n7532), .B1(n7126), .B2(n7525), .ZN(n4459)
         );
  AOI221_X2 U2571 ( .B1(n7488), .B2(REG_FILE_reg_out_27__15_), .C1(n7495), 
        .C2(REG_FILE_reg_out_31__15_), .A(n4462), .ZN(n4461) );
  OAI22_X2 U2572 ( .A1(n6388), .A2(n7550), .B1(n6969), .B2(n7543), .ZN(n4462)
         );
  AOI221_X2 U2573 ( .B1(n7504), .B2(REG_FILE_reg_out_26__15_), .C1(n7513), 
        .C2(REG_FILE_reg_out_30__15_), .A(n4463), .ZN(n4460) );
  OAI22_X2 U2574 ( .A1(n6597), .A2(n7532), .B1(n7125), .B2(n7521), .ZN(n4463)
         );
  AOI221_X2 U2576 ( .B1(n7488), .B2(REG_FILE_reg_out_3__15_), .C1(n7495), .C2(
        REG_FILE_reg_out_7__15_), .A(n4466), .ZN(n4465) );
  OAI22_X2 U2577 ( .A1(n6456), .A2(n7549), .B1(n6984), .B2(n7542), .ZN(n4466)
         );
  AOI221_X2 U2578 ( .B1(n7504), .B2(REG_FILE_reg_out_2__15_), .C1(n7513), .C2(
        REG_FILE_reg_out_6__15_), .A(n4467), .ZN(n4464) );
  OAI22_X2 U2579 ( .A1(n6596), .A2(n7530), .B1(n7086), .B2(n7521), .ZN(n4467)
         );
  OAI22_X2 U2581 ( .A1(n6595), .A2(n7530), .B1(n7085), .B2(n7525), .ZN(n4471)
         );
  OAI22_X2 U2582 ( .A1(n6073), .A2(n7515), .B1(n6968), .B2(n7507), .ZN(n4470)
         );
  OAI22_X2 U2583 ( .A1(n6387), .A2(n7549), .B1(n6921), .B2(n7542), .ZN(n4469)
         );
  OAI22_X2 U2584 ( .A1(n6594), .A2(n7499), .B1(n7124), .B2(n7491), .ZN(n4468)
         );
  AOI221_X2 U2589 ( .B1(n7488), .B2(REG_FILE_reg_out_11__16_), .C1(n7495), 
        .C2(REG_FILE_reg_out_15__16_), .A(n4480), .ZN(n4479) );
  OAI22_X2 U2590 ( .A1(n6945), .A2(n7549), .B1(n6441), .B2(n7542), .ZN(n4480)
         );
  AOI221_X2 U2591 ( .B1(n7504), .B2(REG_FILE_reg_out_10__16_), .C1(n7513), 
        .C2(REG_FILE_reg_out_14__16_), .A(n4481), .ZN(n4478) );
  OAI22_X2 U2592 ( .A1(n7072), .A2(n7530), .B1(n6683), .B2(n7521), .ZN(n4481)
         );
  AOI221_X2 U2594 ( .B1(n7488), .B2(REG_FILE_reg_out_27__16_), .C1(n7495), 
        .C2(REG_FILE_reg_out_31__16_), .A(n4484), .ZN(n4483) );
  OAI22_X2 U2595 ( .A1(n6072), .A2(n7549), .B1(n6440), .B2(n7542), .ZN(n4484)
         );
  AOI221_X2 U2596 ( .B1(n7504), .B2(REG_FILE_reg_out_26__16_), .C1(n7513), 
        .C2(REG_FILE_reg_out_30__16_), .A(n4485), .ZN(n4482) );
  OAI22_X2 U2597 ( .A1(n5987), .A2(n7530), .B1(n6682), .B2(n7521), .ZN(n4485)
         );
  AOI221_X2 U2599 ( .B1(n7488), .B2(REG_FILE_reg_out_3__16_), .C1(n7495), .C2(
        REG_FILE_reg_out_7__16_), .A(n4488), .ZN(n4487) );
  OAI22_X2 U2600 ( .A1(n6455), .A2(n7549), .B1(n6983), .B2(n7542), .ZN(n4488)
         );
  AOI221_X2 U2601 ( .B1(n7504), .B2(REG_FILE_reg_out_2__16_), .C1(n7513), .C2(
        REG_FILE_reg_out_6__16_), .A(n4489), .ZN(n4486) );
  OAI22_X2 U2602 ( .A1(n6593), .A2(n7530), .B1(n7084), .B2(n7521), .ZN(n4489)
         );
  OAI22_X2 U2604 ( .A1(n6592), .A2(n7530), .B1(n7083), .B2(n7525), .ZN(n4493)
         );
  OAI22_X2 U2605 ( .A1(n6944), .A2(n7515), .B1(n6104), .B2(n7507), .ZN(n4492)
         );
  OAI22_X2 U2606 ( .A1(n6943), .A2(n7549), .B1(n6056), .B2(n7542), .ZN(n4491)
         );
  OAI22_X2 U2607 ( .A1(n7071), .A2(n7499), .B1(n6681), .B2(n7491), .ZN(n4490)
         );
  AOI221_X2 U2612 ( .B1(n7488), .B2(REG_FILE_reg_out_11__17_), .C1(n7494), 
        .C2(REG_FILE_reg_out_15__17_), .A(n4502), .ZN(n4501) );
  OAI22_X2 U2613 ( .A1(n6942), .A2(n7549), .B1(n6439), .B2(n7542), .ZN(n4502)
         );
  AOI221_X2 U2614 ( .B1(n7504), .B2(REG_FILE_reg_out_10__17_), .C1(n7510), 
        .C2(REG_FILE_reg_out_14__17_), .A(n4503), .ZN(n4500) );
  OAI22_X2 U2615 ( .A1(n7070), .A2(n7530), .B1(n6680), .B2(n7525), .ZN(n4503)
         );
  AOI221_X2 U2617 ( .B1(n7488), .B2(REG_FILE_reg_out_27__17_), .C1(n7496), 
        .C2(REG_FILE_reg_out_31__17_), .A(n4506), .ZN(n4505) );
  OAI22_X2 U2618 ( .A1(n6071), .A2(n7549), .B1(n6438), .B2(n7542), .ZN(n4506)
         );
  AOI221_X2 U2619 ( .B1(n7504), .B2(REG_FILE_reg_out_26__17_), .C1(n7512), 
        .C2(REG_FILE_reg_out_30__17_), .A(n4507), .ZN(n4504) );
  OAI22_X2 U2620 ( .A1(n5986), .A2(n7530), .B1(n6679), .B2(n7523), .ZN(n4507)
         );
  AOI221_X2 U2622 ( .B1(n7488), .B2(REG_FILE_reg_out_3__17_), .C1(n7496), .C2(
        REG_FILE_reg_out_7__17_), .A(n4510), .ZN(n4509) );
  OAI22_X2 U2623 ( .A1(n6122), .A2(n7549), .B1(n6474), .B2(n7542), .ZN(n4510)
         );
  AOI221_X2 U2624 ( .B1(n7504), .B2(REG_FILE_reg_out_2__17_), .C1(n7513), .C2(
        REG_FILE_reg_out_6__17_), .A(n4511), .ZN(n4508) );
  OAI22_X2 U2625 ( .A1(n6591), .A2(n7530), .B1(n7123), .B2(n7523), .ZN(n4511)
         );
  OAI22_X2 U2627 ( .A1(n6590), .A2(n7530), .B1(n7122), .B2(n7523), .ZN(n4515)
         );
  OAI22_X2 U2628 ( .A1(n6941), .A2(n7515), .B1(n6437), .B2(n7507), .ZN(n4514)
         );
  OAI22_X2 U2629 ( .A1(n6940), .A2(n7549), .B1(n6436), .B2(n7542), .ZN(n4513)
         );
  OAI22_X2 U2630 ( .A1(n7069), .A2(n7499), .B1(n6678), .B2(n7491), .ZN(n4512)
         );
  AOI221_X2 U2635 ( .B1(n7488), .B2(REG_FILE_reg_out_11__18_), .C1(n7496), 
        .C2(REG_FILE_reg_out_15__18_), .A(n4525), .ZN(n4524) );
  OAI22_X2 U2636 ( .A1(n6939), .A2(n7549), .B1(n6435), .B2(n7542), .ZN(n4525)
         );
  AOI221_X2 U2637 ( .B1(n7504), .B2(REG_FILE_reg_out_10__18_), .C1(n7512), 
        .C2(REG_FILE_reg_out_14__18_), .A(n4526), .ZN(n4523) );
  OAI22_X2 U2638 ( .A1(n7068), .A2(n7530), .B1(n6677), .B2(n7523), .ZN(n4526)
         );
  AOI221_X2 U2640 ( .B1(n7488), .B2(REG_FILE_reg_out_27__18_), .C1(n7496), 
        .C2(REG_FILE_reg_out_31__18_), .A(n4529), .ZN(n4528) );
  OAI22_X2 U2641 ( .A1(n5939), .A2(n7548), .B1(n6434), .B2(n7540), .ZN(n4529)
         );
  AOI221_X2 U2642 ( .B1(n7504), .B2(REG_FILE_reg_out_26__18_), .C1(n7512), 
        .C2(REG_FILE_reg_out_30__18_), .A(n4530), .ZN(n4527) );
  OAI22_X2 U2643 ( .A1(n6224), .A2(n7531), .B1(n6676), .B2(n7523), .ZN(n4530)
         );
  AOI221_X2 U2645 ( .B1(n7488), .B2(REG_FILE_reg_out_3__18_), .C1(n7496), .C2(
        REG_FILE_reg_out_7__18_), .A(n4533), .ZN(n4532) );
  OAI22_X2 U2646 ( .A1(n5951), .A2(n7548), .B1(n6473), .B2(n7540), .ZN(n4533)
         );
  AOI221_X2 U2647 ( .B1(n7504), .B2(REG_FILE_reg_out_2__18_), .C1(n7512), .C2(
        REG_FILE_reg_out_6__18_), .A(n4534), .ZN(n4531) );
  OAI22_X2 U2648 ( .A1(n6223), .A2(n7531), .B1(n6675), .B2(n7523), .ZN(n4534)
         );
  OAI22_X2 U2650 ( .A1(n7067), .A2(n7531), .B1(n6674), .B2(n7523), .ZN(n4538)
         );
  OAI22_X2 U2651 ( .A1(n6938), .A2(n7515), .B1(n6433), .B2(n7507), .ZN(n4537)
         );
  OAI22_X2 U2652 ( .A1(n6937), .A2(n7548), .B1(n6432), .B2(n7540), .ZN(n4536)
         );
  OAI22_X2 U2653 ( .A1(n7066), .A2(n7499), .B1(n6673), .B2(n7491), .ZN(n4535)
         );
  AOI221_X2 U2658 ( .B1(n7488), .B2(REG_FILE_reg_out_11__19_), .C1(n7496), 
        .C2(REG_FILE_reg_out_15__19_), .A(n4547), .ZN(n4546) );
  OAI22_X2 U2659 ( .A1(n5938), .A2(n7548), .B1(n6431), .B2(n7540), .ZN(n4547)
         );
  AOI221_X2 U2660 ( .B1(n7504), .B2(REG_FILE_reg_out_10__19_), .C1(n7512), 
        .C2(REG_FILE_reg_out_14__19_), .A(n4548), .ZN(n4545) );
  OAI22_X2 U2661 ( .A1(n6589), .A2(n7531), .B1(n7121), .B2(n7523), .ZN(n4548)
         );
  AOI221_X2 U2663 ( .B1(n7488), .B2(REG_FILE_reg_out_27__19_), .C1(n7496), 
        .C2(REG_FILE_reg_out_31__19_), .A(n4551), .ZN(n4550) );
  OAI22_X2 U2664 ( .A1(n5937), .A2(n7548), .B1(n6430), .B2(n7540), .ZN(n4551)
         );
  AOI221_X2 U2665 ( .B1(n7504), .B2(REG_FILE_reg_out_26__19_), .C1(n7512), 
        .C2(REG_FILE_reg_out_30__19_), .A(n4552), .ZN(n4549) );
  OAI22_X2 U2666 ( .A1(n6222), .A2(n7531), .B1(n6672), .B2(n7523), .ZN(n4552)
         );
  AOI221_X2 U2668 ( .B1(n7488), .B2(REG_FILE_reg_out_3__19_), .C1(n7496), .C2(
        REG_FILE_reg_out_7__19_), .A(n4555), .ZN(n4554) );
  OAI22_X2 U2669 ( .A1(n6454), .A2(n7548), .B1(n6987), .B2(n7540), .ZN(n4555)
         );
  AOI221_X2 U2670 ( .B1(n7504), .B2(REG_FILE_reg_out_2__19_), .C1(n7510), .C2(
        REG_FILE_reg_out_6__19_), .A(n4556), .ZN(n4553) );
  OAI22_X2 U2671 ( .A1(n6588), .A2(n7531), .B1(n7120), .B2(n7523), .ZN(n4556)
         );
  OAI22_X2 U2673 ( .A1(n6587), .A2(n7531), .B1(n7119), .B2(n7523), .ZN(n4560)
         );
  OAI22_X2 U2674 ( .A1(n6386), .A2(n7515), .B1(n6967), .B2(n7507), .ZN(n4559)
         );
  OAI22_X2 U2675 ( .A1(n6385), .A2(n7548), .B1(n6966), .B2(n7540), .ZN(n4558)
         );
  OAI22_X2 U2676 ( .A1(n6586), .A2(n7499), .B1(n7118), .B2(n7491), .ZN(n4557)
         );
  AOI221_X2 U2681 ( .B1(n7488), .B2(REG_FILE_reg_out_11__20_), .C1(n7496), 
        .C2(REG_FILE_reg_out_15__20_), .A(n4569), .ZN(n4568) );
  OAI22_X2 U2682 ( .A1(n6936), .A2(n7548), .B1(n6429), .B2(n7540), .ZN(n4569)
         );
  AOI221_X2 U2683 ( .B1(n7504), .B2(REG_FILE_reg_out_10__20_), .C1(n7512), 
        .C2(REG_FILE_reg_out_14__20_), .A(n4570), .ZN(n4567) );
  OAI22_X2 U2684 ( .A1(n7065), .A2(n7531), .B1(n6671), .B2(n7523), .ZN(n4570)
         );
  AOI221_X2 U2686 ( .B1(n7488), .B2(REG_FILE_reg_out_27__20_), .C1(n7496), 
        .C2(REG_FILE_reg_out_31__20_), .A(n4573), .ZN(n4572) );
  OAI22_X2 U2687 ( .A1(n5936), .A2(n7548), .B1(n6428), .B2(n7540), .ZN(n4573)
         );
  AOI221_X2 U2688 ( .B1(n7504), .B2(REG_FILE_reg_out_26__20_), .C1(n7512), 
        .C2(REG_FILE_reg_out_30__20_), .A(n4574), .ZN(n4571) );
  OAI22_X2 U2689 ( .A1(n6221), .A2(n7531), .B1(n6670), .B2(n7523), .ZN(n4574)
         );
  AOI221_X2 U2691 ( .B1(n7488), .B2(REG_FILE_reg_out_3__20_), .C1(n7496), .C2(
        REG_FILE_reg_out_7__20_), .A(n4577), .ZN(n4576) );
  OAI22_X2 U2692 ( .A1(n5950), .A2(n7548), .B1(n6472), .B2(n7540), .ZN(n4577)
         );
  AOI221_X2 U2693 ( .B1(n7504), .B2(REG_FILE_reg_out_2__20_), .C1(n7512), .C2(
        REG_FILE_reg_out_6__20_), .A(n4578), .ZN(n4575) );
  OAI22_X2 U2694 ( .A1(n6220), .A2(n7531), .B1(n6669), .B2(n7523), .ZN(n4578)
         );
  OAI22_X2 U2696 ( .A1(n7064), .A2(n7531), .B1(n6668), .B2(n7523), .ZN(n4582)
         );
  OAI22_X2 U2697 ( .A1(n6935), .A2(n7515), .B1(n6427), .B2(n7507), .ZN(n4581)
         );
  OAI22_X2 U2698 ( .A1(n6934), .A2(n7548), .B1(n6426), .B2(n7540), .ZN(n4580)
         );
  OAI22_X2 U2699 ( .A1(n7063), .A2(n7499), .B1(n6667), .B2(n7491), .ZN(n4579)
         );
  AOI221_X2 U2704 ( .B1(n7487), .B2(REG_FILE_reg_out_11__21_), .C1(n7497), 
        .C2(REG_FILE_reg_out_15__21_), .A(n4591), .ZN(n4590) );
  OAI22_X2 U2705 ( .A1(n6933), .A2(n7547), .B1(n6425), .B2(n7541), .ZN(n4591)
         );
  AOI221_X2 U2706 ( .B1(n7503), .B2(REG_FILE_reg_out_10__21_), .C1(n7513), 
        .C2(REG_FILE_reg_out_14__21_), .A(n4592), .ZN(n4589) );
  OAI22_X2 U2707 ( .A1(n7062), .A2(n7530), .B1(n6666), .B2(n7523), .ZN(n4592)
         );
  AOI221_X2 U2709 ( .B1(n7487), .B2(REG_FILE_reg_out_27__21_), .C1(n7497), 
        .C2(REG_FILE_reg_out_31__21_), .A(n4595), .ZN(n4594) );
  OAI22_X2 U2710 ( .A1(n6070), .A2(n7547), .B1(n6424), .B2(n7541), .ZN(n4595)
         );
  AOI221_X2 U2711 ( .B1(n7503), .B2(REG_FILE_reg_out_26__21_), .C1(n7513), 
        .C2(REG_FILE_reg_out_30__21_), .A(n4596), .ZN(n4593) );
  OAI22_X2 U2712 ( .A1(n6219), .A2(n7530), .B1(n6665), .B2(n7523), .ZN(n4596)
         );
  AOI221_X2 U2714 ( .B1(n7486), .B2(REG_FILE_reg_out_3__21_), .C1(n7497), .C2(
        REG_FILE_reg_out_7__21_), .A(n4599), .ZN(n4598) );
  OAI22_X2 U2715 ( .A1(n6121), .A2(n7547), .B1(n6471), .B2(n7541), .ZN(n4599)
         );
  AOI221_X2 U2716 ( .B1(n7502), .B2(REG_FILE_reg_out_2__21_), .C1(n7513), .C2(
        REG_FILE_reg_out_6__21_), .A(n4600), .ZN(n4597) );
  OAI22_X2 U2717 ( .A1(n6218), .A2(n7530), .B1(n6664), .B2(n7523), .ZN(n4600)
         );
  OAI22_X2 U2719 ( .A1(n7061), .A2(n7530), .B1(n6663), .B2(n7524), .ZN(n4604)
         );
  OAI22_X2 U2720 ( .A1(n6932), .A2(n7515), .B1(n6423), .B2(n7507), .ZN(n4603)
         );
  OAI22_X2 U2721 ( .A1(n6931), .A2(n7547), .B1(n6422), .B2(n7541), .ZN(n4602)
         );
  OAI22_X2 U2722 ( .A1(n7060), .A2(n7499), .B1(n6662), .B2(n7491), .ZN(n4601)
         );
  AOI221_X2 U2727 ( .B1(n7487), .B2(REG_FILE_reg_out_11__22_), .C1(n7497), 
        .C2(REG_FILE_reg_out_15__22_), .A(n4614), .ZN(n4613) );
  OAI22_X2 U2728 ( .A1(n6930), .A2(n7547), .B1(n6421), .B2(n7541), .ZN(n4614)
         );
  AOI221_X2 U2729 ( .B1(n7503), .B2(REG_FILE_reg_out_10__22_), .C1(n7513), 
        .C2(REG_FILE_reg_out_14__22_), .A(n4615), .ZN(n4612) );
  OAI22_X2 U2730 ( .A1(n7059), .A2(n7530), .B1(n6661), .B2(n7524), .ZN(n4615)
         );
  AOI221_X2 U2732 ( .B1(n7487), .B2(REG_FILE_reg_out_27__22_), .C1(n7497), 
        .C2(REG_FILE_reg_out_31__22_), .A(n4618), .ZN(n4617) );
  OAI22_X2 U2733 ( .A1(n6069), .A2(n7547), .B1(n6420), .B2(n7541), .ZN(n4618)
         );
  AOI221_X2 U2734 ( .B1(n7503), .B2(REG_FILE_reg_out_26__22_), .C1(n7513), 
        .C2(REG_FILE_reg_out_30__22_), .A(n4619), .ZN(n4616) );
  OAI22_X2 U2735 ( .A1(n6217), .A2(n7530), .B1(n6660), .B2(n7524), .ZN(n4619)
         );
  AOI221_X2 U2737 ( .B1(n7487), .B2(REG_FILE_reg_out_3__22_), .C1(n7497), .C2(
        REG_FILE_reg_out_7__22_), .A(n4622), .ZN(n4621) );
  OAI22_X2 U2738 ( .A1(n6120), .A2(n7547), .B1(n6470), .B2(n7541), .ZN(n4622)
         );
  AOI221_X2 U2739 ( .B1(n7503), .B2(REG_FILE_reg_out_2__22_), .C1(n7513), .C2(
        REG_FILE_reg_out_6__22_), .A(n4623), .ZN(n4620) );
  OAI22_X2 U2740 ( .A1(n6216), .A2(n7530), .B1(n6659), .B2(n7524), .ZN(n4623)
         );
  OAI22_X2 U2742 ( .A1(n7058), .A2(n7530), .B1(n6658), .B2(n7524), .ZN(n4627)
         );
  OAI22_X2 U2743 ( .A1(n6929), .A2(n7515), .B1(n6419), .B2(n7507), .ZN(n4626)
         );
  OAI22_X2 U2744 ( .A1(n6928), .A2(n7547), .B1(n6418), .B2(n7541), .ZN(n4625)
         );
  OAI22_X2 U2745 ( .A1(n7057), .A2(n7499), .B1(n6657), .B2(n7491), .ZN(n4624)
         );
  AOI221_X2 U2751 ( .B1(n7486), .B2(REG_FILE_reg_out_11__23_), .C1(n7497), 
        .C2(REG_FILE_reg_out_15__23_), .A(n4637), .ZN(n4636) );
  OAI22_X2 U2752 ( .A1(n6384), .A2(n7547), .B1(n6965), .B2(n7541), .ZN(n4637)
         );
  AOI221_X2 U2753 ( .B1(n7502), .B2(REG_FILE_reg_out_10__23_), .C1(n7513), 
        .C2(REG_FILE_reg_out_14__23_), .A(n4638), .ZN(n4635) );
  OAI22_X2 U2754 ( .A1(n7056), .A2(n7530), .B1(n6656), .B2(n7524), .ZN(n4638)
         );
  AOI221_X2 U2756 ( .B1(n7486), .B2(REG_FILE_reg_out_27__23_), .C1(n7497), 
        .C2(REG_FILE_reg_out_31__23_), .A(n4641), .ZN(n4640) );
  OAI22_X2 U2757 ( .A1(n6068), .A2(n7547), .B1(n6417), .B2(n7541), .ZN(n4641)
         );
  AOI221_X2 U2758 ( .B1(n7502), .B2(REG_FILE_reg_out_26__23_), .C1(n7513), 
        .C2(REG_FILE_reg_out_30__23_), .A(n4642), .ZN(n4639) );
  OAI22_X2 U2759 ( .A1(n6215), .A2(n7530), .B1(n6655), .B2(n7524), .ZN(n4642)
         );
  AOI221_X2 U2761 ( .B1(n7486), .B2(REG_FILE_reg_out_3__23_), .C1(n7497), .C2(
        REG_FILE_reg_out_7__23_), .A(n4645), .ZN(n4644) );
  OAI22_X2 U2762 ( .A1(n6453), .A2(n7547), .B1(n6982), .B2(n7541), .ZN(n4645)
         );
  AOI221_X2 U2763 ( .B1(n7502), .B2(REG_FILE_reg_out_2__23_), .C1(n7513), .C2(
        REG_FILE_reg_out_6__23_), .A(n4646), .ZN(n4643) );
  OAI22_X2 U2764 ( .A1(n6214), .A2(n7530), .B1(n6654), .B2(n7524), .ZN(n4646)
         );
  OAI22_X2 U2766 ( .A1(n7055), .A2(n7529), .B1(n6653), .B2(n7524), .ZN(n4650)
         );
  OAI22_X2 U2767 ( .A1(n6927), .A2(n7515), .B1(n6416), .B2(n7507), .ZN(n4649)
         );
  OAI22_X2 U2768 ( .A1(n6383), .A2(n7550), .B1(n6055), .B2(n7537), .ZN(n4648)
         );
  OAI22_X2 U2769 ( .A1(n7054), .A2(n7499), .B1(n6652), .B2(n7491), .ZN(n4647)
         );
  AOI221_X2 U2774 ( .B1(n7486), .B2(REG_FILE_reg_out_11__24_), .C1(n7497), 
        .C2(REG_FILE_reg_out_15__24_), .A(n4659), .ZN(n4658) );
  OAI22_X2 U2775 ( .A1(n6067), .A2(n7550), .B1(n6415), .B2(n7537), .ZN(n4659)
         );
  AOI221_X2 U2776 ( .B1(n7502), .B2(REG_FILE_reg_out_10__24_), .C1(n7513), 
        .C2(REG_FILE_reg_out_14__24_), .A(n4660), .ZN(n4657) );
  OAI22_X2 U2777 ( .A1(n6585), .A2(n7529), .B1(n7117), .B2(n7524), .ZN(n4660)
         );
  AOI221_X2 U2779 ( .B1(n7486), .B2(REG_FILE_reg_out_27__24_), .C1(n7497), 
        .C2(REG_FILE_reg_out_31__24_), .A(n4663), .ZN(n4662) );
  OAI22_X2 U2780 ( .A1(n6066), .A2(n7551), .B1(n6414), .B2(n7537), .ZN(n4663)
         );
  AOI221_X2 U2781 ( .B1(n7502), .B2(REG_FILE_reg_out_26__24_), .C1(n7513), 
        .C2(REG_FILE_reg_out_30__24_), .A(n4664), .ZN(n4661) );
  OAI22_X2 U2782 ( .A1(n6584), .A2(n7529), .B1(n7116), .B2(n7524), .ZN(n4664)
         );
  AOI221_X2 U2784 ( .B1(n7487), .B2(REG_FILE_reg_out_3__24_), .C1(n7496), .C2(
        REG_FILE_reg_out_7__24_), .A(n4667), .ZN(n4666) );
  OAI22_X2 U2785 ( .A1(n6119), .A2(n7551), .B1(n6469), .B2(n7537), .ZN(n4667)
         );
  AOI221_X2 U2786 ( .B1(n7503), .B2(REG_FILE_reg_out_2__24_), .C1(n7512), .C2(
        REG_FILE_reg_out_6__24_), .A(n4668), .ZN(n4665) );
  OAI22_X2 U2787 ( .A1(n7053), .A2(n7529), .B1(n6651), .B2(n7524), .ZN(n4668)
         );
  OAI22_X2 U2789 ( .A1(n6213), .A2(n7529), .B1(n6650), .B2(n7524), .ZN(n4672)
         );
  OAI22_X2 U2790 ( .A1(n6382), .A2(n7515), .B1(n6964), .B2(n7507), .ZN(n4671)
         );
  OAI22_X2 U2791 ( .A1(n6065), .A2(n7550), .B1(n6413), .B2(n7537), .ZN(n4670)
         );
  OAI22_X2 U2792 ( .A1(n6583), .A2(n7499), .B1(n7115), .B2(n7491), .ZN(n4669)
         );
  AOI221_X2 U2797 ( .B1(n7487), .B2(REG_FILE_reg_out_11__25_), .C1(n7496), 
        .C2(REG_FILE_reg_out_15__25_), .A(n4682), .ZN(n4681) );
  OAI22_X2 U2798 ( .A1(n6064), .A2(n7550), .B1(n6412), .B2(n7539), .ZN(n4682)
         );
  AOI221_X2 U2799 ( .B1(n7503), .B2(REG_FILE_reg_out_10__25_), .C1(n7512), 
        .C2(REG_FILE_reg_out_14__25_), .A(n4683), .ZN(n4680) );
  OAI22_X2 U2800 ( .A1(n6582), .A2(n7533), .B1(n7114), .B2(n7524), .ZN(n4683)
         );
  AOI221_X2 U2802 ( .B1(n7487), .B2(REG_FILE_reg_out_27__25_), .C1(n7496), 
        .C2(REG_FILE_reg_out_31__25_), .A(n4686), .ZN(n4685) );
  OAI22_X2 U2803 ( .A1(n5895), .A2(n7551), .B1(n6103), .B2(n7537), .ZN(n4686)
         );
  AOI221_X2 U2804 ( .B1(n7503), .B2(REG_FILE_reg_out_26__25_), .C1(n7512), 
        .C2(REG_FILE_reg_out_30__25_), .A(n4687), .ZN(n4684) );
  OAI22_X2 U2805 ( .A1(n6212), .A2(n7528), .B1(n7113), .B2(n7524), .ZN(n4687)
         );
  AOI221_X2 U2807 ( .B1(n7487), .B2(REG_FILE_reg_out_3__25_), .C1(n7496), .C2(
        REG_FILE_reg_out_7__25_), .A(n4690), .ZN(n4689) );
  OAI22_X2 U2808 ( .A1(n6452), .A2(n7550), .B1(n6125), .B2(n7537), .ZN(n4690)
         );
  AOI221_X2 U2809 ( .B1(n7503), .B2(REG_FILE_reg_out_2__25_), .C1(n7512), .C2(
        REG_FILE_reg_out_6__25_), .A(n4691), .ZN(n4688) );
  OAI22_X2 U2810 ( .A1(n6581), .A2(n7528), .B1(n7082), .B2(n7524), .ZN(n4691)
         );
  OAI22_X2 U2812 ( .A1(n6580), .A2(n7528), .B1(n7081), .B2(n7524), .ZN(n4695)
         );
  OAI22_X2 U2813 ( .A1(n6381), .A2(n7515), .B1(n6963), .B2(n7507), .ZN(n4694)
         );
  OAI22_X2 U2814 ( .A1(n6380), .A2(n7551), .B1(n6054), .B2(n7537), .ZN(n4693)
         );
  OAI22_X2 U2815 ( .A1(n6579), .A2(n7499), .B1(n7112), .B2(n7491), .ZN(n4692)
         );
  AOI221_X2 U2820 ( .B1(n7487), .B2(REG_FILE_reg_out_11__26_), .C1(n7496), 
        .C2(REG_FILE_reg_out_15__26_), .A(n4705), .ZN(n4704) );
  OAI22_X2 U2821 ( .A1(n6063), .A2(n7551), .B1(n6411), .B2(n7537), .ZN(n4705)
         );
  AOI221_X2 U2822 ( .B1(n7503), .B2(REG_FILE_reg_out_10__26_), .C1(n7512), 
        .C2(REG_FILE_reg_out_14__26_), .A(n4706), .ZN(n4703) );
  OAI22_X2 U2823 ( .A1(n7052), .A2(n7533), .B1(n6649), .B2(n7524), .ZN(n4706)
         );
  AOI221_X2 U2825 ( .B1(n7487), .B2(REG_FILE_reg_out_27__26_), .C1(n7496), 
        .C2(REG_FILE_reg_out_31__26_), .A(n4709), .ZN(n4708) );
  OAI22_X2 U2826 ( .A1(n5875), .A2(n7550), .B1(n5896), .B2(n7537), .ZN(n4709)
         );
  AOI221_X2 U2827 ( .B1(n7503), .B2(REG_FILE_reg_out_26__26_), .C1(n7512), 
        .C2(REG_FILE_reg_out_30__26_), .A(n4710), .ZN(n4707) );
  OAI22_X2 U2828 ( .A1(n6211), .A2(n7528), .B1(n7111), .B2(n7525), .ZN(n4710)
         );
  AOI221_X2 U2830 ( .B1(n7487), .B2(REG_FILE_reg_out_3__26_), .C1(n7496), .C2(
        REG_FILE_reg_out_7__26_), .A(n4713), .ZN(n4712) );
  OAI22_X2 U2831 ( .A1(n6451), .A2(n7549), .B1(n6981), .B2(n7540), .ZN(n4713)
         );
  AOI221_X2 U2832 ( .B1(n7503), .B2(REG_FILE_reg_out_2__26_), .C1(n7512), .C2(
        REG_FILE_reg_out_6__26_), .A(n4714), .ZN(n4711) );
  OAI22_X2 U2833 ( .A1(n6578), .A2(n7529), .B1(n7080), .B2(n7525), .ZN(n4714)
         );
  OAI22_X2 U2835 ( .A1(n6577), .A2(n7529), .B1(n7079), .B2(n7525), .ZN(n4718)
         );
  OAI22_X2 U2836 ( .A1(n6926), .A2(n7515), .B1(n6410), .B2(n7507), .ZN(n4717)
         );
  OAI22_X2 U2837 ( .A1(n6925), .A2(n7549), .B1(n5933), .B2(n7540), .ZN(n4716)
         );
  OAI22_X2 U2838 ( .A1(n7051), .A2(n7499), .B1(n6648), .B2(n7491), .ZN(n4715)
         );
  AOI221_X2 U2845 ( .B1(n7487), .B2(REG_FILE_reg_out_11__27_), .C1(n7496), 
        .C2(REG_FILE_reg_out_15__27_), .A(n4728), .ZN(n4727) );
  OAI22_X2 U2846 ( .A1(n6924), .A2(n7547), .B1(n5947), .B2(n7540), .ZN(n4728)
         );
  AOI221_X2 U2847 ( .B1(n7503), .B2(REG_FILE_reg_out_10__27_), .C1(n7512), 
        .C2(REG_FILE_reg_out_14__27_), .A(n4729), .ZN(n4726) );
  OAI22_X2 U2848 ( .A1(n7050), .A2(n7529), .B1(n6647), .B2(n7525), .ZN(n4729)
         );
  AOI221_X2 U2850 ( .B1(n7487), .B2(REG_FILE_reg_out_27__27_), .C1(n7496), 
        .C2(REG_FILE_reg_out_31__27_), .A(n4732), .ZN(n4731) );
  OAI22_X2 U2851 ( .A1(n5874), .A2(n7547), .B1(n5946), .B2(n7540), .ZN(n4732)
         );
  AOI221_X2 U2852 ( .B1(n7503), .B2(REG_FILE_reg_out_26__27_), .C1(n7512), 
        .C2(REG_FILE_reg_out_30__27_), .A(n4733), .ZN(n4730) );
  OAI22_X2 U2853 ( .A1(n6210), .A2(n7529), .B1(n6646), .B2(n7525), .ZN(n4733)
         );
  AOI221_X2 U2855 ( .B1(n7487), .B2(REG_FILE_reg_out_3__27_), .C1(n7496), .C2(
        REG_FILE_reg_out_7__27_), .A(n4736), .ZN(n4735) );
  OAI22_X2 U2856 ( .A1(n5949), .A2(n7547), .B1(n6131), .B2(n7540), .ZN(n4736)
         );
  AOI221_X2 U2857 ( .B1(n7503), .B2(REG_FILE_reg_out_2__27_), .C1(n7512), .C2(
        REG_FILE_reg_out_6__27_), .A(n4737), .ZN(n4734) );
  OAI22_X2 U2858 ( .A1(n6576), .A2(n7529), .B1(n7110), .B2(n7525), .ZN(n4737)
         );
  OAI22_X2 U2860 ( .A1(n6575), .A2(n7529), .B1(n7109), .B2(n7525), .ZN(n4741)
         );
  OAI22_X2 U2861 ( .A1(n6923), .A2(n7515), .B1(n6409), .B2(n7507), .ZN(n4740)
         );
  OAI22_X2 U2862 ( .A1(n5935), .A2(n7547), .B1(n6962), .B2(n7540), .ZN(n4739)
         );
  OAI22_X2 U2863 ( .A1(n7049), .A2(n7499), .B1(n6645), .B2(n7491), .ZN(n4738)
         );
  AOI221_X2 U2869 ( .B1(n7487), .B2(REG_FILE_reg_out_11__28_), .C1(n7496), 
        .C2(REG_FILE_reg_out_15__28_), .A(n4750), .ZN(n4749) );
  OAI22_X2 U2870 ( .A1(n5873), .A2(n7549), .B1(n6961), .B2(n7540), .ZN(n4750)
         );
  AOI221_X2 U2871 ( .B1(n7503), .B2(REG_FILE_reg_out_10__28_), .C1(n7512), 
        .C2(REG_FILE_reg_out_14__28_), .A(n4751), .ZN(n4748) );
  OAI22_X2 U2872 ( .A1(n6574), .A2(n7529), .B1(n7108), .B2(n7525), .ZN(n4751)
         );
  AOI221_X2 U2874 ( .B1(n7486), .B2(REG_FILE_reg_out_27__28_), .C1(n7495), 
        .C2(REG_FILE_reg_out_31__28_), .A(n4754), .ZN(n4753) );
  OAI22_X2 U2875 ( .A1(n5934), .A2(n7549), .B1(n6960), .B2(n7540), .ZN(n4754)
         );
  AOI221_X2 U2876 ( .B1(n7502), .B2(REG_FILE_reg_out_26__28_), .C1(n7511), 
        .C2(REG_FILE_reg_out_30__28_), .A(n4755), .ZN(n4752) );
  OAI22_X2 U2877 ( .A1(n6573), .A2(n7529), .B1(n7107), .B2(n7525), .ZN(n4755)
         );
  AOI221_X2 U2879 ( .B1(n7486), .B2(REG_FILE_reg_out_3__28_), .C1(n7495), .C2(
        REG_FILE_reg_out_7__28_), .A(n4758), .ZN(n4757) );
  OAI22_X2 U2880 ( .A1(n5882), .A2(n7547), .B1(n6124), .B2(n7540), .ZN(n4758)
         );
  AOI221_X2 U2881 ( .B1(n7502), .B2(REG_FILE_reg_out_2__28_), .C1(n7511), .C2(
        REG_FILE_reg_out_6__28_), .A(n4759), .ZN(n4756) );
  OAI22_X2 U2882 ( .A1(n6572), .A2(n7529), .B1(n7078), .B2(n7525), .ZN(n4759)
         );
  OAI22_X2 U2884 ( .A1(n6571), .A2(n7529), .B1(n7077), .B2(n7525), .ZN(n4763)
         );
  OAI22_X2 U2885 ( .A1(n6379), .A2(n7515), .B1(n6959), .B2(n7507), .ZN(n4762)
         );
  OAI22_X2 U2886 ( .A1(n5872), .A2(n7549), .B1(n6920), .B2(n7540), .ZN(n4761)
         );
  OAI22_X2 U2887 ( .A1(n6570), .A2(n7499), .B1(n7106), .B2(n7491), .ZN(n4760)
         );
  AOI221_X2 U2893 ( .B1(n7486), .B2(REG_FILE_reg_out_11__29_), .C1(n7495), 
        .C2(REG_FILE_reg_out_15__29_), .A(n4772), .ZN(n4771) );
  OAI22_X2 U2894 ( .A1(n5871), .A2(n7549), .B1(n6958), .B2(n7540), .ZN(n4772)
         );
  AOI221_X2 U2895 ( .B1(n7502), .B2(REG_FILE_reg_out_10__29_), .C1(n7511), 
        .C2(REG_FILE_reg_out_14__29_), .A(n4773), .ZN(n4770) );
  OAI22_X2 U2896 ( .A1(n6569), .A2(n7529), .B1(n7105), .B2(n7525), .ZN(n4773)
         );
  AOI221_X2 U2898 ( .B1(n7486), .B2(REG_FILE_reg_out_27__29_), .C1(n7495), 
        .C2(REG_FILE_reg_out_31__29_), .A(n4776), .ZN(n4775) );
  OAI22_X2 U2899 ( .A1(n6378), .A2(n7546), .B1(n6957), .B2(n7539), .ZN(n4776)
         );
  AOI221_X2 U2900 ( .B1(n7502), .B2(REG_FILE_reg_out_26__29_), .C1(n7511), 
        .C2(REG_FILE_reg_out_30__29_), .A(n4777), .ZN(n4774) );
  OAI22_X2 U2901 ( .A1(n6568), .A2(n7528), .B1(n7104), .B2(n7525), .ZN(n4777)
         );
  AOI221_X2 U2903 ( .B1(n7486), .B2(REG_FILE_reg_out_3__29_), .C1(n7495), .C2(
        REG_FILE_reg_out_7__29_), .A(n4780), .ZN(n4779) );
  OAI22_X2 U2904 ( .A1(n5899), .A2(n7546), .B1(n6123), .B2(n7539), .ZN(n4780)
         );
  AOI221_X2 U2905 ( .B1(n7502), .B2(REG_FILE_reg_out_2__29_), .C1(n7511), .C2(
        REG_FILE_reg_out_6__29_), .A(n4781), .ZN(n4778) );
  OAI22_X2 U2906 ( .A1(n6567), .A2(n7528), .B1(n7076), .B2(n7525), .ZN(n4781)
         );
  OAI22_X2 U2908 ( .A1(n6566), .A2(n7528), .B1(n7075), .B2(n7525), .ZN(n4785)
         );
  OAI22_X2 U2909 ( .A1(n6377), .A2(n7515), .B1(n6956), .B2(n7507), .ZN(n4784)
         );
  OAI22_X2 U2910 ( .A1(n6376), .A2(n7546), .B1(n6919), .B2(n7539), .ZN(n4783)
         );
  OAI22_X2 U2911 ( .A1(n6565), .A2(n7499), .B1(n7103), .B2(n7491), .ZN(n4782)
         );
  AOI221_X2 U2917 ( .B1(n7486), .B2(REG_FILE_reg_out_11__30_), .C1(n7495), 
        .C2(REG_FILE_reg_out_15__30_), .A(n4794), .ZN(n4793) );
  OAI22_X2 U2918 ( .A1(n6375), .A2(n7546), .B1(n6955), .B2(n7539), .ZN(n4794)
         );
  AOI221_X2 U2919 ( .B1(n7502), .B2(REG_FILE_reg_out_10__30_), .C1(n7511), 
        .C2(REG_FILE_reg_out_14__30_), .A(n4795), .ZN(n4792) );
  OAI22_X2 U2920 ( .A1(n6564), .A2(n7528), .B1(n7102), .B2(n7525), .ZN(n4795)
         );
  AOI221_X2 U2922 ( .B1(n7486), .B2(REG_FILE_reg_out_27__30_), .C1(n7495), 
        .C2(REG_FILE_reg_out_31__30_), .A(n4798), .ZN(n4797) );
  OAI22_X2 U2923 ( .A1(n6374), .A2(n7546), .B1(n6954), .B2(n7539), .ZN(n4798)
         );
  AOI221_X2 U2924 ( .B1(n7502), .B2(REG_FILE_reg_out_26__30_), .C1(n7511), 
        .C2(REG_FILE_reg_out_30__30_), .A(n4799), .ZN(n4796) );
  OAI22_X2 U2925 ( .A1(n6563), .A2(n7528), .B1(n7101), .B2(n7525), .ZN(n4799)
         );
  AOI221_X2 U2927 ( .B1(n7486), .B2(REG_FILE_reg_out_3__30_), .C1(n7495), .C2(
        REG_FILE_reg_out_7__30_), .A(n4802), .ZN(n4801) );
  OAI22_X2 U2928 ( .A1(n5898), .A2(n7546), .B1(n6130), .B2(n7539), .ZN(n4802)
         );
  AOI221_X2 U2929 ( .B1(n7502), .B2(REG_FILE_reg_out_2__30_), .C1(n7511), .C2(
        REG_FILE_reg_out_6__30_), .A(n4803), .ZN(n4800) );
  OAI22_X2 U2930 ( .A1(n7048), .A2(n7528), .B1(n6644), .B2(n7525), .ZN(n4803)
         );
  OAI22_X2 U2932 ( .A1(n6209), .A2(n7528), .B1(n6643), .B2(n7522), .ZN(n4807)
         );
  OAI22_X2 U2933 ( .A1(n6373), .A2(n7515), .B1(n6953), .B2(n7507), .ZN(n4806)
         );
  OAI22_X2 U2934 ( .A1(n6062), .A2(n7546), .B1(n6408), .B2(n7539), .ZN(n4805)
         );
  OAI22_X2 U2935 ( .A1(n6562), .A2(n7499), .B1(n7100), .B2(n7491), .ZN(n4804)
         );
  OR2_X2 U2939 ( .A1(n3368), .A2(n6346), .ZN(n3351) );
  OR2_X2 U2940 ( .A1(n3363), .A2(IF_ID_OUT[33]), .ZN(n3368) );
  NOR4_X2 U2948 ( .A1(n4812), .A2(n4813), .A3(ID_STAGE_imm16_aluA[23]), .A4(
        ID_STAGE_imm16_aluA[22]), .ZN(n4811) );
  OR3_X2 U2949 ( .A1(ID_STAGE_imm16_aluA[25]), .A2(ID_STAGE_imm16_aluA[29]), 
        .A3(ID_STAGE_imm16_aluA[24]), .ZN(n4813) );
  NAND4_X2 U2950 ( .A1(n6347), .A2(n6886), .A3(n6011), .A4(n4814), .ZN(n4812)
         );
  NOR4_X2 U2952 ( .A1(n4815), .A2(ID_STAGE_imm16_aluA[16]), .A3(
        ID_STAGE_imm16_aluA[18]), .A4(ID_STAGE_imm16_aluA[17]), .ZN(n4810) );
  NOR3_X4 U2954 ( .A1(n3366), .A2(n4449), .A3(n3364), .ZN(n4809) );
  NAND2_X2 U2955 ( .A1(n6864), .A2(n6346), .ZN(n3364) );
  NAND2_X2 U2956 ( .A1(n3329), .A2(n6343), .ZN(n4449) );
  NAND2_X2 U2957 ( .A1(n3375), .A2(n6012), .ZN(n3366) );
  NAND2_X2 U2960 ( .A1(n4089), .A2(n5857), .ZN(n4090) );
  AOI221_X2 U2967 ( .B1(n7486), .B2(REG_FILE_reg_out_11__31_), .C1(n7495), 
        .C2(REG_FILE_reg_out_15__31_), .A(n4824), .ZN(n4822) );
  OAI22_X2 U2968 ( .A1(n6061), .A2(n7546), .B1(n6407), .B2(n7539), .ZN(n4824)
         );
  AOI221_X2 U2969 ( .B1(n7502), .B2(REG_FILE_reg_out_10__31_), .C1(n7511), 
        .C2(REG_FILE_reg_out_14__31_), .A(n4825), .ZN(n4821) );
  OAI22_X2 U2970 ( .A1(n6208), .A2(n7528), .B1(n6642), .B2(n7522), .ZN(n4825)
         );
  AND2_X2 U2973 ( .A1(offset_26_id[6]), .A2(n4100), .ZN(n4823) );
  AOI221_X2 U2974 ( .B1(n7486), .B2(REG_FILE_reg_out_27__31_), .C1(n7495), 
        .C2(REG_FILE_reg_out_31__31_), .A(n4828), .ZN(n4827) );
  OAI22_X2 U2975 ( .A1(n6372), .A2(n7546), .B1(n6952), .B2(n7539), .ZN(n4828)
         );
  AOI221_X2 U2976 ( .B1(n7502), .B2(REG_FILE_reg_out_26__31_), .C1(n7511), 
        .C2(REG_FILE_reg_out_30__31_), .A(n4829), .ZN(n4826) );
  OAI22_X2 U2977 ( .A1(n6207), .A2(n7528), .B1(n6641), .B2(n7522), .ZN(n4829)
         );
  AOI221_X2 U2980 ( .B1(n7486), .B2(REG_FILE_reg_out_3__31_), .C1(n7495), .C2(
        REG_FILE_reg_out_7__31_), .A(n4833), .ZN(n4831) );
  OAI22_X2 U2981 ( .A1(n6118), .A2(n7546), .B1(n6468), .B2(n7539), .ZN(n4833)
         );
  AOI221_X2 U2982 ( .B1(n7502), .B2(REG_FILE_reg_out_2__31_), .C1(n7511), .C2(
        REG_FILE_reg_out_6__31_), .A(n4834), .ZN(n4830) );
  OAI22_X2 U2983 ( .A1(n5985), .A2(n7528), .B1(n6640), .B2(n7522), .ZN(n4834)
         );
  NAND2_X2 U2984 ( .A1(n4832), .A2(offset_26_id[5]), .ZN(n4099) );
  AND2_X2 U2985 ( .A1(n4100), .A2(n6351), .ZN(n4832) );
  OAI22_X2 U2994 ( .A1(n5906), .A2(n7528), .B1(n6639), .B2(n7524), .ZN(n4844)
         );
  OAI22_X2 U2997 ( .A1(n6371), .A2(n7515), .B1(n6951), .B2(n7507), .ZN(n4843)
         );
  NAND2_X2 U2998 ( .A1(n4845), .A2(n1641), .ZN(n4129) );
  OAI22_X2 U3001 ( .A1(n6060), .A2(n7546), .B1(n6406), .B2(n7539), .ZN(n4842)
         );
  NAND2_X2 U3002 ( .A1(n4846), .A2(n1641), .ZN(n4110) );
  OAI22_X2 U3005 ( .A1(n6561), .A2(n7499), .B1(n7099), .B2(n7491), .ZN(n4841)
         );
  NAND2_X2 U3006 ( .A1(n4847), .A2(n1641), .ZN(n4131) );
  NAND2_X2 U3012 ( .A1(ID_STAGE_imm16_aluA[18]), .A2(n7305), .ZN(n4516) );
  NAND2_X2 U3016 ( .A1(ID_STAGE_imm16_aluA[22]), .A2(n7774), .ZN(n4605) );
  NAND2_X2 U3017 ( .A1(ID_STAGE_imm16_aluA[23]), .A2(n7774), .ZN(n4628) );
  NAND2_X2 U3019 ( .A1(ID_STAGE_imm16_aluA[25]), .A2(n7774), .ZN(n4673) );
  NAND2_X2 U3020 ( .A1(ID_STAGE_imm16_aluA[26]), .A2(n7774), .ZN(n4696) );
  AND2_X2 U3327 ( .A1(EXEC_MEM_IN[101]), .A2(n7774), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N81) );
  AND2_X2 U3328 ( .A1(EXEC_MEM_IN[103]), .A2(n7774), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N79) );
  AND2_X2 U3329 ( .A1(EXEC_MEM_IN[104]), .A2(n7774), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N78) );
  AND2_X2 U3331 ( .A1(EXEC_MEM_IN[106]), .A2(n7774), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N76) );
  AND2_X2 U3332 ( .A1(DSize_ex_out[0]), .A2(n7774), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N75) );
  AND2_X2 U3333 ( .A1(DSize_ex_out[1]), .A2(n7774), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N74) );
  XOR2_X2 U3491 ( .A(n5400), .B(ID_EXEC_OUT[147]), .Z(n5399) );
  OAI221_X2 U3503 ( .B1(n6817), .B2(n5908), .C1(n5888), .C2(n7483), .A(n5411), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N40) );
  NAND2_X2 U3504 ( .A1(ID_EXEC_OUT[160]), .A2(n10300), .ZN(n5411) );
  OAI221_X2 U3505 ( .B1(n7034), .B2(n5908), .C1(n5948), .C2(n7484), .A(n5412), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N39) );
  NAND2_X2 U3506 ( .A1(ID_EXEC_OUT[161]), .A2(n10300), .ZN(n5412) );
  OAI221_X2 U3507 ( .B1(n6827), .B2(n5908), .C1(n5926), .C2(n7483), .A(n5413), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N38) );
  NAND2_X2 U3508 ( .A1(ID_EXEC_OUT[162]), .A2(n10300), .ZN(n5413) );
  OAI221_X2 U3509 ( .B1(n6826), .B2(n5908), .C1(n5952), .C2(n7484), .A(n5414), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N37) );
  NAND2_X2 U3510 ( .A1(ID_EXEC_OUT[163]), .A2(n10300), .ZN(n5414) );
  OAI221_X2 U3511 ( .B1(n6816), .B2(n5908), .C1(n5925), .C2(n7483), .A(n5415), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N36) );
  NAND2_X2 U3512 ( .A1(ID_EXEC_OUT[164]), .A2(n10300), .ZN(n5415) );
  OAI221_X2 U3513 ( .B1(n6815), .B2(n5908), .C1(n5914), .C2(n7484), .A(n5416), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N35) );
  NAND2_X2 U3514 ( .A1(ID_EXEC_OUT[165]), .A2(n10300), .ZN(n5416) );
  OAI221_X2 U3515 ( .B1(n6814), .B2(n5908), .C1(n5921), .C2(n7483), .A(n5417), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N34) );
  NAND2_X2 U3516 ( .A1(ID_EXEC_OUT[166]), .A2(n10300), .ZN(n5417) );
  OAI221_X2 U3517 ( .B1(n6825), .B2(n5908), .C1(n5920), .C2(n7484), .A(n5418), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N33) );
  NAND2_X2 U3518 ( .A1(ID_EXEC_OUT[167]), .A2(n10300), .ZN(n5418) );
  OAI221_X2 U3519 ( .B1(n7033), .B2(n5908), .C1(n5922), .C2(n7484), .A(n5419), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N32) );
  NAND2_X2 U3520 ( .A1(ID_EXEC_OUT[168]), .A2(n10300), .ZN(n5419) );
  OAI221_X2 U3521 ( .B1(n6824), .B2(n5908), .C1(n5953), .C2(n7484), .A(n5420), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N31) );
  NAND2_X2 U3522 ( .A1(ID_EXEC_OUT[169]), .A2(n10300), .ZN(n5420) );
  OAI221_X2 U3523 ( .B1(n6823), .B2(n5908), .C1(n5923), .C2(n7484), .A(n5421), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N30) );
  NAND2_X2 U3524 ( .A1(ID_EXEC_OUT[170]), .A2(n10300), .ZN(n5421) );
  AND2_X2 U3561 ( .A1(destReg_ex_out[0]), .A2(n7774), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N118) );
  AND2_X2 U3562 ( .A1(destReg_ex_out[1]), .A2(n7774), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N117) );
  AND2_X2 U3563 ( .A1(destReg_ex_out[2]), .A2(n7774), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N116) );
  AND2_X2 U3564 ( .A1(destReg_ex_out[3]), .A2(n7774), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N115) );
  AND2_X2 U3565 ( .A1(destReg_ex_out[4]), .A2(n7774), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N114) );
  INV_X4 U4160 ( .A(n3188), .ZN(n1543) );
  INV_X4 U4161 ( .A(n3190), .ZN(n1544) );
  INV_X4 U4162 ( .A(n3192), .ZN(n1545) );
  INV_X4 U4163 ( .A(n3194), .ZN(n1546) );
  INV_X4 U4164 ( .A(n3196), .ZN(n1547) );
  INV_X4 U4165 ( .A(n3198), .ZN(n1548) );
  INV_X4 U4166 ( .A(n3200), .ZN(n1549) );
  INV_X4 U4167 ( .A(n3202), .ZN(n1550) );
  INV_X4 U4168 ( .A(n3204), .ZN(n1551) );
  INV_X4 U4169 ( .A(n3206), .ZN(n1552) );
  INV_X4 U4170 ( .A(n3210), .ZN(n1553) );
  INV_X4 U4171 ( .A(n3212), .ZN(n1554) );
  INV_X4 U4172 ( .A(n3214), .ZN(n1555) );
  INV_X4 U4173 ( .A(n3216), .ZN(n1556) );
  INV_X4 U4174 ( .A(n3218), .ZN(n1557) );
  INV_X4 U4175 ( .A(n3220), .ZN(n1558) );
  INV_X4 U4176 ( .A(n3222), .ZN(n1559) );
  INV_X4 U4177 ( .A(n3224), .ZN(n1560) );
  INV_X4 U4178 ( .A(n3226), .ZN(n1561) );
  INV_X4 U4179 ( .A(n3228), .ZN(n1562) );
  INV_X4 U4180 ( .A(n3170), .ZN(n1563) );
  INV_X4 U4181 ( .A(n3172), .ZN(n1564) );
  INV_X4 U4182 ( .A(n3174), .ZN(n1565) );
  INV_X4 U4183 ( .A(n3176), .ZN(n1566) );
  INV_X4 U4184 ( .A(n3178), .ZN(n1567) );
  INV_X4 U4185 ( .A(n3180), .ZN(n1568) );
  INV_X4 U4186 ( .A(n3182), .ZN(n1569) );
  INV_X4 U4187 ( .A(n3186), .ZN(n1570) );
  INV_X4 U4188 ( .A(n3208), .ZN(n1571) );
  INV_X4 U4189 ( .A(n3230), .ZN(n1572) );
  INV_X4 U4190 ( .A(n3303), .ZN(n1573) );
  INV_X4 U4191 ( .A(IMEM_BUS_IN[0]), .ZN(n1574) );
  INV_X4 U4192 ( .A(IMEM_BUS_IN[2]), .ZN(n1575) );
  INV_X4 U4193 ( .A(IMEM_BUS_IN[5]), .ZN(n1576) );
  INV_X4 U4194 ( .A(n3344), .ZN(n1577) );
  INV_X4 U4205 ( .A(n4447), .ZN(n1588) );
  INV_X4 U4206 ( .A(n3355), .ZN(n1589) );
  INV_X4 U4207 ( .A(n3370), .ZN(n1590) );
  INV_X4 U4210 ( .A(n3317), .ZN(n1593) );
  INV_X4 U4211 ( .A(n3366), .ZN(n1594) );
  INV_X4 U4215 ( .A(n3328), .ZN(n1598) );
  INV_X4 U4218 ( .A(n4696), .ZN(n1601) );
  INV_X4 U4219 ( .A(n4673), .ZN(n1602) );
  INV_X4 U4221 ( .A(n4628), .ZN(n1604) );
  INV_X4 U4222 ( .A(n4605), .ZN(n1605) );
  INV_X4 U4226 ( .A(n4516), .ZN(n1609) );
  INV_X4 U4269 ( .A(ID_EX_REG_ID_EX_REG_N94), .ZN(n1652) );
  INV_X4 U4271 ( .A(n3353), .ZN(n1654) );
  INV_X4 U4273 ( .A(ID_EX_REG_ID_EX_REG_N61), .ZN(n1656) );
  INV_X4 U4276 ( .A(n4449), .ZN(n1659) );
  INV_X4 U4277 ( .A(n3354), .ZN(n1660) );
  OAI33_X1 U5659 ( .A1(n3341), .A2(IF_ID_OUT[36]), .A3(n6347), .B1(n3347), 
        .B2(ID_STAGE_imm16_aluA[29]), .B3(n6012), .ZN(n3346) );
  OAI33_X1 U5660 ( .A1(n3347), .A2(n6867), .A3(n6012), .B1(n3362), .B2(n6343), 
        .B3(n3363), .ZN(n3340) );
  OAI33_X1 U5661 ( .A1(n3357), .A2(n6346), .A3(n6864), .B1(n3374), .B2(n6012), 
        .B3(n3358), .ZN(n3339) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_146_ ( .D(n1593), .CK(clk), .RN(n7779), 
        .QN(n7323) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_103_ ( .D(MEM_WB_REG_MEM_WB_REG_N7), 
        .CK(clk), .RN(n7791), .QN(n7223) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_105_ ( .D(DMEM_BUS_OUT[65]), .CK(clk), 
        .RN(n7789), .QN(n7308) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_106_ ( .D(DMEM_BUS_OUT[66]), .CK(clk), 
        .RN(n7792), .Q(MEM_WB_OUT[106]), .QN(n7329) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_157_ ( .D(ID_EX_REG_ID_EX_REG_N49), .CK(
        clk), .RN(n7780), .Q(ID_EXEC_OUT[157]), .QN(n6883) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_158_ ( .D(ID_EX_REG_ID_EX_REG_N48), .CK(
        clk), .RN(n7780), .Q(ID_EXEC_OUT[158]), .QN(n6013) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_159_ ( .D(ID_EX_REG_ID_EX_REG_N47), .CK(
        clk), .RN(n7780), .Q(ID_EXEC_OUT[159]), .QN(n7307) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_68_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N114), .CK(clk), .RN(n7790), .Q(
        MEM_WB_REG_MEM_WB_REG_N74), .QN(n7331) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_65_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N117), .CK(clk), .RN(n7790), .Q(
        MEM_WB_REG_MEM_WB_REG_N77), .QN(n7349) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_66_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N116), .CK(clk), .RN(n7790), .Q(
        MEM_WB_REG_MEM_WB_REG_N76), .QN(n7333) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_64_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N118), .CK(clk), .RN(n7790), .Q(
        MEM_WB_REG_MEM_WB_REG_N78) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_67_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N115), .CK(clk), .RN(n7790), .Q(
        MEM_WB_REG_MEM_WB_REG_N75) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_199_ ( .D(ID_EX_REG_ID_EX_REG_N88), .CK(
        clk), .RN(n7791), .Q(ID_EXEC_OUT[199]) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_63_ ( .D(IF_ID_REG_IF_ID_REG_N3), .CK(
        clk), .RN(n7787), .Q(ID_STAGE_imm16_aluA[31]), .QN(n6012) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_36_ ( .D(IF_ID_REG_IF_ID_REG_N30), .CK(
        clk), .RN(n7786), .Q(IF_ID_OUT[36]), .QN(n6864) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_34_ ( .D(MEM_WB_REG_MEM_WB_REG_N76), 
        .CK(clk), .RN(n7790), .Q(destReg_wb_out[2]), .QN(n7320) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_32_ ( .D(MEM_WB_REG_MEM_WB_REG_N78), 
        .CK(clk), .RN(n7790), .Q(destReg_wb_out[0]), .QN(n6349) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_33_ ( .D(MEM_WB_REG_MEM_WB_REG_N77), 
        .CK(clk), .RN(n7790), .QN(n6900) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_35_ ( .D(MEM_WB_REG_MEM_WB_REG_N75), 
        .CK(clk), .RN(n7790), .QN(n6345) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_192_ ( .D(ID_EX_REG_ID_EX_REG_N14), .CK(
        clk), .RN(n7778), .Q(ID_EXEC_OUT[192]), .QN(n6889) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_198_ ( .D(ID_EX_REG_ID_EX_REG_N89), .CK(
        clk), .RN(n7791), .Q(ID_EXEC_OUT[198]) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_101_ ( .D(MEM_WB_REG_MEM_WB_REG_N9), 
        .CK(clk), .RN(n7791), .QN(n7239) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_141_ ( .D(
        EX_MEM_REGISTER_EX_MEM_REG_N41), .CK(clk), .RN(n7793), .Q(
        EXEC_MEM_OUT_141), .QN(n7305) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_37_ ( .D(IF_ID_REG_IF_ID_REG_N29), .CK(
        clk), .RN(n7782), .Q(IF_ID_OUT[37]), .QN(n6346) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_61_ ( .D(IF_ID_REG_IF_ID_REG_N5), .CK(
        clk), .RN(n7780), .Q(ID_STAGE_imm16_aluA[29]), .QN(n6867) );
  NOR2_X4 U5663 ( .A1(n7993), .A2(n7034), .ZN(n9210) );
  INV_X4 U5664 ( .A(n7973), .ZN(n8095) );
  INV_X4 U5665 ( .A(n8005), .ZN(n9224) );
  OAI21_X4 U5666 ( .B1(n8075), .B2(n8074), .A(n8073), .ZN(n9260) );
  NOR2_X4 U5667 ( .A1(n7993), .A2(n7033), .ZN(n9239) );
  INV_X4 U5668 ( .A(n7999), .ZN(n8850) );
  OAI21_X4 U5671 ( .B1(n8075), .B2(n8060), .A(n8059), .ZN(n9290) );
  INV_X4 U5672 ( .A(n7907), .ZN(n8843) );
  NAND2_X2 U5675 ( .A1(n8016), .A2(n8015), .ZN(n8017) );
  NAND2_X2 U5676 ( .A1(MEM_WB_OUT[37]), .A2(n7941), .ZN(n8033) );
  NAND2_X2 U5677 ( .A1(MEM_WB_OUT[41]), .A2(n7363), .ZN(n8052) );
  NAND2_X2 U5678 ( .A1(MEM_WB_OUT[42]), .A2(n7855), .ZN(n7988) );
  NAND2_X2 U5679 ( .A1(MEM_WB_OUT[43]), .A2(n7889), .ZN(n7981) );
  NAND2_X2 U5680 ( .A1(MEM_WB_OUT[53]), .A2(n7357), .ZN(n7913) );
  NAND2_X2 U5681 ( .A1(MEM_WB_OUT[54]), .A2(n7363), .ZN(n7875) );
  NAND2_X2 U5682 ( .A1(MEM_WB_OUT[55]), .A2(n7363), .ZN(n7869) );
  NAND2_X2 U5683 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[19]), .A2(n7931), 
        .ZN(n7891) );
  NAND2_X2 U5684 ( .A1(MEM_WB_OUT[57]), .A2(n7364), .ZN(n7881) );
  NAND2_X2 U5685 ( .A1(MEM_WB_OUT[58]), .A2(n7941), .ZN(n7960) );
  NAND2_X2 U5686 ( .A1(MEM_WB_OUT[59]), .A2(n7361), .ZN(n7952) );
  INV_X4 U5687 ( .A(n7958), .ZN(n7935) );
  NAND2_X2 U5688 ( .A1(n7941), .A2(MEM_WB_OUT[61]), .ZN(n7949) );
  NAND2_X2 U5689 ( .A1(MEM_WB_OUT[62]), .A2(n7361), .ZN(n7844) );
  NAND2_X2 U5690 ( .A1(MEM_WB_OUT[63]), .A2(n7360), .ZN(n7837) );
  NAND2_X2 U5691 ( .A1(n7855), .A2(MEM_WB_OUT[64]), .ZN(n7861) );
  NAND2_X2 U5692 ( .A1(MEM_WB_OUT[65]), .A2(n7360), .ZN(n7851) );
  NAND2_X2 U5693 ( .A1(MEM_WB_OUT[66]), .A2(n7358), .ZN(n8029) );
  NAND2_X2 U5694 ( .A1(n8038), .A2(MEM_WB_OUT[68]), .ZN(n8040) );
  INV_X8 U5695 ( .A(n10050), .ZN(n10037) );
  NAND2_X1 U5696 ( .A1(n6893), .A2(n8590), .ZN(n8583) );
  NAND3_X1 U5697 ( .A1(ID_EXEC_OUT[90]), .A2(n8493), .A3(n7469), .ZN(n8472) );
  NAND3_X1 U5698 ( .A1(ID_EXEC_OUT[85]), .A2(n8493), .A3(n7384), .ZN(n8495) );
  NAND2_X2 U5699 ( .A1(n8446), .A2(n9668), .ZN(n8650) );
  NOR2_X4 U5700 ( .A1(n8649), .A2(n8478), .ZN(n7344) );
  XNOR2_X2 U5701 ( .A(n9871), .B(n7449), .ZN(n8446) );
  NAND3_X2 U5702 ( .A1(DMEM_BUS_OUT[8]), .A2(n7463), .A3(n8070), .ZN(n7980) );
  NAND3_X2 U5703 ( .A1(ID_EXEC_OUT[91]), .A2(n7384), .A3(n5853), .ZN(n8468) );
  NAND3_X2 U5704 ( .A1(ID_EXEC_OUT[51]), .A2(n7311), .A3(n7337), .ZN(n7895) );
  INV_X4 U5705 ( .A(n8216), .ZN(n5844) );
  INV_X4 U5706 ( .A(n5844), .ZN(n5845) );
  INV_X4 U5707 ( .A(n5844), .ZN(n5846) );
  INV_X16 U5708 ( .A(n3184), .ZN(n1541) );
  INV_X4 U5709 ( .A(n3299), .ZN(n5847) );
  INV_X8 U5710 ( .A(n5847), .ZN(n5848) );
  XOR2_X1 U5711 ( .A(IMEM_BUS_IN[9]), .B(n3306), .Z(n3302) );
  XOR2_X1 U5712 ( .A(IMEM_BUS_IN[14]), .B(n3306), .Z(n3312) );
  NOR2_X1 U5713 ( .A1(n7773), .A2(n3306), .ZN(ID_EX_REG_ID_EX_REG_N65) );
  AOI221_X4 U5714 ( .B1(n5850), .B2(offset_26_id[9]), .C1(n1591), .C2(
        ID_STAGE_imm16_aluA[20]), .A(n3316), .ZN(n3305) );
  INV_X16 U5715 ( .A(n7465), .ZN(n7462) );
  NAND3_X2 U5716 ( .A1(DMEM_BUS_OUT[29]), .A2(n8070), .A3(n7337), .ZN(n8032)
         );
  NAND3_X1 U5717 ( .A1(n9900), .A2(n9842), .A3(n9901), .ZN(n9848) );
  INV_X16 U5718 ( .A(n5850), .ZN(n1591) );
  INV_X16 U5719 ( .A(n5849), .ZN(n5850) );
  OAI221_X2 U5720 ( .B1(n8854), .B2(n9239), .C1(n9239), .C2(n7314), .A(n7465), 
        .ZN(n7979) );
  INV_X4 U5721 ( .A(n3315), .ZN(n5849) );
  NAND3_X1 U5722 ( .A1(n3329), .A2(n6346), .A3(n3324), .ZN(n3315) );
  XOR2_X1 U5723 ( .A(IMEM_BUS_IN[10]), .B(n3305), .Z(n3304) );
  XOR2_X1 U5724 ( .A(IMEM_BUS_IN[15]), .B(n3305), .Z(n3313) );
  NOR2_X1 U5725 ( .A1(n7773), .A2(n3305), .ZN(ID_EX_REG_ID_EX_REG_N64) );
  NAND3_X1 U5726 ( .A1(ID_STAGE_imm16_aluA[29]), .A2(n6862), .A3(n3373), .ZN(
        n3370) );
  NAND2_X1 U5727 ( .A1(ID_STAGE_imm16_aluA[29]), .A2(n7305), .ZN(n3328) );
  NAND2_X1 U5728 ( .A1(ID_STAGE_imm16_aluA[29]), .A2(n1591), .ZN(n3358) );
  OR3_X1 U5729 ( .A1(ID_STAGE_imm16_aluA[29]), .A2(ID_STAGE_imm16_aluA[31]), 
        .A3(n3347), .ZN(n3372) );
  INV_X32 U5730 ( .A(n7460), .ZN(n7465) );
  OAI22_X2 U5731 ( .A1(n8693), .A2(n7389), .B1(n9060), .B2(n9164), .ZN(n9063)
         );
  NAND3_X2 U5732 ( .A1(n9858), .A2(n9856), .A3(n9857), .ZN(n9893) );
  OAI21_X2 U5733 ( .B1(n9147), .B2(n9855), .A(n9854), .ZN(n9856) );
  INV_X4 U5734 ( .A(n10162), .ZN(n10004) );
  NOR2_X2 U5735 ( .A1(n10010), .A2(n10041), .ZN(n10021) );
  NOR2_X2 U5736 ( .A1(n9185), .A2(n9184), .ZN(n9414) );
  NOR2_X2 U5737 ( .A1(n9183), .A2(n9182), .ZN(n9184) );
  OAI221_X2 U5738 ( .B1(n9818), .B2(n7392), .C1(n9817), .C2(n7393), .A(n9816), 
        .ZN(n9837) );
  NAND3_X1 U5739 ( .A1(n9862), .A2(n7366), .A3(n9815), .ZN(n9816) );
  AOI211_X2 U5740 ( .C1(n9814), .C2(n9813), .A(n9812), .B(n9811), .ZN(n9817)
         );
  INV_X16 U5741 ( .A(n7467), .ZN(n7466) );
  NOR2_X1 U5742 ( .A1(n9919), .A2(n9930), .ZN(n7898) );
  NAND3_X1 U5743 ( .A1(n8356), .A2(n8334), .A3(n6356), .ZN(n8325) );
  OAI21_X2 U5744 ( .B1(n8391), .B2(n8165), .A(n7036), .ZN(n8376) );
  OAI21_X2 U5745 ( .B1(n8701), .B2(n7383), .A(n8700), .ZN(n8725) );
  NAND3_X1 U5746 ( .A1(ID_STAGE_imm16_aluA[28]), .A2(n6011), .A3(n3373), .ZN(
        n3347) );
  NAND3_X2 U5747 ( .A1(n7954), .A2(n7953), .A3(n7952), .ZN(n8891) );
  AOI21_X2 U5748 ( .B1(MEM_WB_OUT[91]), .B2(n7951), .A(n7958), .ZN(n7954) );
  NAND3_X2 U5749 ( .A1(n7949), .A2(n7948), .A3(n7947), .ZN(n8902) );
  AOI21_X2 U5750 ( .B1(n7946), .B2(n8037), .A(n7945), .ZN(n7947) );
  INV_X16 U5751 ( .A(n7461), .ZN(n7460) );
  NAND3_X2 U5752 ( .A1(n7871), .A2(n7870), .A3(n7869), .ZN(n9079) );
  AOI21_X2 U5753 ( .B1(MEM_WB_OUT[87]), .B2(n7951), .A(n7958), .ZN(n7871) );
  OAI21_X2 U5754 ( .B1(n8075), .B2(n8053), .A(n8052), .ZN(n9230) );
  NOR2_X2 U5755 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[20]), .A2(n8072), 
        .ZN(n8053) );
  NOR2_X2 U5756 ( .A1(n9877), .A2(n9182), .ZN(n9019) );
  NAND2_X2 U5757 ( .A1(n9893), .A2(n9860), .ZN(n9892) );
  NOR2_X2 U5758 ( .A1(n9160), .A2(n9159), .ZN(n9438) );
  NOR2_X1 U5759 ( .A1(n9148), .A2(n7391), .ZN(n9149) );
  NOR2_X2 U5760 ( .A1(n8533), .A2(n8532), .ZN(n9531) );
  NAND3_X2 U5761 ( .A1(n8531), .A2(n9154), .A3(n8637), .ZN(n8532) );
  NAND3_X2 U5762 ( .A1(n9372), .A2(n9371), .A3(n9370), .ZN(n9698) );
  NAND2_X2 U5763 ( .A1(n7380), .A2(n7384), .ZN(n9293) );
  NAND3_X2 U5764 ( .A1(DMEM_BUS_OUT[31]), .A2(n7384), .A3(n7380), .ZN(n8435)
         );
  NAND3_X2 U5765 ( .A1(ID_EXEC_OUT[95]), .A2(n7384), .A3(n7381), .ZN(n8436) );
  NOR3_X2 U5766 ( .A1(n8409), .A2(MEM_WB_REG_MEM_WB_REG_N7), .A3(n6461), .ZN(
        n8413) );
  NAND2_X2 U5767 ( .A1(MEM_WB_REG_MEM_WB_REG_N8), .A2(n6889), .ZN(n8409) );
  NOR2_X2 U5768 ( .A1(n8083), .A2(n7000), .ZN(n8084) );
  NOR2_X1 U5769 ( .A1(n9894), .A2(n9853), .ZN(n7866) );
  OAI21_X2 U5770 ( .B1(n8293), .B2(n8295), .A(n6357), .ZN(n8215) );
  OAI21_X1 U5771 ( .B1(EXEC_STAGE_imm26_32[9]), .B2(n8151), .A(n5846), .ZN(
        n8211) );
  OAI21_X1 U5772 ( .B1(EXEC_STAGE_imm26_32[10]), .B2(n8133), .A(n5846), .ZN(
        n8210) );
  NOR2_X1 U5773 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[27]), .A2(n8072), 
        .ZN(n8066) );
  OAI21_X1 U5774 ( .B1(EXEC_STAGE_imm26_32[12]), .B2(n8135), .A(n5846), .ZN(
        n8150) );
  NOR3_X2 U5775 ( .A1(n8377), .A2(n8185), .A3(n8184), .ZN(n8200) );
  AOI21_X2 U5776 ( .B1(n8181), .B2(n8367), .A(n8180), .ZN(n8202) );
  AOI21_X2 U5777 ( .B1(n8376), .B2(n8380), .A(n8381), .ZN(n8368) );
  OAI21_X2 U5778 ( .B1(n8552), .B2(n8554), .A(n6918), .ZN(n8162) );
  AOI22_X2 U5779 ( .A1(MEM_WB_OUT[94]), .A2(n7841), .B1(n7834), .B2(
        WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[17]), .ZN(n7842) );
  NOR3_X2 U5780 ( .A1(n8697), .A2(n8696), .A3(n8695), .ZN(n8726) );
  NOR2_X2 U5781 ( .A1(n7388), .A2(n8693), .ZN(n8696) );
  NOR2_X2 U5782 ( .A1(n10246), .A2(n8694), .ZN(n8695) );
  OAI21_X2 U5783 ( .B1(n3368), .B2(n3353), .A(n3369), .ZN(n3345) );
  NAND3_X2 U5784 ( .A1(ID_STAGE_imm16_aluA[30]), .A2(n6012), .A3(n1590), .ZN(
        n3369) );
  AOI21_X2 U5785 ( .B1(MEM_WB_OUT[89]), .B2(n7951), .A(n7958), .ZN(n7883) );
  AOI21_X2 U5786 ( .B1(MEM_WB_OUT[90]), .B2(n7959), .A(n7958), .ZN(n7962) );
  NOR2_X1 U5787 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[30]), .A2(n8072), 
        .ZN(n7903) );
  NOR2_X1 U5788 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[22]), .A2(n8072), 
        .ZN(n7982) );
  NOR2_X1 U5789 ( .A1(n6881), .A2(IF_ID_OUT[32]), .ZN(n3323) );
  NOR3_X2 U5790 ( .A1(n9311), .A2(n9626), .A3(n9388), .ZN(n9312) );
  NAND3_X2 U5791 ( .A1(n9416), .A2(n9415), .A3(n7214), .ZN(n9433) );
  NAND3_X2 U5792 ( .A1(n7877), .A2(n7876), .A3(n7875), .ZN(n9086) );
  AOI21_X2 U5793 ( .B1(MEM_WB_OUT[86]), .B2(n7951), .A(n7958), .ZN(n7877) );
  NOR2_X1 U5794 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[31]), .A2(n8072), 
        .ZN(n7922) );
  NOR2_X1 U5795 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[21]), .A2(n8072), 
        .ZN(n7989) );
  NAND3_X2 U5796 ( .A1(ID_EXEC_OUT[156]), .A2(ID_EXEC_OUT[157]), .A3(
        ID_EXEC_OUT[158]), .ZN(n9742) );
  NOR2_X1 U5797 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[23]), .A2(n8072), 
        .ZN(n8074) );
  NOR3_X2 U5798 ( .A1(n8733), .A2(n8732), .A3(n8731), .ZN(n9755) );
  NOR2_X1 U5799 ( .A1(n9032), .A2(n7386), .ZN(n8732) );
  INV_X8 U5800 ( .A(n7382), .ZN(n7383) );
  NOR2_X1 U5801 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[26]), .A2(n8072), 
        .ZN(n7968) );
  NOR3_X2 U5802 ( .A1(n9298), .A2(n9297), .A3(n9495), .ZN(n9302) );
  NAND2_X2 U5803 ( .A1(n9862), .A2(n6013), .ZN(n10255) );
  NOR2_X1 U5804 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[28]), .A2(n8072), 
        .ZN(n8060) );
  NAND2_X2 U5805 ( .A1(n6799), .A2(n9173), .ZN(n10281) );
  NAND2_X2 U5806 ( .A1(n9753), .A2(n9173), .ZN(n10274) );
  OAI21_X2 U5807 ( .B1(IF_ID_OUT[36]), .B2(n3351), .A(n3352), .ZN(n3343) );
  NAND3_X2 U5808 ( .A1(ID_STAGE_imm16_aluA[31]), .A2(n6011), .A3(n1590), .ZN(
        n3352) );
  OAI21_X2 U5809 ( .B1(n8122), .B2(n8121), .A(n8123), .ZN(n8229) );
  NAND2_X1 U5810 ( .A1(n7465), .A2(n8850), .ZN(n8000) );
  OAI21_X2 U5811 ( .B1(n8309), .B2(n8308), .A(n8307), .ZN(n8314) );
  NAND3_X2 U5812 ( .A1(DMEM_BUS_OUT[19]), .A2(n8070), .A3(n7462), .ZN(n7894)
         );
  NAND3_X1 U5813 ( .A1(DMEM_BUS_OUT[22]), .A2(n8070), .A3(n7462), .ZN(n7957)
         );
  OAI21_X2 U5814 ( .B1(n8577), .B2(n6999), .A(n8568), .ZN(n8574) );
  OAI21_X2 U5815 ( .B1(n7940), .B2(n7939), .A(n7460), .ZN(n7950) );
  OAI21_X2 U5816 ( .B1(n3364), .B2(n3354), .A(n3372), .ZN(n3334) );
  NAND3_X1 U5817 ( .A1(DMEM_BUS_OUT[18]), .A2(n8070), .A3(n7462), .ZN(n7872)
         );
  NAND3_X2 U5818 ( .A1(n8056), .A2(n8055), .A3(n8054), .ZN(n9964) );
  NAND3_X1 U5819 ( .A1(n7356), .A2(n7337), .A3(ID_EXEC_OUT[40]), .ZN(n7978) );
  AOI21_X2 U5820 ( .B1(n9940), .B2(n9939), .A(n6450), .ZN(n9942) );
  NOR2_X2 U5821 ( .A1(n9920), .A2(n6450), .ZN(n9921) );
  NOR2_X2 U5822 ( .A1(n9866), .A2(n9865), .ZN(n9867) );
  NAND3_X2 U5823 ( .A1(n10048), .A2(n10017), .A3(n10062), .ZN(n10018) );
  NOR2_X2 U5824 ( .A1(n10034), .A2(n10033), .ZN(n10035) );
  NOR3_X2 U5825 ( .A1(n8104), .A2(n4087), .A3(n8103), .ZN(n10299) );
  NAND3_X1 U5826 ( .A1(n4084), .A2(RegWrite_wb_out), .A3(n4083), .ZN(n8103) );
  NOR2_X2 U5827 ( .A1(MEM_WB_OUT[106]), .A2(n7451), .ZN(n8014) );
  NOR2_X2 U5828 ( .A1(n7771), .A2(n7223), .ZN(n7833) );
  OAI21_X2 U5829 ( .B1(n10008), .B2(n10007), .A(n10006), .ZN(n10027) );
  AOI21_X1 U5830 ( .B1(n10005), .B2(n10170), .A(n10004), .ZN(n10006) );
  NOR2_X2 U5831 ( .A1(n9779), .A2(n9778), .ZN(n9795) );
  INV_X4 U5832 ( .A(n7223), .ZN(n7452) );
  NOR2_X2 U5833 ( .A1(n9531), .A2(n10246), .ZN(n8618) );
  NOR2_X2 U5834 ( .A1(n8983), .A2(n7386), .ZN(n8619) );
  NAND3_X2 U5835 ( .A1(n7868), .A2(n7452), .A3(n7867), .ZN(n7915) );
  NOR2_X1 U5836 ( .A1(n7451), .A2(n6913), .ZN(n7868) );
  NOR3_X2 U5837 ( .A1(n6352), .A2(MEM_WB_OUT[106]), .A3(n7771), .ZN(n7867) );
  NAND2_X1 U5838 ( .A1(n9588), .A2(n9909), .ZN(n9633) );
  INV_X4 U5839 ( .A(n9804), .ZN(n9189) );
  NAND3_X2 U5840 ( .A1(n9375), .A2(n9374), .A3(n9373), .ZN(n10177) );
  NAND3_X2 U5841 ( .A1(ID_EXEC_OUT[156]), .A2(n6013), .A3(n7450), .ZN(n5665)
         );
  NOR2_X1 U5842 ( .A1(n10163), .A2(n7351), .ZN(n7987) );
  NOR2_X1 U5843 ( .A1(n9318), .A2(n7366), .ZN(n8047) );
  OAI21_X1 U5844 ( .B1(EXEC_STAGE_imm26_32[6]), .B2(n8120), .A(n5846), .ZN(
        n8225) );
  NAND3_X2 U5845 ( .A1(n3247), .A2(IMEM_BUS_OUT[8]), .A3(IMEM_BUS_OUT[7]), 
        .ZN(n3243) );
  OAI21_X1 U5846 ( .B1(EXEC_STAGE_imm26_32[7]), .B2(n8120), .A(n5846), .ZN(
        n8218) );
  OAI21_X1 U5847 ( .B1(EXEC_STAGE_imm26_32[8]), .B2(n8151), .A(n5846), .ZN(
        n8214) );
  NAND4_X2 U5848 ( .A1(n8207), .A2(n8206), .A3(n8205), .A4(n8204), .ZN(n8292)
         );
  NOR2_X2 U5849 ( .A1(n8308), .A2(n8153), .ZN(n8207) );
  NOR2_X2 U5850 ( .A1(n8346), .A2(n8323), .ZN(n8206) );
  NOR3_X2 U5851 ( .A1(n3251), .A2(n6907), .A3(n1996), .ZN(n3247) );
  NAND3_X2 U5852 ( .A1(IMEM_BUS_OUT[11]), .A2(n3255), .A3(IMEM_BUS_OUT[12]), 
        .ZN(n3251) );
  NOR3_X2 U5853 ( .A1(n6040), .A2(n3259), .A3(n5909), .ZN(n3255) );
  OAI21_X1 U5854 ( .B1(EXEC_STAGE_imm26_32[14]), .B2(n8138), .A(n5846), .ZN(
        n8144) );
  NAND3_X2 U5855 ( .A1(IMEM_BUS_OUT[15]), .A2(n3263), .A3(IMEM_BUS_OUT[16]), 
        .ZN(n3259) );
  NOR3_X2 U5856 ( .A1(n6041), .A2(n3267), .A3(n6877), .ZN(n3263) );
  NAND3_X2 U5857 ( .A1(IMEM_BUS_OUT[19]), .A2(n3271), .A3(IMEM_BUS_OUT[20]), 
        .ZN(n3267) );
  AOI21_X2 U5858 ( .B1(n4545), .B2(n4546), .A(n7554), .ZN(n4544) );
  AOI21_X2 U5859 ( .B1(n4549), .B2(n4550), .A(n7520), .ZN(n4543) );
  AOI21_X2 U5860 ( .B1(n4553), .B2(n4554), .A(n7518), .ZN(n4542) );
  NOR3_X2 U5861 ( .A1(n6914), .A2(n3275), .A3(n2008), .ZN(n3271) );
  NAND3_X2 U5862 ( .A1(IMEM_BUS_OUT[23]), .A2(n3279), .A3(IMEM_BUS_OUT[24]), 
        .ZN(n3275) );
  NOR3_X2 U5863 ( .A1(n6915), .A2(n3283), .A3(n2012), .ZN(n3279) );
  AOI21_X2 U5864 ( .B1(n4680), .B2(n4681), .A(n7553), .ZN(n4679) );
  AOI21_X2 U5865 ( .B1(n4684), .B2(n4685), .A(n7519), .ZN(n4678) );
  AOI21_X2 U5866 ( .B1(n4688), .B2(n4689), .A(n7517), .ZN(n4677) );
  NAND3_X2 U5867 ( .A1(IMEM_BUS_OUT[28]), .A2(IMEM_BUS_OUT[27]), .A3(
        IMEM_BUS_OUT[29]), .ZN(n3283) );
  NAND3_X2 U5868 ( .A1(n8564), .A2(n8560), .A3(n8197), .ZN(n8590) );
  AOI21_X2 U5869 ( .B1(n4703), .B2(n4704), .A(n7553), .ZN(n4702) );
  AOI21_X2 U5870 ( .B1(n4707), .B2(n4708), .A(n7519), .ZN(n4701) );
  AOI21_X2 U5871 ( .B1(n4711), .B2(n4712), .A(n7517), .ZN(n4700) );
  INV_X8 U5872 ( .A(n9894), .ZN(n9179) );
  NAND2_X2 U5873 ( .A1(n7618), .A2(n7796), .ZN(n3168) );
  INV_X8 U5874 ( .A(n7618), .ZN(n7616) );
  AOI21_X2 U5875 ( .B1(n4478), .B2(n4479), .A(n7554), .ZN(n4477) );
  AOI21_X2 U5876 ( .B1(n4482), .B2(n4483), .A(n7520), .ZN(n4476) );
  AOI21_X2 U5877 ( .B1(n4486), .B2(n4487), .A(n7518), .ZN(n4475) );
  AOI21_X2 U5878 ( .B1(n4504), .B2(n4505), .A(n7520), .ZN(n4498) );
  AOI21_X2 U5879 ( .B1(n4508), .B2(n4509), .A(n7518), .ZN(n4497) );
  AOI21_X2 U5880 ( .B1(n4500), .B2(n4501), .A(n7554), .ZN(n4499) );
  AOI21_X2 U5881 ( .B1(n4523), .B2(n4524), .A(n7554), .ZN(n4522) );
  AOI21_X2 U5882 ( .B1(n4527), .B2(n4528), .A(n7520), .ZN(n4521) );
  AOI21_X2 U5883 ( .B1(n4531), .B2(n4532), .A(n7518), .ZN(n4520) );
  AOI21_X2 U5884 ( .B1(n4567), .B2(n4568), .A(n7553), .ZN(n4566) );
  AOI21_X2 U5885 ( .B1(n4571), .B2(n4572), .A(n7519), .ZN(n4565) );
  AOI21_X2 U5886 ( .B1(n4575), .B2(n4576), .A(n7517), .ZN(n4564) );
  AOI21_X2 U5887 ( .B1(n4589), .B2(n4590), .A(n7553), .ZN(n4588) );
  AOI21_X2 U5888 ( .B1(n4593), .B2(n4594), .A(n7519), .ZN(n4587) );
  AOI21_X2 U5889 ( .B1(n4597), .B2(n4598), .A(n7517), .ZN(n4586) );
  AOI21_X2 U5890 ( .B1(n4612), .B2(n4613), .A(n7553), .ZN(n4611) );
  AOI21_X2 U5891 ( .B1(n4616), .B2(n4617), .A(n7519), .ZN(n4610) );
  AOI21_X2 U5892 ( .B1(n4620), .B2(n4621), .A(n7517), .ZN(n4609) );
  AOI21_X2 U5893 ( .B1(n4635), .B2(n4636), .A(n7553), .ZN(n4634) );
  AOI21_X2 U5894 ( .B1(n4639), .B2(n4640), .A(n7519), .ZN(n4633) );
  AOI21_X2 U5895 ( .B1(n4643), .B2(n4644), .A(n7517), .ZN(n4632) );
  AOI21_X2 U5896 ( .B1(n4408), .B2(n4409), .A(n7554), .ZN(n4407) );
  AOI21_X2 U5897 ( .B1(n4412), .B2(n4413), .A(n7520), .ZN(n4406) );
  AOI21_X2 U5898 ( .B1(n4416), .B2(n4417), .A(n7518), .ZN(n4405) );
  AOI21_X2 U5899 ( .B1(n4431), .B2(n4432), .A(n7554), .ZN(n4430) );
  AOI21_X2 U5900 ( .B1(n4435), .B2(n4436), .A(n7520), .ZN(n4429) );
  AOI21_X2 U5901 ( .B1(n4439), .B2(n4440), .A(n7518), .ZN(n4428) );
  AOI21_X2 U5902 ( .B1(n4460), .B2(n4461), .A(n7520), .ZN(n4454) );
  AOI21_X2 U5903 ( .B1(n4464), .B2(n4465), .A(n7518), .ZN(n4453) );
  AOI21_X2 U5904 ( .B1(n4456), .B2(n4457), .A(n7554), .ZN(n4455) );
  AOI21_X2 U5905 ( .B1(n4657), .B2(n4658), .A(n7553), .ZN(n4656) );
  AOI21_X2 U5906 ( .B1(n4661), .B2(n4662), .A(n7519), .ZN(n4655) );
  AOI21_X2 U5907 ( .B1(n4665), .B2(n4666), .A(n7517), .ZN(n4654) );
  AOI21_X2 U5908 ( .B1(n4748), .B2(n4749), .A(n7553), .ZN(n4747) );
  AOI21_X2 U5909 ( .B1(n4752), .B2(n4753), .A(n7519), .ZN(n4746) );
  AOI21_X2 U5910 ( .B1(n4756), .B2(n4757), .A(n7517), .ZN(n4745) );
  AOI21_X2 U5911 ( .B1(n4770), .B2(n4771), .A(n7553), .ZN(n4769) );
  AOI21_X2 U5912 ( .B1(n4774), .B2(n4775), .A(n7519), .ZN(n4768) );
  AOI21_X2 U5913 ( .B1(n4778), .B2(n4779), .A(n7517), .ZN(n4767) );
  AOI21_X2 U5914 ( .B1(n4792), .B2(n4793), .A(n7553), .ZN(n4791) );
  AOI21_X2 U5915 ( .B1(n4796), .B2(n4797), .A(n7519), .ZN(n4790) );
  AOI21_X2 U5916 ( .B1(n4800), .B2(n4801), .A(n7517), .ZN(n4789) );
  AOI21_X2 U5917 ( .B1(n4273), .B2(n4274), .A(n7553), .ZN(n4272) );
  AOI21_X2 U5918 ( .B1(n4277), .B2(n4278), .A(n7519), .ZN(n4271) );
  AOI21_X2 U5919 ( .B1(n4281), .B2(n4282), .A(n7517), .ZN(n4270) );
  AOI21_X2 U5920 ( .B1(n4119), .B2(n4120), .A(n7518), .ZN(n4102) );
  AOI21_X2 U5921 ( .B1(n4105), .B2(n4106), .A(n7554), .ZN(n4104) );
  AOI21_X2 U5922 ( .B1(n4114), .B2(n4115), .A(n7520), .ZN(n4103) );
  AOI21_X2 U5923 ( .B1(n4146), .B2(n4147), .A(n7517), .ZN(n4135) );
  AOI21_X2 U5924 ( .B1(n4138), .B2(n4139), .A(n7553), .ZN(n4137) );
  AOI21_X2 U5925 ( .B1(n4142), .B2(n4143), .A(n7519), .ZN(n4136) );
  AOI21_X2 U5926 ( .B1(n4318), .B2(n4319), .A(n7554), .ZN(n4317) );
  AOI21_X2 U5927 ( .B1(n4322), .B2(n4323), .A(n7520), .ZN(n4316) );
  AOI21_X2 U5928 ( .B1(n4326), .B2(n4327), .A(n7518), .ZN(n4315) );
  AOI21_X2 U5929 ( .B1(n4183), .B2(n4184), .A(n7553), .ZN(n4182) );
  AOI21_X2 U5930 ( .B1(n4187), .B2(n4188), .A(n7519), .ZN(n4181) );
  AOI21_X2 U5931 ( .B1(n4191), .B2(n4192), .A(n7517), .ZN(n4180) );
  AOI21_X2 U5932 ( .B1(n4363), .B2(n4364), .A(n7554), .ZN(n4362) );
  AOI21_X2 U5933 ( .B1(n4367), .B2(n4368), .A(n7520), .ZN(n4361) );
  AOI21_X2 U5934 ( .B1(n4371), .B2(n4372), .A(n7518), .ZN(n4360) );
  AOI21_X2 U5935 ( .B1(n4228), .B2(n4229), .A(n7553), .ZN(n4227) );
  AOI21_X2 U5936 ( .B1(n4232), .B2(n4233), .A(n7519), .ZN(n4226) );
  AOI21_X2 U5937 ( .B1(n4236), .B2(n4237), .A(n7517), .ZN(n4225) );
  AOI21_X2 U5938 ( .B1(n4251), .B2(n4252), .A(n7554), .ZN(n4250) );
  AOI21_X2 U5939 ( .B1(n4255), .B2(n4256), .A(n7520), .ZN(n4249) );
  AOI21_X2 U5940 ( .B1(n4259), .B2(n4260), .A(n7518), .ZN(n4248) );
  AOI21_X2 U5941 ( .B1(n4296), .B2(n4297), .A(n7554), .ZN(n4295) );
  AOI21_X2 U5942 ( .B1(n4300), .B2(n4301), .A(n7520), .ZN(n4294) );
  AOI21_X2 U5943 ( .B1(n4304), .B2(n4305), .A(n7518), .ZN(n4293) );
  AOI21_X2 U5944 ( .B1(n4161), .B2(n4162), .A(n7554), .ZN(n4160) );
  AOI21_X2 U5945 ( .B1(n4165), .B2(n4166), .A(n7520), .ZN(n4159) );
  AOI21_X2 U5946 ( .B1(n4169), .B2(n4170), .A(n7518), .ZN(n4158) );
  AOI21_X2 U5947 ( .B1(n4341), .B2(n4342), .A(n7554), .ZN(n4340) );
  AOI21_X2 U5948 ( .B1(n4345), .B2(n4346), .A(n7520), .ZN(n4339) );
  AOI21_X2 U5949 ( .B1(n4349), .B2(n4350), .A(n7518), .ZN(n4338) );
  AOI21_X2 U5950 ( .B1(n4206), .B2(n4207), .A(n7554), .ZN(n4205) );
  AOI21_X2 U5951 ( .B1(n4210), .B2(n4211), .A(n7520), .ZN(n4204) );
  AOI21_X2 U5952 ( .B1(n4214), .B2(n4215), .A(n7518), .ZN(n4203) );
  AOI21_X2 U5953 ( .B1(n4386), .B2(n4387), .A(n7554), .ZN(n4385) );
  AOI21_X2 U5954 ( .B1(n4390), .B2(n4391), .A(n7520), .ZN(n4384) );
  AOI21_X2 U5955 ( .B1(n4394), .B2(n4395), .A(n7518), .ZN(n4383) );
  NOR3_X2 U5956 ( .A1(n8986), .A2(n8985), .A3(n8984), .ZN(n8998) );
  NOR2_X2 U5957 ( .A1(n8982), .A2(n7385), .ZN(n8985) );
  NOR2_X1 U5958 ( .A1(n8983), .A2(n7388), .ZN(n8984) );
  NOR2_X2 U5959 ( .A1(n8526), .A2(n8525), .ZN(n8527) );
  NOR2_X1 U5960 ( .A1(n9539), .A2(n9806), .ZN(n8526) );
  OAI21_X2 U5961 ( .B1(n9468), .B2(n10274), .A(n9467), .ZN(n9476) );
  OAI21_X2 U5962 ( .B1(n9967), .B2(n10230), .A(n10229), .ZN(n9478) );
  NOR2_X2 U5963 ( .A1(n9534), .A2(n9533), .ZN(n9535) );
  NOR2_X2 U5964 ( .A1(n9531), .A2(n7386), .ZN(n9534) );
  NOR2_X2 U5965 ( .A1(n9541), .A2(n9540), .ZN(n9542) );
  NOR2_X2 U5966 ( .A1(n9539), .A2(n7386), .ZN(n9540) );
  NOR2_X2 U5967 ( .A1(n8538), .A2(n8537), .ZN(n8539) );
  NOR2_X2 U5968 ( .A1(n9532), .A2(n7385), .ZN(n8537) );
  NAND2_X2 U5969 ( .A1(n9308), .A2(n9307), .ZN(n9389) );
  AOI21_X2 U5970 ( .B1(n9653), .B2(n9304), .A(n9663), .ZN(n9308) );
  NOR3_X2 U5971 ( .A1(n9305), .A2(n9660), .A3(n9654), .ZN(n9306) );
  NOR3_X2 U5972 ( .A1(n9357), .A2(n9356), .A3(n9355), .ZN(n9645) );
  NOR2_X1 U5973 ( .A1(n9721), .A2(n9806), .ZN(n9356) );
  NOR2_X2 U5974 ( .A1(n9722), .A2(n7385), .ZN(n9355) );
  NOR3_X2 U5975 ( .A1(n9644), .A2(n9643), .A3(n9642), .ZN(n9681) );
  OAI21_X2 U5976 ( .B1(n9640), .B2(n7386), .A(n9639), .ZN(n9644) );
  NOR2_X1 U5977 ( .A1(n9707), .A2(n9806), .ZN(n9643) );
  NOR3_X2 U5978 ( .A1(n9680), .A2(n9679), .A3(n9678), .ZN(n9745) );
  NOR2_X1 U5979 ( .A1(n9719), .A2(n7388), .ZN(n9679) );
  NOR2_X2 U5980 ( .A1(n9721), .A2(n7386), .ZN(n9678) );
  NOR3_X2 U5981 ( .A1(n9710), .A2(n9709), .A3(n9708), .ZN(n9746) );
  NOR2_X1 U5982 ( .A1(n7388), .A2(n9706), .ZN(n9709) );
  NOR2_X2 U5983 ( .A1(n9707), .A2(n7385), .ZN(n9708) );
  NOR3_X2 U5984 ( .A1(n9725), .A2(n9724), .A3(n9723), .ZN(n10143) );
  NOR2_X2 U5985 ( .A1(n9722), .A2(n10246), .ZN(n9723) );
  NAND2_X2 U5986 ( .A1(n6800), .A2(n9173), .ZN(n10279) );
  AOI21_X2 U5987 ( .B1(n4821), .B2(n4822), .A(n7553), .ZN(n4820) );
  AOI21_X2 U5988 ( .B1(n4826), .B2(n4827), .A(n7519), .ZN(n4819) );
  AOI21_X2 U5989 ( .B1(n4830), .B2(n4831), .A(n7517), .ZN(n4818) );
  OAI211_X2 U5990 ( .C1(n3290), .C2(n3291), .A(n3292), .B(n3293), .ZN(n3232)
         );
  NOR4_X2 U5991 ( .A1(n3295), .A2(n3296), .A3(n3297), .A4(n3298), .ZN(n3291)
         );
  NAND3_X2 U5992 ( .A1(ID_STAGE_imm16_aluA[30]), .A2(n6867), .A3(n3373), .ZN(
        n3355) );
  OAI21_X2 U5993 ( .B1(n3347), .B2(ID_STAGE_imm16_aluA[31]), .A(n3371), .ZN(
        n3367) );
  NOR2_X2 U5994 ( .A1(n8129), .A2(n8229), .ZN(n8130) );
  NOR2_X2 U5995 ( .A1(n8245), .A2(n8228), .ZN(n8125) );
  NAND4_X2 U5996 ( .A1(n8232), .A2(n8231), .A3(n8230), .A4(n8269), .ZN(n8233)
         );
  NOR2_X2 U5997 ( .A1(n8228), .A2(n8245), .ZN(n8232) );
  NAND2_X2 U5998 ( .A1(n7464), .A2(n9234), .ZN(n7990) );
  OAI21_X2 U5999 ( .B1(n5915), .B2(n8212), .A(n6189), .ZN(n8213) );
  OAI21_X2 U6000 ( .B1(n8325), .B2(n8306), .A(n8305), .ZN(n8319) );
  NOR2_X2 U6001 ( .A1(n8323), .A2(n8329), .ZN(n8303) );
  OAI21_X2 U6002 ( .B1(n8370), .B2(n8369), .A(n8368), .ZN(n8386) );
  NAND3_X2 U6003 ( .A1(n8550), .A2(n8390), .A3(n6892), .ZN(n8369) );
  NAND3_X2 U6004 ( .A1(n8379), .A2(n8551), .A3(n8378), .ZN(n8384) );
  AOI21_X2 U6005 ( .B1(n3811), .B2(n7612), .A(n8400), .ZN(n8401) );
  NAND3_X2 U6006 ( .A1(n3812), .A2(n3813), .A3(n3814), .ZN(n3811) );
  OAI21_X2 U6007 ( .B1(n6185), .B2(n10274), .A(n8517), .ZN(n8546) );
  OAI21_X2 U6008 ( .B1(n8393), .B2(n8392), .A(n8391), .ZN(n8555) );
  OAI21_X2 U6009 ( .B1(n8185), .B2(n6036), .A(n6520), .ZN(n8160) );
  NOR2_X2 U6010 ( .A1(n8562), .A2(n8561), .ZN(n8563) );
  AOI21_X2 U6011 ( .B1(n3938), .B2(n7612), .A(n8598), .ZN(n8599) );
  NAND3_X2 U6012 ( .A1(n3939), .A2(n3940), .A3(n3941), .ZN(n3938) );
  NAND3_X1 U6013 ( .A1(DMEM_BUS_OUT[25]), .A2(n8070), .A3(n7462), .ZN(n7845)
         );
  AOI21_X2 U6014 ( .B1(n3959), .B2(n7612), .A(n8670), .ZN(n8671) );
  NAND3_X2 U6015 ( .A1(n3960), .A2(n3961), .A3(n3962), .ZN(n3959) );
  NOR2_X2 U6016 ( .A1(n8705), .A2(n10155), .ZN(n8706) );
  OAI21_X2 U6017 ( .B1(n8687), .B2(n7392), .A(n8686), .ZN(n8704) );
  OAI21_X2 U6018 ( .B1(n8726), .B2(n7393), .A(n8702), .ZN(n8703) );
  NOR2_X2 U6019 ( .A1(n9179), .A2(n8683), .ZN(n8707) );
  AOI21_X1 U6020 ( .B1(n10264), .B2(n8682), .A(n6844), .ZN(n8683) );
  AOI21_X2 U6021 ( .B1(n3980), .B2(n7612), .A(n8718), .ZN(n8719) );
  NAND3_X2 U6022 ( .A1(n3981), .A2(n3982), .A3(n3983), .ZN(n3980) );
  NOR3_X2 U6023 ( .A1(n4723), .A2(n4724), .A3(n4725), .ZN(n4722) );
  OAI21_X2 U6024 ( .B1(n8751), .B2(n6998), .A(n8711), .ZN(n8748) );
  AOI21_X2 U6025 ( .B1(n3916), .B2(n7612), .A(n8771), .ZN(n8772) );
  NAND3_X2 U6026 ( .A1(n3917), .A2(n3918), .A3(n3919), .ZN(n3916) );
  AOI21_X2 U6027 ( .B1(n3853), .B2(n7612), .A(n8779), .ZN(n8780) );
  NAND3_X2 U6028 ( .A1(n3854), .A2(n3855), .A3(n3856), .ZN(n3853) );
  AOI21_X2 U6029 ( .B1(n3832), .B2(n7612), .A(n8787), .ZN(n8788) );
  NAND3_X2 U6030 ( .A1(n3833), .A2(n3834), .A3(n3835), .ZN(n3832) );
  AOI21_X2 U6031 ( .B1(n3769), .B2(n7612), .A(n8795), .ZN(n8796) );
  NAND3_X2 U6032 ( .A1(n3770), .A2(n3771), .A3(n3772), .ZN(n3769) );
  AOI21_X2 U6033 ( .B1(n3748), .B2(n7612), .A(n8803), .ZN(n8804) );
  NAND3_X2 U6034 ( .A1(n3749), .A2(n3750), .A3(n3751), .ZN(n3748) );
  AOI21_X2 U6035 ( .B1(n4064), .B2(n7612), .A(n8807), .ZN(n8808) );
  NAND3_X2 U6036 ( .A1(n4065), .A2(n4066), .A3(n4067), .ZN(n4064) );
  AOI21_X2 U6037 ( .B1(n4043), .B2(n7612), .A(n8815), .ZN(n8816) );
  NAND3_X2 U6038 ( .A1(n4044), .A2(n4045), .A3(n4046), .ZN(n4043) );
  AOI21_X2 U6039 ( .B1(n4001), .B2(n7612), .A(n8823), .ZN(n8824) );
  NAND3_X2 U6040 ( .A1(n4002), .A2(n4003), .A3(n4004), .ZN(n4001) );
  AOI21_X2 U6041 ( .B1(n4022), .B2(n7612), .A(n8827), .ZN(n8828) );
  NAND3_X2 U6042 ( .A1(n4023), .A2(n4024), .A3(n4025), .ZN(n4022) );
  AOI21_X2 U6043 ( .B1(n3895), .B2(n7612), .A(n8831), .ZN(n8832) );
  NAND3_X2 U6044 ( .A1(n3896), .A2(n3897), .A3(n3898), .ZN(n3895) );
  AOI21_X2 U6045 ( .B1(n3874), .B2(n7612), .A(n8835), .ZN(n8836) );
  NAND3_X2 U6046 ( .A1(n3875), .A2(n3876), .A3(n3877), .ZN(n3874) );
  AOI21_X2 U6047 ( .B1(n3790), .B2(n7612), .A(n8839), .ZN(n8840) );
  NAND3_X2 U6048 ( .A1(n3791), .A2(n3792), .A3(n3793), .ZN(n3790) );
  AOI21_X2 U6049 ( .B1(n3725), .B2(n7612), .A(n7237), .ZN(n8841) );
  NAND3_X2 U6050 ( .A1(n3726), .A2(n3727), .A3(n3728), .ZN(n3725) );
  AOI21_X2 U6051 ( .B1(n3703), .B2(n7612), .A(n7238), .ZN(n8842) );
  NAND3_X2 U6052 ( .A1(n3704), .A2(n3705), .A3(n3706), .ZN(n3703) );
  AOI21_X2 U6053 ( .B1(n3681), .B2(n7612), .A(n7284), .ZN(n8846) );
  NAND3_X2 U6054 ( .A1(n3682), .A2(n3683), .A3(n3684), .ZN(n3681) );
  AOI21_X2 U6055 ( .B1(n3660), .B2(n7612), .A(n7285), .ZN(n8847) );
  NAND3_X2 U6056 ( .A1(n3661), .A2(n3662), .A3(n3663), .ZN(n3660) );
  AOI21_X2 U6057 ( .B1(n3638), .B2(n7612), .A(n7269), .ZN(n8848) );
  NAND3_X2 U6058 ( .A1(n3639), .A2(n3640), .A3(n3641), .ZN(n3638) );
  AOI21_X2 U6059 ( .B1(n3617), .B2(n7612), .A(n7235), .ZN(n8849) );
  NAND3_X2 U6060 ( .A1(n3618), .A2(n3619), .A3(n3620), .ZN(n3617) );
  AOI21_X2 U6061 ( .B1(n3595), .B2(n7612), .A(n7287), .ZN(n8853) );
  NAND3_X2 U6062 ( .A1(n3596), .A2(n3597), .A3(n3598), .ZN(n3595) );
  AOI21_X2 U6063 ( .B1(n3574), .B2(n3390), .A(n7286), .ZN(n8856) );
  NAND3_X2 U6064 ( .A1(n3575), .A2(n3576), .A3(n3577), .ZN(n3574) );
  NAND3_X2 U6065 ( .A1(n3553), .A2(n3554), .A3(n3555), .ZN(n3552) );
  NAND3_X2 U6066 ( .A1(n3532), .A2(n3533), .A3(n3534), .ZN(n3531) );
  NAND3_X2 U6067 ( .A1(n3510), .A2(n3511), .A3(n3512), .ZN(n3509) );
  NAND3_X2 U6068 ( .A1(n3489), .A2(n3490), .A3(n3491), .ZN(n3488) );
  NAND3_X2 U6069 ( .A1(n3467), .A2(n3468), .A3(n3469), .ZN(n3466) );
  NAND3_X2 U6070 ( .A1(n3446), .A2(n3447), .A3(n3448), .ZN(n3445) );
  NAND3_X2 U6071 ( .A1(n3424), .A2(n3425), .A3(n3426), .ZN(n3423) );
  NAND3_X2 U6072 ( .A1(n3392), .A2(n3393), .A3(n3394), .ZN(n3391) );
  NAND3_X2 U6073 ( .A1(n6343), .A2(n6881), .A3(IF_ID_OUT[32]), .ZN(n3326) );
  NOR2_X2 U6074 ( .A1(IF_ID_OUT[32]), .A2(IF_ID_OUT[35]), .ZN(n3329) );
  NOR2_X2 U6075 ( .A1(n4090), .A2(n4113), .ZN(n3378) );
  NAND3_X2 U6076 ( .A1(n3329), .A2(n6347), .A3(IF_ID_OUT[36]), .ZN(n3322) );
  NOR3_X2 U6077 ( .A1(n3326), .A2(n1654), .A3(n6347), .ZN(n3319) );
  NOR2_X2 U6078 ( .A1(n3322), .A2(n6346), .ZN(n3316) );
  OAI21_X2 U6079 ( .B1(n8963), .B2(n10230), .A(n10229), .ZN(n8965) );
  AOI21_X2 U6080 ( .B1(n9010), .B2(n10229), .A(n9009), .ZN(n9011) );
  OAI21_X2 U6081 ( .B1(n9026), .B2(n7392), .A(n9025), .ZN(n9043) );
  AOI21_X2 U6082 ( .B1(n9049), .B2(n10229), .A(n9872), .ZN(n9050) );
  OAI21_X2 U6083 ( .B1(n9134), .B2(n7393), .A(n9133), .ZN(n9135) );
  OAI21_X2 U6084 ( .B1(n6482), .B2(n7392), .A(n9118), .ZN(n9136) );
  AOI21_X2 U6085 ( .B1(n9141), .B2(n10229), .A(n9140), .ZN(n9142) );
  AOI21_X2 U6086 ( .B1(n9322), .B2(n9321), .A(n7479), .ZN(n9323) );
  NAND3_X2 U6087 ( .A1(n9207), .A2(n9206), .A3(n9205), .ZN(n9209) );
  AOI21_X2 U6088 ( .B1(n9517), .B2(n9204), .A(n9203), .ZN(n9205) );
  AOI21_X2 U6089 ( .B1(n10277), .B2(n9410), .A(n9172), .ZN(n9207) );
  OAI21_X2 U6090 ( .B1(n9338), .B2(n10230), .A(n10229), .ZN(n9339) );
  AOI21_X1 U6091 ( .B1(n9618), .B2(n9433), .A(n9420), .ZN(n9421) );
  OAI21_X2 U6092 ( .B1(n9971), .B2(n10230), .A(n10229), .ZN(n9425) );
  NAND3_X2 U6093 ( .A1(n9489), .A2(n9488), .A3(n7236), .ZN(n9490) );
  OAI21_X2 U6094 ( .B1(n9646), .B2(n9515), .A(n9514), .ZN(n9520) );
  OAI21_X1 U6095 ( .B1(n9506), .B2(n9505), .A(n9504), .ZN(n9507) );
  NAND3_X1 U6096 ( .A1(DMEM_BUS_OUT[17]), .A2(n8070), .A3(n7462), .ZN(n7880)
         );
  OAI21_X2 U6097 ( .B1(n9509), .B2(n10230), .A(n10229), .ZN(n9510) );
  AOI21_X2 U6098 ( .B1(n9556), .B2(n10229), .A(n9555), .ZN(n9557) );
  AOI21_X2 U6099 ( .B1(n9574), .B2(n10229), .A(n9573), .ZN(n9575) );
  AOI21_X2 U6100 ( .B1(n9583), .B2(n9582), .A(n9581), .ZN(n9585) );
  OAI21_X1 U6101 ( .B1(n9586), .B2(n10230), .A(n10229), .ZN(n9587) );
  AOI21_X2 U6102 ( .B1(n9621), .B2(n10229), .A(n9620), .ZN(n9622) );
  OAI21_X2 U6103 ( .B1(n9630), .B2(n10274), .A(n9629), .ZN(n9648) );
  AOI21_X2 U6104 ( .B1(n9662), .B2(n9661), .A(n9660), .ZN(n9664) );
  AOI21_X2 U6105 ( .B1(n9685), .B2(n9684), .A(n10155), .ZN(n9686) );
  NOR2_X2 U6106 ( .A1(n9683), .A2(n9682), .ZN(n9684) );
  NOR2_X2 U6107 ( .A1(n9676), .A2(n9675), .ZN(n9685) );
  NOR2_X2 U6108 ( .A1(n9681), .A2(n7392), .ZN(n9682) );
  OAI21_X1 U6109 ( .B1(n9980), .B2(n10230), .A(n10229), .ZN(n9697) );
  NOR2_X2 U6110 ( .A1(n9735), .A2(n9734), .ZN(n9738) );
  OAI21_X2 U6111 ( .B1(n9740), .B2(n10230), .A(n10229), .ZN(n9741) );
  OAI21_X2 U6112 ( .B1(n9755), .B2(n7392), .A(n9754), .ZN(n9759) );
  NOR2_X2 U6113 ( .A1(n9757), .A2(n6860), .ZN(n9758) );
  NAND3_X2 U6114 ( .A1(DMEM_BUS_OUT[28]), .A2(n7380), .A3(n7469), .ZN(n8477)
         );
  NOR2_X2 U6115 ( .A1(n9762), .A2(n7479), .ZN(n9766) );
  NOR2_X2 U6116 ( .A1(ID_EXEC_OUT[157]), .A2(n9838), .ZN(n9799) );
  NOR2_X2 U6117 ( .A1(n10268), .A2(n10098), .ZN(n10101) );
  AOI21_X2 U6118 ( .B1(n10122), .B2(n10121), .A(n10155), .ZN(n10123) );
  NOR2_X2 U6119 ( .A1(n10120), .A2(n10119), .ZN(n10121) );
  AOI21_X2 U6120 ( .B1(n6799), .B2(n10275), .A(n10118), .ZN(n10122) );
  NOR2_X2 U6121 ( .A1(n7138), .A2(n7393), .ZN(n10120) );
  AOI21_X2 U6122 ( .B1(n10106), .B2(n10229), .A(n10105), .ZN(n10124) );
  AOI21_X2 U6123 ( .B1(n10157), .B2(n10156), .A(n10155), .ZN(n10158) );
  NOR2_X2 U6124 ( .A1(n10145), .A2(n10144), .ZN(n10157) );
  NOR2_X2 U6125 ( .A1(n10154), .A2(n10153), .ZN(n10156) );
  NOR2_X2 U6126 ( .A1(n10143), .A2(n7392), .ZN(n10144) );
  AOI21_X2 U6127 ( .B1(n10137), .B2(n10229), .A(n10136), .ZN(n10159) );
  OAI21_X2 U6128 ( .B1(n6917), .B2(n10274), .A(n10171), .ZN(n10182) );
  AOI21_X2 U6129 ( .B1(n10188), .B2(n10189), .A(n10167), .ZN(n10169) );
  OAI21_X2 U6130 ( .B1(n10193), .B2(n10274), .A(n10192), .ZN(n10213) );
  NOR2_X2 U6131 ( .A1(n10225), .A2(n10224), .ZN(n10227) );
  OAI21_X1 U6132 ( .B1(n10269), .B2(n10222), .A(n10221), .ZN(n10225) );
  OAI21_X2 U6133 ( .B1(n10231), .B2(n10230), .A(n10229), .ZN(n10235) );
  NOR2_X2 U6134 ( .A1(ID_EXEC_OUT[156]), .A2(ID_EXEC_OUT[157]), .ZN(n8505) );
  OAI21_X2 U6135 ( .B1(n6188), .B2(n10274), .A(n10273), .ZN(n10284) );
  AOI21_X2 U6136 ( .B1(n10268), .B2(n10267), .A(n10266), .ZN(n10270) );
  INV_X4 U6137 ( .A(n10230), .ZN(n10264) );
  NOR2_X2 U6138 ( .A1(EXEC_MEM_OUT_141), .A2(n5398), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N41) );
  NOR2_X2 U6139 ( .A1(n7773), .A2(n3332), .ZN(ID_EX_REG_ID_EX_REG_N50) );
  NOR2_X2 U6140 ( .A1(n9862), .A2(n9861), .ZN(n9870) );
  NOR3_X2 U6141 ( .A1(n9030), .A2(n9029), .A3(n9028), .ZN(n9031) );
  NOR2_X2 U6142 ( .A1(n9652), .A2(n9804), .ZN(n9028) );
  NOR2_X2 U6143 ( .A1(n10289), .A2(n7391), .ZN(n9030) );
  NOR3_X2 U6144 ( .A1(n10004), .A2(n10271), .A3(n7348), .ZN(n9952) );
  NOR2_X2 U6145 ( .A1(n10271), .A2(n9954), .ZN(n9957) );
  AOI21_X2 U6146 ( .B1(n9949), .B2(n9948), .A(n9947), .ZN(n9960) );
  AOI21_X2 U6147 ( .B1(n9942), .B2(n9945), .A(n9941), .ZN(n9949) );
  NOR3_X2 U6148 ( .A1(n9933), .A2(n9932), .A3(n9931), .ZN(n9934) );
  OAI21_X2 U6149 ( .B1(n9907), .B2(n9906), .A(n9905), .ZN(n9935) );
  INV_X4 U6150 ( .A(n9893), .ZN(n9907) );
  NOR3_X2 U6151 ( .A1(n9904), .A2(n9903), .A3(n9902), .ZN(n9905) );
  NOR3_X2 U6152 ( .A1(n9848), .A2(n9847), .A3(n9904), .ZN(n9884) );
  AOI21_X2 U6153 ( .B1(n9882), .B2(n9881), .A(n9880), .ZN(n9883) );
  NOR2_X2 U6154 ( .A1(n9846), .A2(n9845), .ZN(n9847) );
  INV_X4 U6155 ( .A(n10067), .ZN(n10010) );
  NOR2_X2 U6156 ( .A1(n9776), .A2(n7338), .ZN(n9777) );
  NOR2_X2 U6157 ( .A1(n9773), .A2(n9772), .ZN(n9774) );
  NAND2_X2 U6158 ( .A1(n9844), .A2(n9764), .ZN(n9195) );
  NAND2_X2 U6159 ( .A1(n7943), .A2(n8014), .ZN(n8024) );
  NOR2_X2 U6160 ( .A1(n6348), .A2(n6868), .ZN(n4093) );
  NOR2_X2 U6161 ( .A1(n6348), .A2(offset_26_id[3]), .ZN(n4094) );
  NOR2_X2 U6162 ( .A1(n5861), .A2(offset_26_id[8]), .ZN(n4846) );
  NOR2_X2 U6163 ( .A1(n5856), .A2(offset_26_id[9]), .ZN(n4845) );
  NOR2_X2 U6164 ( .A1(n5861), .A2(n5856), .ZN(n4847) );
  NOR3_X2 U6165 ( .A1(n10055), .A2(n10054), .A3(n10053), .ZN(n10057) );
  INV_X4 U6166 ( .A(n10028), .ZN(n10074) );
  NOR2_X2 U6167 ( .A1(n10062), .A2(n10061), .ZN(n10065) );
  NOR2_X2 U6168 ( .A1(n9611), .A2(n9094), .ZN(n9095) );
  NAND2_X2 U6169 ( .A1(n7900), .A2(n8025), .ZN(n9223) );
  NOR2_X2 U6170 ( .A1(n6352), .A2(n6913), .ZN(n7899) );
  OAI21_X2 U6171 ( .B1(EXEC_STAGE_imm26_32[11]), .B2(n8135), .A(n5846), .ZN(
        n8137) );
  OAI21_X2 U6172 ( .B1(EXEC_STAGE_imm26_32[13]), .B2(n8133), .A(n5846), .ZN(
        n8147) );
  NOR3_X2 U6173 ( .A1(n8177), .A2(n8186), .A3(n6912), .ZN(n8181) );
  NOR2_X2 U6174 ( .A1(n8368), .A2(n8184), .ZN(n8300) );
  NAND2_X2 U6175 ( .A1(n7453), .A2(n6334), .ZN(n8216) );
  OAI21_X2 U6176 ( .B1(EXEC_STAGE_imm26_32[15]), .B2(n8138), .A(n5845), .ZN(
        n8141) );
  BUF_X4 U6177 ( .A(n8653), .Z(n7322) );
  NAND3_X2 U6178 ( .A1(n8711), .A2(n8712), .A3(n8751), .ZN(n8560) );
  OAI21_X2 U6179 ( .B1(n8623), .B2(n7383), .A(n8622), .ZN(n8685) );
  NOR2_X2 U6180 ( .A1(n6991), .A2(n8024), .ZN(n7857) );
  NOR2_X2 U6181 ( .A1(n7942), .A2(n7856), .ZN(n7858) );
  NAND3_X2 U6182 ( .A1(DMEM_BUS_OUT[31]), .A2(n8070), .A3(n7462), .ZN(n9770)
         );
  NOR2_X2 U6183 ( .A1(n6868), .A2(offset_26_id[4]), .ZN(n4091) );
  NOR3_X2 U6184 ( .A1(n7447), .A2(n10299), .A3(n1652), .ZN(n4077) );
  NOR3_X2 U6185 ( .A1(n10299), .A2(offset_26_id[0]), .A3(n3747), .ZN(n4069) );
  INV_X4 U6186 ( .A(n7944), .ZN(n7945) );
  NOR3_X2 U6187 ( .A1(n6996), .A2(n7329), .A3(n7771), .ZN(n7946) );
  INV_X4 U6188 ( .A(n6900), .ZN(n7312) );
  NAND3_X2 U6189 ( .A1(n3092), .A2(n6349), .A3(n8114), .ZN(n8118) );
  NOR2_X2 U6190 ( .A1(offset_26_id[3]), .A2(offset_26_id[4]), .ZN(n4089) );
  NOR3_X2 U6191 ( .A1(n7888), .A2(n7771), .A3(n7223), .ZN(n7959) );
  OAI21_X2 U6192 ( .B1(n7380), .B2(n7227), .A(n8447), .ZN(n8450) );
  INV_X4 U6193 ( .A(n9055), .ZN(n8439) );
  NOR2_X2 U6194 ( .A1(n7449), .A2(n9786), .ZN(n8438) );
  NAND3_X2 U6195 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[22]), .A2(n7943), 
        .A3(n8014), .ZN(n8015) );
  NAND3_X2 U6196 ( .A1(MEM_WB_OUT[67]), .A2(n7223), .A3(n7772), .ZN(n8016) );
  NAND3_X2 U6197 ( .A1(n8617), .A2(n8637), .A3(n8616), .ZN(n9036) );
  NOR2_X2 U6198 ( .A1(n8615), .A2(n8614), .ZN(n8616) );
  NOR2_X2 U6199 ( .A1(n9538), .A2(n7385), .ZN(n8525) );
  NAND3_X2 U6200 ( .A1(n8536), .A2(n8637), .A3(n8535), .ZN(n9340) );
  NOR2_X2 U6201 ( .A1(n8534), .A2(n6911), .ZN(n8535) );
  NAND2_X2 U6202 ( .A1(n8957), .A2(n8681), .ZN(n8653) );
  NAND2_X2 U6203 ( .A1(n8491), .A2(n8490), .ZN(n9090) );
  INV_X4 U6204 ( .A(n7915), .ZN(n7958) );
  OAI21_X2 U6205 ( .B1(n8648), .B2(n8478), .A(n6895), .ZN(n8954) );
  NAND3_X2 U6206 ( .A1(n8523), .A2(n8637), .A3(n8522), .ZN(n8977) );
  NOR2_X2 U6207 ( .A1(n8521), .A2(n8520), .ZN(n8522) );
  NAND3_X2 U6208 ( .A1(n8632), .A2(n8637), .A3(n8631), .ZN(n9537) );
  NOR2_X2 U6209 ( .A1(n8630), .A2(n8629), .ZN(n8631) );
  NOR2_X2 U6210 ( .A1(n9531), .A2(n9806), .ZN(n8538) );
  NAND2_X2 U6211 ( .A1(n9294), .A2(n9296), .ZN(n9655) );
  NOR2_X2 U6212 ( .A1(n7450), .A2(ID_EXEC_OUT[158]), .ZN(n10084) );
  NAND2_X2 U6213 ( .A1(n7340), .A2(n10027), .ZN(n10023) );
  NOR3_X2 U6214 ( .A1(n9791), .A2(n9790), .A3(n9789), .ZN(n9792) );
  NOR3_X2 U6215 ( .A1(n9785), .A2(n9996), .A3(n9784), .ZN(n9793) );
  NAND3_X2 U6216 ( .A1(n9366), .A2(n9365), .A3(n9364), .ZN(n10138) );
  NAND2_X2 U6217 ( .A1(n9656), .A2(n9655), .ZN(n9690) );
  NAND3_X2 U6218 ( .A1(n9635), .A2(n9634), .A3(n9633), .ZN(n10203) );
  INV_X4 U6219 ( .A(n7451), .ZN(n8072) );
  NAND3_X2 U6220 ( .A1(n9801), .A2(n9590), .A3(n9589), .ZN(n10236) );
  NAND3_X2 U6221 ( .A1(n9671), .A2(n9670), .A3(n9669), .ZN(n10237) );
  NAND2_X2 U6222 ( .A1(n10100), .A2(n10099), .ZN(n9301) );
  INV_X4 U6223 ( .A(n7308), .ZN(n7451) );
  NOR2_X2 U6224 ( .A1(IMEM_BUS_IN[1]), .A2(IMEM_BUS_IN[3]), .ZN(n3294) );
  NOR3_X2 U6225 ( .A1(ID_STAGE_imm16_aluA[27]), .A2(ID_STAGE_imm16_aluA[28]), 
        .A3(ID_STAGE_imm16_aluA[26]), .ZN(n3375) );
  NOR2_X2 U6226 ( .A1(n7806), .A2(n7805), .ZN(n7809) );
  NOR3_X2 U6227 ( .A1(n7807), .A2(n5869), .A3(n6908), .ZN(n7808) );
  NOR2_X2 U6228 ( .A1(n3237), .A2(n6894), .ZN(n3235) );
  OAI21_X2 U6229 ( .B1(n8264), .B2(n8239), .A(n8238), .ZN(n8240) );
  NAND3_X2 U6230 ( .A1(n3239), .A2(IMEM_BUS_OUT[4]), .A3(IMEM_BUS_OUT[3]), 
        .ZN(n3237) );
  NOR3_X2 U6231 ( .A1(n3243), .A2(n6015), .A3(n6906), .ZN(n3239) );
  OAI22_X2 U6232 ( .A1(n8150), .A2(n7211), .B1(n8324), .B2(n8329), .ZN(n8304)
         );
  OAI21_X2 U6233 ( .B1(n8196), .B2(n6037), .A(n6521), .ZN(n8561) );
  OAI21_X2 U6234 ( .B1(n6912), .B2(n8586), .A(n8366), .ZN(n8559) );
  NOR2_X2 U6235 ( .A1(n8612), .A2(n8611), .ZN(n8621) );
  NOR2_X2 U6236 ( .A1(n8619), .A2(n8618), .ZN(n8620) );
  NOR2_X2 U6237 ( .A1(n9032), .A2(n7388), .ZN(n8611) );
  NAND3_X2 U6238 ( .A1(n8473), .A2(n8472), .A3(n8471), .ZN(n8682) );
  AOI21_X2 U6239 ( .B1(n4726), .B2(n4727), .A(n7553), .ZN(n4725) );
  AOI21_X2 U6240 ( .B1(n4730), .B2(n4731), .A(n7519), .ZN(n4724) );
  AOI21_X2 U6241 ( .B1(n4734), .B2(n4735), .A(n7517), .ZN(n4723) );
  NOR2_X2 U6242 ( .A1(n9245), .A2(n7803), .ZN(n7437) );
  INV_X4 U6243 ( .A(reset), .ZN(n7804) );
  INV_X4 U6244 ( .A(n7803), .ZN(n7795) );
  INV_X4 U6245 ( .A(reset), .ZN(n7803) );
  NOR3_X2 U6246 ( .A1(n8112), .A2(n8114), .A3(n6349), .ZN(n8113) );
  INV_X4 U6247 ( .A(n7800), .ZN(n7796) );
  NOR3_X2 U6248 ( .A1(offset_26_id[1]), .A2(offset_26_id[6]), .A3(
        offset_26_id[5]), .ZN(n4814) );
  NAND3_X2 U6249 ( .A1(n6353), .A2(n6899), .A3(n6022), .ZN(n4815) );
  OAI21_X2 U6250 ( .B1(n7450), .B2(n9786), .A(n7366), .ZN(n9055) );
  OAI211_X2 U6251 ( .C1(n9293), .C2(n6030), .A(n9138), .B(n9137), .ZN(n9926)
         );
  OAI21_X2 U6252 ( .B1(n6350), .B2(n9202), .A(n9201), .ZN(n9203) );
  OAI21_X2 U6253 ( .B1(n9199), .B2(n9417), .A(n9198), .ZN(n9200) );
  AOI21_X2 U6254 ( .B1(n7478), .B2(n9413), .A(n9192), .ZN(n9193) );
  OAI21_X2 U6255 ( .B1(n9077), .B2(n9076), .A(n6990), .ZN(n9330) );
  NOR3_X2 U6256 ( .A1(n6911), .A2(n9150), .A3(n9149), .ZN(n9168) );
  AOI21_X2 U6257 ( .B1(n7478), .B2(n9436), .A(n9166), .ZN(n9167) );
  NOR2_X2 U6258 ( .A1(n9147), .A2(n9804), .ZN(n9150) );
  NOR2_X2 U6259 ( .A1(n9419), .A2(n7392), .ZN(n9420) );
  OAI21_X2 U6260 ( .B1(n6350), .B2(n7388), .A(n9417), .ZN(n9418) );
  OAI21_X2 U6261 ( .B1(n9444), .B2(n9443), .A(n10282), .ZN(n9455) );
  OAI21_X2 U6262 ( .B1(n10281), .B2(n9435), .A(n9434), .ZN(n9444) );
  OAI21_X2 U6263 ( .B1(n9969), .B2(n10230), .A(n10229), .ZN(n9446) );
  OAI21_X2 U6264 ( .B1(n9864), .B2(n9346), .A(n9345), .ZN(n9511) );
  INV_X4 U6265 ( .A(n10046), .ZN(n10044) );
  NAND3_X2 U6266 ( .A1(n9378), .A2(n9377), .A3(n9376), .ZN(n9628) );
  NOR2_X2 U6267 ( .A1(n7224), .A2(n6860), .ZN(n9675) );
  NOR2_X2 U6268 ( .A1(n7035), .A2(n10255), .ZN(n9676) );
  NOR2_X2 U6269 ( .A1(n9745), .A2(n7393), .ZN(n9683) );
  INV_X16 U6270 ( .A(n7464), .ZN(n7463) );
  INV_X4 U6271 ( .A(n10255), .ZN(n9753) );
  NOR2_X2 U6272 ( .A1(n8635), .A2(n8634), .ZN(n8636) );
  NOR2_X2 U6273 ( .A1(n9665), .A2(n7391), .ZN(n8634) );
  INV_X16 U6274 ( .A(n7470), .ZN(n7469) );
  NAND2_X2 U6275 ( .A1(n9819), .A2(n9837), .ZN(n9820) );
  NOR2_X2 U6276 ( .A1(n9841), .A2(n9840), .ZN(n10083) );
  NOR2_X2 U6277 ( .A1(n9839), .A2(n9838), .ZN(n9840) );
  NAND3_X2 U6278 ( .A1(n7449), .A2(n7366), .A3(n6799), .ZN(n9836) );
  NOR2_X2 U6279 ( .A1(n10117), .A2(n10255), .ZN(n10118) );
  NOR2_X2 U6280 ( .A1(n7225), .A2(n6860), .ZN(n10119) );
  NOR2_X2 U6281 ( .A1(n7208), .A2(n10255), .ZN(n10153) );
  NOR2_X2 U6282 ( .A1(n7139), .A2(n7393), .ZN(n10154) );
  NOR2_X2 U6283 ( .A1(n6917), .A2(n6860), .ZN(n10145) );
  NOR3_X2 U6284 ( .A1(n7930), .A2(n7929), .A3(n7928), .ZN(n8082) );
  NOR3_X2 U6285 ( .A1(n8051), .A2(n8050), .A3(n8049), .ZN(n8080) );
  NAND3_X2 U6286 ( .A1(n7814), .A2(n7774), .A3(n6869), .ZN(n8119) );
  INV_X4 U6287 ( .A(n8119), .ZN(n10300) );
  NAND3_X2 U6288 ( .A1(n7814), .A2(n7774), .A3(n6869), .ZN(n7354) );
  NOR3_X2 U6289 ( .A1(n7374), .A2(n8245), .A3(n8244), .ZN(n8247) );
  NOR2_X2 U6290 ( .A1(n8249), .A2(n7374), .ZN(n8242) );
  NOR3_X2 U6291 ( .A1(n7374), .A2(n8249), .A3(n8248), .ZN(n8250) );
  INV_X4 U6292 ( .A(n8263), .ZN(n8269) );
  NOR2_X2 U6293 ( .A1(n6015), .A2(n3243), .ZN(n3245) );
  OAI21_X2 U6294 ( .B1(n8222), .B2(n8221), .A(n8220), .ZN(n8281) );
  OAI21_X2 U6295 ( .B1(n8284), .B2(n8217), .A(n6190), .ZN(n8221) );
  NOR3_X2 U6296 ( .A1(n8285), .A2(n8217), .A3(n8286), .ZN(n8222) );
  NAND2_X2 U6297 ( .A1(n6186), .A2(n8281), .ZN(n8280) );
  NOR2_X2 U6298 ( .A1(n3251), .A2(n1996), .ZN(n3253) );
  NOR2_X2 U6299 ( .A1(n3259), .A2(n5909), .ZN(n3261) );
  NOR2_X2 U6300 ( .A1(n3267), .A2(n6877), .ZN(n3269) );
  NOR3_X2 U6301 ( .A1(n4542), .A2(n4543), .A3(n4544), .ZN(n4541) );
  NOR2_X2 U6302 ( .A1(n3275), .A2(n2008), .ZN(n3277) );
  NOR2_X2 U6303 ( .A1(n3283), .A2(n2012), .ZN(n3285) );
  NOR3_X2 U6304 ( .A1(n4677), .A2(n4678), .A3(n4679), .ZN(n4676) );
  AOI21_X2 U6305 ( .B1(n8654), .B2(n8951), .A(n7479), .ZN(n8657) );
  OAI21_X2 U6306 ( .B1(n7352), .B2(n10230), .A(n10229), .ZN(n8647) );
  NOR3_X2 U6307 ( .A1(n4700), .A2(n4701), .A3(n4702), .ZN(n4699) );
  OAI21_X2 U6308 ( .B1(n9844), .B2(n10230), .A(n10229), .ZN(n8737) );
  OAI21_X2 U6309 ( .B1(n8736), .B2(n8735), .A(n10257), .ZN(n8746) );
  NAND3_X2 U6310 ( .A1(n7616), .A2(n7775), .A3(n7773), .ZN(n3184) );
  NOR3_X2 U6311 ( .A1(n4475), .A2(n4476), .A3(n4477), .ZN(n4474) );
  NOR3_X2 U6312 ( .A1(n4497), .A2(n4498), .A3(n4499), .ZN(n4496) );
  NOR3_X2 U6313 ( .A1(n4520), .A2(n4521), .A3(n4522), .ZN(n4519) );
  NOR3_X2 U6314 ( .A1(n4564), .A2(n4565), .A3(n4566), .ZN(n4563) );
  NOR3_X2 U6315 ( .A1(n4586), .A2(n4587), .A3(n4588), .ZN(n4585) );
  NOR3_X2 U6316 ( .A1(n4609), .A2(n4610), .A3(n4611), .ZN(n4608) );
  NOR3_X2 U6317 ( .A1(n4632), .A2(n4633), .A3(n4634), .ZN(n4631) );
  NOR3_X2 U6318 ( .A1(n4405), .A2(n4406), .A3(n4407), .ZN(n4404) );
  NOR3_X2 U6319 ( .A1(n4428), .A2(n4429), .A3(n4430), .ZN(n4427) );
  NOR3_X2 U6320 ( .A1(n4453), .A2(n4454), .A3(n4455), .ZN(n4452) );
  NOR3_X2 U6321 ( .A1(n4654), .A2(n4655), .A3(n4656), .ZN(n4653) );
  NOR3_X2 U6322 ( .A1(n4745), .A2(n4746), .A3(n4747), .ZN(n4744) );
  NOR3_X2 U6323 ( .A1(n4767), .A2(n4768), .A3(n4769), .ZN(n4766) );
  NOR3_X2 U6324 ( .A1(n4789), .A2(n4790), .A3(n4791), .ZN(n4788) );
  NAND2_X2 U6325 ( .A1(n7794), .A2(n8909), .ZN(n8910) );
  NAND2_X2 U6326 ( .A1(n7794), .A2(n8909), .ZN(n7435) );
  NAND2_X2 U6327 ( .A1(n7794), .A2(n8909), .ZN(n7436) );
  NOR3_X2 U6328 ( .A1(n4270), .A2(n4271), .A3(n4272), .ZN(n4269) );
  AOI211_X2 U6329 ( .C1(n9169), .C2(n7457), .A(n7245), .B(n8102), .ZN(n1634)
         );
  NOR2_X2 U6330 ( .A1(n4098), .A2(n4099), .ZN(n8102) );
  AOI211_X2 U6331 ( .C1(n8106), .C2(n7457), .A(n7244), .B(n8101), .ZN(n1633)
         );
  NOR2_X2 U6332 ( .A1(n4133), .A2(n4099), .ZN(n8101) );
  NOR3_X2 U6333 ( .A1(n4315), .A2(n4316), .A3(n4317), .ZN(n4314) );
  AOI211_X2 U6334 ( .C1(n8109), .C2(n7457), .A(n7242), .B(n8094), .ZN(n1631)
         );
  NOR2_X2 U6335 ( .A1(n4178), .A2(n4099), .ZN(n8094) );
  NOR3_X2 U6336 ( .A1(n4360), .A2(n4361), .A3(n4362), .ZN(n4359) );
  AOI211_X2 U6337 ( .C1(n9234), .C2(n7457), .A(n7240), .B(n8090), .ZN(n1629)
         );
  NOR2_X2 U6338 ( .A1(n4223), .A2(n4099), .ZN(n8090) );
  NOR3_X2 U6339 ( .A1(n4248), .A2(n4249), .A3(n4250), .ZN(n4247) );
  NOR3_X2 U6340 ( .A1(n4293), .A2(n4294), .A3(n4295), .ZN(n4292) );
  AOI211_X2 U6341 ( .C1(n9215), .C2(n7457), .A(n7243), .B(n8098), .ZN(n1632)
         );
  NOR2_X2 U6342 ( .A1(n4155), .A2(n4099), .ZN(n8098) );
  NOR3_X2 U6343 ( .A1(n4338), .A2(n4339), .A3(n4340), .ZN(n4337) );
  AOI211_X2 U6344 ( .C1(n9230), .C2(n7457), .A(n7241), .B(n8091), .ZN(n1630)
         );
  NOR2_X2 U6345 ( .A1(n4200), .A2(n4099), .ZN(n8091) );
  NOR3_X2 U6346 ( .A1(n4383), .A2(n4384), .A3(n4385), .ZN(n4382) );
  OAI21_X2 U6347 ( .B1(n6865), .B2(n1592), .A(n3325), .ZN(n3292) );
  NAND2_X2 U6348 ( .A1(n8043), .A2(n8909), .ZN(n8021) );
  OAI21_X2 U6349 ( .B1(n9067), .B2(n9066), .A(n10257), .ZN(n9072) );
  NOR2_X2 U6350 ( .A1(n9818), .A2(n7393), .ZN(n9067) );
  OAI21_X2 U6351 ( .B1(n9965), .B2(n10230), .A(n10229), .ZN(n9386) );
  AOI21_X2 U6352 ( .B1(n9387), .B2(n9449), .A(n7479), .ZN(n9395) );
  NAND3_X2 U6353 ( .A1(n9460), .A2(n9459), .A3(n6916), .ZN(n9461) );
  NOR2_X2 U6354 ( .A1(n7324), .A2(n9450), .ZN(n9462) );
  NAND3_X2 U6355 ( .A1(n9453), .A2(n9449), .A3(n9480), .ZN(n9450) );
  NOR2_X2 U6356 ( .A1(n1591), .A2(n7447), .ZN(n4447) );
  NOR3_X2 U6357 ( .A1(n4818), .A2(n4819), .A3(n4820), .ZN(n4817) );
  NOR2_X2 U6358 ( .A1(EXEC_MEM_OUT_141), .A2(n3360), .ZN(
        ID_EX_REG_ID_EX_REG_N47) );
  AOI21_X2 U6359 ( .B1(n3348), .B2(n3349), .A(EXEC_MEM_OUT_141), .ZN(
        ID_EX_REG_ID_EX_REG_N48) );
  NOR2_X2 U6360 ( .A1(n3335), .A2(n3356), .ZN(n3348) );
  NOR2_X2 U6361 ( .A1(ID_STAGE_imm16_aluA[31]), .A2(n6862), .ZN(n3350) );
  NOR2_X2 U6362 ( .A1(n7773), .A2(n3337), .ZN(ID_EX_REG_ID_EX_REG_N49) );
  OAI21_X2 U6363 ( .B1(n6347), .B2(n3341), .A(n3342), .ZN(n3338) );
  NAND3_X2 U6364 ( .A1(ID_STAGE_imm16_aluA[31]), .A2(ID_STAGE_imm16_aluA[28]), 
        .A3(n1589), .ZN(n3342) );
  NAND3_X2 U6365 ( .A1(n8125), .A2(n8229), .A3(n8124), .ZN(n8237) );
  OAI21_X2 U6366 ( .B1(n8132), .B2(n8131), .A(n8130), .ZN(n8236) );
  NOR3_X2 U6367 ( .A1(n8267), .A2(n8266), .A3(n8265), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N71) );
  NOR2_X2 U6368 ( .A1(n8759), .A2(n8258), .ZN(n8266) );
  AOI21_X2 U6369 ( .B1(n8264), .B2(n8263), .A(n8262), .ZN(n8265) );
  NOR2_X2 U6370 ( .A1(n8257), .A2(n8256), .ZN(n8267) );
  OAI21_X2 U6371 ( .B1(n8279), .B2(n7374), .A(n8278), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N68) );
  OAI21_X2 U6372 ( .B1(n7374), .B2(n8290), .A(n8289), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N66) );
  AOI211_X2 U6373 ( .C1(n8295), .C2(n8294), .A(n8293), .B(n6357), .ZN(n8299)
         );
  OAI21_X2 U6374 ( .B1(n7374), .B2(n8313), .A(n8312), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N64) );
  NAND2_X2 U6375 ( .A1(EXEC_MEM_OUT_119), .A2(n1541), .ZN(n3229) );
  OAI21_X2 U6376 ( .B1(n8318), .B2(n8317), .A(n8316), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N63) );
  NOR2_X2 U6377 ( .A1(n5915), .A2(n8314), .ZN(n8318) );
  OAI21_X2 U6378 ( .B1(n8322), .B2(n7374), .A(n8321), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N62) );
  OAI21_X2 U6379 ( .B1(n8333), .B2(n8332), .A(n8331), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N61) );
  NOR2_X2 U6380 ( .A1(n8327), .A2(n8328), .ZN(n8333) );
  OAI21_X2 U6381 ( .B1(n8330), .B2(n8329), .A(n8759), .ZN(n8332) );
  OAI21_X2 U6382 ( .B1(n8341), .B2(n7374), .A(n8340), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N60) );
  OAI21_X2 U6383 ( .B1(n8350), .B2(n8349), .A(n8348), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N59) );
  NOR2_X2 U6384 ( .A1(n8344), .A2(n8345), .ZN(n8350) );
  OAI21_X2 U6385 ( .B1(n8347), .B2(n8346), .A(n8759), .ZN(n8349) );
  OAI21_X2 U6386 ( .B1(n8358), .B2(n7374), .A(n8357), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N58) );
  OAI21_X2 U6387 ( .B1(n8364), .B2(n8363), .A(n8362), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N57) );
  NOR2_X2 U6388 ( .A1(n8360), .A2(n8359), .ZN(n8364) );
  OAI21_X2 U6389 ( .B1(n7374), .B2(n8375), .A(n8374), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N56) );
  OAI21_X2 U6390 ( .B1(n8389), .B2(n8388), .A(n8387), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N55) );
  AOI211_X2 U6391 ( .C1(n8385), .C2(n8384), .A(n8383), .B(n8382), .ZN(n8389)
         );
  OAI21_X2 U6392 ( .B1(n8397), .B2(n7374), .A(n8396), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N54) );
  OAI21_X2 U6393 ( .B1(n3816), .B2(n3817), .A(n7575), .ZN(n3809) );
  OAI21_X2 U6394 ( .B1(n3820), .B2(n3821), .A(n7558), .ZN(n3808) );
  OAI21_X2 U6395 ( .B1(n3824), .B2(n3825), .A(n7556), .ZN(n3807) );
  AOI21_X2 U6396 ( .B1(n10264), .B2(n9915), .A(n6844), .ZN(n8549) );
  OAI21_X2 U6397 ( .B1(n8546), .B2(n8545), .A(n10282), .ZN(n8547) );
  OAI21_X2 U6398 ( .B1(n8558), .B2(n8557), .A(n8556), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N53) );
  AOI211_X2 U6399 ( .C1(n8554), .C2(n8553), .A(n8552), .B(n6918), .ZN(n8558)
         );
  OAI21_X2 U6400 ( .B1(n7374), .B2(n8572), .A(n8571), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N52) );
  OAI21_X2 U6401 ( .B1(n8579), .B2(n7374), .A(n8578), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N50) );
  OAI21_X2 U6402 ( .B1(n8589), .B2(n8588), .A(n8587), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N49) );
  AOI211_X2 U6403 ( .C1(n8584), .C2(n8583), .A(n8582), .B(n8581), .ZN(n8589)
         );
  OAI21_X2 U6404 ( .B1(n7234), .B2(n8586), .A(n8759), .ZN(n8588) );
  OAI21_X2 U6405 ( .B1(n8595), .B2(n7374), .A(n8594), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N48) );
  OAI21_X2 U6406 ( .B1(n3943), .B2(n3944), .A(n7574), .ZN(n3936) );
  OAI21_X2 U6407 ( .B1(n3947), .B2(n3948), .A(n7557), .ZN(n3935) );
  OAI21_X2 U6408 ( .B1(n3951), .B2(n3952), .A(n7555), .ZN(n3934) );
  OAI21_X2 U6409 ( .B1(n8667), .B2(n8666), .A(n8665), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N47) );
  NOR2_X2 U6410 ( .A1(n8663), .A2(n8662), .ZN(n8667) );
  OAI21_X2 U6411 ( .B1(n3964), .B2(n3965), .A(n7574), .ZN(n3957) );
  OAI21_X2 U6412 ( .B1(n3968), .B2(n3969), .A(n7557), .ZN(n3956) );
  OAI21_X2 U6413 ( .B1(n3972), .B2(n3973), .A(n7555), .ZN(n3955) );
  NOR2_X2 U6414 ( .A1(n8707), .A2(n8706), .ZN(n8708) );
  OAI21_X2 U6415 ( .B1(n7374), .B2(n8715), .A(n8714), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N46) );
  OAI21_X2 U6416 ( .B1(n3985), .B2(n3986), .A(n7574), .ZN(n3978) );
  OAI21_X2 U6417 ( .B1(n3989), .B2(n3990), .A(n7557), .ZN(n3977) );
  OAI21_X2 U6418 ( .B1(n3993), .B2(n3994), .A(n7555), .ZN(n3976) );
  AOI21_X2 U6419 ( .B1(n7448), .B2(n7305), .A(ID_EX_REG_ID_EX_REG_N99), .ZN(
        n4719) );
  OAI21_X2 U6420 ( .B1(n8753), .B2(n7374), .A(n8752), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N44) );
  NOR2_X2 U6421 ( .A1(n7618), .A2(n6476), .ZN(IF_ID_REG_IF_ID_REG_N36) );
  INV_X4 U6422 ( .A(n7797), .ZN(n7775) );
  NOR2_X2 U6423 ( .A1(n7618), .A2(n6477), .ZN(IF_ID_REG_IF_ID_REG_N35) );
  NOR2_X2 U6424 ( .A1(n7773), .A2(n5869), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N77)
         );
  NOR2_X2 U6425 ( .A1(n6868), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N91) );
  OAI21_X2 U6426 ( .B1(n3921), .B2(n3922), .A(n7574), .ZN(n3914) );
  OAI21_X2 U6427 ( .B1(n3925), .B2(n3926), .A(n7557), .ZN(n3913) );
  OAI21_X2 U6428 ( .B1(n3929), .B2(n3930), .A(n7555), .ZN(n3912) );
  NOR2_X2 U6429 ( .A1(n7216), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N76) );
  OAI21_X2 U6430 ( .B1(n3858), .B2(n3859), .A(n7574), .ZN(n3851) );
  OAI21_X2 U6431 ( .B1(n3862), .B2(n3863), .A(n7557), .ZN(n3850) );
  OAI21_X2 U6432 ( .B1(n3866), .B2(n3867), .A(n7555), .ZN(n3849) );
  NOR2_X2 U6433 ( .A1(n6899), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N79) );
  OAI21_X2 U6434 ( .B1(n3837), .B2(n3838), .A(n7574), .ZN(n3830) );
  OAI21_X2 U6435 ( .B1(n3841), .B2(n3842), .A(n7557), .ZN(n3829) );
  OAI21_X2 U6436 ( .B1(n3845), .B2(n3846), .A(n7555), .ZN(n3828) );
  NOR2_X2 U6437 ( .A1(n6353), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N80) );
  NOR2_X2 U6438 ( .A1(n6022), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N81) );
  OAI21_X2 U6439 ( .B1(n3774), .B2(n3775), .A(n7575), .ZN(n3767) );
  OAI21_X2 U6440 ( .B1(n3778), .B2(n3779), .A(n7558), .ZN(n3766) );
  OAI21_X2 U6441 ( .B1(n3782), .B2(n3783), .A(n7556), .ZN(n3765) );
  NOR2_X2 U6442 ( .A1(n6992), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N83) );
  NOR2_X2 U6443 ( .A1(n5857), .A2(EXEC_MEM_OUT_141), .ZN(
        ID_EX_REG_ID_EX_REG_N92) );
  OAI21_X2 U6444 ( .B1(n3753), .B2(n3754), .A(n7575), .ZN(n3745) );
  OAI21_X2 U6445 ( .B1(n3757), .B2(n3758), .A(n7558), .ZN(n3744) );
  OAI21_X2 U6446 ( .B1(n3761), .B2(n3762), .A(n7556), .ZN(n3743) );
  NOR2_X2 U6447 ( .A1(n6891), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N84) );
  OAI21_X2 U6448 ( .B1(n4071), .B2(n4072), .A(n7574), .ZN(n4062) );
  OAI21_X2 U6449 ( .B1(n4075), .B2(n4076), .A(n7557), .ZN(n4061) );
  OAI21_X2 U6450 ( .B1(n4080), .B2(n4081), .A(n7555), .ZN(n4060) );
  NOR2_X2 U6451 ( .A1(n6012), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N95) );
  OAI21_X2 U6452 ( .B1(n4048), .B2(n4049), .A(n7574), .ZN(n4041) );
  OAI21_X2 U6453 ( .B1(n4052), .B2(n4053), .A(n7557), .ZN(n4040) );
  OAI21_X2 U6454 ( .B1(n4056), .B2(n4057), .A(n7555), .ZN(n4039) );
  NOR2_X2 U6455 ( .A1(n6011), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N96) );
  OAI21_X2 U6456 ( .B1(n4006), .B2(n4007), .A(n7574), .ZN(n3999) );
  OAI21_X2 U6457 ( .B1(n4010), .B2(n4011), .A(n7557), .ZN(n3998) );
  OAI21_X2 U6458 ( .B1(n4014), .B2(n4015), .A(n7555), .ZN(n3997) );
  NOR2_X2 U6459 ( .A1(n6862), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N98) );
  NOR2_X2 U6460 ( .A1(n6898), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N99) );
  OAI21_X2 U6461 ( .B1(n4027), .B2(n4028), .A(n7574), .ZN(n4020) );
  OAI21_X2 U6462 ( .B1(n4031), .B2(n4032), .A(n7557), .ZN(n4019) );
  OAI21_X2 U6463 ( .B1(n4035), .B2(n4036), .A(n7555), .ZN(n4018) );
  OAI21_X2 U6464 ( .B1(n3900), .B2(n3901), .A(n7574), .ZN(n3893) );
  OAI21_X2 U6465 ( .B1(n3904), .B2(n3905), .A(n7557), .ZN(n3892) );
  OAI21_X2 U6466 ( .B1(n3908), .B2(n3909), .A(n7555), .ZN(n3891) );
  OAI21_X2 U6467 ( .B1(n3879), .B2(n3880), .A(n7574), .ZN(n3872) );
  OAI21_X2 U6468 ( .B1(n3883), .B2(n3884), .A(n7557), .ZN(n3871) );
  OAI21_X2 U6469 ( .B1(n3887), .B2(n3888), .A(n7555), .ZN(n3870) );
  OAI21_X2 U6470 ( .B1(n3795), .B2(n3796), .A(n7575), .ZN(n3788) );
  OAI21_X2 U6471 ( .B1(n3799), .B2(n3800), .A(n7558), .ZN(n3787) );
  OAI21_X2 U6472 ( .B1(n3803), .B2(n3804), .A(n7556), .ZN(n3786) );
  OAI21_X2 U6473 ( .B1(n3731), .B2(n3732), .A(n7575), .ZN(n3723) );
  OAI21_X2 U6474 ( .B1(n3735), .B2(n3736), .A(n7558), .ZN(n3722) );
  OAI21_X2 U6475 ( .B1(n3739), .B2(n3740), .A(n7556), .ZN(n3721) );
  OAI21_X2 U6476 ( .B1(n3708), .B2(n3709), .A(n7575), .ZN(n3701) );
  OAI21_X2 U6477 ( .B1(n3712), .B2(n3713), .A(n7558), .ZN(n3700) );
  OAI21_X2 U6478 ( .B1(n3716), .B2(n3717), .A(n7556), .ZN(n3699) );
  OAI21_X2 U6479 ( .B1(n3687), .B2(n3688), .A(n7575), .ZN(n3679) );
  OAI21_X2 U6480 ( .B1(n3691), .B2(n3692), .A(n7558), .ZN(n3678) );
  OAI21_X2 U6481 ( .B1(n3695), .B2(n3696), .A(n7556), .ZN(n3677) );
  OAI21_X2 U6482 ( .B1(n3665), .B2(n3666), .A(n7575), .ZN(n3658) );
  OAI21_X2 U6483 ( .B1(n3669), .B2(n3670), .A(n7558), .ZN(n3657) );
  OAI21_X2 U6484 ( .B1(n3673), .B2(n3674), .A(n7556), .ZN(n3656) );
  OAI21_X2 U6485 ( .B1(n3644), .B2(n3645), .A(n7575), .ZN(n3636) );
  OAI21_X2 U6486 ( .B1(n3648), .B2(n3649), .A(n7558), .ZN(n3635) );
  OAI21_X2 U6487 ( .B1(n3652), .B2(n3653), .A(n7556), .ZN(n3634) );
  OAI21_X2 U6488 ( .B1(n3622), .B2(n3623), .A(n7575), .ZN(n3615) );
  OAI21_X2 U6489 ( .B1(n3626), .B2(n3627), .A(n7558), .ZN(n3614) );
  OAI21_X2 U6490 ( .B1(n3630), .B2(n3631), .A(n7556), .ZN(n3613) );
  OAI21_X2 U6491 ( .B1(n3601), .B2(n3602), .A(n7575), .ZN(n3593) );
  OAI21_X2 U6492 ( .B1(n3605), .B2(n3606), .A(n7558), .ZN(n3592) );
  OAI21_X2 U6493 ( .B1(n3609), .B2(n3610), .A(n7556), .ZN(n3591) );
  OAI21_X2 U6494 ( .B1(n3579), .B2(n3580), .A(n7575), .ZN(n3572) );
  OAI21_X2 U6495 ( .B1(n3583), .B2(n3584), .A(n7558), .ZN(n3571) );
  OAI21_X2 U6496 ( .B1(n3587), .B2(n3588), .A(n7556), .ZN(n3570) );
  OAI21_X2 U6497 ( .B1(n3558), .B2(n3559), .A(n7575), .ZN(n3550) );
  OAI21_X2 U6498 ( .B1(n3566), .B2(n3567), .A(n7556), .ZN(n3548) );
  OAI21_X2 U6499 ( .B1(n3562), .B2(n3563), .A(n7558), .ZN(n3549) );
  OAI21_X2 U6500 ( .B1(n3536), .B2(n3537), .A(n7574), .ZN(n3529) );
  OAI21_X2 U6501 ( .B1(n3544), .B2(n3545), .A(n7555), .ZN(n3527) );
  OAI21_X2 U6502 ( .B1(n3540), .B2(n3541), .A(n7557), .ZN(n3528) );
  OAI21_X2 U6503 ( .B1(n3515), .B2(n3516), .A(n7575), .ZN(n3507) );
  OAI21_X2 U6504 ( .B1(n3523), .B2(n3524), .A(n7556), .ZN(n3505) );
  OAI21_X2 U6505 ( .B1(n3519), .B2(n3520), .A(n7558), .ZN(n3506) );
  OAI21_X2 U6506 ( .B1(n3493), .B2(n3494), .A(n7574), .ZN(n3486) );
  OAI21_X2 U6507 ( .B1(n3501), .B2(n3502), .A(n7555), .ZN(n3484) );
  OAI21_X2 U6508 ( .B1(n3497), .B2(n3498), .A(n7557), .ZN(n3485) );
  OAI21_X2 U6509 ( .B1(n3472), .B2(n3473), .A(n7575), .ZN(n3464) );
  OAI21_X2 U6510 ( .B1(n3480), .B2(n3481), .A(n7556), .ZN(n3462) );
  OAI21_X2 U6511 ( .B1(n3476), .B2(n3477), .A(n7558), .ZN(n3463) );
  OAI21_X2 U6512 ( .B1(n3450), .B2(n3451), .A(n7574), .ZN(n3443) );
  OAI21_X2 U6513 ( .B1(n3458), .B2(n3459), .A(n7555), .ZN(n3441) );
  OAI21_X2 U6514 ( .B1(n3454), .B2(n3455), .A(n7557), .ZN(n3442) );
  OAI21_X2 U6515 ( .B1(n3429), .B2(n3430), .A(n7575), .ZN(n3421) );
  OAI21_X2 U6516 ( .B1(n3437), .B2(n3438), .A(n7556), .ZN(n3419) );
  OAI21_X2 U6517 ( .B1(n3433), .B2(n3434), .A(n7558), .ZN(n3420) );
  OAI21_X2 U6518 ( .B1(n3402), .B2(n3403), .A(n7574), .ZN(n3387) );
  OAI21_X2 U6519 ( .B1(n3414), .B2(n3415), .A(n7555), .ZN(n3385) );
  OAI21_X2 U6520 ( .B1(n3409), .B2(n3410), .A(n7557), .ZN(n3386) );
  NOR2_X2 U6521 ( .A1(n6016), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N93) );
  NOR2_X2 U6522 ( .A1(n6886), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N94) );
  NOR2_X2 U6523 ( .A1(n1656), .A2(n6343), .ZN(ID_EX_REG_ID_EX_REG_N62) );
  NOR2_X2 U6524 ( .A1(n3322), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N61) );
  NOR2_X2 U6525 ( .A1(EXEC_MEM_OUT_141), .A2(n6354), .ZN(
        ID_EX_REG_ID_EX_REG_N39) );
  NOR2_X2 U6526 ( .A1(n5861), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N85) );
  NOR2_X2 U6527 ( .A1(n7773), .A2(n6355), .ZN(ID_EX_REG_ID_EX_REG_N40) );
  NOR2_X2 U6528 ( .A1(EXEC_MEM_OUT_141), .A2(n1629), .ZN(
        ID_EX_REG_ID_EX_REG_N41) );
  NOR2_X2 U6529 ( .A1(n7773), .A2(n1630), .ZN(ID_EX_REG_ID_EX_REG_N42) );
  NOR2_X2 U6530 ( .A1(EXEC_MEM_OUT_141), .A2(n1631), .ZN(
        ID_EX_REG_ID_EX_REG_N43) );
  NOR2_X2 U6531 ( .A1(EXEC_MEM_OUT_141), .A2(n1632), .ZN(
        ID_EX_REG_ID_EX_REG_N44) );
  NOR2_X2 U6532 ( .A1(n7773), .A2(n1633), .ZN(ID_EX_REG_ID_EX_REG_N45) );
  NOR2_X2 U6533 ( .A1(n7773), .A2(n1634), .ZN(ID_EX_REG_ID_EX_REG_N46) );
  NOR2_X2 U6534 ( .A1(n5856), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N86) );
  OAI21_X2 U6535 ( .B1(n6354), .B2(n7445), .A(n4096), .ZN(
        ID_EX_REG_ID_EX_REG_N135) );
  OAI21_X2 U6536 ( .B1(n1634), .B2(n7445), .A(n4096), .ZN(
        ID_EX_REG_ID_EX_REG_N142) );
  OAI21_X2 U6537 ( .B1(n1633), .B2(n7445), .A(n4096), .ZN(
        ID_EX_REG_ID_EX_REG_N141) );
  OAI21_X2 U6538 ( .B1(n1631), .B2(n7445), .A(n4096), .ZN(
        ID_EX_REG_ID_EX_REG_N139) );
  OAI21_X2 U6539 ( .B1(n1629), .B2(n7445), .A(n4096), .ZN(
        ID_EX_REG_ID_EX_REG_N137) );
  OAI21_X2 U6540 ( .B1(n6355), .B2(n7445), .A(n4096), .ZN(
        ID_EX_REG_ID_EX_REG_N136) );
  OAI21_X2 U6541 ( .B1(n1632), .B2(n7445), .A(n4096), .ZN(
        ID_EX_REG_ID_EX_REG_N140) );
  OAI21_X2 U6542 ( .B1(n1630), .B2(n7445), .A(n4096), .ZN(
        ID_EX_REG_ID_EX_REG_N138) );
  NOR2_X2 U6543 ( .A1(n1641), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N87) );
  NOR2_X2 U6544 ( .A1(n7773), .A2(n5848), .ZN(ID_EX_REG_ID_EX_REG_N66) );
  NOR2_X2 U6545 ( .A1(n7773), .A2(n3301), .ZN(ID_EX_REG_ID_EX_REG_N67) );
  NOR2_X2 U6546 ( .A1(n7773), .A2(n3300), .ZN(ID_EX_REG_ID_EX_REG_N68) );
  NOR2_X2 U6547 ( .A1(n6348), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N90) );
  AOI21_X2 U6548 ( .B1(n3322), .B2(n7774), .A(ID_EX_REG_ID_EX_REG_N63), .ZN(
        n3321) );
  INV_X4 U6549 ( .A(n7802), .ZN(n7794) );
  NOR2_X2 U6550 ( .A1(IF_ID_OUT[37]), .A2(n3317), .ZN(ID_EX_REG_ID_EX_REG_N59)
         );
  OAI21_X2 U6551 ( .B1(n8988), .B2(n8987), .A(n10257), .ZN(n8989) );
  OAI21_X2 U6552 ( .B1(n9001), .B2(n9000), .A(n10257), .ZN(n9013) );
  NAND3_X2 U6553 ( .A1(n9053), .A2(n9052), .A3(n9051), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N84) );
  AOI21_X2 U6554 ( .B1(n9143), .B2(n7338), .A(n9050), .ZN(n9051) );
  OAI21_X2 U6555 ( .B1(n9043), .B2(n9042), .A(n10257), .ZN(n9053) );
  OAI21_X2 U6556 ( .B1(n9136), .B2(n9135), .A(n10257), .ZN(n9145) );
  AOI21_X2 U6557 ( .B1(n10282), .B2(n9209), .A(n9208), .ZN(n9329) );
  NOR2_X2 U6558 ( .A1(n10034), .A2(n10229), .ZN(n9208) );
  OAI21_X2 U6559 ( .B1(n9349), .B2(n9348), .A(n10282), .ZN(n9350) );
  OAI21_X2 U6560 ( .B1(n9409), .B2(n9405), .A(n7480), .ZN(n9431) );
  AOI21_X2 U6561 ( .B1(n10257), .B2(n9428), .A(n9427), .ZN(n9429) );
  NOR3_X2 U6562 ( .A1(n9465), .A2(n9464), .A3(n9463), .ZN(n10295) );
  NOR2_X2 U6563 ( .A1(n9458), .A2(n9451), .ZN(n9465) );
  NOR2_X2 U6564 ( .A1(n9462), .A2(n9461), .ZN(n9463) );
  OAI21_X2 U6565 ( .B1(n9458), .B2(n9460), .A(n9457), .ZN(n9464) );
  OAI21_X2 U6566 ( .B1(n9487), .B2(n9489), .A(n9486), .ZN(n9493) );
  OAI21_X2 U6567 ( .B1(n9520), .B2(n9519), .A(n7379), .ZN(n9521) );
  AOI21_X2 U6568 ( .B1(n10257), .B2(n9558), .A(n9557), .ZN(n9559) );
  AOI21_X2 U6569 ( .B1(n10257), .B2(n9576), .A(n9575), .ZN(n9577) );
  AOI21_X2 U6570 ( .B1(n9567), .B2(n9566), .A(n9565), .ZN(n9569) );
  OAI21_X2 U6571 ( .B1(n9607), .B2(n9606), .A(n7379), .ZN(n9608) );
  AOI21_X2 U6572 ( .B1(n10257), .B2(n9623), .A(n9622), .ZN(n9624) );
  AOI21_X2 U6573 ( .B1(n9613), .B2(n9612), .A(n9611), .ZN(n9615) );
  OAI21_X2 U6574 ( .B1(n9648), .B2(n9647), .A(n7379), .ZN(n9649) );
  NOR2_X2 U6575 ( .A1(n9687), .A2(n9686), .ZN(n9688) );
  AOI21_X2 U6576 ( .B1(n9666), .B2(n10229), .A(n9665), .ZN(n9687) );
  OAI21_X2 U6577 ( .B1(n9728), .B2(n9727), .A(n10257), .ZN(n9729) );
  OAI21_X2 U6578 ( .B1(n9748), .B2(n9747), .A(n7379), .ZN(n9749) );
  AOI21_X2 U6579 ( .B1(n9766), .B2(n7281), .A(n9765), .ZN(n9767) );
  AOI211_X2 U6580 ( .C1(n6800), .C2(n9760), .A(n9759), .B(n9758), .ZN(n9768)
         );
  OAI221_X2 U6581 ( .B1(n10097), .B2(n10096), .C1(n10095), .C2(n10094), .A(
        n10093), .ZN(n10293) );
  AOI21_X2 U6582 ( .B1(n9799), .B2(n9798), .A(n9797), .ZN(n10096) );
  NOR2_X2 U6583 ( .A1(n10124), .A2(n10123), .ZN(n10125) );
  OAI21_X2 U6584 ( .B1(n10101), .B2(n10100), .A(n10099), .ZN(n10102) );
  NOR2_X2 U6585 ( .A1(n10159), .A2(n10158), .ZN(n10160) );
  AOI21_X2 U6586 ( .B1(n10131), .B2(n10130), .A(n10129), .ZN(n10133) );
  OAI21_X2 U6587 ( .B1(n10182), .B2(n10181), .A(n7379), .ZN(n10183) );
  OAI21_X2 U6588 ( .B1(n10213), .B2(n10212), .A(n7379), .ZN(n10214) );
  OAI21_X2 U6589 ( .B1(n10259), .B2(n10258), .A(n10257), .ZN(n10260) );
  OAI21_X2 U6590 ( .B1(n10284), .B2(n10283), .A(n7379), .ZN(n10285) );
  INV_X4 U6591 ( .A(n7799), .ZN(n7786) );
  INV_X4 U6592 ( .A(n7801), .ZN(n7789) );
  INV_X4 U6593 ( .A(n7798), .ZN(n7783) );
  INV_X4 U6594 ( .A(n7801), .ZN(n7791) );
  INV_X4 U6595 ( .A(n7801), .ZN(n7790) );
  INV_X4 U6596 ( .A(n7799), .ZN(n7785) );
  NOR2_X2 U6597 ( .A1(n7618), .A2(n1575), .ZN(IF_ID_REG_IF_ID_REG_N32) );
  INV_X4 U6598 ( .A(n7799), .ZN(n7787) );
  NOR2_X2 U6599 ( .A1(n7618), .A2(n1574), .ZN(IF_ID_REG_IF_ID_REG_N34) );
  XOR2_X1 U6600 ( .A(destReg_wb_out[2]), .B(n1641), .Z(n4835) );
  INV_X4 U6601 ( .A(n9408), .ZN(n9407) );
  NOR2_X2 U6602 ( .A1(n9424), .A2(n9165), .ZN(n7336) );
  INV_X2 U6603 ( .A(n9970), .ZN(n9165) );
  INV_X4 U6604 ( .A(n7477), .ZN(n5851) );
  INV_X4 U6605 ( .A(n7477), .ZN(n5852) );
  INV_X4 U6606 ( .A(n9598), .ZN(n9588) );
  INV_X4 U6607 ( .A(n7477), .ZN(n7475) );
  NAND2_X2 U6608 ( .A1(n9844), .A2(n9876), .ZN(n9598) );
  INV_X4 U6609 ( .A(n9588), .ZN(n7477) );
  OAI221_X2 U6610 ( .B1(n10073), .B2(n10021), .C1(n10019), .C2(n10020), .A(
        n10018), .ZN(n10022) );
  NAND2_X2 U6611 ( .A1(n6479), .A2(n8422), .ZN(n5853) );
  INV_X8 U6612 ( .A(n7380), .ZN(n7381) );
  INV_X8 U6613 ( .A(n9270), .ZN(n7380) );
  INV_X4 U6614 ( .A(n8493), .ZN(n8492) );
  NOR2_X2 U6615 ( .A1(n6351), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N88) );
  XNOR2_X1 U6616 ( .A(n10187), .B(n9989), .ZN(n7319) );
  BUF_X16 U6617 ( .A(n10187), .Z(n7315) );
  OAI21_X2 U6618 ( .B1(n10024), .B2(n10023), .A(n10022), .ZN(n10025) );
  NAND4_X1 U6619 ( .A1(n10031), .A2(n10030), .A3(n10043), .A4(n10029), .ZN(
        n10042) );
  NAND2_X4 U6620 ( .A1(n9975), .A2(n9974), .ZN(n10043) );
  INV_X1 U6621 ( .A(n8408), .ZN(n7805) );
  AND2_X4 U6622 ( .A1(n8408), .A2(n8407), .ZN(n6479) );
  NAND2_X2 U6623 ( .A1(n9252), .A2(n9989), .ZN(n10128) );
  OAI211_X4 U6624 ( .C1(n10081), .C2(n10080), .A(n10079), .B(n6013), .ZN(
        n10082) );
  INV_X1 U6625 ( .A(n10164), .ZN(n9990) );
  OAI211_X4 U6626 ( .C1(n5923), .C2(n7313), .A(n9248), .B(n9247), .ZN(n10164)
         );
  NAND3_X2 U6627 ( .A1(n7809), .A2(n8412), .A3(n7808), .ZN(n7814) );
  NOR2_X1 U6628 ( .A1(n7618), .A2(n1576), .ZN(IF_ID_REG_IF_ID_REG_N29) );
  INV_X8 U6629 ( .A(n6878), .ZN(n5854) );
  INV_X16 U6630 ( .A(n5854), .ZN(n5855) );
  NOR2_X1 U6631 ( .A1(n7771), .A2(n7452), .ZN(n7357) );
  INV_X4 U6632 ( .A(n7799), .ZN(n7782) );
  AND2_X4 U6633 ( .A1(n4846), .A2(offset_26_id[7]), .ZN(n5858) );
  NAND2_X2 U6634 ( .A1(offset_26_id[2]), .A2(n4089), .ZN(n5859) );
  NAND2_X2 U6635 ( .A1(n4093), .A2(n5857), .ZN(n5860) );
  INV_X4 U6636 ( .A(n5865), .ZN(n7593) );
  NOR2_X1 U6637 ( .A1(n7771), .A2(n7452), .ZN(n7358) );
  INV_X4 U6638 ( .A(n7509), .ZN(n7507) );
  INV_X4 U6639 ( .A(n7493), .ZN(n7491) );
  INV_X4 U6640 ( .A(n7516), .ZN(n7515) );
  INV_X4 U6641 ( .A(n7500), .ZN(n7499) );
  INV_X4 U6642 ( .A(n7590), .ZN(n7584) );
  INV_X4 U6643 ( .A(n7798), .ZN(n7784) );
  INV_X4 U6644 ( .A(n7509), .ZN(n7508) );
  INV_X4 U6645 ( .A(n7493), .ZN(n7492) );
  INV_X4 U6646 ( .A(n5858), .ZN(n7552) );
  INV_X4 U6647 ( .A(n4090), .ZN(n7764) );
  INV_X4 U6648 ( .A(n7535), .ZN(n7534) );
  INV_X4 U6649 ( .A(n4110), .ZN(n7538) );
  INV_X4 U6650 ( .A(n5865), .ZN(n7596) );
  INV_X4 U6651 ( .A(n5865), .ZN(n7592) );
  INV_X4 U6652 ( .A(n7798), .ZN(n7781) );
  NAND2_X4 U6653 ( .A1(n7794), .A2(n9246), .ZN(n5862) );
  NAND2_X4 U6654 ( .A1(n7794), .A2(n9290), .ZN(n5863) );
  AND2_X2 U6655 ( .A1(n9180), .A2(n7383), .ZN(n5864) );
  INV_X4 U6656 ( .A(EXEC_MEM_OUT_141), .ZN(n7774) );
  INV_X4 U6657 ( .A(n6333), .ZN(n7604) );
  INV_X4 U6658 ( .A(n7507), .ZN(n7502) );
  INV_X4 U6659 ( .A(n7507), .ZN(n7503) );
  INV_X4 U6660 ( .A(n7491), .ZN(n7486) );
  INV_X4 U6661 ( .A(n7491), .ZN(n7487) );
  INV_X4 U6662 ( .A(n7590), .ZN(n7588) );
  INV_X4 U6663 ( .A(n7358), .ZN(n7362) );
  NOR2_X1 U6664 ( .A1(n7771), .A2(n7452), .ZN(n8038) );
  AND2_X4 U6665 ( .A1(n4094), .A2(offset_26_id[2]), .ZN(n5865) );
  OR2_X4 U6666 ( .A1(n8108), .A2(n7803), .ZN(n5866) );
  NAND2_X4 U6667 ( .A1(n7796), .A2(n9230), .ZN(n5867) );
  NAND2_X4 U6668 ( .A1(n7795), .A2(n9266), .ZN(n5868) );
  INV_X4 U6669 ( .A(n6844), .ZN(n10229) );
  INV_X4 U6670 ( .A(n6897), .ZN(n7750) );
  INV_X4 U6671 ( .A(n6897), .ZN(n7749) );
  INV_X4 U6672 ( .A(n7771), .ZN(n7772) );
  INV_X4 U6673 ( .A(n5859), .ZN(n7577) );
  INV_X4 U6674 ( .A(n5859), .ZN(n7578) );
  INV_X4 U6675 ( .A(n7797), .ZN(n7776) );
  AND2_X4 U6676 ( .A1(n9864), .A2(n9871), .ZN(n5884) );
  INV_X4 U6677 ( .A(n6904), .ZN(n7754) );
  INV_X4 U6678 ( .A(n6904), .ZN(n7753) );
  INV_X4 U6679 ( .A(n6903), .ZN(n7752) );
  INV_X4 U6680 ( .A(n6903), .ZN(n7751) );
  AND2_X2 U6681 ( .A1(n7795), .A2(n8676), .ZN(n6335) );
  INV_X4 U6682 ( .A(n7526), .ZN(n7521) );
  INV_X4 U6683 ( .A(n7526), .ZN(n7525) );
  INV_X4 U6684 ( .A(n6896), .ZN(n7756) );
  INV_X4 U6685 ( .A(n6896), .ZN(n7755) );
  INV_X4 U6686 ( .A(n6866), .ZN(n7758) );
  INV_X4 U6687 ( .A(n6866), .ZN(n7757) );
  INV_X4 U6688 ( .A(n6993), .ZN(n7423) );
  INV_X4 U6689 ( .A(n6993), .ZN(n7422) );
  INV_X4 U6690 ( .A(n6870), .ZN(n7424) );
  INV_X4 U6691 ( .A(n6870), .ZN(n7425) );
  INV_X4 U6692 ( .A(n6871), .ZN(n7426) );
  INV_X4 U6693 ( .A(n6871), .ZN(n7427) );
  INV_X4 U6694 ( .A(n6876), .ZN(n7443) );
  INV_X4 U6695 ( .A(n6876), .ZN(n7444) );
  INV_X4 U6696 ( .A(n5858), .ZN(n7549) );
  INV_X4 U6697 ( .A(n5858), .ZN(n7547) );
  INV_X4 U6698 ( .A(n7566), .ZN(n7559) );
  INV_X4 U6699 ( .A(n7565), .ZN(n7560) );
  INV_X4 U6700 ( .A(n6333), .ZN(n7602) );
  INV_X4 U6701 ( .A(n6333), .ZN(n7603) );
  INV_X4 U6702 ( .A(n7515), .ZN(n7511) );
  INV_X4 U6703 ( .A(n7499), .ZN(n7497) );
  INV_X4 U6704 ( .A(n5860), .ZN(n7606) );
  INV_X4 U6705 ( .A(n7538), .ZN(n7544) );
  INV_X4 U6706 ( .A(n7535), .ZN(n7529) );
  INV_X4 U6707 ( .A(n7535), .ZN(n7528) );
  INV_X4 U6708 ( .A(n3405), .ZN(n7573) );
  INV_X4 U6709 ( .A(n4090), .ZN(n7765) );
  INV_X4 U6710 ( .A(n7437), .ZN(n7438) );
  INV_X4 U6711 ( .A(n7357), .ZN(n7359) );
  NOR2_X1 U6712 ( .A1(n7771), .A2(n7452), .ZN(n7889) );
  INV_X4 U6713 ( .A(reset), .ZN(n7797) );
  INV_X4 U6714 ( .A(n7801), .ZN(n7780) );
  NAND3_X4 U6715 ( .A1(n7813), .A2(n7774), .A3(n7814), .ZN(n5908) );
  INV_X4 U6716 ( .A(ID_EXEC_OUT[159]), .ZN(n7449) );
  INV_X8 U6717 ( .A(n7389), .ZN(n7478) );
  INV_X4 U6718 ( .A(n6338), .ZN(n7408) );
  INV_X4 U6719 ( .A(n6338), .ZN(n7409) );
  INV_X4 U6720 ( .A(n6339), .ZN(n7411) );
  INV_X4 U6721 ( .A(n6339), .ZN(n7412) );
  AND2_X4 U6722 ( .A1(n7795), .A2(n8423), .ZN(n5910) );
  AND2_X2 U6723 ( .A1(n7795), .A2(n8604), .ZN(n5911) );
  AND3_X4 U6724 ( .A1(RegWrite_wb_out), .A2(n7827), .A3(n6889), .ZN(n5913) );
  INV_X4 U6725 ( .A(n6336), .ZN(n7400) );
  XOR2_X2 U6726 ( .A(n8210), .B(n6801), .Z(n5915) );
  INV_X4 U6727 ( .A(n6880), .ZN(n7759) );
  INV_X4 U6728 ( .A(n6880), .ZN(n7760) );
  INV_X4 U6729 ( .A(n6872), .ZN(n7404) );
  INV_X4 U6730 ( .A(n6872), .ZN(n7403) );
  AND2_X2 U6731 ( .A1(n7794), .A2(n8902), .ZN(n6342) );
  INV_X4 U6732 ( .A(n6342), .ZN(n7428) );
  INV_X4 U6733 ( .A(n6335), .ZN(n7398) );
  INV_X4 U6734 ( .A(n6337), .ZN(n7405) );
  INV_X4 U6735 ( .A(n6340), .ZN(n7414) );
  INV_X4 U6736 ( .A(n6341), .ZN(n7417) );
  INV_X4 U6737 ( .A(n6874), .ZN(n7421) );
  INV_X4 U6738 ( .A(n6874), .ZN(n7420) );
  NOR2_X2 U6739 ( .A1(n6326), .A2(n7803), .ZN(n6003) );
  NOR2_X2 U6740 ( .A1(n6327), .A2(n7803), .ZN(n6004) );
  NOR2_X2 U6741 ( .A1(n6328), .A2(n7803), .ZN(n6005) );
  NOR2_X2 U6742 ( .A1(n6329), .A2(n7803), .ZN(n6006) );
  NOR2_X2 U6743 ( .A1(n6331), .A2(n7803), .ZN(n6007) );
  NOR2_X2 U6744 ( .A1(n6332), .A2(n7803), .ZN(n6008) );
  INV_X4 U6745 ( .A(n6333), .ZN(n7601) );
  INV_X4 U6746 ( .A(n6333), .ZN(n7600) );
  INV_X4 U6747 ( .A(n5865), .ZN(n7598) );
  INV_X4 U6748 ( .A(n7515), .ZN(n7513) );
  INV_X4 U6749 ( .A(n7499), .ZN(n7495) );
  AND2_X4 U6750 ( .A1(n4091), .A2(offset_26_id[2]), .ZN(n6009) );
  INV_X4 U6751 ( .A(n7538), .ZN(n7543) );
  INV_X4 U6752 ( .A(n5860), .ZN(n7609) );
  INV_X4 U6753 ( .A(n7590), .ZN(n7585) );
  INV_X4 U6754 ( .A(n7590), .ZN(n7586) );
  NOR2_X1 U6755 ( .A1(n7771), .A2(n7452), .ZN(n7941) );
  INV_X4 U6756 ( .A(n7438), .ZN(n7439) );
  NAND3_X2 U6757 ( .A1(n5856), .A2(n5861), .A3(offset_26_id[7]), .ZN(n4112) );
  INV_X4 U6758 ( .A(reset), .ZN(n7802) );
  INV_X4 U6759 ( .A(n7798), .ZN(n7779) );
  INV_X4 U6760 ( .A(n7801), .ZN(n7778) );
  INV_X4 U6761 ( .A(n7798), .ZN(n7777) );
  AND2_X2 U6762 ( .A1(n1591), .A2(n7774), .ZN(n6010) );
  INV_X4 U6763 ( .A(n7466), .ZN(n7472) );
  INV_X4 U6764 ( .A(n6336), .ZN(n7402) );
  INV_X4 U6765 ( .A(n6336), .ZN(n7401) );
  AND3_X4 U6766 ( .A1(ID_EXEC_OUT[156]), .A2(n10084), .A3(n6883), .ZN(n6023)
         );
  AND3_X4 U6767 ( .A1(n3092), .A2(n7312), .A3(n6349), .ZN(n6027) );
  AND3_X4 U6768 ( .A1(n7317), .A2(n8111), .A3(n8114), .ZN(n6028) );
  AND3_X4 U6769 ( .A1(n7317), .A2(n3092), .A3(n8114), .ZN(n6029) );
  AND3_X4 U6770 ( .A1(n8111), .A2(n6349), .A3(n8114), .ZN(n6034) );
  INV_X4 U6771 ( .A(n7305), .ZN(n7773) );
  AND3_X4 U6772 ( .A1(n7312), .A2(n8111), .A3(n6349), .ZN(n6035) );
  XOR2_X2 U6773 ( .A(nextPC_ex_out[22]), .B(n8158), .Z(n6036) );
  XOR2_X2 U6774 ( .A(nextPC_ex_out[28]), .B(n8194), .Z(n6037) );
  INV_X4 U6775 ( .A(n6335), .ZN(n7397) );
  INV_X4 U6776 ( .A(n6335), .ZN(n7399) );
  INV_X4 U6777 ( .A(n6342), .ZN(n7429) );
  INV_X4 U6778 ( .A(n6342), .ZN(n7430) );
  INV_X4 U6779 ( .A(n6337), .ZN(n7407) );
  INV_X4 U6780 ( .A(n6337), .ZN(n7406) );
  INV_X4 U6781 ( .A(n6338), .ZN(n7410) );
  INV_X4 U6782 ( .A(n6339), .ZN(n7413) );
  INV_X4 U6783 ( .A(n6340), .ZN(n7415) );
  INV_X4 U6784 ( .A(n6340), .ZN(n7416) );
  INV_X4 U6785 ( .A(n6341), .ZN(n7418) );
  INV_X4 U6786 ( .A(n6341), .ZN(n7419) );
  OAI21_X2 U6787 ( .B1(n7038), .B2(n6023), .A(n10282), .ZN(n10230) );
  INV_X4 U6788 ( .A(n6873), .ZN(n7433) );
  INV_X4 U6789 ( .A(n6873), .ZN(n7434) );
  AND2_X2 U6790 ( .A1(n7794), .A2(n8904), .ZN(n6875) );
  INV_X4 U6791 ( .A(n6875), .ZN(n7431) );
  INV_X4 U6792 ( .A(n6875), .ZN(n7432) );
  AND2_X4 U6793 ( .A1(n3110), .A2(n7796), .ZN(n6044) );
  AND2_X4 U6794 ( .A1(n3107), .A2(n7796), .ZN(n6045) );
  AND2_X4 U6795 ( .A1(n3099), .A2(n7796), .ZN(n6046) );
  INV_X4 U6796 ( .A(n6879), .ZN(n7367) );
  INV_X4 U6797 ( .A(n6879), .ZN(n7368) );
  AND2_X4 U6798 ( .A1(n6027), .A2(n3080), .ZN(n6134) );
  AND2_X4 U6799 ( .A1(n6029), .A2(n3080), .ZN(n6135) );
  AND2_X4 U6800 ( .A1(n6027), .A2(n3077), .ZN(n6136) );
  AND2_X4 U6801 ( .A1(n6029), .A2(n3077), .ZN(n6137) );
  AND2_X4 U6802 ( .A1(n8115), .A2(n3077), .ZN(n6138) );
  AND2_X4 U6803 ( .A1(n7795), .A2(n3131), .ZN(n6139) );
  AND2_X4 U6804 ( .A1(n7795), .A2(n3128), .ZN(n6140) );
  AND2_X4 U6805 ( .A1(n7795), .A2(n3148), .ZN(n6141) );
  AND2_X4 U6806 ( .A1(n7795), .A2(n3146), .ZN(n6142) );
  AND4_X4 U6807 ( .A1(n8512), .A2(n8511), .A3(n8510), .A4(n8509), .ZN(n6185)
         );
  XOR2_X2 U6808 ( .A(n8225), .B(n6699), .Z(n6186) );
  XOR2_X2 U6809 ( .A(n8225), .B(n7220), .Z(n6187) );
  AND4_X4 U6810 ( .A1(n10243), .A2(n10242), .A3(n10241), .A4(n10240), .ZN(
        n6188) );
  XOR2_X2 U6811 ( .A(n8211), .B(n6802), .Z(n6189) );
  XOR2_X2 U6812 ( .A(n8218), .B(n6803), .Z(n6190) );
  AND2_X4 U6813 ( .A1(n3105), .A2(n7796), .ZN(n6191) );
  AND2_X4 U6814 ( .A1(n3103), .A2(n7796), .ZN(n6192) );
  INV_X4 U6815 ( .A(n5910), .ZN(n7377) );
  AND2_X4 U6816 ( .A1(n7795), .A2(n3135), .ZN(n6267) );
  INV_X4 U6817 ( .A(n5911), .ZN(n7394) );
  AND2_X4 U6818 ( .A1(n3114), .A2(n7796), .ZN(n6301) );
  AND2_X4 U6819 ( .A1(n3112), .A2(n7796), .ZN(n6303) );
  AND2_X4 U6820 ( .A1(n7795), .A2(n3133), .ZN(n6304) );
  NAND3_X2 U6821 ( .A1(n5856), .A2(n5861), .A3(n1641), .ZN(n4113) );
  INV_X4 U6822 ( .A(n7526), .ZN(n7523) );
  INV_X4 U6823 ( .A(n7526), .ZN(n7524) );
  AND2_X4 U6824 ( .A1(n7795), .A2(n3078), .ZN(n6305) );
  AND2_X4 U6825 ( .A1(n3096), .A2(n7796), .ZN(n6306) );
  NOR2_X2 U6826 ( .A1(n6134), .A2(n7803), .ZN(n6307) );
  NOR2_X2 U6827 ( .A1(n6136), .A2(n7803), .ZN(n6308) );
  NOR2_X2 U6828 ( .A1(n6135), .A2(n7803), .ZN(n6309) );
  NOR2_X2 U6829 ( .A1(n6137), .A2(n7803), .ZN(n6310) );
  NOR2_X2 U6830 ( .A1(n7731), .A2(n7803), .ZN(n6311) );
  NOR2_X2 U6831 ( .A1(n6138), .A2(n7803), .ZN(n6312) );
  AND2_X4 U6832 ( .A1(n7795), .A2(n3101), .ZN(n6313) );
  AND2_X4 U6833 ( .A1(n7795), .A2(n3093), .ZN(n6314) );
  AND2_X4 U6834 ( .A1(n7796), .A2(n3150), .ZN(n6315) );
  AND2_X4 U6835 ( .A1(n7795), .A2(n3126), .ZN(n6316) );
  AND2_X4 U6836 ( .A1(n9543), .A2(n9542), .ZN(n6317) );
  AND2_X4 U6837 ( .A1(n6027), .A2(n3087), .ZN(n6326) );
  AND2_X4 U6838 ( .A1(n6027), .A2(n3084), .ZN(n6327) );
  AND2_X4 U6839 ( .A1(n6029), .A2(n3087), .ZN(n6328) );
  AND2_X4 U6840 ( .A1(n6029), .A2(n3084), .ZN(n6329) );
  NOR2_X2 U6841 ( .A1(n8118), .A2(n8116), .ZN(n6331) );
  NOR2_X2 U6842 ( .A1(n8118), .A2(n8117), .ZN(n6332) );
  INV_X4 U6843 ( .A(n4090), .ZN(n7768) );
  INV_X4 U6844 ( .A(n4090), .ZN(n7767) );
  INV_X4 U6845 ( .A(n4090), .ZN(n7766) );
  INV_X4 U6846 ( .A(n7538), .ZN(n7540) );
  INV_X4 U6847 ( .A(n4129), .ZN(n7504) );
  INV_X4 U6848 ( .A(n4131), .ZN(n7488) );
  INV_X4 U6849 ( .A(n5860), .ZN(n7607) );
  INV_X4 U6850 ( .A(n5860), .ZN(n7608) );
  NOR2_X2 U6851 ( .A1(n7773), .A2(n6031), .ZN(n7369) );
  NOR2_X2 U6852 ( .A1(n7773), .A2(n6031), .ZN(n8762) );
  INV_X4 U6853 ( .A(n7590), .ZN(n7587) );
  NAND2_X2 U6854 ( .A1(n4093), .A2(offset_26_id[2]), .ZN(n6333) );
  NAND2_X1 U6855 ( .A1(n4845), .A2(offset_26_id[7]), .ZN(n4128) );
  NAND2_X1 U6856 ( .A1(n4847), .A2(offset_26_id[7]), .ZN(n4130) );
  NAND2_X4 U6857 ( .A1(EXEC_STAGE_imm16_32_16_), .A2(n7453), .ZN(n6334) );
  INV_X4 U6858 ( .A(n5859), .ZN(n7580) );
  INV_X4 U6859 ( .A(n5864), .ZN(n7385) );
  INV_X4 U6860 ( .A(n4112), .ZN(n7535) );
  INV_X4 U6861 ( .A(n7535), .ZN(n7530) );
  INV_X4 U6862 ( .A(n7438), .ZN(n7440) );
  INV_X4 U6863 ( .A(n6009), .ZN(n7567) );
  INV_X4 U6864 ( .A(reset), .ZN(n7799) );
  INV_X4 U6865 ( .A(reset), .ZN(n7798) );
  AND2_X2 U6866 ( .A1(n7795), .A2(n8724), .ZN(n6336) );
  AND2_X4 U6867 ( .A1(n7795), .A2(n9086), .ZN(n6337) );
  AND2_X4 U6868 ( .A1(n7795), .A2(n9079), .ZN(n6338) );
  AND2_X4 U6869 ( .A1(n7795), .A2(n8886), .ZN(n6339) );
  AND2_X4 U6870 ( .A1(n7795), .A2(n8888), .ZN(n6340) );
  AND2_X4 U6871 ( .A1(n7795), .A2(n8891), .ZN(n6341) );
  AND2_X4 U6872 ( .A1(n9980), .A2(n9979), .ZN(n6344) );
  INV_X4 U6873 ( .A(n9361), .ZN(n7474) );
  INV_X4 U6874 ( .A(n9195), .ZN(n9361) );
  INV_X16 U6875 ( .A(n7474), .ZN(n7473) );
  AND2_X4 U6876 ( .A1(n9196), .A2(n9704), .ZN(n6350) );
  INV_X4 U6877 ( .A(n7613), .ZN(n7612) );
  AND3_X4 U6878 ( .A1(n4269), .A2(n8087), .A3(n8086), .ZN(n6354) );
  AND3_X4 U6879 ( .A1(n4247), .A2(n8089), .A3(n8088), .ZN(n6355) );
  AND2_X4 U6880 ( .A1(n8301), .A2(n8373), .ZN(n6356) );
  XOR2_X2 U6881 ( .A(n8214), .B(n7222), .Z(n6357) );
  AND2_X4 U6882 ( .A1(n9338), .A2(n9919), .ZN(n6450) );
  XNOR2_X1 U6883 ( .A(offset_26_id[8]), .B(n7310), .ZN(n6467) );
  AND3_X4 U6884 ( .A1(n8417), .A2(n8416), .A3(n8415), .ZN(n6478) );
  INV_X1 U6885 ( .A(n9855), .ZN(n7352) );
  AND2_X4 U6886 ( .A1(n4823), .A2(offset_26_id[5]), .ZN(n6480) );
  AND4_X4 U6887 ( .A1(n9111), .A2(n9110), .A3(n9109), .A4(n9108), .ZN(n6482)
         );
  XOR2_X2 U6888 ( .A(nextPC_ex_out[21]), .B(n8159), .Z(n6520) );
  XOR2_X2 U6889 ( .A(nextPC_ex_out[27]), .B(n8195), .Z(n6521) );
  NOR2_X2 U6890 ( .A1(n8940), .A2(n7803), .ZN(n8941) );
  AND2_X4 U6891 ( .A1(n7794), .A2(n8948), .ZN(n6700) );
  AND2_X4 U6892 ( .A1(n4823), .A2(n6014), .ZN(n6791) );
  NAND2_X2 U6893 ( .A1(n4077), .A2(offset_26_id[1]), .ZN(n6792) );
  NAND2_X2 U6894 ( .A1(n4077), .A2(n6016), .ZN(n6793) );
  NAND2_X2 U6895 ( .A1(ID_EX_REG_ID_EX_REG_N93), .A2(n4069), .ZN(n6794) );
  AND2_X4 U6896 ( .A1(n4832), .A2(n6014), .ZN(n6795) );
  AND2_X4 U6897 ( .A1(n7795), .A2(n7759), .ZN(n6796) );
  AND2_X4 U6898 ( .A1(n7815), .A2(n7305), .ZN(n6797) );
  AND2_X4 U6899 ( .A1(n9482), .A2(n9448), .ZN(n6798) );
  AND2_X4 U6900 ( .A1(n9786), .A2(ID_EXEC_OUT[158]), .ZN(n6799) );
  AND2_X4 U6901 ( .A1(n9862), .A2(ID_EXEC_OUT[158]), .ZN(n6800) );
  AND4_X4 U6902 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n6804) );
  AND2_X4 U6903 ( .A1(n8528), .A2(n8527), .ZN(n6805) );
  AND2_X4 U6904 ( .A1(n9536), .A2(n9535), .ZN(n6806) );
  INV_X4 U6905 ( .A(n3168), .ZN(n7623) );
  INV_X4 U6906 ( .A(n7623), .ZN(n7621) );
  AND4_X4 U6907 ( .A1(n9344), .A2(n9343), .A3(n9342), .A4(n9341), .ZN(n6807)
         );
  INV_X4 U6908 ( .A(n7615), .ZN(n7614) );
  INV_X4 U6909 ( .A(n3232), .ZN(n7615) );
  INV_X8 U6910 ( .A(n7614), .ZN(n7618) );
  AND4_X4 U6911 ( .A1(n9795), .A2(n9794), .A3(n9793), .A4(n9792), .ZN(n6828)
         );
  INV_X4 U6912 ( .A(n8024), .ZN(n7834) );
  NOR2_X2 U6913 ( .A1(ID_EXEC_OUT[153]), .A2(EXEC_MEM_OUT_141), .ZN(n10282) );
  INV_X8 U6914 ( .A(n7239), .ZN(n7771) );
  OR4_X4 U6915 ( .A1(n4285), .A2(n4286), .A3(n4287), .A4(n4288), .ZN(n6829) );
  OR4_X4 U6916 ( .A1(n4557), .A2(n4558), .A3(n4559), .A4(n4560), .ZN(n6830) );
  OR4_X4 U6917 ( .A1(n4692), .A2(n4693), .A3(n4694), .A4(n4695), .ZN(n6831) );
  OR4_X4 U6918 ( .A1(n4263), .A2(n4264), .A3(n4265), .A4(n4266), .ZN(n6832) );
  INV_X4 U6919 ( .A(n4113), .ZN(n7526) );
  INV_X4 U6920 ( .A(n6306), .ZN(n7720) );
  INV_X4 U6921 ( .A(n6306), .ZN(n7721) );
  NAND3_X2 U6922 ( .A1(n8085), .A2(n6467), .A3(n8084), .ZN(n4100) );
  NOR2_X2 U6923 ( .A1(n7773), .A2(n6481), .ZN(n6844) );
  INV_X4 U6924 ( .A(n5865), .ZN(n7597) );
  INV_X4 U6925 ( .A(n5865), .ZN(n7594) );
  INV_X4 U6926 ( .A(n5865), .ZN(n7595) );
  INV_X4 U6927 ( .A(n7567), .ZN(n7566) );
  INV_X4 U6928 ( .A(n7566), .ZN(n7561) );
  INV_X4 U6929 ( .A(n7566), .ZN(n7562) );
  INV_X4 U6930 ( .A(n3405), .ZN(n7572) );
  INV_X4 U6931 ( .A(n7572), .ZN(n7568) );
  INV_X4 U6932 ( .A(n7572), .ZN(n7569) );
  INV_X4 U6933 ( .A(n5859), .ZN(n7581) );
  INV_X4 U6934 ( .A(n5859), .ZN(n7582) );
  INV_X4 U6935 ( .A(n5859), .ZN(n7579) );
  INV_X4 U6936 ( .A(n5858), .ZN(n7550) );
  INV_X4 U6937 ( .A(n5858), .ZN(n7551) );
  INV_X4 U6938 ( .A(n5858), .ZN(n7548) );
  INV_X4 U6939 ( .A(n9806), .ZN(n7387) );
  INV_X4 U6940 ( .A(n7387), .ZN(n7388) );
  INV_X4 U6941 ( .A(n7535), .ZN(n7532) );
  INV_X4 U6942 ( .A(n7535), .ZN(n7531) );
  NAND2_X2 U6943 ( .A1(n9786), .A2(n6013), .ZN(n6860) );
  NAND2_X2 U6944 ( .A1(n10272), .A2(n10282), .ZN(n6861) );
  NOR2_X1 U6945 ( .A1(n7771), .A2(n7452), .ZN(n7855) );
  INV_X4 U6946 ( .A(n7449), .ZN(n7450) );
  INV_X4 U6947 ( .A(n7371), .ZN(n7373) );
  INV_X4 U6948 ( .A(n7371), .ZN(n7372) );
  INV_X4 U6949 ( .A(n5864), .ZN(n7386) );
  INV_X4 U6950 ( .A(n4128), .ZN(n7510) );
  INV_X4 U6951 ( .A(n7515), .ZN(n7512) );
  INV_X4 U6952 ( .A(n4130), .ZN(n7494) );
  INV_X4 U6953 ( .A(n7499), .ZN(n7496) );
  INV_X4 U6954 ( .A(n4129), .ZN(n7501) );
  INV_X4 U6955 ( .A(n4131), .ZN(n7485) );
  INV_X4 U6956 ( .A(n7438), .ZN(n7441) );
  INV_X4 U6957 ( .A(n4090), .ZN(n7769) );
  INV_X4 U6958 ( .A(n4090), .ZN(n7770) );
  INV_X4 U6959 ( .A(n7538), .ZN(n7536) );
  INV_X4 U6960 ( .A(n7538), .ZN(n7541) );
  INV_X4 U6961 ( .A(n7538), .ZN(n7542) );
  INV_X4 U6962 ( .A(n5884), .ZN(n7389) );
  INV_X4 U6963 ( .A(n3399), .ZN(n7590) );
  INV_X4 U6964 ( .A(n7590), .ZN(n7589) );
  INV_X4 U6965 ( .A(n6134), .ZN(n7638) );
  INV_X4 U6966 ( .A(n6135), .ZN(n7674) );
  INV_X4 U6967 ( .A(n3090), .ZN(n7731) );
  INV_X4 U6968 ( .A(n6136), .ZN(n7642) );
  INV_X4 U6969 ( .A(n6137), .ZN(n7678) );
  INV_X4 U6970 ( .A(n6138), .ZN(n7735) );
  INV_X4 U6971 ( .A(n6326), .ZN(n7646) );
  INV_X4 U6972 ( .A(n6327), .ZN(n7650) );
  INV_X4 U6973 ( .A(n6328), .ZN(n7682) );
  INV_X4 U6974 ( .A(n6329), .ZN(n7686) );
  INV_X4 U6975 ( .A(n6331), .ZN(n7739) );
  INV_X4 U6976 ( .A(n6332), .ZN(n7743) );
  INV_X4 U6977 ( .A(reset), .ZN(n7801) );
  INV_X8 U6978 ( .A(n9632), .ZN(n9877) );
  AND2_X4 U6979 ( .A1(n7795), .A2(n9260), .ZN(n6866) );
  OR3_X4 U6980 ( .A1(n7812), .A2(n7811), .A3(n7810), .ZN(n6869) );
  AND2_X4 U6981 ( .A1(n7794), .A2(n9275), .ZN(n6870) );
  AND2_X4 U6982 ( .A1(n7794), .A2(n9280), .ZN(n6871) );
  AND2_X4 U6983 ( .A1(n7794), .A2(n9101), .ZN(n6872) );
  AND2_X4 U6984 ( .A1(n7794), .A2(n8907), .ZN(n6873) );
  AND2_X4 U6985 ( .A1(n7795), .A2(n8894), .ZN(n6874) );
  AND2_X4 U6986 ( .A1(n7794), .A2(n7316), .ZN(n6876) );
  AND2_X4 U6987 ( .A1(n7384), .A2(n5853), .ZN(n6878) );
  OR2_X4 U6988 ( .A1(n7447), .A2(n8105), .ZN(n6879) );
  AND2_X4 U6989 ( .A1(n3077), .A2(n6035), .ZN(n6880) );
  INV_X16 U6990 ( .A(n7390), .ZN(n7391) );
  INV_X8 U6991 ( .A(n9802), .ZN(n7390) );
  INV_X4 U6992 ( .A(n10155), .ZN(n10257) );
  INV_X4 U6993 ( .A(n9995), .ZN(n10271) );
  AND2_X4 U6994 ( .A1(n8569), .A2(n8568), .ZN(n6892) );
  AND2_X4 U6995 ( .A1(n8592), .A2(n8591), .ZN(n6893) );
  XOR2_X2 U6996 ( .A(n8482), .B(n9632), .Z(n6895) );
  AND2_X4 U6997 ( .A1(n7796), .A2(n9234), .ZN(n6896) );
  AND2_X4 U6998 ( .A1(n7795), .A2(n9169), .ZN(n6897) );
  NOR2_X2 U6999 ( .A1(n8107), .A2(n7803), .ZN(n6903) );
  NOR2_X2 U7000 ( .A1(n8110), .A2(n7804), .ZN(n6904) );
  AND2_X4 U7001 ( .A1(n7476), .A2(n10135), .ZN(n6911) );
  AND2_X4 U7002 ( .A1(n6893), .A2(n8585), .ZN(n6912) );
  AND2_X4 U7003 ( .A1(n9455), .A2(n9456), .ZN(n6916) );
  AND4_X4 U7004 ( .A1(n10142), .A2(n10141), .A3(n10140), .A4(n10139), .ZN(
        n6917) );
  XOR2_X2 U7005 ( .A(nextPC_ex_out[20]), .B(n8163), .Z(n6918) );
  OR2_X4 U7006 ( .A1(ID_EXEC_OUT[156]), .A2(n10097), .ZN(n6988) );
  XOR2_X2 U7007 ( .A(n9265), .B(n9977), .Z(n6989) );
  XOR2_X2 U7008 ( .A(n9078), .B(n9916), .Z(n6990) );
  AND2_X4 U7009 ( .A1(n7795), .A2(n9269), .ZN(n6993) );
  AND2_X4 U7010 ( .A1(n8967), .A2(n9864), .ZN(n6994) );
  INV_X4 U7011 ( .A(n9871), .ZN(n9180) );
  AND2_X4 U7012 ( .A1(n8710), .A2(n8756), .ZN(n6998) );
  AND2_X4 U7013 ( .A1(n8567), .A2(n8566), .ZN(n6999) );
  XNOR2_X2 U7014 ( .A(n6014), .B(n7317), .ZN(n7000) );
  AND2_X4 U7015 ( .A1(n8967), .A2(n7383), .ZN(n7001) );
  AND3_X4 U7016 ( .A1(n9638), .A2(n9637), .A3(n9636), .ZN(n7035) );
  XOR2_X2 U7017 ( .A(nextPC_ex_out[19]), .B(n8166), .Z(n7036) );
  XOR2_X2 U7018 ( .A(nextPC_ex_out[25]), .B(n8174), .Z(n7037) );
  AND2_X4 U7019 ( .A1(ID_EXEC_OUT[157]), .A2(n9197), .ZN(n7038) );
  AND4_X4 U7020 ( .A1(n9603), .A2(n9602), .A3(n9601), .A4(n9600), .ZN(n7138)
         );
  NAND4_X2 U7021 ( .A1(n4447), .A2(ID_STAGE_imm16_aluA[16]), .A3(n4448), .A4(
        n7774), .ZN(n4096) );
  AND4_X4 U7022 ( .A1(n10152), .A2(n10151), .A3(n10150), .A4(n10149), .ZN(
        n7139) );
  AND4_X4 U7023 ( .A1(n9702), .A2(n9701), .A3(n9700), .A4(n9699), .ZN(n7208)
         );
  AND2_X4 U7024 ( .A1(n8677), .A2(n8679), .ZN(n7209) );
  AND2_X4 U7025 ( .A1(MEM_WB_OUT[106]), .A2(n8072), .ZN(n7210) );
  INV_X4 U7026 ( .A(n5910), .ZN(n7376) );
  INV_X4 U7027 ( .A(n5910), .ZN(n7375) );
  INV_X4 U7028 ( .A(n5911), .ZN(n7395) );
  INV_X4 U7029 ( .A(n5911), .ZN(n7396) );
  XNOR2_X2 U7030 ( .A(offset_26_id[4]), .B(n7335), .ZN(n7213) );
  OR2_X4 U7031 ( .A1(n9414), .A2(n7383), .ZN(n7214) );
  AND3_X4 U7032 ( .A1(n9674), .A2(n9673), .A3(n9672), .ZN(n7224) );
  AND4_X4 U7033 ( .A1(n9595), .A2(n9594), .A3(n9593), .A4(n9592), .ZN(n7225)
         );
  AND2_X4 U7034 ( .A1(n8959), .A2(n8489), .ZN(n7226) );
  XNOR2_X2 U7035 ( .A(offset_26_id[9]), .B(n7335), .ZN(n7228) );
  AND2_X4 U7036 ( .A1(n8310), .A2(n8307), .ZN(n7229) );
  AND2_X4 U7037 ( .A1(n8540), .A2(n8539), .ZN(n7230) );
  AND4_X4 U7038 ( .A1(n8981), .A2(n8980), .A3(n8979), .A4(n8978), .ZN(n7231)
         );
  AND4_X4 U7039 ( .A1(n10254), .A2(n10253), .A3(n10252), .A4(n10251), .ZN(
        n7232) );
  AND4_X4 U7040 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n7233) );
  AND3_X4 U7041 ( .A1(n8585), .A2(n8590), .A3(n6893), .ZN(n7234) );
  AND2_X4 U7042 ( .A1(n7368), .A2(n9246), .ZN(n7235) );
  AND2_X4 U7043 ( .A1(n9484), .A2(n9485), .ZN(n7236) );
  AND2_X4 U7044 ( .A1(n7368), .A2(n9280), .ZN(n7237) );
  AND2_X4 U7045 ( .A1(n7368), .A2(n9275), .ZN(n7238) );
  NAND3_X2 U7046 ( .A1(n9082), .A2(n9081), .A3(n9080), .ZN(n9918) );
  NAND3_X2 U7047 ( .A1(n9089), .A2(n9088), .A3(n9087), .ZN(n9929) );
  INV_X4 U7048 ( .A(n6480), .ZN(n7520) );
  INV_X4 U7049 ( .A(n6480), .ZN(n7519) );
  INV_X4 U7050 ( .A(n6795), .ZN(n7518) );
  INV_X4 U7051 ( .A(n6795), .ZN(n7517) );
  INV_X4 U7052 ( .A(n6791), .ZN(n7554) );
  INV_X4 U7053 ( .A(n6791), .ZN(n7553) );
  INV_X4 U7054 ( .A(n6797), .ZN(n7484) );
  INV_X4 U7055 ( .A(n6797), .ZN(n7483) );
  OR3_X4 U7056 ( .A1(n4225), .A2(n4226), .A3(n4227), .ZN(n7240) );
  OR3_X4 U7057 ( .A1(n4203), .A2(n4204), .A3(n4205), .ZN(n7241) );
  OR3_X4 U7058 ( .A1(n4180), .A2(n4181), .A3(n4182), .ZN(n7242) );
  OR3_X4 U7059 ( .A1(n4158), .A2(n4159), .A3(n4160), .ZN(n7243) );
  OR3_X4 U7060 ( .A1(n4135), .A2(n4136), .A3(n4137), .ZN(n7244) );
  OR3_X4 U7061 ( .A1(n4102), .A2(n4103), .A3(n4104), .ZN(n7245) );
  AND2_X4 U7062 ( .A1(n8344), .A2(n8302), .ZN(n7246) );
  INV_X4 U7063 ( .A(n3114), .ZN(n7691) );
  INV_X4 U7064 ( .A(n7691), .ZN(n7690) );
  INV_X4 U7065 ( .A(n3112), .ZN(n7695) );
  INV_X4 U7066 ( .A(n7695), .ZN(n7694) );
  INV_X4 U7067 ( .A(n3105), .ZN(n7707) );
  INV_X4 U7068 ( .A(n7707), .ZN(n7706) );
  INV_X4 U7069 ( .A(n3103), .ZN(n7711) );
  INV_X4 U7070 ( .A(n7711), .ZN(n7710) );
  INV_X4 U7071 ( .A(n3150), .ZN(n7627) );
  INV_X4 U7072 ( .A(n7627), .ZN(n7626) );
  INV_X4 U7073 ( .A(n3135), .ZN(n7655) );
  INV_X4 U7074 ( .A(n7655), .ZN(n7654) );
  INV_X4 U7075 ( .A(n3133), .ZN(n7659) );
  INV_X4 U7076 ( .A(n7659), .ZN(n7658) );
  INV_X4 U7077 ( .A(n3126), .ZN(n7671) );
  INV_X4 U7078 ( .A(n7671), .ZN(n7670) );
  INV_X4 U7079 ( .A(n3131), .ZN(n7663) );
  INV_X4 U7080 ( .A(n7663), .ZN(n7662) );
  INV_X4 U7081 ( .A(n3128), .ZN(n7667) );
  INV_X4 U7082 ( .A(n7667), .ZN(n7666) );
  INV_X4 U7083 ( .A(n3110), .ZN(n7699) );
  INV_X4 U7084 ( .A(n7699), .ZN(n7698) );
  INV_X4 U7085 ( .A(n3107), .ZN(n7703) );
  INV_X4 U7086 ( .A(n7703), .ZN(n7702) );
  INV_X4 U7087 ( .A(n3101), .ZN(n7715) );
  INV_X4 U7088 ( .A(n7715), .ZN(n7714) );
  INV_X4 U7089 ( .A(n3099), .ZN(n7719) );
  INV_X4 U7090 ( .A(n7719), .ZN(n7718) );
  INV_X4 U7091 ( .A(n3093), .ZN(n7728) );
  INV_X4 U7092 ( .A(n7728), .ZN(n7727) );
  INV_X4 U7093 ( .A(n3148), .ZN(n7631) );
  INV_X4 U7094 ( .A(n7631), .ZN(n7630) );
  INV_X4 U7095 ( .A(n3146), .ZN(n7635) );
  INV_X4 U7096 ( .A(n7635), .ZN(n7634) );
  INV_X4 U7097 ( .A(n3078), .ZN(n7748) );
  INV_X4 U7098 ( .A(n7748), .ZN(n7747) );
  INV_X4 U7099 ( .A(n6792), .ZN(n7557) );
  INV_X4 U7100 ( .A(n6792), .ZN(n7558) );
  INV_X4 U7101 ( .A(n6793), .ZN(n7555) );
  INV_X4 U7102 ( .A(n6793), .ZN(n7556) );
  INV_X4 U7103 ( .A(n6794), .ZN(n7574) );
  INV_X4 U7104 ( .A(n6794), .ZN(n7575) );
  INV_X4 U7105 ( .A(n3096), .ZN(n7724) );
  INV_X4 U7106 ( .A(n7724), .ZN(n7722) );
  INV_X4 U7107 ( .A(n7724), .ZN(n7723) );
  OR4_X4 U7108 ( .A1(n4715), .A2(n4716), .A3(n4717), .A4(n4718), .ZN(n7247) );
  OR4_X4 U7109 ( .A1(n4738), .A2(n4739), .A3(n4740), .A4(n4741), .ZN(n7248) );
  OR4_X4 U7110 ( .A1(n4669), .A2(n4670), .A3(n4671), .A4(n4672), .ZN(n7249) );
  OR4_X4 U7111 ( .A1(n4601), .A2(n4602), .A3(n4603), .A4(n4604), .ZN(n7250) );
  OR4_X4 U7112 ( .A1(n4579), .A2(n4580), .A3(n4581), .A4(n4582), .ZN(n7251) );
  OR4_X4 U7113 ( .A1(n4512), .A2(n4513), .A3(n4514), .A4(n4515), .ZN(n7252) );
  OR4_X4 U7114 ( .A1(n4490), .A2(n4491), .A3(n4492), .A4(n4493), .ZN(n7253) );
  OR4_X4 U7115 ( .A1(n4804), .A2(n4805), .A3(n4806), .A4(n4807), .ZN(n7254) );
  OR4_X4 U7116 ( .A1(n4760), .A2(n4761), .A3(n4762), .A4(n4763), .ZN(n7255) );
  OR4_X4 U7117 ( .A1(n4782), .A2(n4783), .A3(n4784), .A4(n4785), .ZN(n7256) );
  OR4_X4 U7118 ( .A1(n4647), .A2(n4648), .A3(n4649), .A4(n4650), .ZN(n7257) );
  OR4_X4 U7119 ( .A1(n4624), .A2(n4625), .A3(n4626), .A4(n4627), .ZN(n7258) );
  OR4_X4 U7120 ( .A1(n4535), .A2(n4536), .A3(n4537), .A4(n4538), .ZN(n7259) );
  OR4_X4 U7121 ( .A1(n4468), .A2(n4469), .A3(n4470), .A4(n4471), .ZN(n7260) );
  OR4_X4 U7122 ( .A1(n4443), .A2(n4444), .A3(n4445), .A4(n4446), .ZN(n7261) );
  OR4_X4 U7123 ( .A1(n4420), .A2(n4421), .A3(n4422), .A4(n4423), .ZN(n7262) );
  OR4_X4 U7124 ( .A1(n4398), .A2(n4399), .A3(n4400), .A4(n4401), .ZN(n7263) );
  OR4_X4 U7125 ( .A1(n4375), .A2(n4376), .A3(n4377), .A4(n4378), .ZN(n7264) );
  OR4_X4 U7126 ( .A1(n4353), .A2(n4354), .A3(n4355), .A4(n4356), .ZN(n7265) );
  OR4_X4 U7127 ( .A1(n4330), .A2(n4331), .A3(n4332), .A4(n4333), .ZN(n7266) );
  OR4_X4 U7128 ( .A1(n4308), .A2(n4309), .A3(n4310), .A4(n4311), .ZN(n7267) );
  OR4_X4 U7129 ( .A1(n4841), .A2(n4842), .A3(n4843), .A4(n4844), .ZN(n7268) );
  INV_X16 U7130 ( .A(n7467), .ZN(n7384) );
  INV_X4 U7131 ( .A(n3747), .ZN(n7446) );
  NOR2_X2 U7132 ( .A1(n3351), .A2(n6864), .ZN(n3747) );
  INV_X4 U7133 ( .A(n7446), .ZN(n7447) );
  INV_X4 U7134 ( .A(n7446), .ZN(n7448) );
  INV_X4 U7135 ( .A(n6311), .ZN(n7730) );
  INV_X4 U7136 ( .A(n6311), .ZN(n7729) );
  INV_X4 U7137 ( .A(n6312), .ZN(n7734) );
  INV_X4 U7138 ( .A(n6312), .ZN(n7733) );
  INV_X4 U7139 ( .A(n6007), .ZN(n7738) );
  INV_X4 U7140 ( .A(n6007), .ZN(n7737) );
  INV_X4 U7141 ( .A(n6008), .ZN(n7742) );
  INV_X4 U7142 ( .A(n6008), .ZN(n7741) );
  INV_X4 U7143 ( .A(n6307), .ZN(n7637) );
  INV_X4 U7144 ( .A(n6307), .ZN(n7636) );
  INV_X4 U7145 ( .A(n6308), .ZN(n7641) );
  INV_X4 U7146 ( .A(n6308), .ZN(n7640) );
  INV_X4 U7147 ( .A(n6003), .ZN(n7645) );
  INV_X4 U7148 ( .A(n6003), .ZN(n7644) );
  INV_X4 U7149 ( .A(n6004), .ZN(n7649) );
  INV_X4 U7150 ( .A(n6004), .ZN(n7648) );
  INV_X4 U7151 ( .A(n6309), .ZN(n7673) );
  INV_X4 U7152 ( .A(n6309), .ZN(n7672) );
  INV_X4 U7153 ( .A(n6310), .ZN(n7677) );
  INV_X4 U7154 ( .A(n6310), .ZN(n7676) );
  INV_X4 U7155 ( .A(n6005), .ZN(n7681) );
  INV_X4 U7156 ( .A(n6005), .ZN(n7680) );
  INV_X4 U7157 ( .A(n6006), .ZN(n7685) );
  INV_X4 U7158 ( .A(n6006), .ZN(n7684) );
  AND2_X4 U7159 ( .A1(n7367), .A2(n7316), .ZN(n7269) );
  INV_X4 U7160 ( .A(n6796), .ZN(n7761) );
  INV_X4 U7161 ( .A(n6796), .ZN(n7762) );
  INV_X4 U7162 ( .A(n6141), .ZN(n7629) );
  INV_X4 U7163 ( .A(n6141), .ZN(n7628) );
  INV_X4 U7164 ( .A(n6142), .ZN(n7633) );
  INV_X4 U7165 ( .A(n6142), .ZN(n7632) );
  INV_X4 U7166 ( .A(n6139), .ZN(n7661) );
  INV_X4 U7167 ( .A(n6139), .ZN(n7660) );
  INV_X4 U7168 ( .A(n6140), .ZN(n7665) );
  INV_X4 U7169 ( .A(n6140), .ZN(n7664) );
  INV_X4 U7170 ( .A(n6301), .ZN(n7688) );
  INV_X4 U7171 ( .A(n6301), .ZN(n7689) );
  INV_X4 U7172 ( .A(n6303), .ZN(n7692) );
  INV_X4 U7173 ( .A(n6303), .ZN(n7693) );
  INV_X4 U7174 ( .A(n6044), .ZN(n7697) );
  INV_X4 U7175 ( .A(n6044), .ZN(n7696) );
  INV_X4 U7176 ( .A(n6045), .ZN(n7701) );
  INV_X4 U7177 ( .A(n6045), .ZN(n7700) );
  INV_X4 U7178 ( .A(n6191), .ZN(n7704) );
  INV_X4 U7179 ( .A(n6191), .ZN(n7705) );
  INV_X4 U7180 ( .A(n6192), .ZN(n7708) );
  INV_X4 U7181 ( .A(n6192), .ZN(n7709) );
  INV_X4 U7182 ( .A(n6313), .ZN(n7712) );
  INV_X4 U7183 ( .A(n6313), .ZN(n7713) );
  INV_X4 U7184 ( .A(n6046), .ZN(n7717) );
  INV_X4 U7185 ( .A(n6046), .ZN(n7716) );
  INV_X4 U7186 ( .A(n6314), .ZN(n7725) );
  INV_X4 U7187 ( .A(n6314), .ZN(n7726) );
  INV_X4 U7188 ( .A(n6305), .ZN(n7745) );
  INV_X4 U7189 ( .A(n6305), .ZN(n7746) );
  INV_X4 U7190 ( .A(n6700), .ZN(n7481) );
  INV_X4 U7191 ( .A(n6700), .ZN(n7482) );
  INV_X4 U7192 ( .A(n6315), .ZN(n7625) );
  INV_X4 U7193 ( .A(n6315), .ZN(n7624) );
  INV_X4 U7194 ( .A(n6267), .ZN(n7653) );
  INV_X4 U7195 ( .A(n6267), .ZN(n7652) );
  INV_X4 U7196 ( .A(n6304), .ZN(n7657) );
  INV_X4 U7197 ( .A(n6304), .ZN(n7656) );
  INV_X4 U7198 ( .A(n6316), .ZN(n7669) );
  INV_X4 U7199 ( .A(n6316), .ZN(n7668) );
  OR2_X4 U7200 ( .A1(n6895), .A2(n9763), .ZN(n7281) );
  AND2_X4 U7201 ( .A1(n7367), .A2(n9269), .ZN(n7284) );
  AND2_X4 U7202 ( .A1(n7368), .A2(n9290), .ZN(n7285) );
  INV_X4 U7203 ( .A(n4100), .ZN(n7457) );
  INV_X4 U7204 ( .A(n3169), .ZN(n7620) );
  INV_X4 U7205 ( .A(n7620), .ZN(n7619) );
  INV_X8 U7206 ( .A(n7365), .ZN(n7366) );
  INV_X4 U7207 ( .A(n9835), .ZN(n7365) );
  AND2_X4 U7208 ( .A1(n7368), .A2(n8939), .ZN(n7286) );
  AND2_X4 U7209 ( .A1(n7367), .A2(n8913), .ZN(n7287) );
  AND3_X4 U7210 ( .A1(n9403), .A2(n9316), .A3(n9452), .ZN(n7288) );
  INV_X4 U7211 ( .A(n3390), .ZN(n7613) );
  INV_X4 U7212 ( .A(n4129), .ZN(n7509) );
  INV_X4 U7213 ( .A(n4129), .ZN(n7506) );
  INV_X4 U7214 ( .A(n7508), .ZN(n7505) );
  INV_X4 U7215 ( .A(n4131), .ZN(n7493) );
  INV_X4 U7216 ( .A(n4131), .ZN(n7490) );
  INV_X4 U7217 ( .A(n7492), .ZN(n7489) );
  INV_X4 U7218 ( .A(n8759), .ZN(n7374) );
  NOR2_X2 U7219 ( .A1(EXEC_MEM_IN[102]), .A2(EXEC_MEM_OUT_141), .ZN(n8759) );
  INV_X4 U7220 ( .A(n7567), .ZN(n7565) );
  INV_X4 U7221 ( .A(n7565), .ZN(n7564) );
  INV_X4 U7222 ( .A(n7565), .ZN(n7563) );
  INV_X4 U7223 ( .A(n7590), .ZN(n7583) );
  INV_X4 U7224 ( .A(n6333), .ZN(n7599) );
  INV_X4 U7225 ( .A(n6333), .ZN(n7605) );
  INV_X4 U7226 ( .A(n4090), .ZN(n7763) );
  AND2_X4 U7227 ( .A1(ID_EXEC_OUT[80]), .A2(n8493), .ZN(n7306) );
  INV_X4 U7228 ( .A(n7538), .ZN(n7539) );
  INV_X4 U7229 ( .A(n7538), .ZN(n7537) );
  INV_X4 U7230 ( .A(n8941), .ZN(n7456) );
  INV_X4 U7231 ( .A(n8941), .ZN(n7455) );
  INV_X4 U7232 ( .A(n8941), .ZN(n7454) );
  INV_X4 U7233 ( .A(n10286), .ZN(n7480) );
  INV_X4 U7234 ( .A(n7480), .ZN(n7479) );
  NAND3_X2 U7235 ( .A1(n7379), .A2(n6013), .A3(n8505), .ZN(n10286) );
  INV_X4 U7236 ( .A(n6010), .ZN(n7445) );
  INV_X4 U7237 ( .A(n6134), .ZN(n7639) );
  INV_X4 U7238 ( .A(n6136), .ZN(n7643) );
  INV_X4 U7239 ( .A(n6135), .ZN(n7675) );
  INV_X4 U7240 ( .A(n6137), .ZN(n7679) );
  INV_X4 U7241 ( .A(n7731), .ZN(n7732) );
  INV_X4 U7242 ( .A(n6138), .ZN(n7736) );
  INV_X4 U7243 ( .A(n6326), .ZN(n7647) );
  INV_X4 U7244 ( .A(n6327), .ZN(n7651) );
  INV_X4 U7245 ( .A(n6328), .ZN(n7683) );
  INV_X4 U7246 ( .A(n6329), .ZN(n7687) );
  INV_X4 U7247 ( .A(n6331), .ZN(n7740) );
  INV_X4 U7248 ( .A(n6332), .ZN(n7744) );
  INV_X4 U7249 ( .A(n7572), .ZN(n7570) );
  INV_X4 U7250 ( .A(n7572), .ZN(n7571) );
  INV_X4 U7251 ( .A(n4128), .ZN(n7516) );
  INV_X4 U7252 ( .A(n7515), .ZN(n7514) );
  INV_X4 U7253 ( .A(n4130), .ZN(n7500) );
  INV_X4 U7254 ( .A(n7499), .ZN(n7498) );
  INV_X4 U7255 ( .A(n5860), .ZN(n7610) );
  INV_X4 U7256 ( .A(n5860), .ZN(n7611) );
  INV_X4 U7257 ( .A(n7438), .ZN(n7442) );
  INV_X4 U7258 ( .A(n7371), .ZN(n7370) );
  INV_X4 U7259 ( .A(n8762), .ZN(n7371) );
  INV_X4 U7260 ( .A(n5859), .ZN(n7576) );
  INV_X4 U7261 ( .A(n5858), .ZN(n7545) );
  INV_X4 U7262 ( .A(n5858), .ZN(n7546) );
  INV_X4 U7263 ( .A(n6799), .ZN(n7392) );
  INV_X4 U7264 ( .A(n7535), .ZN(n7527) );
  INV_X4 U7265 ( .A(n7535), .ZN(n7533) );
  INV_X4 U7266 ( .A(n6800), .ZN(n7393) );
  INV_X4 U7267 ( .A(n4099), .ZN(n7458) );
  INV_X4 U7268 ( .A(n4099), .ZN(n7459) );
  INV_X4 U7269 ( .A(n6860), .ZN(n9618) );
  INV_X4 U7270 ( .A(n7378), .ZN(n7379) );
  INV_X4 U7271 ( .A(n10282), .ZN(n7378) );
  INV_X4 U7272 ( .A(n7615), .ZN(n7617) );
  INV_X4 U7273 ( .A(n5865), .ZN(n7591) );
  INV_X4 U7274 ( .A(n7526), .ZN(n7522) );
  INV_X4 U7275 ( .A(reset), .ZN(n7800) );
  INV_X4 U7276 ( .A(n7798), .ZN(n7788) );
  INV_X4 U7277 ( .A(n7802), .ZN(n7793) );
  INV_X4 U7278 ( .A(n7801), .ZN(n7792) );
  NAND2_X4 U7283 ( .A1(ID_EXEC_OUT[71]), .A2(n5855), .ZN(n9262) );
  NAND2_X2 U7284 ( .A1(n9361), .A2(n9850), .ZN(n8624) );
  XNOR2_X2 U7285 ( .A(ID_EXEC_OUT[194]), .B(n7312), .ZN(n7823) );
  XNOR2_X1 U7286 ( .A(n8962), .B(n8961), .ZN(n8991) );
  NOR2_X2 U7287 ( .A1(n6014), .A2(n7773), .ZN(ID_EX_REG_ID_EX_REG_N89) );
  NAND3_X2 U7288 ( .A1(n7380), .A2(DMEM_BUS_OUT[19]), .A3(n7468), .ZN(n8426)
         );
  NAND2_X1 U7289 ( .A1(n8407), .A2(n8410), .ZN(n7807) );
  AOI21_X2 U7290 ( .B1(n9981), .B2(n10135), .A(n6344), .ZN(n10031) );
  NAND2_X1 U7291 ( .A1(n7473), .A2(n10135), .ZN(n9371) );
  NAND2_X1 U7292 ( .A1(n9246), .A2(n8947), .ZN(n8876) );
  NAND2_X2 U7293 ( .A1(n8043), .A2(n8902), .ZN(n9003) );
  INV_X2 U7294 ( .A(n8411), .ZN(n7806) );
  XNOR2_X1 U7295 ( .A(n9424), .B(n7449), .ZN(n9220) );
  INV_X1 U7296 ( .A(n9424), .ZN(n9971) );
  NAND2_X2 U7297 ( .A1(n7465), .A2(n9275), .ZN(n7904) );
  OAI211_X4 U7298 ( .C1(n6017), .C2(n9293), .A(n9277), .B(n9276), .ZN(n10104)
         );
  NAND3_X2 U7299 ( .A1(n9214), .A2(n9213), .A3(n9212), .ZN(n9424) );
  OAI221_X2 U7300 ( .B1(n9211), .B2(n9210), .C1(n7314), .C2(n9210), .A(n7472), 
        .ZN(n9212) );
  NAND2_X4 U7301 ( .A1(n9984), .A2(n10052), .ZN(n9985) );
  NOR2_X2 U7302 ( .A1(ID_EXEC_OUT[192]), .A2(n6461), .ZN(n8420) );
  NAND3_X2 U7303 ( .A1(ID_EXEC_OUT[62]), .A2(n7311), .A3(n7337), .ZN(n8022) );
  INV_X32 U7304 ( .A(n7356), .ZN(n8070) );
  NAND2_X4 U7305 ( .A1(n7460), .A2(n7356), .ZN(n7828) );
  NAND2_X1 U7306 ( .A1(n10264), .A2(n10134), .ZN(n10137) );
  INV_X1 U7307 ( .A(n10134), .ZN(n9981) );
  NAND4_X4 U7308 ( .A1(n7851), .A2(n7850), .A3(n7849), .A4(n7848), .ZN(n8904)
         );
  NAND2_X1 U7309 ( .A1(n10272), .A2(n10044), .ZN(n9629) );
  OAI21_X2 U7310 ( .B1(n9877), .B2(n9876), .A(n9875), .ZN(n9878) );
  AOI21_X2 U7311 ( .B1(n7336), .B2(n10051), .A(n10035), .ZN(n10040) );
  NAND2_X1 U7312 ( .A1(n6828), .A2(n10051), .ZN(n9826) );
  NOR2_X1 U7313 ( .A1(n10051), .A2(n9742), .ZN(n9172) );
  NOR2_X2 U7314 ( .A1(n10004), .A2(n7348), .ZN(n9955) );
  NAND3_X2 U7315 ( .A1(n10043), .A2(n10030), .A3(n10031), .ZN(n10063) );
  NAND3_X2 U7316 ( .A1(n7915), .A2(n7891), .A3(n7890), .ZN(n8423) );
  INV_X4 U7317 ( .A(n6345), .ZN(n7310) );
  NOR4_X1 U7318 ( .A1(n9783), .A2(n9782), .A3(n9941), .A4(n9951), .ZN(n9794)
         );
  AOI21_X2 U7319 ( .B1(n9143), .B2(n9941), .A(n9142), .ZN(n9144) );
  AOI211_X4 U7320 ( .C1(n7209), .C2(n8651), .A(n9568), .B(n8953), .ZN(n8483)
         );
  NAND3_X2 U7321 ( .A1(n9655), .A2(n10165), .A3(n9306), .ZN(n9307) );
  NAND2_X1 U7322 ( .A1(n10264), .A2(n9926), .ZN(n9141) );
  INV_X1 U7323 ( .A(n9926), .ZN(n9928) );
  NAND2_X1 U7324 ( .A1(n8057), .A2(DMEM_BUS_OUT[4]), .ZN(n8056) );
  NAND2_X1 U7325 ( .A1(DMEM_BUS_OUT[15]), .A2(n8057), .ZN(n7925) );
  INV_X4 U7326 ( .A(n7355), .ZN(n7311) );
  BUF_X4 U7327 ( .A(n9249), .Z(n7316) );
  NAND2_X1 U7328 ( .A1(n8907), .A2(n8947), .ZN(n8858) );
  NAND2_X1 U7329 ( .A1(n7367), .A2(n8907), .ZN(n8825) );
  INV_X1 U7330 ( .A(n7348), .ZN(n10127) );
  NAND2_X1 U7331 ( .A1(n9101), .A2(n7457), .ZN(n8798) );
  NAND2_X1 U7332 ( .A1(n7464), .A2(n9101), .ZN(n7917) );
  NAND2_X4 U7333 ( .A1(n9098), .A2(n9099), .ZN(n9299) );
  NAND2_X4 U7334 ( .A1(ID_EXEC_OUT[37]), .A2(n8058), .ZN(n7991) );
  NAND2_X4 U7335 ( .A1(n9225), .A2(n7314), .ZN(n8092) );
  NAND2_X1 U7336 ( .A1(n7370), .A2(n10234), .ZN(n8331) );
  AOI21_X1 U7337 ( .B1(n10235), .B2(n10234), .A(n10233), .ZN(n10261) );
  NOR4_X1 U7338 ( .A1(n9964), .A2(n10234), .A3(n9989), .A4(n9977), .ZN(n8079)
         );
  NAND2_X1 U7339 ( .A1(n9303), .A2(n10234), .ZN(n9656) );
  NAND2_X1 U7340 ( .A1(n7473), .A2(n10234), .ZN(n9634) );
  NAND2_X1 U7341 ( .A1(n5851), .A2(n10234), .ZN(n9186) );
  XNOR2_X1 U7342 ( .A(n9303), .B(n10234), .ZN(n10226) );
  INV_X1 U7343 ( .A(n10234), .ZN(n9016) );
  NAND2_X1 U7344 ( .A1(n7372), .A2(n9927), .ZN(n8362) );
  INV_X1 U7345 ( .A(n9927), .ZN(n9140) );
  NOR2_X1 U7346 ( .A1(n9927), .A2(n9925), .ZN(n7926) );
  NAND2_X1 U7347 ( .A1(n7473), .A2(n9927), .ZN(n9127) );
  NAND2_X1 U7348 ( .A1(n9279), .A2(n9927), .ZN(n9580) );
  XNOR2_X1 U7349 ( .A(n9279), .B(n9927), .ZN(n9579) );
  NAND2_X1 U7350 ( .A1(n9928), .A2(n9927), .ZN(n9946) );
  INV_X1 U7351 ( .A(n9976), .ZN(n9740) );
  OAI211_X4 U7352 ( .C1(n5920), .C2(n9293), .A(n9262), .B(n9261), .ZN(n9976)
         );
  OAI211_X4 U7353 ( .C1(n5921), .C2(n9293), .A(n9268), .B(n9267), .ZN(n9973)
         );
  OAI221_X2 U7354 ( .B1(n9016), .B2(n7391), .C1(n9015), .C2(n9804), .A(n9633), 
        .ZN(n9017) );
  NAND3_X2 U7355 ( .A1(DMEM_BUS_OUT[1]), .A2(n8070), .A3(n7337), .ZN(n7995) );
  XOR2_X2 U7356 ( .A(ID_EXEC_OUT[194]), .B(n7350), .Z(n7819) );
  INV_X2 U7357 ( .A(n9837), .ZN(n9839) );
  OAI22_X1 U7358 ( .A1(n9781), .A2(n9742), .B1(n7225), .B2(n10274), .ZN(n9607)
         );
  XNOR2_X2 U7359 ( .A(n9924), .B(n9925), .ZN(n9781) );
  NAND2_X1 U7360 ( .A1(n7373), .A2(n9987), .ZN(n8278) );
  NAND2_X1 U7361 ( .A1(n7475), .A2(n9987), .ZN(n8530) );
  XNOR2_X1 U7362 ( .A(n9309), .B(n9987), .ZN(n9626) );
  NAND2_X1 U7363 ( .A1(n7390), .A2(n9987), .ZN(n8605) );
  NAND2_X1 U7364 ( .A1(n7473), .A2(n9987), .ZN(n9641) );
  INV_X1 U7365 ( .A(n9987), .ZN(n9652) );
  NAND2_X1 U7366 ( .A1(n9988), .A2(n9987), .ZN(n10029) );
  NAND2_X2 U7367 ( .A1(n7382), .A2(n9863), .ZN(n9869) );
  NOR2_X1 U7368 ( .A1(n10232), .A2(n6861), .ZN(n10233) );
  NAND2_X1 U7369 ( .A1(n10232), .A2(n9995), .ZN(n10001) );
  NAND2_X4 U7370 ( .A1(n8492), .A2(n7384), .ZN(n7313) );
  NOR2_X2 U7371 ( .A1(IF_ID_OUT[33]), .A2(n1656), .ZN(ID_EX_REG_ID_EX_REG_N14)
         );
  NAND3_X2 U7372 ( .A1(IF_ID_OUT[33]), .A2(n6347), .A3(n3323), .ZN(n3357) );
  NAND3_X2 U7373 ( .A1(n3329), .A2(IF_ID_OUT[37]), .A3(IF_ID_OUT[33]), .ZN(
        n3341) );
  NOR4_X4 U7374 ( .A1(n3320), .A2(IF_ID_OUT[33]), .A3(IF_ID_OUT[34]), .A4(
        IF_ID_OUT[36]), .ZN(n3324) );
  INV_X4 U7375 ( .A(n8075), .ZN(n7314) );
  NAND2_X1 U7376 ( .A1(n7465), .A2(n9249), .ZN(n8068) );
  INV_X4 U7377 ( .A(n6349), .ZN(n7317) );
  XNOR2_X2 U7378 ( .A(n10187), .B(n9989), .ZN(n7318) );
  XNOR2_X1 U7379 ( .A(n10187), .B(n9989), .ZN(n9992) );
  OAI211_X4 U7380 ( .C1(n7313), .C2(n6019), .A(n9251), .B(n9250), .ZN(n10187)
         );
  INV_X4 U7381 ( .A(n7320), .ZN(n7321) );
  NOR2_X1 U7382 ( .A1(n8983), .A2(n7389), .ZN(n8731) );
  OAI21_X1 U7383 ( .B1(n6350), .B2(n7389), .A(n9639), .ZN(n9357) );
  NOR2_X1 U7384 ( .A1(n9721), .A2(n7389), .ZN(n9724) );
  NOR2_X1 U7385 ( .A1(n8982), .A2(n7389), .ZN(n8612) );
  OAI22_X1 U7386 ( .A1(n9532), .A2(n10246), .B1(n9531), .B2(n7389), .ZN(n8986)
         );
  NOR2_X1 U7387 ( .A1(n9703), .A2(n7389), .ZN(n9642) );
  INV_X1 U7388 ( .A(n7389), .ZN(n10146) );
  OAI22_X1 U7389 ( .A1(n9640), .A2(n7389), .B1(n9703), .B2(n10246), .ZN(n9710)
         );
  NOR2_X2 U7390 ( .A1(n9538), .A2(n7389), .ZN(n9541) );
  OAI22_X1 U7391 ( .A1(n6350), .A2(n10246), .B1(n9722), .B2(n7389), .ZN(n9680)
         );
  NOR2_X1 U7392 ( .A1(n9532), .A2(n7389), .ZN(n9533) );
  NOR2_X1 U7393 ( .A1(n9810), .A2(n7389), .ZN(n9811) );
  INV_X1 U7394 ( .A(n10265), .ZN(n10267) );
  INV_X8 U7395 ( .A(n9470), .ZN(n9473) );
  INV_X1 U7396 ( .A(n9966), .ZN(n9158) );
  OAI21_X2 U7397 ( .B1(n8271), .B2(n7374), .A(n8270), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N70) );
  NAND3_X2 U7398 ( .A1(n9485), .A2(n7479), .A3(n9484), .ZN(n9486) );
  NOR2_X1 U7399 ( .A1(n9158), .A2(n7391), .ZN(n8533) );
  NOR2_X2 U7400 ( .A1(n9158), .A2(n9182), .ZN(n9159) );
  INV_X1 U7401 ( .A(n10066), .ZN(n10070) );
  NOR2_X2 U7402 ( .A1(n9879), .A2(n9878), .ZN(n9880) );
  INV_X1 U7403 ( .A(n9878), .ZN(n9881) );
  OAI21_X2 U7404 ( .B1(n9738), .B2(n9737), .A(n9736), .ZN(n9739) );
  NAND3_X1 U7405 ( .A1(n8958), .A2(n8957), .A3(n8956), .ZN(n9563) );
  INV_X8 U7406 ( .A(n8019), .ZN(n8909) );
  INV_X1 U7407 ( .A(n9863), .ZN(n9060) );
  INV_X1 U7408 ( .A(n9866), .ZN(n9776) );
  OAI21_X2 U7409 ( .B1(n9065), .B2(n7393), .A(n9041), .ZN(n9042) );
  NAND3_X2 U7410 ( .A1(n9713), .A2(n9712), .A3(n9711), .ZN(n10204) );
  OAI21_X2 U7411 ( .B1(n9060), .B2(n7371), .A(n8757), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N43) );
  OAI22_X1 U7412 ( .A1(n9060), .A2(n8971), .B1(n9179), .B2(n9182), .ZN(n8972)
         );
  INV_X4 U7413 ( .A(n7460), .ZN(n8043) );
  NAND2_X4 U7414 ( .A1(DMEM_BUS_OUT[24]), .A2(n7380), .ZN(n8447) );
  NAND3_X1 U7415 ( .A1(n9712), .A2(n9596), .A3(n8518), .ZN(n9599) );
  NAND3_X1 U7416 ( .A1(n9107), .A2(n9596), .A3(n9374), .ZN(n10197) );
  NAND3_X2 U7417 ( .A1(n9119), .A2(n9596), .A3(n9365), .ZN(n10249) );
  NAND3_X2 U7418 ( .A1(n8530), .A2(n9596), .A3(n9670), .ZN(n10107) );
  NAND3_X2 U7419 ( .A1(n8519), .A2(n9596), .A3(n9634), .ZN(n10250) );
  NAND3_X2 U7420 ( .A1(n9106), .A2(n9596), .A3(n9371), .ZN(n10198) );
  NAND3_X2 U7421 ( .A1(n9590), .A2(n9596), .A3(n8529), .ZN(n9529) );
  NAND3_X2 U7422 ( .A1(n3302), .A2(n3303), .A3(n3304), .ZN(n3295) );
  NAND4_X4 U7423 ( .A1(n9302), .A2(n9301), .A3(n9300), .A4(n9299), .ZN(n10165)
         );
  NAND2_X4 U7424 ( .A1(n9301), .A2(n10103), .ZN(n10265) );
  INV_X2 U7425 ( .A(n9627), .ZN(n9391) );
  NAND3_X1 U7426 ( .A1(n9456), .A2(n7479), .A3(n9455), .ZN(n9457) );
  NAND2_X1 U7427 ( .A1(n9813), .A2(n9631), .ZN(n9638) );
  NAND3_X1 U7428 ( .A1(n9176), .A2(n8637), .A3(n8636), .ZN(n9021) );
  NAND2_X1 U7429 ( .A1(n10147), .A2(n9631), .ZN(n9369) );
  NOR2_X4 U7430 ( .A1(n9627), .A2(n9387), .ZN(n7324) );
  NAND2_X1 U7431 ( .A1(n9309), .A2(n9987), .ZN(n9448) );
  AOI22_X1 U7432 ( .A1(n6334), .A2(n7304), .B1(n7453), .B2(n6833), .ZN(n8139)
         );
  AOI21_X1 U7433 ( .B1(n5399), .B2(n7453), .A(ID_EXEC_OUT[145]), .ZN(n5398) );
  NAND3_X1 U7434 ( .A1(n8292), .A2(n8291), .A3(n7229), .ZN(n8294) );
  OAI211_X1 U7435 ( .C1(n6186), .C2(n8281), .A(n8280), .B(n8759), .ZN(n8283)
         );
  AND4_X4 U7436 ( .A1(n3378), .A2(n4809), .A3(n4810), .A4(n4811), .ZN(n3320)
         );
  INV_X4 U7437 ( .A(n7329), .ZN(n7325) );
  NAND2_X4 U7438 ( .A1(n7229), .A2(n8291), .ZN(n8285) );
  AOI21_X4 U7439 ( .B1(n9732), .B2(n9256), .A(n10132), .ZN(n7326) );
  NAND2_X1 U7440 ( .A1(n9254), .A2(n10163), .ZN(n9732) );
  INV_X2 U7441 ( .A(n9256), .ZN(n10131) );
  XNOR2_X1 U7442 ( .A(n9257), .B(n10135), .ZN(n10132) );
  NAND3_X2 U7443 ( .A1(n8451), .A2(n7450), .A3(n7468), .ZN(n8452) );
  NAND4_X4 U7444 ( .A1(n8413), .A2(n8412), .A3(n8411), .A4(n8410), .ZN(n8414)
         );
  NOR2_X2 U7445 ( .A1(n9483), .A2(n9487), .ZN(n9494) );
  NAND2_X4 U7446 ( .A1(n7236), .A2(n9479), .ZN(n9487) );
  OAI221_X4 U7447 ( .B1(n9474), .B2(n10279), .C1(n9473), .C2(n9646), .A(n9472), 
        .ZN(n9475) );
  NAND3_X2 U7448 ( .A1(DMEM_BUS_OUT[25]), .A2(n8492), .A3(n7469), .ZN(n8429)
         );
  NAND3_X2 U7449 ( .A1(DMEM_BUS_OUT[22]), .A2(n8492), .A3(n7469), .ZN(n8464)
         );
  NAND3_X1 U7450 ( .A1(ID_EXEC_OUT[83]), .A2(n8493), .A3(n7469), .ZN(n8425) );
  NAND3_X1 U7451 ( .A1(DMEM_BUS_OUT[18]), .A2(n8492), .A3(n7469), .ZN(n9082)
         );
  NAND3_X1 U7452 ( .A1(ID_EXEC_OUT[73]), .A2(n5853), .A3(n7468), .ZN(n9243) );
  AOI21_X1 U7453 ( .B1(n10264), .B2(n10263), .A(n6844), .ZN(n10288) );
  INV_X1 U7454 ( .A(n10263), .ZN(n9999) );
  NAND3_X2 U7455 ( .A1(n9228), .A2(n9227), .A3(n9226), .ZN(n9477) );
  NAND3_X2 U7456 ( .A1(n9242), .A2(n9241), .A3(n9240), .ZN(n9978) );
  NOR2_X1 U7457 ( .A1(n7329), .A2(n7223), .ZN(n7328) );
  INV_X16 U7458 ( .A(n7470), .ZN(n7468) );
  NAND2_X4 U7459 ( .A1(n9284), .A2(n9283), .ZN(n10100) );
  NAND2_X1 U7460 ( .A1(n7373), .A2(n9850), .ZN(n8587) );
  NAND2_X1 U7461 ( .A1(n7475), .A2(n9850), .ZN(n9128) );
  AOI22_X1 U7462 ( .A1(n9189), .A2(n9850), .B1(n7390), .B2(n9927), .ZN(n9191)
         );
  INV_X2 U7463 ( .A(n9850), .ZN(n9009) );
  AOI22_X1 U7464 ( .A1(n10112), .A2(n9180), .B1(n8967), .B2(n9850), .ZN(n9346)
         );
  NAND2_X1 U7465 ( .A1(n7390), .A2(n9850), .ZN(n9362) );
  OAI21_X1 U7466 ( .B1(n8503), .B2(n9075), .A(n9500), .ZN(n8504) );
  XNOR2_X1 U7467 ( .A(n9528), .B(n9527), .ZN(n9560) );
  INV_X16 U7468 ( .A(n7323), .ZN(n7453) );
  XOR2_X2 U7469 ( .A(n7330), .B(n7331), .Z(n7820) );
  XNOR2_X2 U7470 ( .A(n7332), .B(n7333), .ZN(n7816) );
  NAND2_X2 U7471 ( .A1(n7465), .A2(n8894), .ZN(n7937) );
  NAND2_X2 U7472 ( .A1(n7465), .A2(n8904), .ZN(n7852) );
  OAI211_X1 U7473 ( .C1(n9164), .C2(n9069), .A(n9068), .B(n10229), .ZN(n9070)
         );
  OAI22_X1 U7474 ( .A1(n9800), .A2(n9164), .B1(n9065), .B2(n7392), .ZN(n9066)
         );
  NAND2_X1 U7475 ( .A1(n10264), .A2(n9871), .ZN(n9049) );
  OAI22_X1 U7476 ( .A1(n9872), .A2(n9164), .B1(n7365), .B2(n9024), .ZN(n9756)
         );
  OAI22_X1 U7477 ( .A1(n9877), .A2(n9164), .B1(n9060), .B2(n9024), .ZN(n9752)
         );
  NOR2_X1 U7478 ( .A1(n9165), .A2(n9164), .ZN(n9166) );
  INV_X2 U7479 ( .A(n9164), .ZN(n9815) );
  NAND2_X1 U7480 ( .A1(n9412), .A2(n9871), .ZN(n9440) );
  NAND2_X1 U7481 ( .A1(n7473), .A2(n9871), .ZN(n8971) );
  NOR2_X1 U7482 ( .A1(n9872), .A2(n9871), .ZN(n9873) );
  NAND2_X2 U7483 ( .A1(n7383), .A2(n9871), .ZN(n10246) );
  NAND2_X2 U7484 ( .A1(n9180), .A2(n7382), .ZN(n9806) );
  NOR4_X2 U7485 ( .A1(n10056), .A2(n10070), .A3(n10061), .A4(n10069), .ZN(
        n10059) );
  INV_X4 U7486 ( .A(n7334), .ZN(n7335) );
  INV_X4 U7487 ( .A(n7336), .ZN(n10032) );
  INV_X8 U7488 ( .A(n7461), .ZN(n7337) );
  INV_X16 U7489 ( .A(n7466), .ZN(n7471) );
  NAND3_X2 U7490 ( .A1(n9004), .A2(n9003), .A3(n9002), .ZN(n9005) );
  AOI21_X2 U7491 ( .B1(n9335), .B2(n9334), .A(n9333), .ZN(n9337) );
  NOR2_X2 U7492 ( .A1(n9524), .A2(n9331), .ZN(n8503) );
  NOR3_X2 U7493 ( .A1(n9503), .A2(n9502), .A3(n9501), .ZN(n9506) );
  INV_X2 U7494 ( .A(n9568), .ZN(n8465) );
  OAI221_X1 U7495 ( .B1(n9900), .B2(n6861), .C1(n9578), .C2(n7479), .A(n9577), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N91) );
  BUF_X16 U7496 ( .A(n9868), .Z(n7338) );
  NAND2_X1 U7497 ( .A1(n9045), .A2(n9044), .ZN(n9046) );
  NAND2_X1 U7498 ( .A1(n9425), .A2(n9970), .ZN(n9426) );
  NAND2_X1 U7499 ( .A1(n7473), .A2(n9970), .ZN(n9359) );
  XNOR2_X1 U7500 ( .A(n9220), .B(n9970), .ZN(n9400) );
  NAND2_X1 U7501 ( .A1(n9220), .A2(n9970), .ZN(n9221) );
  NAND2_X1 U7502 ( .A1(n7475), .A2(n9970), .ZN(n9106) );
  NAND2_X1 U7503 ( .A1(n9189), .A2(n9970), .ZN(n8609) );
  NAND2_X1 U7504 ( .A1(n7390), .A2(n9970), .ZN(n8536) );
  AOI21_X1 U7505 ( .B1(n7370), .B2(n9970), .A(n8250), .ZN(n8251) );
  NOR2_X1 U7506 ( .A1(n9987), .A2(n9970), .ZN(n8011) );
  AOI21_X1 U7507 ( .B1(n10264), .B2(n10164), .A(n6844), .ZN(n10185) );
  XNOR2_X1 U7508 ( .A(n10169), .B(n10168), .ZN(n10184) );
  XNOR2_X1 U7509 ( .A(n9615), .B(n9614), .ZN(n9625) );
  NAND2_X1 U7510 ( .A1(n10264), .A2(n9908), .ZN(n9621) );
  INV_X2 U7511 ( .A(n9908), .ZN(n9910) );
  NAND2_X1 U7512 ( .A1(n8502), .A2(n9909), .ZN(n9500) );
  INV_X1 U7513 ( .A(n8953), .ZN(n8951) );
  NOR3_X2 U7514 ( .A1(n10071), .A2(n10070), .A3(n10069), .ZN(n10072) );
  NAND2_X4 U7515 ( .A1(n10009), .A2(n10018), .ZN(n7339) );
  INV_X4 U7516 ( .A(n7339), .ZN(n7340) );
  OR2_X1 U7517 ( .A1(n10217), .A2(n7315), .ZN(n7341) );
  OR2_X2 U7518 ( .A1(n10228), .A2(n9991), .ZN(n7342) );
  NAND3_X4 U7519 ( .A1(n7341), .A2(n7342), .A3(n10005), .ZN(n10008) );
  NOR3_X2 U7520 ( .A1(n10041), .A2(n10010), .A3(n10063), .ZN(n10009) );
  OAI211_X4 U7521 ( .C1(n7313), .C2(n6024), .A(n9292), .B(n9291), .ZN(n10228)
         );
  BUF_X4 U7522 ( .A(n10073), .Z(n7346) );
  NAND4_X4 U7523 ( .A1(n8202), .A2(n8201), .A3(n8200), .A4(n8550), .ZN(n8334)
         );
  NAND2_X1 U7524 ( .A1(n7372), .A2(n9916), .ZN(n8396) );
  NOR2_X1 U7525 ( .A1(n9909), .A2(n9916), .ZN(n7897) );
  NAND2_X1 U7526 ( .A1(n7473), .A2(n9916), .ZN(n8531) );
  NAND2_X1 U7527 ( .A1(n7476), .A2(n9916), .ZN(n9373) );
  INV_X2 U7528 ( .A(n9916), .ZN(n9155) );
  NAND2_X1 U7529 ( .A1(n9078), .A2(n9916), .ZN(n9499) );
  NAND2_X1 U7530 ( .A1(n9917), .A2(n9916), .ZN(n9938) );
  NOR2_X2 U7531 ( .A1(n10057), .A2(n10056), .ZN(n10058) );
  NOR3_X2 U7532 ( .A1(n10042), .A2(n10041), .A3(n10056), .ZN(n10060) );
  NAND2_X4 U7533 ( .A1(n10040), .A2(n10039), .ZN(n10056) );
  XNOR2_X1 U7534 ( .A(n9888), .B(n7449), .ZN(n7343) );
  NOR2_X1 U7535 ( .A1(n8141), .A2(n7215), .ZN(n8142) );
  OAI21_X1 U7536 ( .B1(n8343), .B2(n8353), .A(n8342), .ZN(n8345) );
  AOI21_X1 U7537 ( .B1(n10264), .B2(n9876), .A(n6844), .ZN(n9769) );
  OAI211_X1 U7538 ( .C1(n9061), .C2(n7383), .A(n9023), .B(n9022), .ZN(n9760)
         );
  OAI211_X1 U7539 ( .C1(n10034), .C2(n9598), .A(n9597), .B(n9596), .ZN(n10245)
         );
  NOR2_X2 U7540 ( .A1(n9864), .A2(n9061), .ZN(n9062) );
  INV_X4 U7541 ( .A(n7477), .ZN(n7476) );
  INV_X4 U7542 ( .A(n7623), .ZN(n7622) );
  NOR2_X2 U7543 ( .A1(n7344), .A2(n8953), .ZN(n8480) );
  NAND3_X1 U7544 ( .A1(n9562), .A2(n8959), .A3(n9563), .ZN(n8992) );
  NAND2_X4 U7545 ( .A1(n9984), .A2(n9972), .ZN(n10067) );
  INV_X4 U7546 ( .A(n8649), .ZN(n9045) );
  XNOR2_X2 U7547 ( .A(n10187), .B(n7307), .ZN(n9252) );
  NAND2_X1 U7548 ( .A1(n9280), .A2(n8947), .ZN(n8866) );
  XNOR2_X1 U7549 ( .A(n9585), .B(n9584), .ZN(n9610) );
  NOR2_X1 U7550 ( .A1(n9690), .A2(n9657), .ZN(n9658) );
  INV_X4 U7551 ( .A(n9690), .ZN(n10166) );
  NAND2_X1 U7552 ( .A1(n9285), .A2(n9925), .ZN(n10099) );
  NAND2_X1 U7553 ( .A1(n7472), .A2(n9280), .ZN(n9281) );
  AOI21_X1 U7554 ( .B1(n8992), .B2(n8993), .A(n8960), .ZN(n8962) );
  NAND2_X1 U7555 ( .A1(n10264), .A2(n9849), .ZN(n9010) );
  NAND2_X4 U7556 ( .A1(n8485), .A2(n8465), .ZN(n8466) );
  INV_X2 U7557 ( .A(n9849), .ZN(n9851) );
  NAND3_X2 U7558 ( .A1(DMEM_BUS_OUT[30]), .A2(n8070), .A3(n7337), .ZN(n8020)
         );
  OAI21_X1 U7559 ( .B1(n10016), .B2(n10047), .A(n10048), .ZN(n10020) );
  OAI21_X2 U7560 ( .B1(n10002), .B2(n10001), .A(n10000), .ZN(n10007) );
  AOI21_X1 U7561 ( .B1(n9979), .B2(n9697), .A(n9696), .ZN(n9730) );
  NAND2_X1 U7562 ( .A1(n7473), .A2(n9979), .ZN(n9597) );
  XNOR2_X1 U7563 ( .A(n9258), .B(n9979), .ZN(n9694) );
  NAND2_X1 U7564 ( .A1(n9258), .A2(n9979), .ZN(n9736) );
  NAND2_X1 U7565 ( .A1(n5852), .A2(n9979), .ZN(n9190) );
  NAND2_X1 U7566 ( .A1(n7373), .A2(n9979), .ZN(n8297) );
  NOR2_X1 U7567 ( .A1(n9979), .A2(n9974), .ZN(n7986) );
  OAI21_X2 U7568 ( .B1(n10012), .B2(n6344), .A(n10011), .ZN(n10015) );
  NOR2_X2 U7569 ( .A1(n10012), .A2(n6861), .ZN(n9696) );
  NAND3_X2 U7570 ( .A1(n9363), .A2(n9597), .A3(n9362), .ZN(n9714) );
  AOI21_X1 U7571 ( .B1(n9191), .B2(n9190), .A(n9806), .ZN(n9192) );
  NAND4_X1 U7572 ( .A1(n8637), .A2(n9127), .A3(n9190), .A4(n8524), .ZN(n9120)
         );
  OAI21_X2 U7573 ( .B1(n8299), .B2(n8298), .A(n8297), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N65) );
  XNOR2_X1 U7574 ( .A(n9569), .B(n9568), .ZN(n9578) );
  NAND2_X1 U7575 ( .A1(n8488), .A2(n9853), .ZN(n8959) );
  NAND4_X1 U7576 ( .A1(n9901), .A2(n9900), .A3(n9780), .A4(n9913), .ZN(n9783)
         );
  NAND2_X1 U7577 ( .A1(n7373), .A2(n9632), .ZN(n8749) );
  NOR2_X1 U7578 ( .A1(n9632), .A2(n9843), .ZN(n7865) );
  NAND2_X1 U7579 ( .A1(n8699), .A2(n9632), .ZN(n8622) );
  NAND2_X1 U7580 ( .A1(n7390), .A2(n9632), .ZN(n9635) );
  NAND2_X1 U7581 ( .A1(n9189), .A2(n9632), .ZN(n9187) );
  NAND2_X1 U7582 ( .A1(n8482), .A2(n9632), .ZN(n8677) );
  OAI21_X1 U7583 ( .B1(n7322), .B2(n9761), .A(n8652), .ZN(n8654) );
  OAI21_X1 U7584 ( .B1(n7209), .B2(n7322), .A(n8651), .ZN(n8952) );
  OAI221_X1 U7585 ( .B1(n10013), .B2(n6861), .C1(n9689), .C2(n7479), .A(n9688), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N107) );
  NAND2_X1 U7586 ( .A1(n10264), .A2(n9973), .ZN(n9666) );
  NAND2_X1 U7587 ( .A1(n10046), .A2(n10013), .ZN(n9789) );
  XNOR2_X1 U7588 ( .A(n9973), .B(n7449), .ZN(n9310) );
  INV_X2 U7589 ( .A(n9973), .ZN(n9975) );
  NAND3_X2 U7590 ( .A1(n9137), .A2(n9104), .A3(n7450), .ZN(n9103) );
  OAI21_X2 U7591 ( .B1(n7306), .B2(n9102), .A(n7468), .ZN(n9104) );
  NOR2_X1 U7592 ( .A1(n5853), .A2(n6030), .ZN(n9102) );
  XNOR2_X2 U7593 ( .A(n9994), .B(n9993), .ZN(n7348) );
  INV_X2 U7594 ( .A(n7349), .ZN(n7350) );
  NAND2_X2 U7595 ( .A1(n7464), .A2(n9260), .ZN(n8076) );
  INV_X2 U7596 ( .A(n8489), .ZN(n8960) );
  INV_X16 U7597 ( .A(n7460), .ZN(n7464) );
  NAND2_X1 U7598 ( .A1(n7370), .A2(n9668), .ZN(n8752) );
  NAND2_X1 U7599 ( .A1(n8699), .A2(n9668), .ZN(n8700) );
  NAND2_X1 U7600 ( .A1(n7475), .A2(n9668), .ZN(n8506) );
  NAND2_X1 U7601 ( .A1(n7390), .A2(n9668), .ZN(n9671) );
  NAND2_X1 U7602 ( .A1(n9027), .A2(n9668), .ZN(n9034) );
  NAND2_X1 U7603 ( .A1(n9189), .A2(n9668), .ZN(n9161) );
  INV_X2 U7604 ( .A(n9668), .ZN(n9872) );
  NAND2_X1 U7605 ( .A1(n8649), .A2(n8648), .ZN(n9047) );
  NAND2_X4 U7606 ( .A1(n9876), .A2(n8738), .ZN(n9804) );
  NAND4_X2 U7607 ( .A1(n9957), .A2(n9956), .A3(n9955), .A4(n7318), .ZN(n9958)
         );
  NAND2_X4 U7608 ( .A1(n9852), .A2(n9854), .ZN(n9858) );
  AOI21_X1 U7609 ( .B1(n9143), .B2(n9852), .A(n9011), .ZN(n9012) );
  INV_X1 U7610 ( .A(n9852), .ZN(n9775) );
  NAND4_X2 U7611 ( .A1(n7977), .A2(n7976), .A3(n7975), .A4(n7974), .ZN(n7351)
         );
  NAND4_X2 U7612 ( .A1(n7977), .A2(n7976), .A3(n7975), .A4(n7974), .ZN(n9968)
         );
  NAND3_X1 U7613 ( .A1(ID_EXEC_OUT[34]), .A2(n7356), .A3(n7463), .ZN(n7976) );
  NOR2_X1 U7614 ( .A1(n10036), .A2(n10037), .ZN(n10038) );
  INV_X2 U7615 ( .A(n7383), .ZN(n9864) );
  INV_X8 U7616 ( .A(n9497), .ZN(n9091) );
  NAND2_X4 U7617 ( .A1(n8356), .A2(n8302), .ZN(n8343) );
  INV_X8 U7618 ( .A(n8155), .ZN(n8356) );
  NAND4_X4 U7619 ( .A1(n8226), .A2(n8264), .A3(n8263), .A4(n8229), .ZN(n8227)
         );
  INV_X8 U7620 ( .A(n8343), .ZN(n8335) );
  INV_X8 U7621 ( .A(n9498), .ZN(n9097) );
  NAND3_X1 U7622 ( .A1(n9500), .A2(n9499), .A3(n9498), .ZN(n9502) );
  NAND4_X4 U7623 ( .A1(n7912), .A2(n7911), .A3(n7910), .A4(n7909), .ZN(n7353)
         );
  NAND4_X2 U7624 ( .A1(n7912), .A2(n7911), .A3(n7910), .A4(n7909), .ZN(n9998)
         );
  NAND3_X2 U7625 ( .A1(DMEM_BUS_OUT[13]), .A2(n8070), .A3(n7462), .ZN(n7909)
         );
  NAND2_X1 U7626 ( .A1(n7370), .A2(n9966), .ZN(n8270) );
  NAND2_X1 U7627 ( .A1(n9478), .A2(n9966), .ZN(n9485) );
  NOR2_X1 U7628 ( .A1(n10135), .A2(n9966), .ZN(n8010) );
  NAND2_X1 U7629 ( .A1(n5851), .A2(n9966), .ZN(n9107) );
  NAND2_X1 U7630 ( .A1(n9788), .A2(n10048), .ZN(n9790) );
  NAND2_X1 U7631 ( .A1(n9189), .A2(n9966), .ZN(n8730) );
  XNOR2_X1 U7632 ( .A(n9229), .B(n9966), .ZN(n9488) );
  NAND2_X1 U7633 ( .A1(n7473), .A2(n9966), .ZN(n9360) );
  NAND2_X1 U7634 ( .A1(n9967), .A2(n9966), .ZN(n10066) );
  NOR2_X1 U7635 ( .A1(n9879), .A2(n6861), .ZN(n9765) );
  NAND3_X1 U7636 ( .A1(n9846), .A2(n9879), .A3(n9777), .ZN(n9778) );
  NOR2_X1 U7637 ( .A1(n8955), .A2(n8954), .ZN(n8956) );
  NAND3_X1 U7638 ( .A1(DMEM_BUS_OUT[17]), .A2(n8492), .A3(n7468), .ZN(n9089)
         );
  NAND3_X1 U7639 ( .A1(n7381), .A2(n7468), .A3(ID_EXEC_OUT[67]), .ZN(n9227) );
  NAND3_X1 U7640 ( .A1(ID_EXEC_OUT[81]), .A2(n7381), .A3(n7468), .ZN(n9088) );
  NAND3_X1 U7641 ( .A1(DMEM_BUS_OUT[3]), .A2(n7468), .A3(n8492), .ZN(n9226) );
  NAND3_X1 U7642 ( .A1(ID_EXEC_OUT[82]), .A2(n5853), .A3(n7468), .ZN(n9081) );
  NAND3_X1 U7643 ( .A1(n7381), .A2(n7468), .A3(ID_EXEC_OUT[65]), .ZN(n9213) );
  NAND3_X1 U7644 ( .A1(DMEM_BUS_OUT[1]), .A2(n7468), .A3(n8492), .ZN(n9214) );
  NAND3_X1 U7645 ( .A1(n8492), .A2(DMEM_BUS_OUT[8]), .A3(n7468), .ZN(n9242) );
  NAND3_X1 U7646 ( .A1(ID_EXEC_OUT[72]), .A2(n7381), .A3(n7468), .ZN(n9241) );
  NAND3_X1 U7647 ( .A1(n7380), .A2(DMEM_BUS_OUT[9]), .A3(n7468), .ZN(n9244) );
  INV_X1 U7648 ( .A(n10026), .ZN(n10024) );
  OAI21_X1 U7649 ( .B1(n10085), .B2(n7307), .A(n9055), .ZN(n9056) );
  NAND2_X1 U7650 ( .A1(n7372), .A2(n9993), .ZN(n8348) );
  NAND2_X1 U7651 ( .A1(n9275), .A2(n8947), .ZN(n8868) );
  NAND2_X1 U7652 ( .A1(n7473), .A2(n9993), .ZN(n9712) );
  INV_X2 U7653 ( .A(n9993), .ZN(n10105) );
  NAND2_X1 U7654 ( .A1(n9278), .A2(n9993), .ZN(n10219) );
  XNOR2_X1 U7655 ( .A(n9278), .B(n9993), .ZN(n9297) );
  NAND2_X1 U7656 ( .A1(n9588), .A2(n9993), .ZN(n9176) );
  NAND2_X1 U7657 ( .A1(n7471), .A2(n9275), .ZN(n9276) );
  INV_X2 U7658 ( .A(n9653), .ZN(n9662) );
  INV_X8 U7659 ( .A(n9807), .ZN(n7382) );
  OAI21_X1 U7660 ( .B1(n9877), .B2(n9598), .A(n8628), .ZN(n10112) );
  NAND2_X4 U7661 ( .A1(n10037), .A2(n10032), .ZN(n9984) );
  NAND2_X1 U7662 ( .A1(n7372), .A2(n9887), .ZN(n8578) );
  AOI21_X1 U7663 ( .B1(n8965), .B2(n9887), .A(n8964), .ZN(n8990) );
  NOR2_X1 U7664 ( .A1(n9857), .A2(n6861), .ZN(n8964) );
  NOR4_X1 U7665 ( .A1(n9887), .A2(n9850), .A3(n9889), .A4(n9912), .ZN(n8081)
         );
  NAND3_X1 U7666 ( .A1(n9857), .A2(n9775), .A3(n9774), .ZN(n9779) );
  NAND2_X1 U7667 ( .A1(n7476), .A2(n9887), .ZN(n9801) );
  NAND2_X1 U7668 ( .A1(n7473), .A2(n9887), .ZN(n8613) );
  NAND2_X1 U7669 ( .A1(n7390), .A2(n9887), .ZN(n9152) );
  NAND2_X1 U7670 ( .A1(n8963), .A2(n9887), .ZN(n9896) );
  NOR4_X4 U7671 ( .A1(n3307), .A2(n3308), .A3(n3309), .A4(n3310), .ZN(n3290)
         );
  NOR3_X2 U7672 ( .A1(n9494), .A2(n9493), .A3(n9492), .ZN(n10294) );
  NAND2_X1 U7673 ( .A1(n8894), .A2(n8947), .ZN(n8860) );
  NAND2_X1 U7674 ( .A1(n7367), .A2(n8894), .ZN(n8829) );
  NAND2_X1 U7675 ( .A1(n8461), .A2(n9887), .ZN(n9564) );
  NAND3_X2 U7676 ( .A1(n10089), .A2(n6883), .A3(n10090), .ZN(n10091) );
  AOI21_X4 U7677 ( .B1(n10083), .B2(n10082), .A(n6988), .ZN(n10092) );
  INV_X4 U7678 ( .A(n9491), .ZN(n9483) );
  NOR2_X2 U7679 ( .A1(n9491), .A2(n9490), .ZN(n9492) );
  NAND2_X1 U7680 ( .A1(n9070), .A2(n9863), .ZN(n9071) );
  NAND3_X1 U7681 ( .A1(n9815), .A2(n9618), .A3(n9863), .ZN(n9041) );
  NOR2_X1 U7682 ( .A1(n9863), .A2(n9668), .ZN(n8048) );
  NAND2_X1 U7683 ( .A1(n7390), .A2(n9863), .ZN(n9711) );
  NAND2_X1 U7684 ( .A1(n7475), .A2(n9863), .ZN(n8541) );
  NAND2_X1 U7685 ( .A1(n9189), .A2(n9863), .ZN(n9174) );
  NAND2_X1 U7686 ( .A1(n8440), .A2(n9863), .ZN(n8441) );
  NAND2_X4 U7687 ( .A1(n8057), .A2(DMEM_BUS_OUT[5]), .ZN(n7992) );
  AOI211_X2 U7688 ( .C1(n10074), .C2(n10060), .A(n10058), .B(n10059), .ZN(
        n10077) );
  NAND2_X2 U7689 ( .A1(n7288), .A2(n9402), .ZN(n9324) );
  NAND2_X1 U7690 ( .A1(n9229), .A2(n9966), .ZN(n9452) );
  NAND3_X2 U7691 ( .A1(n9956), .A2(n9953), .A3(n9952), .ZN(n9959) );
  INV_X2 U7692 ( .A(n9986), .ZN(n9988) );
  XNOR2_X1 U7693 ( .A(n9986), .B(n7307), .ZN(n9309) );
  AOI21_X1 U7694 ( .B1(n10264), .B2(n9986), .A(n6844), .ZN(n9651) );
  OAI211_X4 U7695 ( .C1(n5914), .C2(n7313), .A(n9236), .B(n9235), .ZN(n9986)
         );
  AOI22_X1 U7696 ( .A1(n7367), .A2(n9260), .B1(n3552), .B2(n3390), .ZN(n3551)
         );
  NAND2_X1 U7697 ( .A1(n9260), .A2(n7457), .ZN(n8087) );
  OAI22_X1 U7698 ( .A1(n10011), .A2(n9742), .B1(n7224), .B2(n10274), .ZN(n9748) );
  XNOR2_X1 U7699 ( .A(n9976), .B(n7307), .ZN(n9265) );
  OAI221_X1 U7700 ( .B1(n9225), .B2(n9224), .C1(n7314), .C2(n9224), .A(n7471), 
        .ZN(n9228) );
  NAND2_X1 U7701 ( .A1(n7471), .A2(n9260), .ZN(n9261) );
  OAI21_X1 U7702 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[18]), .B2(n7308), 
        .A(n9223), .ZN(n8096) );
  NAND2_X1 U7703 ( .A1(n8854), .A2(n9223), .ZN(n9237) );
  NAND2_X1 U7704 ( .A1(n9211), .A2(n9223), .ZN(n8099) );
  OAI21_X2 U7705 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[25]), .B2(n7308), 
        .A(n9223), .ZN(n8851) );
  OAI21_X2 U7706 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[29]), .B2(n7308), 
        .A(n9223), .ZN(n8844) );
  INV_X8 U7707 ( .A(n8071), .ZN(n7355) );
  NAND2_X1 U7708 ( .A1(n7316), .A2(n8947), .ZN(n8874) );
  AOI21_X1 U7709 ( .B1(n10264), .B2(n7315), .A(n6844), .ZN(n10216) );
  NAND2_X4 U7710 ( .A1(n10027), .A2(n10026), .ZN(n10028) );
  NAND2_X1 U7711 ( .A1(n7471), .A2(n9249), .ZN(n9250) );
  AOI22_X4 U7712 ( .A1(n7994), .A2(n7464), .B1(n8043), .B2(n9210), .ZN(n7997)
         );
  NAND2_X4 U7713 ( .A1(n9561), .A2(n9564), .ZN(n8485) );
  NAND2_X4 U7714 ( .A1(n6479), .A2(n8422), .ZN(n8493) );
  INV_X8 U7715 ( .A(n8414), .ZN(n8422) );
  OAI22_X4 U7716 ( .A1(n8225), .A2(n7212), .B1(n8277), .B2(n8276), .ZN(n8273)
         );
  INV_X1 U7717 ( .A(n8304), .ZN(n8305) );
  XNOR2_X1 U7718 ( .A(n8277), .B(n8276), .ZN(n8279) );
  NAND2_X1 U7719 ( .A1(n8904), .A2(n7457), .ZN(n8818) );
  NAND2_X1 U7720 ( .A1(n7367), .A2(n8904), .ZN(n8821) );
  NAND2_X4 U7721 ( .A1(n7471), .A2(n8904), .ZN(n8475) );
  NAND4_X1 U7722 ( .A1(n7772), .A2(n7325), .A3(
        WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[31]), .A4(n8037), .ZN(n8041) );
  NAND3_X1 U7723 ( .A1(n7772), .A2(MEM_WB_OUT[106]), .A3(
        WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[27]), .ZN(n7856) );
  NAND2_X4 U7724 ( .A1(n7451), .A2(MEM_WB_OUT[106]), .ZN(n7888) );
  NAND3_X2 U7725 ( .A1(n9999), .A2(n7353), .A3(n9997), .ZN(n10000) );
  NAND3_X1 U7726 ( .A1(n8419), .A2(EXEC_MEM_IN[105]), .A3(n8415), .ZN(n7812)
         );
  INV_X2 U7727 ( .A(n7312), .ZN(n8114) );
  XOR2_X1 U7728 ( .A(n6016), .B(n7312), .Z(n4084) );
  XOR2_X1 U7729 ( .A(n6351), .B(n7312), .Z(n4837) );
  OAI21_X1 U7730 ( .B1(n8353), .B2(n8337), .A(n8336), .ZN(n8338) );
  OAI21_X1 U7731 ( .B1(n8326), .B2(n8325), .A(n8324), .ZN(n8328) );
  NAND2_X4 U7732 ( .A1(n7471), .A2(n8894), .ZN(n8457) );
  NAND4_X4 U7733 ( .A1(n7935), .A2(n7934), .A3(n7933), .A4(n7932), .ZN(n8894)
         );
  INV_X2 U7734 ( .A(n9924), .ZN(n9586) );
  AOI21_X2 U7735 ( .B1(n7326), .B2(n9693), .A(n9692), .ZN(n9695) );
  NOR3_X1 U7736 ( .A1(n10223), .A2(n10269), .A3(n10265), .ZN(n10224) );
  OAI21_X1 U7737 ( .B1(n10220), .B2(n10265), .A(n10219), .ZN(n10266) );
  NAND3_X1 U7738 ( .A1(RegWrite_wb_out), .A2(n8416), .A3(n8418), .ZN(n7810) );
  XNOR2_X1 U7739 ( .A(ID_EXEC_OUT[197]), .B(destReg_wb_out[4]), .ZN(n7825) );
  AOI21_X1 U7740 ( .B1(n6343), .B2(n6881), .A(n3324), .ZN(n3331) );
  NAND3_X1 U7741 ( .A1(IF_ID_OUT[36]), .A2(n1659), .A3(IF_ID_OUT[34]), .ZN(
        n3376) );
  NAND3_X1 U7742 ( .A1(n1659), .A2(IF_ID_OUT[37]), .A3(IF_ID_OUT[34]), .ZN(
        n4448) );
  NAND3_X1 U7743 ( .A1(IF_ID_OUT[33]), .A2(n3329), .A3(IF_ID_OUT[34]), .ZN(
        n3354) );
  INV_X2 U7744 ( .A(n3324), .ZN(n1592) );
  OR3_X1 U7745 ( .A1(n6346), .A2(IF_ID_OUT[34]), .A3(n3326), .ZN(n3325) );
  NAND2_X1 U7746 ( .A1(IF_ID_OUT[34]), .A2(n3323), .ZN(n3363) );
  XNOR2_X1 U7747 ( .A(n9057), .B(n9056), .ZN(n9058) );
  NAND3_X1 U7748 ( .A1(n9299), .A2(n9508), .A3(n9300), .ZN(n10223) );
  NAND3_X1 U7749 ( .A1(ID_EXEC_OUT[33]), .A2(n7337), .A3(n7356), .ZN(n7996) );
  NAND3_X1 U7750 ( .A1(ID_EXEC_OUT[63]), .A2(n7311), .A3(n9006), .ZN(n8045) );
  NAND2_X4 U7751 ( .A1(n8070), .A2(n7337), .ZN(n7906) );
  INV_X8 U7752 ( .A(n9006), .ZN(n7461) );
  NAND4_X1 U7753 ( .A1(n10162), .A2(n10003), .A3(n10011), .A4(n10012), .ZN(
        n9785) );
  NAND2_X4 U7754 ( .A1(n7829), .A2(n5913), .ZN(n9006) );
  NAND4_X4 U7755 ( .A1(n9404), .A2(n9403), .A3(n9452), .A4(n9402), .ZN(n9408)
         );
  INV_X2 U7756 ( .A(n8025), .ZN(n7841) );
  NAND2_X4 U7757 ( .A1(n7833), .A2(n7832), .ZN(n8025) );
  XNOR2_X2 U7758 ( .A(ID_EXEC_OUT[193]), .B(destReg_wb_out[0]), .ZN(n7827) );
  OAI21_X2 U7759 ( .B1(n9431), .B2(n9430), .A(n9429), .ZN(n10297) );
  NAND4_X4 U7760 ( .A1(n8486), .A2(n8485), .A3(n8484), .A4(n8483), .ZN(n9497)
         );
  INV_X8 U7761 ( .A(n9273), .ZN(n7467) );
  NAND2_X4 U7762 ( .A1(n6478), .A2(n8434), .ZN(n9273) );
  NAND2_X1 U7763 ( .A1(n7373), .A2(n7353), .ZN(n8340) );
  NAND2_X1 U7764 ( .A1(n10088), .A2(ID_EXEC_OUT[158]), .ZN(n10089) );
  NOR2_X1 U7765 ( .A1(n9993), .A2(n7353), .ZN(n7927) );
  NOR2_X1 U7766 ( .A1(n7310), .A2(n7335), .ZN(n3080) );
  NOR2_X1 U7767 ( .A1(n7334), .A2(n7310), .ZN(n3077) );
  NAND2_X1 U7768 ( .A1(n7473), .A2(n7353), .ZN(n9670) );
  NAND2_X1 U7769 ( .A1(n9288), .A2(n7353), .ZN(n10221) );
  NAND2_X1 U7770 ( .A1(n5852), .A2(n7353), .ZN(n9163) );
  XOR2_X1 U7771 ( .A(offset_26_id[3]), .B(n7310), .Z(n4087) );
  OAI21_X1 U7772 ( .B1(n10050), .B2(n6861), .A(n9426), .ZN(n9427) );
  NAND3_X1 U7773 ( .A1(n10050), .A2(n10052), .A3(n9861), .ZN(n9791) );
  AND4_X1 U7774 ( .A1(n10067), .A2(n10066), .A3(n10065), .A4(n10064), .ZN(
        n10075) );
  NAND2_X1 U7775 ( .A1(n10068), .A2(n10067), .ZN(n10071) );
  NAND2_X1 U7776 ( .A1(n10051), .A2(n10050), .ZN(n10055) );
  NAND3_X1 U7777 ( .A1(n9994), .A2(n9993), .A3(n7319), .ZN(n10002) );
  NAND2_X1 U7778 ( .A1(n9992), .A2(n10234), .ZN(n9991) );
  INV_X2 U7779 ( .A(n7319), .ZN(n10191) );
  NAND2_X4 U7780 ( .A1(n7318), .A2(n10232), .ZN(n9996) );
  OAI211_X1 U7781 ( .C1(n6187), .C2(n8273), .A(n8272), .B(n8759), .ZN(n8275)
         );
  NAND3_X1 U7782 ( .A1(n8241), .A2(n8272), .A3(n8259), .ZN(n8254) );
  OAI21_X1 U7783 ( .B1(n8286), .B2(n8285), .A(n8284), .ZN(n8296) );
  NAND2_X4 U7784 ( .A1(n8241), .A2(n8272), .ZN(n8263) );
  NAND2_X4 U7785 ( .A1(n6187), .A2(n8273), .ZN(n8272) );
  NAND2_X4 U7786 ( .A1(n8320), .A2(n8304), .ZN(n8291) );
  NOR3_X1 U7787 ( .A1(n8329), .A2(n8155), .A3(n8365), .ZN(n8205) );
  NAND2_X4 U7788 ( .A1(n10092), .A2(n10091), .ZN(n10093) );
  NAND2_X1 U7789 ( .A1(n10046), .A2(n10017), .ZN(n10019) );
  NAND2_X1 U7790 ( .A1(n8655), .A2(n8953), .ZN(n8656) );
  NAND3_X2 U7791 ( .A1(n9449), .A2(n9390), .A3(n9627), .ZN(n9393) );
  NAND4_X1 U7792 ( .A1(n9498), .A2(n9332), .A3(n9497), .A4(n9500), .ZN(n9334)
         );
  NAND2_X1 U7793 ( .A1(n9497), .A2(n9496), .ZN(n9503) );
  NAND2_X1 U7794 ( .A1(n9498), .A2(n9497), .ZN(n9524) );
  NOR2_X1 U7795 ( .A1(n7344), .A2(n8953), .ZN(n8958) );
  XNOR2_X1 U7796 ( .A(n9390), .B(n9627), .ZN(n9650) );
  NAND3_X1 U7797 ( .A1(n10165), .A2(n9691), .A3(n9732), .ZN(n9693) );
  NAND3_X1 U7798 ( .A1(n9659), .A2(n10165), .A3(n9658), .ZN(n9661) );
  NAND3_X1 U7799 ( .A1(n10128), .A2(n10165), .A3(n10166), .ZN(n10130) );
  NAND3_X1 U7800 ( .A1(n9733), .A2(n9732), .A3(n10165), .ZN(n9735) );
  NAND2_X1 U7801 ( .A1(n10166), .A2(n10165), .ZN(n10188) );
  AND3_X4 U7802 ( .A1(n3092), .A2(n7312), .A3(n7317), .ZN(n3098) );
  XOR2_X1 U7803 ( .A(n6886), .B(n7317), .Z(n4083) );
  INV_X32 U7804 ( .A(n7355), .ZN(n7356) );
  NAND2_X4 U7805 ( .A1(n7893), .A2(n7892), .ZN(n8071) );
  INV_X8 U7806 ( .A(n7906), .ZN(n8057) );
  INV_X8 U7807 ( .A(n7828), .ZN(n8058) );
  INV_X4 U7808 ( .A(n7359), .ZN(n7360) );
  INV_X4 U7809 ( .A(n7359), .ZN(n7361) );
  INV_X4 U7810 ( .A(n7362), .ZN(n7363) );
  INV_X4 U7811 ( .A(n7362), .ZN(n7364) );
  INV_X8 U7812 ( .A(n7831), .ZN(n8023) );
  INV_X16 U7813 ( .A(n9223), .ZN(n8075) );
  OAI211_X4 U7814 ( .C1(n7906), .C2(n6017), .A(n7905), .B(n7904), .ZN(n9993)
         );
  NAND2_X4 U7815 ( .A1(n7950), .A2(n9003), .ZN(n9850) );
  NAND4_X4 U7816 ( .A1(n8003), .A2(n8002), .A3(n8001), .A4(n8000), .ZN(n10135)
         );
  NAND4_X4 U7817 ( .A1(n8009), .A2(n8008), .A3(n8007), .A4(n8006), .ZN(n9966)
         );
  NAND2_X4 U7818 ( .A1(n9771), .A2(n9770), .ZN(n9835) );
  NAND2_X4 U7819 ( .A1(n6479), .A2(n8422), .ZN(n9270) );
  NAND2_X4 U7820 ( .A1(n9764), .A2(n8738), .ZN(n9802) );
  INV_X32 U7821 ( .A(n7466), .ZN(n7470) );
  XNOR2_X2 U7822 ( .A(MEM_WB_REG_MEM_WB_REG_N78), .B(ID_EXEC_OUT[198]), .ZN(
        n8411) );
  XNOR2_X2 U7823 ( .A(ID_EXEC_OUT[201]), .B(MEM_WB_REG_MEM_WB_REG_N75), .ZN(
        n8408) );
  XNOR2_X2 U7824 ( .A(ID_EXEC_OUT[202]), .B(MEM_WB_REG_MEM_WB_REG_N74), .ZN(
        n8412) );
  XNOR2_X2 U7825 ( .A(ID_EXEC_OUT[200]), .B(MEM_WB_REG_MEM_WB_REG_N76), .ZN(
        n8407) );
  XNOR2_X2 U7826 ( .A(MEM_WB_REG_MEM_WB_REG_N77), .B(ID_EXEC_OUT[199]), .ZN(
        n8410) );
  XNOR2_X2 U7827 ( .A(n7312), .B(ID_EXEC_OUT[199]), .ZN(n8419) );
  XNOR2_X2 U7828 ( .A(destReg_wb_out[2]), .B(ID_EXEC_OUT[200]), .ZN(n8415) );
  XNOR2_X2 U7829 ( .A(n7310), .B(ID_EXEC_OUT[201]), .ZN(n8417) );
  INV_X4 U7830 ( .A(n8417), .ZN(n7811) );
  XNOR2_X2 U7831 ( .A(destReg_wb_out[4]), .B(ID_EXEC_OUT[202]), .ZN(n8416) );
  XNOR2_X2 U7832 ( .A(destReg_wb_out[0]), .B(ID_EXEC_OUT[198]), .ZN(n8418) );
  INV_X4 U7833 ( .A(n6869), .ZN(n7813) );
  INV_X4 U7834 ( .A(n7814), .ZN(n7815) );
  NOR4_X2 U7835 ( .A1(n6908), .A2(EXEC_MEM_IN[105]), .A3(
        MEM_WB_REG_MEM_WB_REG_N7), .A4(ID_EXEC_OUT[192]), .ZN(n7893) );
  XNOR2_X2 U7836 ( .A(ID_EXEC_OUT[196]), .B(MEM_WB_REG_MEM_WB_REG_N75), .ZN(
        n7818) );
  XNOR2_X2 U7837 ( .A(ID_EXEC_OUT[193]), .B(MEM_WB_REG_MEM_WB_REG_N78), .ZN(
        n7817) );
  NAND3_X4 U7838 ( .A1(n7818), .A2(n7817), .A3(n7816), .ZN(n7821) );
  NOR3_X4 U7839 ( .A1(n7821), .A2(n7820), .A3(n7819), .ZN(n7892) );
  XNOR2_X2 U7840 ( .A(ID_EXEC_OUT[196]), .B(n7310), .ZN(n7824) );
  XNOR2_X2 U7841 ( .A(ID_EXEC_OUT[195]), .B(destReg_wb_out[2]), .ZN(n7822) );
  NAND4_X2 U7842 ( .A1(n7825), .A2(n7824), .A3(n7823), .A4(n7822), .ZN(n7826)
         );
  INV_X4 U7843 ( .A(n7826), .ZN(n7829) );
  NAND2_X2 U7844 ( .A1(DMEM_BUS_OUT[26]), .A2(n8057), .ZN(n7840) );
  NAND2_X2 U7845 ( .A1(ID_EXEC_OUT[58]), .A2(n8058), .ZN(n7839) );
  NAND2_X2 U7846 ( .A1(n7452), .A2(n7772), .ZN(n7830) );
  INV_X4 U7847 ( .A(n7830), .ZN(n7943) );
  NAND2_X2 U7848 ( .A1(n7210), .A2(n7943), .ZN(n7831) );
  NAND2_X2 U7849 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[26]), .A2(n8023), 
        .ZN(n7836) );
  INV_X4 U7850 ( .A(n7888), .ZN(n7832) );
  AOI22_X2 U7851 ( .A1(MEM_WB_OUT[95]), .A2(n7841), .B1(n7834), .B2(
        WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[18]), .ZN(n7835) );
  NAND3_X4 U7852 ( .A1(n7837), .A2(n7836), .A3(n7835), .ZN(n8676) );
  NAND2_X2 U7853 ( .A1(n7464), .A2(n8676), .ZN(n7838) );
  NAND3_X4 U7854 ( .A1(n7840), .A2(n7839), .A3(n7838), .ZN(n9894) );
  NAND3_X2 U7855 ( .A1(ID_EXEC_OUT[57]), .A2(n7356), .A3(n7463), .ZN(n7847) );
  NAND2_X2 U7856 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[25]), .A2(n8023), 
        .ZN(n7843) );
  NAND3_X4 U7857 ( .A1(n7844), .A2(n7843), .A3(n7842), .ZN(n8604) );
  NAND2_X2 U7858 ( .A1(n7465), .A2(n8604), .ZN(n7846) );
  NAND3_X4 U7859 ( .A1(n7845), .A2(n7846), .A3(n7847), .ZN(n9853) );
  NAND2_X2 U7860 ( .A1(DMEM_BUS_OUT[28]), .A2(n8057), .ZN(n7854) );
  NAND2_X2 U7861 ( .A1(ID_EXEC_OUT[60]), .A2(n8058), .ZN(n7853) );
  NAND2_X2 U7862 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[28]), .A2(n8023), 
        .ZN(n7850) );
  NAND2_X2 U7863 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[20]), .A2(n7834), 
        .ZN(n7849) );
  NAND2_X2 U7864 ( .A1(MEM_WB_OUT[97]), .A2(n7951), .ZN(n7848) );
  NAND3_X4 U7865 ( .A1(n7854), .A2(n7853), .A3(n7852), .ZN(n9632) );
  NAND3_X2 U7866 ( .A1(ID_EXEC_OUT[59]), .A2(n7356), .A3(n7463), .ZN(n7864) );
  NAND4_X2 U7867 ( .A1(n7772), .A2(n7451), .A3(MEM_WB_OUT[96]), .A4(n7328), 
        .ZN(n7860) );
  NAND2_X2 U7868 ( .A1(n7452), .A2(n8072), .ZN(n7942) );
  NOR2_X4 U7869 ( .A1(n7858), .A2(n7857), .ZN(n7859) );
  NAND3_X4 U7870 ( .A1(n7861), .A2(n7860), .A3(n7859), .ZN(n8724) );
  NAND2_X2 U7871 ( .A1(n7464), .A2(n8724), .ZN(n7863) );
  NAND3_X4 U7872 ( .A1(DMEM_BUS_OUT[27]), .A2(n8070), .A3(n7462), .ZN(n7862)
         );
  NAND3_X4 U7873 ( .A1(n7864), .A2(n7863), .A3(n7862), .ZN(n9843) );
  NAND2_X2 U7874 ( .A1(n7866), .A2(n7865), .ZN(n7930) );
  INV_X4 U7875 ( .A(n8025), .ZN(n7951) );
  NAND2_X2 U7876 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[18]), .A2(n8023), 
        .ZN(n7870) );
  NAND2_X2 U7877 ( .A1(n7464), .A2(n9079), .ZN(n7874) );
  NAND3_X2 U7878 ( .A1(ID_EXEC_OUT[50]), .A2(n7356), .A3(n7463), .ZN(n7873) );
  NAND3_X4 U7879 ( .A1(n7874), .A2(n7873), .A3(n7872), .ZN(n9919) );
  NAND3_X2 U7880 ( .A1(ID_EXEC_OUT[49]), .A2(n7356), .A3(n7463), .ZN(n7879) );
  NAND2_X2 U7881 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[17]), .A2(n8023), 
        .ZN(n7876) );
  NAND2_X2 U7882 ( .A1(n7465), .A2(n9086), .ZN(n7878) );
  NAND3_X4 U7883 ( .A1(n7880), .A2(n7879), .A3(n7878), .ZN(n9930) );
  NAND3_X4 U7884 ( .A1(DMEM_BUS_OUT[20]), .A2(n8070), .A3(n7462), .ZN(n7886)
         );
  NAND3_X2 U7885 ( .A1(ID_EXEC_OUT[52]), .A2(n7356), .A3(n7337), .ZN(n7885) );
  NAND2_X2 U7886 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[20]), .A2(n8023), 
        .ZN(n7882) );
  NAND3_X4 U7887 ( .A1(n7883), .A2(n7882), .A3(n7881), .ZN(n8886) );
  NAND2_X2 U7888 ( .A1(n7464), .A2(n8886), .ZN(n7884) );
  NAND3_X4 U7889 ( .A1(n7886), .A2(n7885), .A3(n7884), .ZN(n9909) );
  NAND2_X2 U7890 ( .A1(n7210), .A2(n7943), .ZN(n7887) );
  INV_X4 U7891 ( .A(n7887), .ZN(n7931) );
  AOI22_X2 U7892 ( .A1(n7889), .A2(MEM_WB_OUT[56]), .B1(MEM_WB_OUT[88]), .B2(
        n7959), .ZN(n7890) );
  NAND2_X2 U7893 ( .A1(n8043), .A2(n8423), .ZN(n7896) );
  NAND3_X4 U7894 ( .A1(n7896), .A2(n7894), .A3(n7895), .ZN(n9916) );
  NAND2_X2 U7895 ( .A1(n7898), .A2(n7897), .ZN(n7929) );
  NAND2_X2 U7896 ( .A1(ID_EXEC_OUT[46]), .A2(n8058), .ZN(n7905) );
  NAND4_X2 U7897 ( .A1(n7899), .A2(n8072), .A3(n7452), .A4(n7772), .ZN(n7900)
         );
  NAND2_X2 U7898 ( .A1(MEM_WB_OUT[51]), .A2(n7364), .ZN(n7902) );
  NAND3_X2 U7899 ( .A1(ID_EXEC_OUT[45]), .A2(n7356), .A3(n7462), .ZN(n7912) );
  NAND2_X2 U7900 ( .A1(MEM_WB_OUT[50]), .A2(n7360), .ZN(n7907) );
  NAND2_X2 U7901 ( .A1(n7465), .A2(n8843), .ZN(n7911) );
  INV_X4 U7902 ( .A(n8844), .ZN(n7908) );
  NAND2_X2 U7903 ( .A1(n7908), .A2(n7465), .ZN(n7910) );
  NAND2_X2 U7904 ( .A1(DMEM_BUS_OUT[16]), .A2(n8057), .ZN(n7919) );
  NAND2_X2 U7905 ( .A1(ID_EXEC_OUT[48]), .A2(n8058), .ZN(n7918) );
  NAND2_X2 U7906 ( .A1(n8023), .A2(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[16]), 
        .ZN(n7916) );
  NAND2_X2 U7907 ( .A1(MEM_WB_OUT[85]), .A2(n7951), .ZN(n7914) );
  NAND4_X2 U7908 ( .A1(n7916), .A2(n7915), .A3(n7914), .A4(n7913), .ZN(n9101)
         );
  NAND3_X4 U7909 ( .A1(n7919), .A2(n7918), .A3(n7917), .ZN(n9927) );
  NAND2_X2 U7910 ( .A1(ID_EXEC_OUT[47]), .A2(n8058), .ZN(n7924) );
  NAND2_X2 U7911 ( .A1(MEM_WB_OUT[52]), .A2(n7361), .ZN(n7921) );
  NAND2_X2 U7912 ( .A1(n7464), .A2(n9280), .ZN(n7923) );
  NAND3_X4 U7913 ( .A1(n7925), .A2(n7924), .A3(n7923), .ZN(n9925) );
  NAND2_X2 U7914 ( .A1(n7927), .A2(n7926), .ZN(n7928) );
  NAND3_X2 U7915 ( .A1(ID_EXEC_OUT[55]), .A2(n7356), .A3(n7463), .ZN(n7938) );
  NAND2_X2 U7916 ( .A1(MEM_WB_OUT[60]), .A2(n7361), .ZN(n7934) );
  NAND2_X2 U7917 ( .A1(MEM_WB_OUT[92]), .A2(n7959), .ZN(n7933) );
  NAND2_X2 U7918 ( .A1(n7931), .A2(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[23]), 
        .ZN(n7932) );
  NAND3_X4 U7919 ( .A1(DMEM_BUS_OUT[23]), .A2(n8070), .A3(n7462), .ZN(n7936)
         );
  NAND3_X4 U7920 ( .A1(n7938), .A2(n7937), .A3(n7936), .ZN(n9887) );
  NAND2_X2 U7921 ( .A1(DMEM_BUS_OUT[24]), .A2(n8070), .ZN(n9004) );
  INV_X4 U7922 ( .A(n9004), .ZN(n7940) );
  NAND2_X2 U7923 ( .A1(ID_EXEC_OUT[56]), .A2(n7311), .ZN(n9002) );
  INV_X4 U7924 ( .A(n9002), .ZN(n7939) );
  NAND4_X2 U7925 ( .A1(n7772), .A2(n7451), .A3(MEM_WB_OUT[93]), .A4(n7328), 
        .ZN(n7948) );
  INV_X4 U7926 ( .A(n7942), .ZN(n8037) );
  NAND3_X4 U7927 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[16]), .A2(n8014), 
        .A3(n7943), .ZN(n7944) );
  NAND3_X2 U7928 ( .A1(ID_EXEC_OUT[54]), .A2(n7356), .A3(n7337), .ZN(n7956) );
  NAND2_X2 U7929 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[22]), .A2(n8023), 
        .ZN(n7953) );
  NAND2_X2 U7930 ( .A1(n7464), .A2(n8891), .ZN(n7955) );
  NAND3_X4 U7931 ( .A1(n7957), .A2(n7956), .A3(n7955), .ZN(n9889) );
  NAND3_X4 U7932 ( .A1(DMEM_BUS_OUT[21]), .A2(n8070), .A3(n7463), .ZN(n7965)
         );
  NAND3_X2 U7933 ( .A1(ID_EXEC_OUT[53]), .A2(n7356), .A3(n7337), .ZN(n7964) );
  NAND2_X2 U7934 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[21]), .A2(n8023), 
        .ZN(n7961) );
  NAND3_X4 U7935 ( .A1(n7962), .A2(n7961), .A3(n7960), .ZN(n8888) );
  NAND2_X2 U7936 ( .A1(n7464), .A2(n8888), .ZN(n7963) );
  NAND3_X4 U7937 ( .A1(n7965), .A2(n7964), .A3(n7963), .ZN(n9912) );
  NAND2_X2 U7938 ( .A1(ID_EXEC_OUT[42]), .A2(n8058), .ZN(n7971) );
  NAND2_X2 U7939 ( .A1(MEM_WB_OUT[47]), .A2(n7361), .ZN(n7967) );
  NAND2_X2 U7940 ( .A1(n7464), .A2(n9246), .ZN(n7970) );
  NAND2_X2 U7941 ( .A1(n8057), .A2(DMEM_BUS_OUT[10]), .ZN(n7969) );
  NAND3_X4 U7942 ( .A1(n7971), .A2(n7970), .A3(n7969), .ZN(n10163) );
  NAND3_X2 U7943 ( .A1(n8070), .A2(DMEM_BUS_OUT[2]), .A3(n7460), .ZN(n7977) );
  INV_X4 U7944 ( .A(n8096), .ZN(n7972) );
  NAND2_X2 U7945 ( .A1(n7972), .A2(n7465), .ZN(n7975) );
  NAND2_X2 U7946 ( .A1(MEM_WB_OUT[39]), .A2(n7364), .ZN(n7973) );
  NAND2_X2 U7947 ( .A1(n7465), .A2(n8095), .ZN(n7974) );
  NAND2_X2 U7948 ( .A1(n7451), .A2(n6996), .ZN(n8854) );
  INV_X4 U7949 ( .A(n7889), .ZN(n7993) );
  NAND3_X4 U7950 ( .A1(n7980), .A2(n7978), .A3(n7979), .ZN(n9979) );
  NAND2_X2 U7951 ( .A1(n8057), .A2(DMEM_BUS_OUT[6]), .ZN(n7985) );
  NAND2_X2 U7952 ( .A1(ID_EXEC_OUT[38]), .A2(n8058), .ZN(n7984) );
  OAI21_X4 U7953 ( .B1(n8075), .B2(n7982), .A(n7981), .ZN(n9266) );
  NAND2_X2 U7954 ( .A1(n7464), .A2(n9266), .ZN(n7983) );
  NAND3_X4 U7955 ( .A1(n7985), .A2(n7984), .A3(n7983), .ZN(n9974) );
  NAND2_X2 U7956 ( .A1(n7987), .A2(n7986), .ZN(n8051) );
  OAI21_X4 U7957 ( .B1(n8075), .B2(n7989), .A(n7988), .ZN(n9234) );
  NAND3_X4 U7958 ( .A1(n7992), .A2(n7990), .A3(n7991), .ZN(n9987) );
  NAND2_X2 U7959 ( .A1(n7451), .A2(n6997), .ZN(n9211) );
  INV_X4 U7960 ( .A(n8099), .ZN(n7994) );
  NAND3_X4 U7961 ( .A1(n7997), .A2(n7996), .A3(n7995), .ZN(n9970) );
  NAND3_X2 U7962 ( .A1(n8070), .A2(DMEM_BUS_OUT[9]), .A3(n7463), .ZN(n8003) );
  NAND3_X2 U7963 ( .A1(ID_EXEC_OUT[41]), .A2(n7356), .A3(n7463), .ZN(n8002) );
  INV_X4 U7964 ( .A(n8851), .ZN(n7998) );
  NAND2_X2 U7965 ( .A1(n7998), .A2(n7464), .ZN(n8001) );
  NAND2_X2 U7966 ( .A1(MEM_WB_OUT[46]), .A2(n8038), .ZN(n7999) );
  NAND3_X2 U7967 ( .A1(n8070), .A2(DMEM_BUS_OUT[3]), .A3(n7463), .ZN(n8009) );
  NAND3_X2 U7968 ( .A1(ID_EXEC_OUT[35]), .A2(n7356), .A3(n7337), .ZN(n8008) );
  NAND2_X2 U7969 ( .A1(n7451), .A2(n6991), .ZN(n9225) );
  INV_X4 U7970 ( .A(n8092), .ZN(n8004) );
  NAND2_X2 U7971 ( .A1(n8004), .A2(n7465), .ZN(n8007) );
  NAND2_X2 U7972 ( .A1(MEM_WB_OUT[40]), .A2(n7364), .ZN(n8005) );
  NAND2_X2 U7973 ( .A1(n7464), .A2(n9224), .ZN(n8006) );
  NAND2_X2 U7974 ( .A1(n8011), .A2(n8010), .ZN(n8050) );
  NAND4_X2 U7975 ( .A1(n7772), .A2(n7325), .A3(
        WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[30]), .A4(n8037), .ZN(n8013) );
  NAND4_X2 U7976 ( .A1(n7772), .A2(n7451), .A3(MEM_WB_OUT[99]), .A4(n7328), 
        .ZN(n8012) );
  NAND2_X2 U7977 ( .A1(n8013), .A2(n8012), .ZN(n8018) );
  NOR2_X4 U7978 ( .A1(n8018), .A2(n8017), .ZN(n8019) );
  NAND3_X4 U7979 ( .A1(n8021), .A2(n8022), .A3(n8020), .ZN(n9863) );
  NAND3_X2 U7980 ( .A1(ID_EXEC_OUT[61]), .A2(n7356), .A3(n7463), .ZN(n8031) );
  NAND2_X2 U7981 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[29]), .A2(n8023), 
        .ZN(n8028) );
  NAND2_X2 U7982 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[21]), .A2(n7834), 
        .ZN(n8027) );
  NAND2_X2 U7983 ( .A1(MEM_WB_OUT[98]), .A2(n7841), .ZN(n8026) );
  NAND4_X2 U7984 ( .A1(n8029), .A2(n8028), .A3(n8027), .A4(n8026), .ZN(n8907)
         );
  NAND2_X2 U7985 ( .A1(n7464), .A2(n8907), .ZN(n8030) );
  NAND3_X4 U7986 ( .A1(n8031), .A2(n8032), .A3(n8030), .ZN(n9668) );
  NAND2_X2 U7987 ( .A1(n8057), .A2(DMEM_BUS_OUT[0]), .ZN(n8036) );
  NAND2_X2 U7988 ( .A1(ID_EXEC_OUT[32]), .A2(n8058), .ZN(n8035) );
  OAI21_X4 U7989 ( .B1(n8075), .B2(n6352), .A(n8033), .ZN(n9169) );
  NAND2_X2 U7990 ( .A1(n7464), .A2(n9169), .ZN(n8034) );
  NAND3_X4 U7991 ( .A1(n8036), .A2(n8035), .A3(n8034), .ZN(n9318) );
  NAND4_X2 U7992 ( .A1(n7772), .A2(n7329), .A3(
        WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[23]), .A4(n8037), .ZN(n8042) );
  NAND4_X2 U7993 ( .A1(n7772), .A2(n7451), .A3(MEM_WB_OUT[100]), .A4(n7328), 
        .ZN(n8039) );
  NAND4_X2 U7994 ( .A1(n8042), .A2(n8041), .A3(n8040), .A4(n8039), .ZN(n8948)
         );
  NAND2_X2 U7995 ( .A1(n8043), .A2(n8948), .ZN(n8044) );
  NAND2_X2 U7996 ( .A1(n8045), .A2(n8044), .ZN(n8046) );
  INV_X4 U7997 ( .A(n8046), .ZN(n9771) );
  NAND2_X2 U7998 ( .A1(n8048), .A2(n8047), .ZN(n8049) );
  NAND2_X2 U7999 ( .A1(ID_EXEC_OUT[36]), .A2(n8058), .ZN(n8055) );
  NAND2_X2 U8000 ( .A1(n7464), .A2(n9230), .ZN(n8054) );
  NAND2_X2 U8001 ( .A1(DMEM_BUS_OUT[12]), .A2(n8057), .ZN(n8063) );
  NAND2_X2 U8002 ( .A1(ID_EXEC_OUT[44]), .A2(n8058), .ZN(n8062) );
  NAND2_X2 U8003 ( .A1(MEM_WB_OUT[49]), .A2(n7363), .ZN(n8059) );
  NAND2_X2 U8004 ( .A1(n7465), .A2(n9290), .ZN(n8061) );
  NAND3_X4 U8005 ( .A1(n8063), .A2(n8062), .A3(n8061), .ZN(n10234) );
  NAND3_X2 U8006 ( .A1(ID_EXEC_OUT[43]), .A2(n7356), .A3(n7463), .ZN(n8069) );
  NAND2_X2 U8007 ( .A1(MEM_WB_OUT[48]), .A2(n7364), .ZN(n8065) );
  NAND3_X4 U8008 ( .A1(DMEM_BUS_OUT[11]), .A2(n8070), .A3(n7462), .ZN(n8067)
         );
  NAND3_X4 U8009 ( .A1(n8069), .A2(n8068), .A3(n8067), .ZN(n9989) );
  NAND3_X2 U8010 ( .A1(n8070), .A2(DMEM_BUS_OUT[7]), .A3(n7463), .ZN(n8078) );
  NAND3_X2 U8011 ( .A1(ID_EXEC_OUT[39]), .A2(n7356), .A3(n7337), .ZN(n8077) );
  NAND2_X2 U8012 ( .A1(MEM_WB_OUT[44]), .A2(n7363), .ZN(n8073) );
  NAND3_X4 U8013 ( .A1(n8078), .A2(n8077), .A3(n8076), .ZN(n9977) );
  NAND4_X2 U8014 ( .A1(n8082), .A2(n8081), .A3(n8080), .A4(n8079), .ZN(n5400)
         );
  AND2_X2 U8015 ( .A1(n4835), .A2(n7228), .ZN(n8085) );
  NAND2_X2 U8016 ( .A1(n4837), .A2(RegWrite_wb_out), .ZN(n8083) );
  INV_X4 U8017 ( .A(n4100), .ZN(n8947) );
  NAND2_X2 U8018 ( .A1(n7459), .A2(n6829), .ZN(n8086) );
  NAND2_X2 U8019 ( .A1(n9266), .A2(n7457), .ZN(n8089) );
  NAND2_X2 U8020 ( .A1(n7458), .A2(n6832), .ZN(n8088) );
  INV_X4 U8021 ( .A(n9224), .ZN(n8093) );
  NAND2_X2 U8022 ( .A1(n8093), .A2(n8092), .ZN(n8109) );
  INV_X4 U8023 ( .A(n8095), .ZN(n8097) );
  NAND2_X2 U8024 ( .A1(n8097), .A2(n8096), .ZN(n9215) );
  INV_X4 U8025 ( .A(n9210), .ZN(n8100) );
  NAND2_X2 U8026 ( .A1(n8100), .A2(n8099), .ZN(n8106) );
  NAND2_X2 U8027 ( .A1(n4082), .A2(n7213), .ZN(n8104) );
  NAND2_X2 U8028 ( .A1(n10299), .A2(n7774), .ZN(n8105) );
  AOI22_X2 U8029 ( .A1(n7368), .A2(n9266), .B1(n3531), .B2(n3390), .ZN(n3530)
         );
  AOI22_X2 U8030 ( .A1(n7368), .A2(n9234), .B1(n3509), .B2(n3390), .ZN(n3508)
         );
  AOI22_X2 U8032 ( .A1(n7367), .A2(n8109), .B1(n3466), .B2(n3390), .ZN(n3465)
         );
  AOI22_X2 U8033 ( .A1(n7367), .A2(n9215), .B1(n3445), .B2(n3390), .ZN(n3444)
         );
  AOI22_X2 U8034 ( .A1(n7368), .A2(n8106), .B1(n3423), .B2(n3390), .ZN(n3422)
         );
  AOI22_X2 U8035 ( .A1(n7368), .A2(n9169), .B1(n3391), .B2(n3390), .ZN(n3388)
         );
  NAND2_X2 U8036 ( .A1(RegWrite_wb_out), .A2(n7320), .ZN(n8112) );
  INV_X4 U8037 ( .A(n8112), .ZN(n8111) );
  NAND2_X2 U8038 ( .A1(n6034), .A2(n3080), .ZN(n3150) );
  INV_X4 U8039 ( .A(n8106), .ZN(n8107) );
  INV_X4 U8040 ( .A(n9215), .ZN(n8108) );
  INV_X4 U8041 ( .A(n8109), .ZN(n8110) );
  NAND2_X2 U8042 ( .A1(n3087), .A2(n6035), .ZN(n3148) );
  NAND2_X2 U8043 ( .A1(n3084), .A2(n6035), .ZN(n3146) );
  NAND2_X2 U8044 ( .A1(n6028), .A2(n3080), .ZN(n3135) );
  NAND2_X2 U8045 ( .A1(n6028), .A2(n3077), .ZN(n3133) );
  NAND2_X2 U8046 ( .A1(n6028), .A2(n3087), .ZN(n3131) );
  NAND2_X2 U8047 ( .A1(n6028), .A2(n3084), .ZN(n3128) );
  NAND2_X2 U8048 ( .A1(n6034), .A2(n3077), .ZN(n3126) );
  NAND2_X2 U8049 ( .A1(n8113), .A2(n3080), .ZN(n3114) );
  NAND2_X2 U8050 ( .A1(n8113), .A2(n3077), .ZN(n3112) );
  NAND2_X2 U8051 ( .A1(n8113), .A2(n3087), .ZN(n3110) );
  NAND2_X2 U8052 ( .A1(n8113), .A2(n3084), .ZN(n3107) );
  NAND2_X2 U8053 ( .A1(n6034), .A2(n3087), .ZN(n3101) );
  NAND2_X2 U8054 ( .A1(n6034), .A2(n3084), .ZN(n3093) );
  INV_X4 U8055 ( .A(n8118), .ZN(n8115) );
  NAND2_X2 U8056 ( .A1(n8115), .A2(n3080), .ZN(n3090) );
  INV_X4 U8057 ( .A(n3087), .ZN(n8116) );
  INV_X4 U8058 ( .A(n3084), .ZN(n8117) );
  NAND2_X2 U8059 ( .A1(n3080), .A2(n6035), .ZN(n3078) );
  OAI222_X2 U8060 ( .A1(n6266), .A2(n5908), .B1(n7354), .B2(n6834), .C1(n7484), 
        .C2(n5889), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N10) );
  OAI222_X2 U8061 ( .A1(n6320), .A2(n5908), .B1(n8119), .B2(n6835), .C1(n7484), 
        .C2(n5885), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N11) );
  OAI222_X2 U8062 ( .A1(n6321), .A2(n5908), .B1(n7354), .B2(n6836), .C1(n7484), 
        .C2(n5919), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N12) );
  OAI222_X2 U8063 ( .A1(n6324), .A2(n5908), .B1(n8119), .B2(n6837), .C1(n7484), 
        .C2(n5912), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N13) );
  OAI222_X2 U8064 ( .A1(n6322), .A2(n5908), .B1(n7354), .B2(n6838), .C1(n7484), 
        .C2(n5924), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N14) );
  OAI222_X2 U8065 ( .A1(n6323), .A2(n5908), .B1(n8119), .B2(n6839), .C1(n7484), 
        .C2(n5916), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N15) );
  OAI222_X2 U8066 ( .A1(n6325), .A2(n5908), .B1(n7354), .B2(n6840), .C1(n7484), 
        .C2(n5887), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N16) );
  OAI222_X2 U8067 ( .A1(n6330), .A2(n5908), .B1(n8119), .B2(n6841), .C1(n7484), 
        .C2(n5886), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N17) );
  OAI222_X2 U8068 ( .A1(n6318), .A2(n5908), .B1(n7354), .B2(n6842), .C1(n7484), 
        .C2(n5917), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N18) );
  OAI222_X2 U8069 ( .A1(n6319), .A2(n5908), .B1(n8119), .B2(n6843), .C1(n7483), 
        .C2(n5918), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N19) );
  OAI222_X2 U8070 ( .A1(n6808), .A2(n5908), .B1(n7354), .B2(n7270), .C1(n7483), 
        .C2(n6025), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N20) );
  OAI222_X2 U8071 ( .A1(n6812), .A2(n5908), .B1(n8119), .B2(n7271), .C1(n7483), 
        .C2(n6026), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N21) );
  OAI222_X2 U8072 ( .A1(n6809), .A2(n5908), .B1(n7354), .B2(n7272), .C1(n7483), 
        .C2(n6032), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N22) );
  OAI222_X2 U8073 ( .A1(n6810), .A2(n5908), .B1(n8119), .B2(n7273), .C1(n7483), 
        .C2(n6033), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N23) );
  OAI222_X2 U8074 ( .A1(n6811), .A2(n5908), .B1(n7354), .B2(n7274), .C1(n7483), 
        .C2(n6030), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N24) );
  OAI222_X2 U8075 ( .A1(n6818), .A2(n5908), .B1(n8119), .B2(n7275), .C1(n7483), 
        .C2(n6042), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N25) );
  OAI222_X2 U8076 ( .A1(n6819), .A2(n5908), .B1(n7354), .B2(n7276), .C1(n7483), 
        .C2(n6017), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N26) );
  OAI222_X2 U8077 ( .A1(n6820), .A2(n5908), .B1(n8119), .B2(n7277), .C1(n7483), 
        .C2(n6043), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N27) );
  OAI222_X2 U8078 ( .A1(n6821), .A2(n5908), .B1(n7354), .B2(n7278), .C1(n7483), 
        .C2(n6024), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N28) );
  OAI222_X2 U8079 ( .A1(n6822), .A2(n5908), .B1(n8119), .B2(n7279), .C1(n7483), 
        .C2(n6019), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N29) );
  OAI222_X2 U8080 ( .A1(n6813), .A2(n5908), .B1(n7354), .B2(n7280), .C1(n7483), 
        .C2(n6018), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N9) );
  INV_X4 U8081 ( .A(n6334), .ZN(n8120) );
  INV_X4 U8082 ( .A(n8225), .ZN(n8224) );
  NAND2_X2 U8083 ( .A1(nextPC_ex_out[2]), .A2(n8224), .ZN(n8248) );
  INV_X4 U8084 ( .A(n8248), .ZN(n8245) );
  NAND2_X2 U8085 ( .A1(nextPC_ex_out[1]), .A2(n8224), .ZN(n8127) );
  NAND2_X2 U8086 ( .A1(nextPC_ex_out[3]), .A2(n8224), .ZN(n8259) );
  NAND2_X2 U8087 ( .A1(n8127), .A2(n8259), .ZN(n8228) );
  NAND2_X2 U8088 ( .A1(n7369), .A2(n9318), .ZN(n8231) );
  INV_X4 U8089 ( .A(n8231), .ZN(n8122) );
  XNOR2_X2 U8090 ( .A(n8224), .B(nextPC_ex_out[0]), .ZN(n8121) );
  NAND2_X2 U8091 ( .A1(n8231), .A2(n7374), .ZN(n8123) );
  NAND2_X2 U8092 ( .A1(n8123), .A2(n8231), .ZN(n8132) );
  INV_X4 U8093 ( .A(n8132), .ZN(n8124) );
  INV_X4 U8094 ( .A(n8228), .ZN(n8126) );
  XNOR2_X2 U8095 ( .A(n8225), .B(n7217), .ZN(n8268) );
  NAND2_X2 U8096 ( .A1(n8126), .A2(n8268), .ZN(n8131) );
  XNOR2_X2 U8097 ( .A(n8225), .B(n7218), .ZN(n8244) );
  INV_X4 U8098 ( .A(n8244), .ZN(n8249) );
  XNOR2_X2 U8099 ( .A(n8225), .B(n7219), .ZN(n8261) );
  INV_X4 U8100 ( .A(n8261), .ZN(n8238) );
  NAND2_X2 U8101 ( .A1(n8249), .A2(n8238), .ZN(n8128) );
  NAND4_X2 U8102 ( .A1(n8231), .A2(n8128), .A3(n8127), .A4(n8248), .ZN(n8226)
         );
  INV_X4 U8103 ( .A(n8226), .ZN(n8129) );
  NAND2_X2 U8104 ( .A1(nextPC_ex_out[4]), .A2(n8224), .ZN(n8241) );
  INV_X4 U8105 ( .A(n6334), .ZN(n8133) );
  INV_X4 U8106 ( .A(n8210), .ZN(n8134) );
  NAND2_X2 U8107 ( .A1(nextPC_ex_out[10]), .A2(n8134), .ZN(n8310) );
  INV_X4 U8108 ( .A(n6334), .ZN(n8135) );
  INV_X4 U8109 ( .A(n8137), .ZN(n8136) );
  NAND2_X2 U8110 ( .A1(nextPC_ex_out[11]), .A2(n8136), .ZN(n8307) );
  XNOR2_X2 U8111 ( .A(n8137), .B(n7221), .ZN(n8308) );
  INV_X4 U8112 ( .A(n8308), .ZN(n8320) );
  INV_X4 U8113 ( .A(n8147), .ZN(n8149) );
  INV_X4 U8114 ( .A(n6334), .ZN(n8138) );
  INV_X4 U8115 ( .A(n8144), .ZN(n8146) );
  XNOR2_X2 U8116 ( .A(n8141), .B(n7215), .ZN(n8155) );
  NAND2_X2 U8117 ( .A1(nextPC_ex_out[16]), .A2(n8139), .ZN(n8354) );
  XNOR2_X2 U8118 ( .A(nextPC_ex_out[16]), .B(n8139), .ZN(n8351) );
  NAND2_X2 U8119 ( .A1(n8354), .A2(n8351), .ZN(n8302) );
  MUX2_X2 U8120 ( .A(n6845), .B(n7289), .S(n7453), .Z(n8140) );
  INV_X4 U8121 ( .A(n8140), .ZN(n8154) );
  NAND2_X2 U8122 ( .A1(nextPC_ex_out[17]), .A2(n8154), .ZN(n8352) );
  NAND2_X2 U8123 ( .A1(n8354), .A2(n8352), .ZN(n8143) );
  AOI21_X4 U8124 ( .B1(n8335), .B2(n8143), .A(n8142), .ZN(n8342) );
  XNOR2_X2 U8125 ( .A(n8144), .B(n7136), .ZN(n8346) );
  NOR2_X4 U8126 ( .A1(n8342), .A2(n8346), .ZN(n8145) );
  AOI21_X4 U8127 ( .B1(nextPC_ex_out[14]), .B2(n8146), .A(n8145), .ZN(n8336)
         );
  XNOR2_X2 U8128 ( .A(n8147), .B(n7137), .ZN(n8323) );
  NOR2_X4 U8129 ( .A1(n8336), .A2(n8323), .ZN(n8148) );
  AOI21_X4 U8130 ( .B1(nextPC_ex_out[13]), .B2(n8149), .A(n8148), .ZN(n8324)
         );
  XNOR2_X2 U8131 ( .A(n8150), .B(n7211), .ZN(n8329) );
  INV_X4 U8132 ( .A(n6334), .ZN(n8151) );
  INV_X4 U8133 ( .A(n8214), .ZN(n8152) );
  NAND2_X2 U8134 ( .A1(nextPC_ex_out[8]), .A2(n8152), .ZN(n8287) );
  INV_X4 U8135 ( .A(n8287), .ZN(n8217) );
  INV_X4 U8136 ( .A(n8302), .ZN(n8153) );
  XNOR2_X2 U8137 ( .A(nextPC_ex_out[17]), .B(n8154), .ZN(n8365) );
  MUX2_X2 U8138 ( .A(n6846), .B(n7290), .S(n7453), .Z(n8156) );
  INV_X4 U8139 ( .A(n8156), .ZN(n8159) );
  NAND2_X2 U8140 ( .A1(nextPC_ex_out[21]), .A2(n8159), .ZN(n8390) );
  INV_X4 U8141 ( .A(n8390), .ZN(n8552) );
  MUX2_X2 U8142 ( .A(n6847), .B(n7291), .S(n7453), .Z(n8157) );
  INV_X4 U8143 ( .A(n8157), .ZN(n8158) );
  NAND2_X2 U8144 ( .A1(nextPC_ex_out[22]), .A2(n8158), .ZN(n8569) );
  INV_X4 U8145 ( .A(n8569), .ZN(n8185) );
  INV_X4 U8146 ( .A(n8160), .ZN(n8554) );
  MUX2_X2 U8147 ( .A(n6848), .B(n7292), .S(n7453), .Z(n8161) );
  INV_X4 U8148 ( .A(n8161), .ZN(n8163) );
  INV_X4 U8149 ( .A(n8162), .ZN(n8391) );
  NAND2_X2 U8150 ( .A1(nextPC_ex_out[20]), .A2(n8163), .ZN(n8394) );
  INV_X4 U8151 ( .A(n8394), .ZN(n8165) );
  MUX2_X2 U8152 ( .A(n6849), .B(n7293), .S(n7453), .Z(n8164) );
  INV_X4 U8153 ( .A(n8164), .ZN(n8166) );
  NAND2_X2 U8154 ( .A1(nextPC_ex_out[19]), .A2(n8166), .ZN(n8380) );
  MUX2_X2 U8155 ( .A(n6850), .B(n7294), .S(n7453), .Z(n8167) );
  INV_X4 U8156 ( .A(n8167), .ZN(n8168) );
  XNOR2_X2 U8157 ( .A(nextPC_ex_out[18]), .B(n8168), .ZN(n8381) );
  NAND2_X2 U8158 ( .A1(nextPC_ex_out[18]), .A2(n8168), .ZN(n8371) );
  INV_X4 U8159 ( .A(n8371), .ZN(n8184) );
  MUX2_X2 U8160 ( .A(n6851), .B(n7295), .S(n7453), .Z(n8169) );
  INV_X4 U8161 ( .A(n8169), .ZN(n8170) );
  NAND2_X2 U8162 ( .A1(nextPC_ex_out[26]), .A2(n8170), .ZN(n8592) );
  INV_X4 U8163 ( .A(n8592), .ZN(n8173) );
  XNOR2_X2 U8164 ( .A(nextPC_ex_out[26]), .B(n8170), .ZN(n8171) );
  INV_X4 U8165 ( .A(n8171), .ZN(n8662) );
  MUX2_X2 U8166 ( .A(n6852), .B(n7296), .S(n7453), .Z(n8172) );
  INV_X4 U8167 ( .A(n8172), .ZN(n8174) );
  OAI21_X4 U8168 ( .B1(n8173), .B2(n8662), .A(n7037), .ZN(n8580) );
  NAND2_X2 U8169 ( .A1(nextPC_ex_out[25]), .A2(n8174), .ZN(n8585) );
  NAND2_X2 U8170 ( .A1(n8580), .A2(n8585), .ZN(n8565) );
  INV_X4 U8171 ( .A(n8565), .ZN(n8177) );
  MUX2_X2 U8172 ( .A(n6853), .B(n7297), .S(n7453), .Z(n8175) );
  INV_X4 U8173 ( .A(n8175), .ZN(n8182) );
  XNOR2_X2 U8174 ( .A(nextPC_ex_out[24]), .B(n8182), .ZN(n8186) );
  MUX2_X2 U8175 ( .A(n6854), .B(n7298), .S(n7453), .Z(n8176) );
  INV_X4 U8176 ( .A(n8176), .ZN(n8195) );
  NAND2_X2 U8177 ( .A1(nextPC_ex_out[27]), .A2(n8195), .ZN(n8591) );
  MUX2_X2 U8178 ( .A(n6855), .B(n7299), .S(n7453), .Z(n8178) );
  INV_X4 U8179 ( .A(n8178), .ZN(n8179) );
  XNOR2_X2 U8180 ( .A(nextPC_ex_out[23]), .B(n8179), .ZN(n8577) );
  INV_X4 U8181 ( .A(n8577), .ZN(n8367) );
  NAND2_X2 U8182 ( .A1(nextPC_ex_out[23]), .A2(n8179), .ZN(n8568) );
  NAND2_X2 U8183 ( .A1(n8568), .A2(n8380), .ZN(n8180) );
  NAND2_X2 U8184 ( .A1(nextPC_ex_out[24]), .A2(n8182), .ZN(n8366) );
  INV_X4 U8185 ( .A(n8366), .ZN(n8183) );
  NAND2_X2 U8186 ( .A1(n8183), .A2(n8367), .ZN(n8201) );
  NAND2_X2 U8187 ( .A1(n8394), .A2(n8390), .ZN(n8377) );
  INV_X4 U8188 ( .A(n8186), .ZN(n8581) );
  NAND2_X2 U8189 ( .A1(n8581), .A2(n8565), .ZN(n8586) );
  INV_X4 U8190 ( .A(n8586), .ZN(n8199) );
  MUX2_X2 U8191 ( .A(n6856), .B(n7300), .S(n7453), .Z(n8187) );
  INV_X4 U8192 ( .A(n8187), .ZN(n8189) );
  NAND2_X2 U8193 ( .A1(nextPC_ex_out[30]), .A2(n8189), .ZN(n8710) );
  MUX2_X2 U8194 ( .A(n6857), .B(n7301), .S(n7453), .Z(n8188) );
  INV_X4 U8195 ( .A(n8188), .ZN(n8193) );
  NAND2_X2 U8196 ( .A1(nextPC_ex_out[29]), .A2(n8193), .ZN(n8711) );
  MUX2_X2 U8197 ( .A(n6858), .B(n7302), .S(n7453), .Z(n8758) );
  NAND2_X2 U8198 ( .A1(nextPC_ex_out[31]), .A2(n8761), .ZN(n8760) );
  INV_X4 U8199 ( .A(n8760), .ZN(n8191) );
  XNOR2_X2 U8200 ( .A(nextPC_ex_out[30]), .B(n8189), .ZN(n8754) );
  INV_X4 U8201 ( .A(n8754), .ZN(n8190) );
  NAND2_X2 U8202 ( .A1(n8191), .A2(n8190), .ZN(n8756) );
  MUX2_X2 U8203 ( .A(n6859), .B(n7303), .S(n7453), .Z(n8192) );
  INV_X4 U8204 ( .A(n8192), .ZN(n8194) );
  NAND2_X2 U8205 ( .A1(nextPC_ex_out[28]), .A2(n8194), .ZN(n8712) );
  NAND4_X2 U8206 ( .A1(n8710), .A2(n8711), .A3(n8756), .A4(n8712), .ZN(n8564)
         );
  XNOR2_X2 U8207 ( .A(nextPC_ex_out[29]), .B(n8193), .ZN(n8751) );
  INV_X4 U8208 ( .A(n8712), .ZN(n8196) );
  INV_X4 U8209 ( .A(n8561), .ZN(n8197) );
  INV_X4 U8210 ( .A(n8590), .ZN(n8198) );
  NAND3_X4 U8211 ( .A1(n8199), .A2(n8367), .A3(n8198), .ZN(n8550) );
  INV_X4 U8212 ( .A(n8334), .ZN(n8203) );
  NOR2_X4 U8213 ( .A1(n8300), .A2(n8203), .ZN(n8204) );
  INV_X4 U8214 ( .A(n8211), .ZN(n8208) );
  NAND2_X2 U8215 ( .A1(nextPC_ex_out[9]), .A2(n8208), .ZN(n8209) );
  NAND2_X2 U8216 ( .A1(n8292), .A2(n8209), .ZN(n8286) );
  INV_X4 U8217 ( .A(n8209), .ZN(n8293) );
  INV_X4 U8218 ( .A(n8310), .ZN(n8212) );
  INV_X4 U8219 ( .A(n8213), .ZN(n8295) );
  INV_X4 U8220 ( .A(n8215), .ZN(n8284) );
  INV_X4 U8221 ( .A(n8218), .ZN(n8219) );
  NAND2_X2 U8222 ( .A1(nextPC_ex_out[7]), .A2(n8219), .ZN(n8220) );
  INV_X4 U8223 ( .A(n8280), .ZN(n8223) );
  AOI21_X4 U8224 ( .B1(nextPC_ex_out[6]), .B2(n8224), .A(n8223), .ZN(n8277) );
  XNOR2_X2 U8225 ( .A(n8225), .B(n7212), .ZN(n8276) );
  INV_X4 U8226 ( .A(n8227), .ZN(n8235) );
  INV_X4 U8227 ( .A(n8229), .ZN(n8230) );
  INV_X4 U8228 ( .A(n8233), .ZN(n8234) );
  AOI211_X4 U8229 ( .C1(n8237), .C2(n8236), .A(n8235), .B(n8234), .ZN(n10296)
         );
  INV_X4 U8230 ( .A(n8268), .ZN(n8264) );
  INV_X4 U8231 ( .A(n8259), .ZN(n8239) );
  INV_X4 U8232 ( .A(n8240), .ZN(n8255) );
  NAND2_X2 U8233 ( .A1(n8255), .A2(n8254), .ZN(n8246) );
  INV_X4 U8234 ( .A(n8246), .ZN(n8243) );
  NAND2_X2 U8235 ( .A1(n8243), .A2(n8242), .ZN(n8253) );
  NAND2_X2 U8236 ( .A1(n8247), .A2(n8246), .ZN(n8252) );
  NAND3_X2 U8237 ( .A1(n8253), .A2(n8252), .A3(n8251), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N72) );
  INV_X4 U8238 ( .A(n8254), .ZN(n8257) );
  NAND2_X2 U8239 ( .A1(n8762), .A2(n7351), .ZN(n8260) );
  NAND2_X2 U8240 ( .A1(n8255), .A2(n8260), .ZN(n8256) );
  INV_X4 U8241 ( .A(n8260), .ZN(n8258) );
  NAND3_X2 U8242 ( .A1(n8261), .A2(n8260), .A3(n8259), .ZN(n8262) );
  XNOR2_X2 U8243 ( .A(n8269), .B(n8268), .ZN(n8271) );
  NAND2_X2 U8245 ( .A1(n8275), .A2(n8274), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N69)
         );
  NAND2_X2 U8246 ( .A1(n7372), .A2(n9974), .ZN(n8282) );
  NAND2_X2 U8247 ( .A1(n8283), .A2(n8282), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N67)
         );
  NAND2_X2 U8248 ( .A1(n8296), .A2(n8287), .ZN(n8288) );
  XNOR2_X2 U8249 ( .A(n6190), .B(n8288), .ZN(n8290) );
  NAND2_X2 U8250 ( .A1(n7372), .A2(n9977), .ZN(n8289) );
  NAND2_X2 U8251 ( .A1(n8759), .A2(n8296), .ZN(n8298) );
  INV_X4 U8252 ( .A(n8300), .ZN(n8301) );
  INV_X4 U8253 ( .A(n8346), .ZN(n8344) );
  NAND2_X2 U8254 ( .A1(n8303), .A2(n7246), .ZN(n8306) );
  INV_X4 U8255 ( .A(n8319), .ZN(n8309) );
  NAND2_X2 U8256 ( .A1(n5915), .A2(n8314), .ZN(n8315) );
  NAND2_X2 U8257 ( .A1(n8315), .A2(n8310), .ZN(n8311) );
  XNOR2_X2 U8258 ( .A(n6189), .B(n8311), .ZN(n8313) );
  NAND2_X2 U8259 ( .A1(n7372), .A2(n10135), .ZN(n8312) );
  NAND2_X2 U8260 ( .A1(n8759), .A2(n8315), .ZN(n8317) );
  NAND2_X2 U8261 ( .A1(n7373), .A2(n10163), .ZN(n8316) );
  XNOR2_X2 U8262 ( .A(n8320), .B(n8319), .ZN(n8322) );
  NAND2_X2 U8263 ( .A1(n7370), .A2(n9989), .ZN(n8321) );
  INV_X4 U8264 ( .A(n8329), .ZN(n8327) );
  INV_X4 U8265 ( .A(n8323), .ZN(n8339) );
  NAND2_X2 U8266 ( .A1(n7246), .A2(n8339), .ZN(n8326) );
  INV_X4 U8267 ( .A(n8328), .ZN(n8330) );
  NAND2_X2 U8268 ( .A1(n6356), .A2(n8334), .ZN(n8353) );
  NAND2_X2 U8269 ( .A1(n8344), .A2(n8335), .ZN(n8337) );
  XNOR2_X2 U8270 ( .A(n8339), .B(n8338), .ZN(n8341) );
  INV_X4 U8271 ( .A(n8345), .ZN(n8347) );
  INV_X4 U8272 ( .A(n8351), .ZN(n8360) );
  NAND2_X2 U8273 ( .A1(n8353), .A2(n8352), .ZN(n8359) );
  NAND2_X2 U8274 ( .A1(n8360), .A2(n8359), .ZN(n8361) );
  NAND2_X2 U8275 ( .A1(n8354), .A2(n8361), .ZN(n8355) );
  XNOR2_X2 U8276 ( .A(n8356), .B(n8355), .ZN(n8358) );
  NAND2_X2 U8277 ( .A1(n7373), .A2(n9925), .ZN(n8357) );
  NAND2_X2 U8278 ( .A1(n8759), .A2(n8361), .ZN(n8363) );
  INV_X4 U8279 ( .A(n8365), .ZN(n8373) );
  NAND2_X2 U8280 ( .A1(n8559), .A2(n8367), .ZN(n8551) );
  NAND3_X2 U8281 ( .A1(n8394), .A2(n8551), .A3(n8380), .ZN(n8370) );
  NAND2_X2 U8282 ( .A1(n8386), .A2(n8371), .ZN(n8372) );
  XNOR2_X2 U8283 ( .A(n8373), .B(n8372), .ZN(n8375) );
  NAND2_X2 U8284 ( .A1(n7372), .A2(n9930), .ZN(n8374) );
  INV_X4 U8285 ( .A(n8376), .ZN(n8385) );
  INV_X4 U8286 ( .A(n8377), .ZN(n8379) );
  NAND2_X2 U8287 ( .A1(n6892), .A2(n8550), .ZN(n8392) );
  INV_X4 U8288 ( .A(n8392), .ZN(n8378) );
  INV_X4 U8289 ( .A(n8380), .ZN(n8383) );
  INV_X4 U8290 ( .A(n8381), .ZN(n8382) );
  NAND2_X2 U8291 ( .A1(n8759), .A2(n8386), .ZN(n8388) );
  NAND2_X2 U8292 ( .A1(n7373), .A2(n9919), .ZN(n8387) );
  NAND2_X2 U8293 ( .A1(n8551), .A2(n8390), .ZN(n8393) );
  NAND2_X2 U8294 ( .A1(n8394), .A2(n8555), .ZN(n8395) );
  XNOR2_X2 U8295 ( .A(n7036), .B(n8395), .ZN(n8397) );
  NAND2_X2 U8296 ( .A1(ID_EX_REG_ID_EX_REG_N81), .A2(n7447), .ZN(n8399) );
  NAND2_X2 U8297 ( .A1(n7367), .A2(n8423), .ZN(n8398) );
  NAND2_X2 U8298 ( .A1(n8399), .A2(n8398), .ZN(n8400) );
  NAND4_X2 U8299 ( .A1(n3808), .A2(n3809), .A3(n3807), .A4(n8401), .ZN(
        ID_EX_REG_ID_EX_REG_N155) );
  NAND2_X2 U8300 ( .A1(n8423), .A2(n7457), .ZN(n8403) );
  NAND2_X2 U8301 ( .A1(n7459), .A2(n6830), .ZN(n8402) );
  NAND3_X2 U8302 ( .A1(n4541), .A2(n8403), .A3(n8402), .ZN(n8406) );
  NAND2_X2 U8303 ( .A1(n6010), .A2(n8406), .ZN(n8405) );
  NAND2_X2 U8304 ( .A1(ID_EX_REG_ID_EX_REG_N81), .A2(n4447), .ZN(n8404) );
  NAND2_X2 U8305 ( .A1(n8405), .A2(n8404), .ZN(n1580) );
  AND2_X2 U8306 ( .A1(n8406), .A2(n7305), .ZN(ID_EX_REG_ID_EX_REG_N27) );
  OAI22_X2 U8307 ( .A1(n7626), .A2(n7375), .B1(n7120), .B2(n7624), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8308 ( .A1(n3148), .A2(n7376), .B1(n6167), .B2(n7628), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8309 ( .A1(n3146), .A2(n7375), .B1(n7178), .B2(n7632), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8310 ( .A1(n7639), .A2(n7376), .B1(n6589), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8311 ( .A1(n7643), .A2(n7376), .B1(n5938), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8312 ( .A1(n7647), .A2(n7377), .B1(n7026), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8313 ( .A1(n7651), .A2(n7376), .B1(n6717), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8314 ( .A1(n7654), .A2(n7377), .B1(n7119), .B2(n7652), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8315 ( .A1(n7658), .A2(n7376), .B1(n6966), .B2(n7656), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8316 ( .A1(n3131), .A2(n7377), .B1(n6967), .B2(n7660), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8317 ( .A1(n3128), .A2(n7375), .B1(n7118), .B2(n7664), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8318 ( .A1(n7670), .A2(n7376), .B1(n6987), .B2(n7668), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8319 ( .A1(n7675), .A2(n7375), .B1(n6587), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8320 ( .A1(n7679), .A2(n7375), .B1(n6385), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8321 ( .A1(n7683), .A2(n7375), .B1(n6386), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8322 ( .A1(n7687), .A2(n7377), .B1(n6586), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8323 ( .A1(n7690), .A2(n7375), .B1(n6672), .B2(n7688), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8324 ( .A1(n7694), .A2(n7377), .B1(n6430), .B2(n7692), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8325 ( .A1(n7698), .A2(n7375), .B1(n6166), .B2(n7696), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8326 ( .A1(n7702), .A2(n7376), .B1(n6750), .B2(n7700), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8327 ( .A1(n7706), .A2(n7375), .B1(n6222), .B2(n7704), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8328 ( .A1(n7710), .A2(n7376), .B1(n5937), .B2(n7708), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8329 ( .A1(n7714), .A2(n7376), .B1(n6302), .B2(n7712), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8330 ( .A1(n7718), .A2(n7377), .B1(n6514), .B2(n7716), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8331 ( .A1(n7723), .A2(n7375), .B1(n6718), .B2(n7720), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8332 ( .A1(n7727), .A2(n7377), .B1(n7091), .B2(n7725), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8333 ( .A1(n7732), .A2(n7377), .B1(n6588), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8334 ( .A1(n7736), .A2(n7377), .B1(n6454), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8335 ( .A1(n7739), .A2(n7375), .B1(n6719), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8336 ( .A1(n7744), .A2(n7376), .B1(n6546), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8337 ( .A1(n3078), .A2(n7377), .B1(n7121), .B2(n7745), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8338 ( .A1(n7760), .A2(n7377), .B1(n6431), .B2(n7761), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U8339 ( .A1(ID_EXEC_OUT[158]), .A2(n7307), .ZN(n9823) );
  NAND2_X2 U8340 ( .A1(n5665), .A2(n9823), .ZN(n9197) );
  NAND4_X2 U8341 ( .A1(n8420), .A2(RegWrite_wb_out), .A3(n8419), .A4(n8418), 
        .ZN(n8421) );
  INV_X4 U8342 ( .A(n8421), .ZN(n8434) );
  NAND2_X2 U8343 ( .A1(n7471), .A2(n8423), .ZN(n8424) );
  NAND3_X4 U8344 ( .A1(n8426), .A2(n8425), .A3(n8424), .ZN(n9915) );
  XNOR2_X2 U8345 ( .A(n9915), .B(n7449), .ZN(n9078) );
  NAND3_X2 U8346 ( .A1(ID_EXEC_OUT[89]), .A2(n7381), .A3(n7469), .ZN(n8428) );
  NAND2_X2 U8347 ( .A1(n7471), .A2(n8604), .ZN(n8427) );
  NAND3_X4 U8348 ( .A1(n8429), .A2(n8428), .A3(n8427), .ZN(n9855) );
  XNOR2_X2 U8349 ( .A(n9855), .B(n7449), .ZN(n8488) );
  XNOR2_X2 U8350 ( .A(n8488), .B(n9853), .ZN(n8953) );
  XNOR2_X2 U8351 ( .A(n9863), .B(n7449), .ZN(n8433) );
  NAND3_X2 U8352 ( .A1(DMEM_BUS_OUT[30]), .A2(n7380), .A3(n7468), .ZN(n8432)
         );
  NAND3_X2 U8353 ( .A1(ID_EXEC_OUT[94]), .A2(n8493), .A3(n7469), .ZN(n8431) );
  NAND2_X2 U8354 ( .A1(n7471), .A2(n8909), .ZN(n8430) );
  NAND3_X4 U8355 ( .A1(n8432), .A2(n8431), .A3(n8430), .ZN(n9807) );
  XNOR2_X2 U8356 ( .A(n8433), .B(n7383), .ZN(n9057) );
  NAND2_X2 U8357 ( .A1(n7471), .A2(n8948), .ZN(n8437) );
  NAND3_X4 U8358 ( .A1(n8437), .A2(n8436), .A3(n8435), .ZN(n9786) );
  NOR2_X4 U8359 ( .A1(n8439), .A2(n8438), .ZN(n8442) );
  XNOR2_X2 U8360 ( .A(n9807), .B(n7449), .ZN(n8440) );
  OAI21_X4 U8361 ( .B1(n9057), .B2(n8442), .A(n8441), .ZN(n8649) );
  NAND3_X2 U8362 ( .A1(DMEM_BUS_OUT[29]), .A2(n8492), .A3(n7469), .ZN(n8445)
         );
  NAND3_X2 U8363 ( .A1(ID_EXEC_OUT[93]), .A2(n7381), .A3(n7469), .ZN(n8444) );
  NAND2_X2 U8364 ( .A1(n7471), .A2(n8907), .ZN(n8443) );
  NAND3_X4 U8365 ( .A1(n8445), .A2(n8444), .A3(n8443), .ZN(n9871) );
  NAND2_X2 U8366 ( .A1(n7471), .A2(n8902), .ZN(n8448) );
  NAND2_X2 U8367 ( .A1(n8450), .A2(n7469), .ZN(n8453) );
  NAND2_X2 U8368 ( .A1(n8448), .A2(n8453), .ZN(n9849) );
  XNOR2_X2 U8369 ( .A(n9849), .B(n7449), .ZN(n8449) );
  NAND2_X2 U8370 ( .A1(n8449), .A2(n9850), .ZN(n8489) );
  XNOR2_X2 U8371 ( .A(n7450), .B(n8902), .ZN(n8454) );
  INV_X4 U8372 ( .A(n8450), .ZN(n8451) );
  OAI221_X2 U8373 ( .B1(n8454), .B2(n7468), .C1(n7450), .C2(n8453), .A(n8452), 
        .ZN(n8455) );
  XNOR2_X2 U8374 ( .A(n8455), .B(n9850), .ZN(n8456) );
  INV_X4 U8375 ( .A(n8456), .ZN(n8993) );
  NAND3_X2 U8376 ( .A1(DMEM_BUS_OUT[23]), .A2(n7380), .A3(n7384), .ZN(n8459)
         );
  NAND3_X2 U8377 ( .A1(ID_EXEC_OUT[87]), .A2(n8493), .A3(n7384), .ZN(n8458) );
  NAND3_X4 U8378 ( .A1(n8459), .A2(n8458), .A3(n8457), .ZN(n9886) );
  XNOR2_X2 U8379 ( .A(n9886), .B(n7307), .ZN(n8461) );
  XNOR2_X2 U8380 ( .A(n8461), .B(n9887), .ZN(n8961) );
  INV_X4 U8381 ( .A(n8961), .ZN(n8460) );
  OAI21_X4 U8382 ( .B1(n8960), .B2(n8993), .A(n8460), .ZN(n9561) );
  NAND3_X2 U8383 ( .A1(ID_EXEC_OUT[86]), .A2(n7381), .A3(n7469), .ZN(n8463) );
  NAND2_X2 U8384 ( .A1(n7471), .A2(n8891), .ZN(n8462) );
  NAND3_X4 U8385 ( .A1(n8464), .A2(n8463), .A3(n8462), .ZN(n9888) );
  XNOR2_X2 U8386 ( .A(n9888), .B(n7449), .ZN(n8487) );
  XNOR2_X2 U8387 ( .A(n8487), .B(n9889), .ZN(n9568) );
  INV_X4 U8388 ( .A(n8466), .ZN(n8491) );
  NAND2_X2 U8389 ( .A1(n7470), .A2(n8724), .ZN(n8469) );
  NAND3_X4 U8390 ( .A1(DMEM_BUS_OUT[27]), .A2(n7384), .A3(n7380), .ZN(n8467)
         );
  NAND3_X4 U8391 ( .A1(n8469), .A2(n8468), .A3(n8467), .ZN(n8738) );
  XNOR2_X2 U8392 ( .A(n8738), .B(n7307), .ZN(n8470) );
  XNOR2_X2 U8393 ( .A(n8470), .B(n9843), .ZN(n8678) );
  NAND2_X2 U8394 ( .A1(n8470), .A2(n9843), .ZN(n8679) );
  NAND2_X2 U8395 ( .A1(n8678), .A2(n8679), .ZN(n8957) );
  NAND3_X2 U8396 ( .A1(DMEM_BUS_OUT[26]), .A2(n7380), .A3(n7469), .ZN(n8473)
         );
  NAND2_X2 U8397 ( .A1(n7471), .A2(n8676), .ZN(n8471) );
  XNOR2_X2 U8398 ( .A(n8682), .B(n7449), .ZN(n8481) );
  XNOR2_X2 U8399 ( .A(n8481), .B(n9894), .ZN(n8955) );
  INV_X4 U8400 ( .A(n8955), .ZN(n8681) );
  INV_X4 U8401 ( .A(n8650), .ZN(n8478) );
  XNOR2_X2 U8402 ( .A(n9668), .B(n7307), .ZN(n8474) );
  XNOR2_X2 U8403 ( .A(n8474), .B(n9871), .ZN(n9044) );
  INV_X4 U8404 ( .A(n9044), .ZN(n8648) );
  NAND3_X2 U8405 ( .A1(ID_EXEC_OUT[92]), .A2(n8493), .A3(n7469), .ZN(n8476) );
  NAND3_X4 U8406 ( .A1(n8477), .A2(n8476), .A3(n8475), .ZN(n9876) );
  XNOR2_X2 U8407 ( .A(n9876), .B(n7449), .ZN(n8482) );
  NOR2_X4 U8408 ( .A1(n8653), .A2(n8954), .ZN(n8479) );
  NAND3_X4 U8409 ( .A1(n8480), .A2(n8491), .A3(n8479), .ZN(n9498) );
  NAND2_X2 U8410 ( .A1(n8481), .A2(n9894), .ZN(n8651) );
  NAND3_X2 U8411 ( .A1(n8678), .A2(n8651), .A3(n8679), .ZN(n8486) );
  NAND2_X2 U8412 ( .A1(n8955), .A2(n8651), .ZN(n8484) );
  NAND2_X2 U8413 ( .A1(n7343), .A2(n9889), .ZN(n9093) );
  NAND2_X2 U8414 ( .A1(n7226), .A2(n9564), .ZN(n8490) );
  NAND2_X2 U8415 ( .A1(n9093), .A2(n9090), .ZN(n9501) );
  INV_X4 U8416 ( .A(n9501), .ZN(n9526) );
  NAND3_X2 U8417 ( .A1(DMEM_BUS_OUT[21]), .A2(n7380), .A3(n7384), .ZN(n8496)
         );
  NAND2_X2 U8418 ( .A1(n7471), .A2(n8888), .ZN(n8494) );
  NAND3_X4 U8419 ( .A1(n8496), .A2(n8495), .A3(n8494), .ZN(n9911) );
  XNOR2_X2 U8420 ( .A(n9911), .B(n7449), .ZN(n8497) );
  NAND2_X2 U8421 ( .A1(n8497), .A2(n9912), .ZN(n9496) );
  NAND2_X2 U8422 ( .A1(n9526), .A2(n9496), .ZN(n9331) );
  INV_X4 U8423 ( .A(n9496), .ZN(n9611) );
  XNOR2_X2 U8424 ( .A(n8497), .B(n9912), .ZN(n9527) );
  INV_X4 U8425 ( .A(n9527), .ZN(n9612) );
  NAND3_X2 U8426 ( .A1(DMEM_BUS_OUT[20]), .A2(n8492), .A3(n7469), .ZN(n8500)
         );
  NAND3_X2 U8427 ( .A1(ID_EXEC_OUT[84]), .A2(n7381), .A3(n7469), .ZN(n8499) );
  NAND2_X2 U8428 ( .A1(n7471), .A2(n8886), .ZN(n8498) );
  NAND3_X4 U8429 ( .A1(n8500), .A2(n8499), .A3(n8498), .ZN(n9908) );
  XNOR2_X2 U8430 ( .A(n9908), .B(n7449), .ZN(n8502) );
  XNOR2_X2 U8431 ( .A(n8502), .B(n9909), .ZN(n9614) );
  INV_X4 U8432 ( .A(n9614), .ZN(n8501) );
  OAI21_X4 U8433 ( .B1(n9611), .B2(n9612), .A(n8501), .ZN(n9075) );
  XNOR2_X2 U8434 ( .A(n6990), .B(n8504), .ZN(n8548) );
  INV_X4 U8435 ( .A(n8738), .ZN(n9844) );
  INV_X4 U8436 ( .A(n9876), .ZN(n9764) );
  NAND2_X2 U8437 ( .A1(n7473), .A2(n9912), .ZN(n8606) );
  NAND2_X2 U8438 ( .A1(n8506), .A2(n8606), .ZN(n9591) );
  NAND2_X2 U8439 ( .A1(n5864), .A2(n9591), .ZN(n8512) );
  INV_X4 U8440 ( .A(n8971), .ZN(n8967) );
  NAND2_X2 U8441 ( .A1(n7001), .A2(n9853), .ZN(n8511) );
  NAND2_X2 U8442 ( .A1(n7475), .A2(n9843), .ZN(n8507) );
  NAND2_X2 U8443 ( .A1(n8507), .A2(n8531), .ZN(n10238) );
  NAND2_X2 U8444 ( .A1(n8627), .A2(n10238), .ZN(n8510) );
  NAND2_X2 U8445 ( .A1(n7475), .A2(n7366), .ZN(n8508) );
  NAND2_X2 U8446 ( .A1(n8508), .A2(n8613), .ZN(n9544) );
  NAND2_X2 U8447 ( .A1(n7478), .A2(n9544), .ZN(n8509) );
  INV_X4 U8448 ( .A(n9786), .ZN(n9862) );
  NAND2_X2 U8449 ( .A1(n7450), .A2(n6013), .ZN(n10086) );
  NAND2_X2 U8450 ( .A1(n10086), .A2(n9823), .ZN(n9819) );
  NAND2_X2 U8451 ( .A1(ID_EXEC_OUT[156]), .A2(n9819), .ZN(n8515) );
  NAND2_X2 U8452 ( .A1(n7450), .A2(ID_EXEC_OUT[158]), .ZN(n9838) );
  INV_X4 U8453 ( .A(n9838), .ZN(n8513) );
  NAND2_X2 U8454 ( .A1(n8513), .A2(n6863), .ZN(n8514) );
  MUX2_X2 U8455 ( .A(n8515), .B(n8514), .S(ID_EXEC_OUT[157]), .Z(n8516) );
  INV_X4 U8456 ( .A(n8516), .ZN(n9173) );
  INV_X4 U8457 ( .A(n9742), .ZN(n10272) );
  XNOR2_X2 U8458 ( .A(n9915), .B(n9916), .ZN(n9780) );
  INV_X4 U8459 ( .A(n9780), .ZN(n9937) );
  NAND2_X2 U8460 ( .A1(n10272), .A2(n9937), .ZN(n8517) );
  NAND2_X2 U8461 ( .A1(ID_EXEC_OUT[157]), .A2(n9318), .ZN(n9417) );
  INV_X4 U8462 ( .A(n9417), .ZN(n9412) );
  NAND2_X2 U8463 ( .A1(n9412), .A2(n8738), .ZN(n9596) );
  NAND2_X2 U8464 ( .A1(n5851), .A2(n9974), .ZN(n8518) );
  NAND2_X2 U8465 ( .A1(n7475), .A2(n9964), .ZN(n8519) );
  AOI22_X2 U8466 ( .A1(n7478), .A2(n9599), .B1(n10248), .B2(n10250), .ZN(n8528) );
  NAND2_X2 U8467 ( .A1(n7390), .A2(n7351), .ZN(n8523) );
  NAND2_X2 U8468 ( .A1(n9189), .A2(n9412), .ZN(n8637) );
  NAND2_X2 U8469 ( .A1(n7473), .A2(n9919), .ZN(n9125) );
  INV_X4 U8470 ( .A(n9125), .ZN(n8521) );
  NAND2_X2 U8471 ( .A1(n9588), .A2(n10163), .ZN(n9177) );
  INV_X4 U8472 ( .A(n9177), .ZN(n8520) );
  INV_X4 U8473 ( .A(n8977), .ZN(n9539) );
  NAND2_X2 U8474 ( .A1(n7390), .A2(n9318), .ZN(n8524) );
  INV_X4 U8475 ( .A(n9120), .ZN(n9538) );
  NAND2_X2 U8476 ( .A1(n7473), .A2(n9925), .ZN(n9590) );
  NAND2_X2 U8477 ( .A1(n7475), .A2(n9977), .ZN(n8529) );
  AOI22_X2 U8478 ( .A1(n7478), .A2(n9529), .B1(n10195), .B2(n10107), .ZN(n8540) );
  NAND2_X2 U8479 ( .A1(n5852), .A2(n9989), .ZN(n9154) );
  NAND2_X2 U8480 ( .A1(n7473), .A2(n9930), .ZN(n9112) );
  INV_X4 U8481 ( .A(n9112), .ZN(n8534) );
  INV_X4 U8482 ( .A(n9340), .ZN(n9532) );
  NAND2_X2 U8483 ( .A1(n9618), .A2(n9173), .ZN(n9646) );
  INV_X4 U8484 ( .A(n9646), .ZN(n10277) );
  NAND2_X2 U8485 ( .A1(n7473), .A2(n9889), .ZN(n8633) );
  NAND2_X2 U8486 ( .A1(n8541), .A2(n8633), .ZN(n9550) );
  INV_X4 U8487 ( .A(n9550), .ZN(n8543) );
  NAND2_X2 U8488 ( .A1(n7473), .A2(n9909), .ZN(n8628) );
  NAND2_X2 U8489 ( .A1(n7001), .A2(n9894), .ZN(n8542) );
  OAI221_X2 U8490 ( .B1(n8543), .B2(n7386), .C1(n9346), .C2(n7383), .A(n8542), 
        .ZN(n9616) );
  NAND2_X2 U8491 ( .A1(n10277), .A2(n9616), .ZN(n8544) );
  OAI221_X2 U8492 ( .B1(n6805), .B2(n10281), .C1(n7230), .C2(n10279), .A(n8544), .ZN(n8545) );
  OAI221_X2 U8493 ( .B1(n9155), .B2(n8549), .C1(n8548), .C2(n7479), .A(n8547), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N94) );
  NAND3_X2 U8494 ( .A1(n8551), .A2(n8550), .A3(n6892), .ZN(n8553) );
  NAND2_X2 U8495 ( .A1(n8759), .A2(n8555), .ZN(n8557) );
  NAND2_X2 U8496 ( .A1(n7372), .A2(n9909), .ZN(n8556) );
  INV_X4 U8497 ( .A(n8559), .ZN(n8567) );
  INV_X4 U8498 ( .A(n8560), .ZN(n8562) );
  NAND4_X2 U8499 ( .A1(n8565), .A2(n8564), .A3(n8581), .A4(n8563), .ZN(n8566)
         );
  NAND2_X2 U8500 ( .A1(n8574), .A2(n6036), .ZN(n8573) );
  NAND2_X2 U8501 ( .A1(n8573), .A2(n8569), .ZN(n8570) );
  XNOR2_X2 U8502 ( .A(n6520), .B(n8570), .ZN(n8572) );
  NAND2_X2 U8503 ( .A1(n7370), .A2(n9912), .ZN(n8571) );
  OAI211_X2 U8504 ( .C1(n8574), .C2(n6036), .A(n8573), .B(n8759), .ZN(n8576)
         );
  NAND2_X2 U8505 ( .A1(n7370), .A2(n9889), .ZN(n8575) );
  NAND2_X2 U8506 ( .A1(n8576), .A2(n8575), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N51)
         );
  XNOR2_X2 U8507 ( .A(n6999), .B(n8577), .ZN(n8579) );
  INV_X4 U8508 ( .A(n8580), .ZN(n8584) );
  INV_X4 U8509 ( .A(n8585), .ZN(n8582) );
  NAND2_X2 U8510 ( .A1(n8591), .A2(n8590), .ZN(n8663) );
  NAND2_X2 U8511 ( .A1(n8663), .A2(n8662), .ZN(n8664) );
  NAND2_X2 U8512 ( .A1(n8592), .A2(n8664), .ZN(n8593) );
  XNOR2_X2 U8513 ( .A(n7037), .B(n8593), .ZN(n8595) );
  NAND2_X2 U8514 ( .A1(n7373), .A2(n9853), .ZN(n8594) );
  NAND2_X2 U8515 ( .A1(n1602), .A2(n7448), .ZN(n8597) );
  NAND2_X2 U8516 ( .A1(n7368), .A2(n8604), .ZN(n8596) );
  NAND2_X2 U8517 ( .A1(n8597), .A2(n8596), .ZN(n8598) );
  NAND4_X2 U8518 ( .A1(n3935), .A2(n3936), .A3(n3934), .A4(n8599), .ZN(
        ID_EX_REG_ID_EX_REG_N149) );
  NAND2_X2 U8519 ( .A1(n8604), .A2(n7457), .ZN(n8601) );
  NAND2_X2 U8520 ( .A1(n7458), .A2(n6831), .ZN(n8600) );
  NAND3_X2 U8521 ( .A1(n4676), .A2(n8601), .A3(n8600), .ZN(n8603) );
  INV_X4 U8522 ( .A(n8603), .ZN(n8602) );
  OAI22_X2 U8523 ( .A1(n7445), .A2(n8602), .B1(n4673), .B2(n1588), .ZN(
        ID_EX_REG_ID_EX_REG_N117) );
  AND2_X2 U8524 ( .A1(n8603), .A2(n7305), .ZN(ID_EX_REG_ID_EX_REG_N21) );
  OAI22_X2 U8525 ( .A1(n7082), .A2(n7625), .B1(n7626), .B2(n7394), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8526 ( .A1(n3148), .A2(n7394), .B1(n6161), .B2(n7628), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8527 ( .A1(n3146), .A2(n7395), .B1(n7179), .B2(n7632), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8528 ( .A1(n7639), .A2(n7396), .B1(n6582), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8529 ( .A1(n7643), .A2(n7394), .B1(n6064), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8530 ( .A1(n7647), .A2(n7394), .B1(n7020), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8531 ( .A1(n7651), .A2(n7395), .B1(n7140), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8532 ( .A1(n7081), .A2(n7653), .B1(n7654), .B2(n7396), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8533 ( .A1(n6054), .A2(n7657), .B1(n7658), .B2(n7396), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8534 ( .A1(n3131), .A2(n7394), .B1(n6963), .B2(n7660), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8535 ( .A1(n3128), .A2(n7396), .B1(n7112), .B2(n7664), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8536 ( .A1(n6125), .A2(n7669), .B1(n7670), .B2(n7396), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8537 ( .A1(n7675), .A2(n7394), .B1(n6580), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8538 ( .A1(n7679), .A2(n7395), .B1(n6380), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8539 ( .A1(n7683), .A2(n7394), .B1(n6381), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8540 ( .A1(n7687), .A2(n7396), .B1(n6579), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8541 ( .A1(n7690), .A2(n7396), .B1(n7113), .B2(n7688), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8542 ( .A1(n7694), .A2(n7395), .B1(n6103), .B2(n7692), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8543 ( .A1(n3110), .A2(n7394), .B1(n5963), .B2(n7696), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8544 ( .A1(n3107), .A2(n7396), .B1(n7180), .B2(n7700), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8545 ( .A1(n3105), .A2(n7395), .B1(n6212), .B2(n7704), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8546 ( .A1(n3103), .A2(n7396), .B1(n5895), .B2(n7708), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8547 ( .A1(n3101), .A2(n7394), .B1(n7181), .B2(n7712), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8548 ( .A1(n3099), .A2(n7395), .B1(n7019), .B2(n7716), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8549 ( .A1(n7722), .A2(n7395), .B1(n6720), .B2(n7720), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8550 ( .A1(n3093), .A2(n7395), .B1(n6244), .B2(n7725), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8551 ( .A1(n7732), .A2(n7394), .B1(n6581), .B2(n7730), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8552 ( .A1(n7736), .A2(n7395), .B1(n6452), .B2(n7734), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8553 ( .A1(n7739), .A2(n7394), .B1(n6721), .B2(n7738), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8554 ( .A1(n7744), .A2(n7396), .B1(n6547), .B2(n7742), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8555 ( .A1(n3078), .A2(n7394), .B1(n7114), .B2(n7745), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8556 ( .A1(n7760), .A2(n7395), .B1(n6412), .B2(n7761), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U8557 ( .A1(n7379), .A2(n9173), .ZN(n10155) );
  NAND4_X2 U8558 ( .A1(n8637), .A2(n8606), .A3(n9163), .A4(n8605), .ZN(n9530)
         );
  INV_X4 U8559 ( .A(n9530), .ZN(n8982) );
  NAND2_X2 U8560 ( .A1(n5851), .A2(n9930), .ZN(n9370) );
  NAND2_X2 U8561 ( .A1(n7473), .A2(n9853), .ZN(n8608) );
  NAND2_X2 U8562 ( .A1(n7390), .A2(n10135), .ZN(n8607) );
  NAND4_X2 U8563 ( .A1(n8609), .A2(n9370), .A3(n8608), .A4(n8607), .ZN(n8610)
         );
  INV_X4 U8564 ( .A(n8610), .ZN(n9032) );
  NAND2_X2 U8565 ( .A1(n7390), .A2(n9977), .ZN(n8617) );
  INV_X4 U8566 ( .A(n8613), .ZN(n8615) );
  NAND2_X2 U8567 ( .A1(n7476), .A2(n9925), .ZN(n9153) );
  INV_X4 U8568 ( .A(n9153), .ZN(n8614) );
  INV_X4 U8569 ( .A(n9036), .ZN(n8983) );
  NAND2_X2 U8570 ( .A1(n8621), .A2(n8620), .ZN(n8684) );
  NAND2_X2 U8571 ( .A1(n6800), .A2(n8684), .ZN(n8645) );
  NAND2_X2 U8572 ( .A1(n9180), .A2(n9361), .ZN(n9182) );
  INV_X4 U8573 ( .A(n8972), .ZN(n8623) );
  NAND2_X2 U8574 ( .A1(n8976), .A2(n7473), .ZN(n9024) );
  INV_X4 U8575 ( .A(n9024), .ZN(n8699) );
  NAND2_X2 U8576 ( .A1(n8685), .A2(n9618), .ZN(n8644) );
  INV_X4 U8577 ( .A(n7388), .ZN(n8627) );
  NAND2_X2 U8578 ( .A1(n7390), .A2(n9979), .ZN(n8626) );
  NAND2_X2 U8579 ( .A1(n9189), .A2(n9318), .ZN(n8625) );
  NAND2_X2 U8580 ( .A1(n9588), .A2(n9927), .ZN(n9363) );
  NAND4_X2 U8581 ( .A1(n8626), .A2(n8625), .A3(n9363), .A4(n8624), .ZN(n9018)
         );
  NAND2_X2 U8582 ( .A1(n8627), .A2(n9018), .ZN(n8641) );
  NAND2_X2 U8583 ( .A1(n7390), .A2(n9964), .ZN(n8632) );
  INV_X4 U8584 ( .A(n8628), .ZN(n8630) );
  INV_X4 U8585 ( .A(n9186), .ZN(n8629) );
  NAND2_X2 U8586 ( .A1(n7478), .A2(n9537), .ZN(n8640) );
  INV_X4 U8587 ( .A(n8633), .ZN(n8635) );
  INV_X4 U8588 ( .A(n9974), .ZN(n9665) );
  NAND2_X2 U8589 ( .A1(n8976), .A2(n9021), .ZN(n8639) );
  NAND2_X2 U8590 ( .A1(n10195), .A2(n8977), .ZN(n8638) );
  NAND4_X2 U8591 ( .A1(n8641), .A2(n8640), .A3(n8639), .A4(n8638), .ZN(n8995)
         );
  NAND2_X2 U8592 ( .A1(n6799), .A2(n8995), .ZN(n8643) );
  INV_X4 U8593 ( .A(n9843), .ZN(n9156) );
  OAI22_X2 U8594 ( .A1(n7365), .A2(n8971), .B1(n9156), .B2(n9182), .ZN(n8698)
         );
  INV_X4 U8595 ( .A(n9853), .ZN(n9147) );
  OAI22_X2 U8596 ( .A1(n9872), .A2(n8971), .B1(n9147), .B2(n9182), .ZN(n8966)
         );
  MUX2_X2 U8597 ( .A(n8698), .B(n8966), .S(n9864), .Z(n8994) );
  NAND2_X2 U8598 ( .A1(n9753), .A2(n8994), .ZN(n8642) );
  NAND4_X2 U8599 ( .A1(n8645), .A2(n8644), .A3(n8643), .A4(n8642), .ZN(n8646)
         );
  NAND2_X2 U8600 ( .A1(n10257), .A2(n8646), .ZN(n8661) );
  NAND2_X2 U8601 ( .A1(n8647), .A2(n9853), .ZN(n8660) );
  INV_X4 U8602 ( .A(n6861), .ZN(n9143) );
  XNOR2_X2 U8603 ( .A(n9855), .B(n9853), .ZN(n9859) );
  INV_X4 U8604 ( .A(n9859), .ZN(n9772) );
  NAND2_X2 U8605 ( .A1(n9143), .A2(n9772), .ZN(n8659) );
  NAND2_X2 U8606 ( .A1(n9047), .A2(n8650), .ZN(n9763) );
  NAND2_X2 U8607 ( .A1(n9763), .A2(n6895), .ZN(n9761) );
  INV_X4 U8608 ( .A(n8952), .ZN(n8652) );
  INV_X4 U8609 ( .A(n8654), .ZN(n8655) );
  NAND2_X2 U8610 ( .A1(n8657), .A2(n8656), .ZN(n8658) );
  NAND4_X2 U8611 ( .A1(n8661), .A2(n8660), .A3(n8659), .A4(n8658), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N88) );
  NAND2_X2 U8612 ( .A1(n8759), .A2(n8664), .ZN(n8666) );
  NAND2_X2 U8613 ( .A1(n7373), .A2(n9894), .ZN(n8665) );
  NAND2_X2 U8614 ( .A1(n1601), .A2(n7448), .ZN(n8669) );
  NAND2_X2 U8615 ( .A1(n7367), .A2(n8676), .ZN(n8668) );
  NAND2_X2 U8616 ( .A1(n8669), .A2(n8668), .ZN(n8670) );
  NAND4_X2 U8617 ( .A1(n3956), .A2(n3957), .A3(n3955), .A4(n8671), .ZN(
        ID_EX_REG_ID_EX_REG_N148) );
  NAND2_X2 U8618 ( .A1(n8676), .A2(n7457), .ZN(n8673) );
  NAND2_X2 U8619 ( .A1(n7459), .A2(n7247), .ZN(n8672) );
  NAND3_X2 U8620 ( .A1(n4699), .A2(n8673), .A3(n8672), .ZN(n8675) );
  INV_X4 U8621 ( .A(n8675), .ZN(n8674) );
  OAI22_X2 U8622 ( .A1(n7445), .A2(n8674), .B1(n4696), .B2(n1588), .ZN(
        ID_EX_REG_ID_EX_REG_N116) );
  AND2_X2 U8623 ( .A1(n8675), .A2(n7305), .ZN(ID_EX_REG_ID_EX_REG_N20) );
  OAI22_X2 U8624 ( .A1(n7080), .A2(n7625), .B1(n7626), .B2(n7399), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8625 ( .A1(n7630), .A2(n7398), .B1(n6495), .B2(n7628), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8626 ( .A1(n7634), .A2(n7397), .B1(n6751), .B2(n7632), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8627 ( .A1(n7639), .A2(n7398), .B1(n7052), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8628 ( .A1(n7643), .A2(n7399), .B1(n6063), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8629 ( .A1(n7647), .A2(n7398), .B1(n7018), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8630 ( .A1(n7651), .A2(n7397), .B1(n7141), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8631 ( .A1(n7079), .A2(n7653), .B1(n7654), .B2(n7398), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8632 ( .A1(n5933), .A2(n7657), .B1(n7658), .B2(n7398), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8633 ( .A1(n7662), .A2(n7399), .B1(n6410), .B2(n7660), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8634 ( .A1(n7666), .A2(n7397), .B1(n6648), .B2(n7664), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8635 ( .A1(n6981), .A2(n7669), .B1(n7670), .B2(n7399), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8636 ( .A1(n7675), .A2(n7398), .B1(n6577), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8637 ( .A1(n7679), .A2(n7397), .B1(n6925), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8638 ( .A1(n7683), .A2(n7399), .B1(n6926), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8639 ( .A1(n7687), .A2(n7397), .B1(n7051), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8640 ( .A1(n7690), .A2(n7398), .B1(n7111), .B2(n7688), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8641 ( .A1(n7694), .A2(n7399), .B1(n5896), .B2(n7692), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8642 ( .A1(n3110), .A2(n7397), .B1(n6160), .B2(n7696), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8643 ( .A1(n3107), .A2(n7397), .B1(n7182), .B2(n7700), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8644 ( .A1(n3105), .A2(n7398), .B1(n6211), .B2(n7704), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8645 ( .A1(n3103), .A2(n7399), .B1(n5875), .B2(n7708), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8646 ( .A1(n7714), .A2(n7398), .B1(n6752), .B2(n7712), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8647 ( .A1(n3099), .A2(n7397), .B1(n7017), .B2(n7716), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8648 ( .A1(n7723), .A2(n7398), .B1(n6722), .B2(n7720), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8649 ( .A1(n7727), .A2(n7399), .B1(n6608), .B2(n7725), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8650 ( .A1(n7732), .A2(n7398), .B1(n6578), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8651 ( .A1(n7736), .A2(n7397), .B1(n6451), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8652 ( .A1(n7739), .A2(n7399), .B1(n6723), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8653 ( .A1(n7744), .A2(n7399), .B1(n6548), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8654 ( .A1(n7747), .A2(n7398), .B1(n6649), .B2(n7745), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8655 ( .A1(n7760), .A2(n7397), .B1(n6411), .B2(n7761), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  INV_X4 U8656 ( .A(n8682), .ZN(n9895) );
  XNOR2_X2 U8657 ( .A(n9179), .B(n9895), .ZN(n9842) );
  NAND2_X2 U8658 ( .A1(n9761), .A2(n8677), .ZN(n8741) );
  INV_X4 U8659 ( .A(n8678), .ZN(n8742) );
  NAND2_X2 U8660 ( .A1(n8741), .A2(n8742), .ZN(n8740) );
  NAND2_X2 U8661 ( .A1(n8740), .A2(n8679), .ZN(n8680) );
  XNOR2_X2 U8662 ( .A(n8681), .B(n8680), .ZN(n8709) );
  INV_X4 U8663 ( .A(n8684), .ZN(n8687) );
  NAND2_X2 U8664 ( .A1(n9753), .A2(n8685), .ZN(n8686) );
  INV_X4 U8665 ( .A(n9021), .ZN(n8689) );
  INV_X4 U8666 ( .A(n9018), .ZN(n8688) );
  OAI22_X2 U8667 ( .A1(n7389), .A2(n8689), .B1(n7385), .B2(n8688), .ZN(n8697)
         );
  NAND2_X2 U8668 ( .A1(n9189), .A2(n7351), .ZN(n8692) );
  NAND2_X2 U8669 ( .A1(n7476), .A2(n9919), .ZN(n9364) );
  NAND2_X2 U8670 ( .A1(n7473), .A2(n9894), .ZN(n8691) );
  NAND2_X2 U8671 ( .A1(n7390), .A2(n10163), .ZN(n8690) );
  NAND4_X2 U8672 ( .A1(n8692), .A2(n9364), .A3(n8691), .A4(n8690), .ZN(n9059)
         );
  INV_X4 U8673 ( .A(n9059), .ZN(n8693) );
  INV_X4 U8674 ( .A(n9537), .ZN(n8694) );
  INV_X4 U8675 ( .A(n8698), .ZN(n8701) );
  NAND2_X2 U8676 ( .A1(n9618), .A2(n8725), .ZN(n8702) );
  NOR2_X4 U8677 ( .A1(n8704), .A2(n8703), .ZN(n8705) );
  OAI221_X2 U8678 ( .B1(n9842), .B2(n6861), .C1(n8709), .C2(n7479), .A(n8708), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N87) );
  NAND2_X2 U8679 ( .A1(n8748), .A2(n6037), .ZN(n8747) );
  NAND2_X2 U8680 ( .A1(n8747), .A2(n8712), .ZN(n8713) );
  XNOR2_X2 U8681 ( .A(n6521), .B(n8713), .ZN(n8715) );
  NAND2_X2 U8682 ( .A1(n7372), .A2(n9843), .ZN(n8714) );
  NAND2_X2 U8683 ( .A1(ID_EX_REG_ID_EX_REG_N99), .A2(n7448), .ZN(n8717) );
  NAND2_X2 U8684 ( .A1(n7368), .A2(n8724), .ZN(n8716) );
  NAND2_X2 U8685 ( .A1(n8717), .A2(n8716), .ZN(n8718) );
  NAND4_X2 U8686 ( .A1(n3977), .A2(n3978), .A3(n3976), .A4(n8719), .ZN(
        ID_EX_REG_ID_EX_REG_N147) );
  NAND2_X2 U8687 ( .A1(n8724), .A2(n7457), .ZN(n8721) );
  NAND2_X2 U8688 ( .A1(n7459), .A2(n7248), .ZN(n8720) );
  NAND3_X2 U8689 ( .A1(n4722), .A2(n8721), .A3(n8720), .ZN(n8723) );
  INV_X4 U8690 ( .A(n8723), .ZN(n8722) );
  OAI22_X2 U8691 ( .A1(n7445), .A2(n8722), .B1(n4719), .B2(n1591), .ZN(
        ID_EX_REG_ID_EX_REG_N115) );
  AND2_X2 U8692 ( .A1(n8723), .A2(n7305), .ZN(ID_EX_REG_ID_EX_REG_N19) );
  OAI22_X2 U8693 ( .A1(n7626), .A2(n7400), .B1(n7110), .B2(n7625), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8694 ( .A1(n7630), .A2(n7400), .B1(n6494), .B2(n7628), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8695 ( .A1(n7634), .A2(n7400), .B1(n6753), .B2(n7632), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8696 ( .A1(n7639), .A2(n7400), .B1(n7050), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8697 ( .A1(n7643), .A2(n7401), .B1(n6924), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8698 ( .A1(n7647), .A2(n7402), .B1(n7016), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8699 ( .A1(n7651), .A2(n7401), .B1(n7142), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8700 ( .A1(n7654), .A2(n7402), .B1(n7109), .B2(n7653), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8701 ( .A1(n7658), .A2(n7402), .B1(n6962), .B2(n7657), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8702 ( .A1(n7662), .A2(n7401), .B1(n6409), .B2(n7660), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8703 ( .A1(n7666), .A2(n7400), .B1(n6645), .B2(n7664), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8704 ( .A1(n7670), .A2(n7400), .B1(n6131), .B2(n7669), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8705 ( .A1(n7675), .A2(n7402), .B1(n6575), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8706 ( .A1(n7679), .A2(n7401), .B1(n5935), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8707 ( .A1(n7683), .A2(n7401), .B1(n6923), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8708 ( .A1(n7687), .A2(n7402), .B1(n7049), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8709 ( .A1(n7690), .A2(n7402), .B1(n6646), .B2(n7688), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8710 ( .A1(n7694), .A2(n7401), .B1(n5946), .B2(n7692), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8711 ( .A1(n7698), .A2(n7400), .B1(n6159), .B2(n7696), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8712 ( .A1(n7702), .A2(n7400), .B1(n6754), .B2(n7700), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8713 ( .A1(n7706), .A2(n7400), .B1(n6210), .B2(n7704), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8714 ( .A1(n7710), .A2(n7400), .B1(n5874), .B2(n7708), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8715 ( .A1(n7714), .A2(n7401), .B1(n6755), .B2(n7712), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8716 ( .A1(n7718), .A2(n7402), .B1(n6508), .B2(n7716), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8717 ( .A1(n7723), .A2(n7401), .B1(n7143), .B2(n7720), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8718 ( .A1(n7727), .A2(n7402), .B1(n6609), .B2(n7725), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8719 ( .A1(n7732), .A2(n7401), .B1(n6576), .B2(n7730), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8720 ( .A1(n7736), .A2(n7402), .B1(n5949), .B2(n7734), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8721 ( .A1(n7739), .A2(n7400), .B1(n6724), .B2(n7738), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8722 ( .A1(n7744), .A2(n7400), .B1(n6549), .B2(n7742), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8723 ( .A1(n7747), .A2(n7401), .B1(n6647), .B2(n7745), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8724 ( .A1(n7760), .A2(n7402), .B1(n5947), .B2(n7761), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  INV_X4 U8725 ( .A(n8725), .ZN(n8727) );
  OAI22_X2 U8726 ( .A1(n8727), .A2(n10255), .B1(n8726), .B2(n7392), .ZN(n8736)
         );
  NAND2_X2 U8727 ( .A1(n7387), .A2(n7473), .ZN(n9164) );
  INV_X4 U8728 ( .A(n9752), .ZN(n8734) );
  NAND2_X2 U8729 ( .A1(n7473), .A2(n9843), .ZN(n8729) );
  NAND2_X2 U8730 ( .A1(n7390), .A2(n9989), .ZN(n8728) );
  NAND4_X2 U8731 ( .A1(n8730), .A2(n9373), .A3(n8729), .A4(n8728), .ZN(n9035)
         );
  INV_X4 U8732 ( .A(n9035), .ZN(n9810) );
  OAI22_X2 U8733 ( .A1(n8982), .A2(n10246), .B1(n9810), .B2(n9806), .ZN(n8733)
         );
  OAI22_X2 U8734 ( .A1(n8734), .A2(n6860), .B1(n9755), .B2(n7393), .ZN(n8735)
         );
  NAND2_X2 U8735 ( .A1(n8737), .A2(n9843), .ZN(n8745) );
  XNOR2_X2 U8736 ( .A(n8738), .B(n9843), .ZN(n9846) );
  INV_X4 U8737 ( .A(n9846), .ZN(n8739) );
  NAND2_X2 U8738 ( .A1(n9143), .A2(n8739), .ZN(n8744) );
  OAI211_X2 U8739 ( .C1(n8742), .C2(n8741), .A(n8740), .B(n7480), .ZN(n8743)
         );
  NAND4_X2 U8740 ( .A1(n8746), .A2(n8745), .A3(n8744), .A4(n8743), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N86) );
  OAI211_X2 U8741 ( .C1(n8748), .C2(n6037), .A(n8747), .B(n8759), .ZN(n8750)
         );
  NAND2_X2 U8742 ( .A1(n8750), .A2(n8749), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N45)
         );
  XNOR2_X2 U8743 ( .A(n6998), .B(n8751), .ZN(n8753) );
  NAND2_X2 U8744 ( .A1(n8754), .A2(n8760), .ZN(n8755) );
  NAND3_X2 U8745 ( .A1(n8759), .A2(n8756), .A3(n8755), .ZN(n8757) );
  INV_X4 U8746 ( .A(n8758), .ZN(n8761) );
  OAI211_X2 U8747 ( .C1(nextPC_ex_out[31]), .C2(n8761), .A(n8760), .B(n8759), 
        .ZN(n8764) );
  NAND2_X2 U8748 ( .A1(n7370), .A2(n7366), .ZN(n8763) );
  NAND2_X2 U8749 ( .A1(n8764), .A2(n8763), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N42)
         );
  NAND2_X2 U8750 ( .A1(n8902), .A2(n7457), .ZN(n8766) );
  NAND2_X2 U8751 ( .A1(n7459), .A2(n7249), .ZN(n8765) );
  NAND3_X2 U8752 ( .A1(n4653), .A2(n8766), .A3(n8765), .ZN(n8901) );
  NAND2_X2 U8753 ( .A1(n6010), .A2(n8901), .ZN(n8768) );
  NAND2_X2 U8754 ( .A1(ID_EX_REG_ID_EX_REG_N76), .A2(n4447), .ZN(n8767) );
  NAND2_X2 U8755 ( .A1(n8768), .A2(n8767), .ZN(n1583) );
  NAND2_X2 U8756 ( .A1(ID_EX_REG_ID_EX_REG_N76), .A2(n7447), .ZN(n8770) );
  NAND2_X2 U8757 ( .A1(n7367), .A2(n8902), .ZN(n8769) );
  NAND2_X2 U8758 ( .A1(n8770), .A2(n8769), .ZN(n8771) );
  NAND4_X2 U8759 ( .A1(n3913), .A2(n3914), .A3(n3912), .A4(n8772), .ZN(
        ID_EX_REG_ID_EX_REG_N150) );
  NAND2_X2 U8760 ( .A1(n8888), .A2(n7457), .ZN(n8774) );
  NAND2_X2 U8761 ( .A1(n7459), .A2(n7250), .ZN(n8773) );
  NAND3_X2 U8762 ( .A1(n4585), .A2(n8774), .A3(n8773), .ZN(n8887) );
  NAND2_X2 U8763 ( .A1(n6010), .A2(n8887), .ZN(n8776) );
  NAND2_X2 U8764 ( .A1(ID_EX_REG_ID_EX_REG_N79), .A2(n4447), .ZN(n8775) );
  NAND2_X2 U8765 ( .A1(n8776), .A2(n8775), .ZN(n1582) );
  NAND2_X2 U8766 ( .A1(ID_EX_REG_ID_EX_REG_N79), .A2(n7448), .ZN(n8778) );
  NAND2_X2 U8767 ( .A1(n7368), .A2(n8888), .ZN(n8777) );
  NAND2_X2 U8768 ( .A1(n8778), .A2(n8777), .ZN(n8779) );
  NAND4_X2 U8769 ( .A1(n3850), .A2(n3851), .A3(n3849), .A4(n8780), .ZN(
        ID_EX_REG_ID_EX_REG_N153) );
  NAND2_X2 U8770 ( .A1(n8886), .A2(n7457), .ZN(n8782) );
  NAND2_X2 U8771 ( .A1(n7459), .A2(n7251), .ZN(n8781) );
  NAND3_X2 U8772 ( .A1(n4563), .A2(n8782), .A3(n8781), .ZN(n8885) );
  NAND2_X2 U8773 ( .A1(n6010), .A2(n8885), .ZN(n8784) );
  NAND2_X2 U8774 ( .A1(ID_EX_REG_ID_EX_REG_N80), .A2(n4447), .ZN(n8783) );
  NAND2_X2 U8775 ( .A1(n8784), .A2(n8783), .ZN(n1581) );
  NAND2_X2 U8776 ( .A1(ID_EX_REG_ID_EX_REG_N80), .A2(n7448), .ZN(n8786) );
  NAND2_X2 U8777 ( .A1(n7368), .A2(n8886), .ZN(n8785) );
  NAND2_X2 U8778 ( .A1(n8786), .A2(n8785), .ZN(n8787) );
  NAND4_X2 U8779 ( .A1(n3829), .A2(n3830), .A3(n3828), .A4(n8788), .ZN(
        ID_EX_REG_ID_EX_REG_N154) );
  NAND2_X2 U8780 ( .A1(n9086), .A2(n7457), .ZN(n8790) );
  NAND2_X2 U8781 ( .A1(n7459), .A2(n7252), .ZN(n8789) );
  NAND3_X2 U8782 ( .A1(n4496), .A2(n8790), .A3(n8789), .ZN(n8882) );
  NAND2_X2 U8783 ( .A1(n6010), .A2(n8882), .ZN(n8792) );
  NAND2_X2 U8784 ( .A1(ID_EX_REG_ID_EX_REG_N83), .A2(n4447), .ZN(n8791) );
  NAND2_X2 U8785 ( .A1(n8792), .A2(n8791), .ZN(n1579) );
  NAND2_X2 U8786 ( .A1(ID_EX_REG_ID_EX_REG_N83), .A2(n7448), .ZN(n8794) );
  NAND2_X2 U8787 ( .A1(n7368), .A2(n9086), .ZN(n8793) );
  NAND2_X2 U8788 ( .A1(n8794), .A2(n8793), .ZN(n8795) );
  NAND4_X2 U8789 ( .A1(n3766), .A2(n3767), .A3(n3765), .A4(n8796), .ZN(
        ID_EX_REG_ID_EX_REG_N157) );
  NAND2_X2 U8790 ( .A1(n7459), .A2(n7253), .ZN(n8797) );
  NAND3_X2 U8791 ( .A1(n4474), .A2(n8798), .A3(n8797), .ZN(n8881) );
  NAND2_X2 U8792 ( .A1(n6010), .A2(n8881), .ZN(n8800) );
  NAND2_X2 U8793 ( .A1(ID_EX_REG_ID_EX_REG_N84), .A2(n4447), .ZN(n8799) );
  NAND2_X2 U8794 ( .A1(n8800), .A2(n8799), .ZN(n1578) );
  NAND2_X2 U8795 ( .A1(ID_EX_REG_ID_EX_REG_N84), .A2(n7447), .ZN(n8802) );
  NAND2_X2 U8796 ( .A1(n7368), .A2(n9101), .ZN(n8801) );
  NAND2_X2 U8797 ( .A1(n8802), .A2(n8801), .ZN(n8803) );
  NAND4_X2 U8798 ( .A1(n3744), .A2(n3745), .A3(n3743), .A4(n8804), .ZN(
        ID_EX_REG_ID_EX_REG_N158) );
  NAND2_X2 U8799 ( .A1(n7448), .A2(ID_EX_REG_ID_EX_REG_N95), .ZN(n8806) );
  NAND2_X2 U8800 ( .A1(n7367), .A2(n8948), .ZN(n8805) );
  NAND2_X2 U8801 ( .A1(n8806), .A2(n8805), .ZN(n8807) );
  NAND4_X2 U8802 ( .A1(n4061), .A2(n4062), .A3(n4060), .A4(n8808), .ZN(
        ID_EX_REG_ID_EX_REG_N143) );
  NAND2_X2 U8803 ( .A1(n8909), .A2(n8947), .ZN(n8810) );
  NAND2_X2 U8804 ( .A1(n7459), .A2(n7254), .ZN(n8809) );
  NAND3_X2 U8805 ( .A1(n4788), .A2(n8810), .A3(n8809), .ZN(n8908) );
  NAND2_X2 U8806 ( .A1(n6010), .A2(n8908), .ZN(n8812) );
  NAND2_X2 U8807 ( .A1(ID_EX_REG_ID_EX_REG_N96), .A2(n4447), .ZN(n8811) );
  NAND2_X2 U8808 ( .A1(n8812), .A2(n8811), .ZN(n1585) );
  NAND2_X2 U8809 ( .A1(ID_EX_REG_ID_EX_REG_N96), .A2(n7448), .ZN(n8814) );
  NAND2_X2 U8810 ( .A1(n7368), .A2(n8909), .ZN(n8813) );
  NAND2_X2 U8811 ( .A1(n8814), .A2(n8813), .ZN(n8815) );
  NAND4_X2 U8812 ( .A1(n4040), .A2(n4041), .A3(n4039), .A4(n8816), .ZN(
        ID_EX_REG_ID_EX_REG_N144) );
  NAND2_X2 U8813 ( .A1(n7459), .A2(n7255), .ZN(n8817) );
  NAND3_X2 U8814 ( .A1(n4744), .A2(n8818), .A3(n8817), .ZN(n8903) );
  NAND2_X2 U8815 ( .A1(n6010), .A2(n8903), .ZN(n8820) );
  NAND2_X2 U8816 ( .A1(ID_EX_REG_ID_EX_REG_N98), .A2(n4447), .ZN(n8819) );
  NAND2_X2 U8817 ( .A1(n8820), .A2(n8819), .ZN(n1584) );
  NAND2_X2 U8818 ( .A1(ID_EX_REG_ID_EX_REG_N98), .A2(n7448), .ZN(n8822) );
  NAND2_X2 U8819 ( .A1(n8822), .A2(n8821), .ZN(n8823) );
  NAND4_X2 U8820 ( .A1(n3998), .A2(n3999), .A3(n3997), .A4(n8824), .ZN(
        ID_EX_REG_ID_EX_REG_N146) );
  NAND2_X2 U8821 ( .A1(n1598), .A2(n7448), .ZN(n8826) );
  NAND2_X2 U8822 ( .A1(n8826), .A2(n8825), .ZN(n8827) );
  NAND4_X2 U8823 ( .A1(n4019), .A2(n4020), .A3(n4018), .A4(n8828), .ZN(
        ID_EX_REG_ID_EX_REG_N145) );
  NAND2_X2 U8824 ( .A1(n1604), .A2(n7447), .ZN(n8830) );
  NAND2_X2 U8825 ( .A1(n8830), .A2(n8829), .ZN(n8831) );
  NAND4_X2 U8826 ( .A1(n3892), .A2(n3893), .A3(n3891), .A4(n8832), .ZN(
        ID_EX_REG_ID_EX_REG_N151) );
  NAND2_X2 U8827 ( .A1(n1605), .A2(n7448), .ZN(n8834) );
  NAND2_X2 U8828 ( .A1(n7368), .A2(n8891), .ZN(n8833) );
  NAND2_X2 U8829 ( .A1(n8834), .A2(n8833), .ZN(n8835) );
  NAND4_X2 U8830 ( .A1(n3871), .A2(n3872), .A3(n3870), .A4(n8836), .ZN(
        ID_EX_REG_ID_EX_REG_N152) );
  NAND2_X2 U8831 ( .A1(n1609), .A2(n7448), .ZN(n8838) );
  NAND2_X2 U8832 ( .A1(n7368), .A2(n9079), .ZN(n8837) );
  NAND2_X2 U8833 ( .A1(n8838), .A2(n8837), .ZN(n8839) );
  NAND4_X2 U8834 ( .A1(n3787), .A2(n3788), .A3(n3786), .A4(n8840), .ZN(
        ID_EX_REG_ID_EX_REG_N156) );
  NAND4_X2 U8835 ( .A1(n3722), .A2(n3723), .A3(n3721), .A4(n8841), .ZN(
        ID_EX_REG_ID_EX_REG_N159) );
  NAND4_X2 U8836 ( .A1(n3700), .A2(n3701), .A3(n3699), .A4(n8842), .ZN(
        ID_EX_REG_ID_EX_REG_N160) );
  INV_X4 U8837 ( .A(n8843), .ZN(n8845) );
  NAND2_X2 U8838 ( .A1(n8845), .A2(n8844), .ZN(n9269) );
  NAND4_X2 U8839 ( .A1(n3678), .A2(n3679), .A3(n3677), .A4(n8846), .ZN(
        ID_EX_REG_ID_EX_REG_N161) );
  NAND4_X2 U8840 ( .A1(n3657), .A2(n3658), .A3(n3656), .A4(n8847), .ZN(
        ID_EX_REG_ID_EX_REG_N162) );
  NAND4_X2 U8841 ( .A1(n3635), .A2(n3636), .A3(n3634), .A4(n8848), .ZN(
        ID_EX_REG_ID_EX_REG_N163) );
  NAND4_X2 U8842 ( .A1(n3614), .A2(n3615), .A3(n3613), .A4(n8849), .ZN(
        ID_EX_REG_ID_EX_REG_N164) );
  INV_X4 U8843 ( .A(n8850), .ZN(n8852) );
  NAND2_X2 U8844 ( .A1(n8852), .A2(n8851), .ZN(n8913) );
  NAND4_X2 U8845 ( .A1(n3592), .A2(n3593), .A3(n3591), .A4(n8853), .ZN(
        ID_EX_REG_ID_EX_REG_N165) );
  INV_X4 U8846 ( .A(n9239), .ZN(n8855) );
  NAND2_X2 U8847 ( .A1(n8855), .A2(n9237), .ZN(n8939) );
  NAND4_X2 U8848 ( .A1(n3571), .A2(n3572), .A3(n3570), .A4(n8856), .ZN(
        ID_EX_REG_ID_EX_REG_N166) );
  NAND2_X2 U8849 ( .A1(n7459), .A2(n7256), .ZN(n8857) );
  NAND3_X2 U8850 ( .A1(n4766), .A2(n8858), .A3(n8857), .ZN(n8905) );
  AND2_X2 U8851 ( .A1(n8905), .A2(n7305), .ZN(ID_EX_REG_ID_EX_REG_N17) );
  NAND2_X2 U8852 ( .A1(n7459), .A2(n7257), .ZN(n8859) );
  NAND3_X2 U8853 ( .A1(n4631), .A2(n8860), .A3(n8859), .ZN(n8892) );
  AND2_X2 U8854 ( .A1(n8892), .A2(n7305), .ZN(ID_EX_REG_ID_EX_REG_N23) );
  NAND2_X2 U8855 ( .A1(n8891), .A2(n7457), .ZN(n8862) );
  NAND2_X2 U8856 ( .A1(n7458), .A2(n7258), .ZN(n8861) );
  NAND3_X2 U8857 ( .A1(n4608), .A2(n8862), .A3(n8861), .ZN(n8889) );
  AND2_X2 U8858 ( .A1(n8889), .A2(n7305), .ZN(ID_EX_REG_ID_EX_REG_N24) );
  NAND2_X2 U8859 ( .A1(n9079), .A2(n7457), .ZN(n8864) );
  NAND2_X2 U8860 ( .A1(n7458), .A2(n7259), .ZN(n8863) );
  NAND3_X2 U8861 ( .A1(n4519), .A2(n8864), .A3(n8863), .ZN(n8883) );
  AND2_X2 U8862 ( .A1(n8883), .A2(n7305), .ZN(ID_EX_REG_ID_EX_REG_N28) );
  NAND2_X2 U8863 ( .A1(n7458), .A2(n7260), .ZN(n8865) );
  NAND3_X2 U8864 ( .A1(n4452), .A2(n8866), .A3(n8865), .ZN(n8899) );
  AND2_X2 U8865 ( .A1(n8899), .A2(n7305), .ZN(ID_EX_REG_ID_EX_REG_N31) );
  NAND2_X2 U8866 ( .A1(n7458), .A2(n7261), .ZN(n8867) );
  NAND3_X2 U8867 ( .A1(n4427), .A2(n8868), .A3(n8867), .ZN(n8897) );
  AND2_X2 U8868 ( .A1(n8897), .A2(n7305), .ZN(ID_EX_REG_ID_EX_REG_N32) );
  NAND2_X2 U8869 ( .A1(n9269), .A2(n7457), .ZN(n8870) );
  NAND2_X2 U8870 ( .A1(n7458), .A2(n7262), .ZN(n8869) );
  NAND3_X2 U8871 ( .A1(n4404), .A2(n8870), .A3(n8869), .ZN(n8895) );
  AND2_X2 U8872 ( .A1(n8895), .A2(n7305), .ZN(ID_EX_REG_ID_EX_REG_N33) );
  NAND2_X2 U8873 ( .A1(n9290), .A2(n8947), .ZN(n8872) );
  NAND2_X2 U8874 ( .A1(n7458), .A2(n7263), .ZN(n8871) );
  NAND3_X2 U8875 ( .A1(n4382), .A2(n8872), .A3(n8871), .ZN(n8945) );
  AND2_X2 U8876 ( .A1(n8945), .A2(n7305), .ZN(ID_EX_REG_ID_EX_REG_N34) );
  NAND2_X2 U8877 ( .A1(n7458), .A2(n7264), .ZN(n8873) );
  NAND3_X2 U8878 ( .A1(n4359), .A2(n8874), .A3(n8873), .ZN(n8935) );
  AND2_X2 U8879 ( .A1(n8935), .A2(n7305), .ZN(ID_EX_REG_ID_EX_REG_N35) );
  NAND2_X2 U8880 ( .A1(n7458), .A2(n7265), .ZN(n8875) );
  NAND3_X2 U8881 ( .A1(n4337), .A2(n8876), .A3(n8875), .ZN(n8942) );
  AND2_X2 U8882 ( .A1(n8942), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N36) );
  NAND2_X2 U8883 ( .A1(n8913), .A2(n8947), .ZN(n8878) );
  NAND2_X2 U8884 ( .A1(n7458), .A2(n7266), .ZN(n8877) );
  NAND3_X2 U8885 ( .A1(n4314), .A2(n8878), .A3(n8877), .ZN(n8911) );
  AND2_X2 U8886 ( .A1(n8911), .A2(n7305), .ZN(ID_EX_REG_ID_EX_REG_N37) );
  NAND2_X2 U8887 ( .A1(n8939), .A2(n8947), .ZN(n8880) );
  NAND2_X2 U8888 ( .A1(n7458), .A2(n7267), .ZN(n8879) );
  NAND3_X2 U8889 ( .A1(n4292), .A2(n8880), .A3(n8879), .ZN(n8937) );
  AND2_X2 U8890 ( .A1(n8937), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N38) );
  AND2_X2 U8891 ( .A1(n8881), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N30) );
  OAI22_X2 U8892 ( .A1(n7084), .A2(n7625), .B1(n7626), .B2(n7404), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8893 ( .A1(n7630), .A2(n7404), .B1(n6171), .B2(n7628), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8894 ( .A1(n7634), .A2(n7404), .B1(n6756), .B2(n7632), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8895 ( .A1(n7639), .A2(n7403), .B1(n7072), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8896 ( .A1(n7643), .A2(n7404), .B1(n6945), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8897 ( .A1(n7647), .A2(n7403), .B1(n7029), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8898 ( .A1(n7651), .A2(n7404), .B1(n7144), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8899 ( .A1(n7083), .A2(n7653), .B1(n3135), .B2(n7403), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8900 ( .A1(n6056), .A2(n7657), .B1(n3133), .B2(n7404), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8901 ( .A1(n7662), .A2(n7403), .B1(n6104), .B2(n7660), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8902 ( .A1(n7666), .A2(n7404), .B1(n6681), .B2(n7664), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8903 ( .A1(n6983), .A2(n7669), .B1(n7670), .B2(n7403), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8904 ( .A1(n7675), .A2(n7404), .B1(n6592), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8905 ( .A1(n7679), .A2(n7404), .B1(n6943), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8906 ( .A1(n7683), .A2(n7403), .B1(n6944), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8907 ( .A1(n7687), .A2(n7403), .B1(n7071), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8908 ( .A1(n7690), .A2(n7403), .B1(n6682), .B2(n7688), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8909 ( .A1(n7694), .A2(n7403), .B1(n6440), .B2(n7692), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8910 ( .A1(n7698), .A2(n7404), .B1(n5964), .B2(n7696), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8911 ( .A1(n7702), .A2(n7403), .B1(n6757), .B2(n7700), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8912 ( .A1(n7706), .A2(n7404), .B1(n5987), .B2(n7704), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8913 ( .A1(n7710), .A2(n7404), .B1(n6072), .B2(n7708), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8914 ( .A1(n7714), .A2(n7404), .B1(n6758), .B2(n7712), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8915 ( .A1(n7718), .A2(n7403), .B1(n6174), .B2(n7716), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8916 ( .A1(n7723), .A2(n7403), .B1(n7145), .B2(n7720), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8917 ( .A1(n7727), .A2(n7403), .B1(n6610), .B2(n7725), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8918 ( .A1(n7732), .A2(n7403), .B1(n6593), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8919 ( .A1(n7736), .A2(n7404), .B1(n6455), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8920 ( .A1(n7739), .A2(n7403), .B1(n6725), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8921 ( .A1(n7744), .A2(n7404), .B1(n6550), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8922 ( .A1(n7747), .A2(n7403), .B1(n6683), .B2(n7745), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8923 ( .A1(n7760), .A2(n7404), .B1(n6441), .B2(n7762), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  AND2_X2 U8924 ( .A1(n8882), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N29) );
  OAI22_X2 U8925 ( .A1(n7626), .A2(n7405), .B1(n7123), .B2(n7625), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8926 ( .A1(n7630), .A2(n7405), .B1(n6170), .B2(n7628), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8927 ( .A1(n7634), .A2(n7405), .B1(n6759), .B2(n7632), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8928 ( .A1(n7639), .A2(n7405), .B1(n7070), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8929 ( .A1(n7643), .A2(n7406), .B1(n6942), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8930 ( .A1(n7647), .A2(n7407), .B1(n7028), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8931 ( .A1(n7651), .A2(n7406), .B1(n7146), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8932 ( .A1(n7654), .A2(n7407), .B1(n7122), .B2(n7653), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8933 ( .A1(n7658), .A2(n7406), .B1(n6436), .B2(n7657), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8934 ( .A1(n7662), .A2(n7407), .B1(n6437), .B2(n7660), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8935 ( .A1(n7666), .A2(n7405), .B1(n6678), .B2(n7664), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8936 ( .A1(n7670), .A2(n7405), .B1(n6474), .B2(n7669), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8937 ( .A1(n7675), .A2(n7406), .B1(n6590), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8938 ( .A1(n7679), .A2(n7406), .B1(n6940), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8939 ( .A1(n7683), .A2(n7406), .B1(n6941), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8940 ( .A1(n7687), .A2(n7407), .B1(n7069), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8941 ( .A1(n7690), .A2(n7407), .B1(n6679), .B2(n7688), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8942 ( .A1(n7694), .A2(n7406), .B1(n6438), .B2(n7692), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8943 ( .A1(n7698), .A2(n7405), .B1(n6169), .B2(n7696), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8944 ( .A1(n7702), .A2(n7405), .B1(n6760), .B2(n7700), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8945 ( .A1(n7706), .A2(n7405), .B1(n5986), .B2(n7704), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8946 ( .A1(n7710), .A2(n7405), .B1(n6071), .B2(n7708), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8947 ( .A1(n7714), .A2(n7406), .B1(n6761), .B2(n7712), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8948 ( .A1(n7718), .A2(n7407), .B1(n6516), .B2(n7716), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8949 ( .A1(n7723), .A2(n7406), .B1(n7147), .B2(n7720), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8950 ( .A1(n7727), .A2(n7407), .B1(n6611), .B2(n7725), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8951 ( .A1(n7732), .A2(n7407), .B1(n6591), .B2(n7730), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8952 ( .A1(n7736), .A2(n7407), .B1(n6122), .B2(n7734), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8953 ( .A1(n7739), .A2(n7405), .B1(n6726), .B2(n7738), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8954 ( .A1(n7744), .A2(n7405), .B1(n6551), .B2(n7742), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8955 ( .A1(n7747), .A2(n7407), .B1(n6680), .B2(n7745), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8956 ( .A1(n7760), .A2(n7406), .B1(n6439), .B2(n7761), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  INV_X4 U8957 ( .A(n8883), .ZN(n8884) );
  OAI22_X2 U8958 ( .A1(n7445), .A2(n8884), .B1(n4516), .B2(n1588), .ZN(
        ID_EX_REG_ID_EX_REG_N124) );
  OAI22_X2 U8959 ( .A1(n7626), .A2(n7408), .B1(n6675), .B2(n7625), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8960 ( .A1(n7630), .A2(n7409), .B1(n6501), .B2(n7628), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8961 ( .A1(n7634), .A2(n7408), .B1(n6762), .B2(n7632), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8962 ( .A1(n7639), .A2(n7409), .B1(n7068), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8963 ( .A1(n7643), .A2(n7410), .B1(n6939), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8964 ( .A1(n7647), .A2(n7410), .B1(n7027), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8965 ( .A1(n7651), .A2(n7410), .B1(n7148), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8966 ( .A1(n7654), .A2(n7410), .B1(n6674), .B2(n7653), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8967 ( .A1(n7658), .A2(n7409), .B1(n6432), .B2(n7656), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8968 ( .A1(n7662), .A2(n7410), .B1(n6433), .B2(n7660), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8969 ( .A1(n7666), .A2(n7408), .B1(n6673), .B2(n7664), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8970 ( .A1(n7670), .A2(n7409), .B1(n6473), .B2(n7668), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8971 ( .A1(n7675), .A2(n7409), .B1(n7067), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8972 ( .A1(n7679), .A2(n7409), .B1(n6937), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8973 ( .A1(n7683), .A2(n7410), .B1(n6938), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8974 ( .A1(n7687), .A2(n7408), .B1(n7066), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8975 ( .A1(n7690), .A2(n7409), .B1(n6676), .B2(n7688), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8976 ( .A1(n7694), .A2(n7408), .B1(n6434), .B2(n7692), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8977 ( .A1(n7698), .A2(n7408), .B1(n6168), .B2(n7696), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8978 ( .A1(n7702), .A2(n7409), .B1(n6763), .B2(n7700), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8979 ( .A1(n7706), .A2(n7408), .B1(n6224), .B2(n7704), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8980 ( .A1(n7710), .A2(n7409), .B1(n5939), .B2(n7708), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8981 ( .A1(n7714), .A2(n7410), .B1(n6764), .B2(n7712), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8982 ( .A1(n7718), .A2(n7409), .B1(n6515), .B2(n7716), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8983 ( .A1(n7723), .A2(n7410), .B1(n7149), .B2(n7720), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8984 ( .A1(n7727), .A2(n7410), .B1(n6612), .B2(n7725), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8985 ( .A1(n7732), .A2(n7408), .B1(n6223), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8986 ( .A1(n7736), .A2(n7410), .B1(n5951), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8987 ( .A1(n7739), .A2(n7408), .B1(n6727), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8988 ( .A1(n7744), .A2(n7409), .B1(n6552), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8989 ( .A1(n7747), .A2(n7408), .B1(n6677), .B2(n7745), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8990 ( .A1(n7760), .A2(n7410), .B1(n6435), .B2(n7762), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  AND2_X2 U8991 ( .A1(n8885), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N26) );
  OAI22_X2 U8992 ( .A1(n7626), .A2(n7411), .B1(n6669), .B2(n7624), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8993 ( .A1(n7630), .A2(n7412), .B1(n6500), .B2(n7628), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8994 ( .A1(n7634), .A2(n7411), .B1(n6765), .B2(n7632), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8995 ( .A1(n7639), .A2(n7412), .B1(n7065), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8996 ( .A1(n7643), .A2(n7413), .B1(n6936), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8997 ( .A1(n7647), .A2(n7411), .B1(n7025), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8998 ( .A1(n7651), .A2(n7413), .B1(n7150), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8999 ( .A1(n7654), .A2(n7412), .B1(n6668), .B2(n7652), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9000 ( .A1(n7658), .A2(n7412), .B1(n6426), .B2(n7656), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9001 ( .A1(n7662), .A2(n7413), .B1(n6427), .B2(n7660), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9002 ( .A1(n7666), .A2(n7411), .B1(n6667), .B2(n7664), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9003 ( .A1(n7670), .A2(n7412), .B1(n6472), .B2(n7668), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9004 ( .A1(n7675), .A2(n7412), .B1(n7064), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9005 ( .A1(n7679), .A2(n7413), .B1(n6934), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9006 ( .A1(n7683), .A2(n7413), .B1(n6935), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9007 ( .A1(n7687), .A2(n7412), .B1(n7063), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9008 ( .A1(n7690), .A2(n7412), .B1(n6670), .B2(n7688), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9009 ( .A1(n7694), .A2(n7411), .B1(n6428), .B2(n7692), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9010 ( .A1(n7698), .A2(n7411), .B1(n6165), .B2(n7696), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9011 ( .A1(n7702), .A2(n7412), .B1(n6766), .B2(n7700), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9012 ( .A1(n7706), .A2(n7411), .B1(n6221), .B2(n7704), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9013 ( .A1(n7710), .A2(n7412), .B1(n5936), .B2(n7708), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9014 ( .A1(n7714), .A2(n7413), .B1(n6767), .B2(n7712), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9015 ( .A1(n7718), .A2(n7413), .B1(n6513), .B2(n7716), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9016 ( .A1(n7723), .A2(n7413), .B1(n7151), .B2(n7720), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9017 ( .A1(n7727), .A2(n7413), .B1(n6613), .B2(n7725), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9018 ( .A1(n7732), .A2(n7411), .B1(n6220), .B2(n7730), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9019 ( .A1(n7736), .A2(n7413), .B1(n5950), .B2(n7734), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9020 ( .A1(n7739), .A2(n7411), .B1(n6728), .B2(n7738), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9021 ( .A1(n7744), .A2(n7412), .B1(n6553), .B2(n7742), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9022 ( .A1(n7747), .A2(n7411), .B1(n6671), .B2(n7745), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9023 ( .A1(n7760), .A2(n7413), .B1(n6429), .B2(n7761), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  AND2_X2 U9024 ( .A1(n8887), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N25) );
  OAI22_X2 U9025 ( .A1(n7626), .A2(n7414), .B1(n6664), .B2(n7624), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9026 ( .A1(n7630), .A2(n7414), .B1(n6499), .B2(n7628), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9027 ( .A1(n7634), .A2(n7414), .B1(n6768), .B2(n7632), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9028 ( .A1(n7639), .A2(n7414), .B1(n7062), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9029 ( .A1(n7643), .A2(n7415), .B1(n6933), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9030 ( .A1(n7647), .A2(n7415), .B1(n7024), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9031 ( .A1(n7651), .A2(n7415), .B1(n7152), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9032 ( .A1(n7654), .A2(n7416), .B1(n6663), .B2(n7652), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9033 ( .A1(n7658), .A2(n7415), .B1(n6422), .B2(n7656), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9034 ( .A1(n7662), .A2(n7416), .B1(n6423), .B2(n7660), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9035 ( .A1(n7666), .A2(n7414), .B1(n6662), .B2(n7664), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9036 ( .A1(n7670), .A2(n7414), .B1(n6471), .B2(n7668), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9037 ( .A1(n7675), .A2(n7416), .B1(n7061), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9038 ( .A1(n7679), .A2(n7416), .B1(n6931), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9039 ( .A1(n7683), .A2(n7415), .B1(n6932), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9040 ( .A1(n7687), .A2(n7416), .B1(n7060), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9041 ( .A1(n7690), .A2(n7415), .B1(n6665), .B2(n7688), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9042 ( .A1(n7694), .A2(n7416), .B1(n6424), .B2(n7692), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9043 ( .A1(n7698), .A2(n7414), .B1(n6164), .B2(n7696), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9044 ( .A1(n7702), .A2(n7414), .B1(n6769), .B2(n7700), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9045 ( .A1(n7706), .A2(n7414), .B1(n6219), .B2(n7704), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9046 ( .A1(n7710), .A2(n7414), .B1(n6070), .B2(n7708), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9047 ( .A1(n7714), .A2(n7415), .B1(n6770), .B2(n7712), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9048 ( .A1(n7718), .A2(n7416), .B1(n6512), .B2(n7716), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9049 ( .A1(n7723), .A2(n7415), .B1(n7153), .B2(n7720), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9050 ( .A1(n7727), .A2(n7415), .B1(n6614), .B2(n7725), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9051 ( .A1(n7732), .A2(n7415), .B1(n6218), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9052 ( .A1(n7736), .A2(n7416), .B1(n6121), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9053 ( .A1(n7739), .A2(n7414), .B1(n6729), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9054 ( .A1(n7744), .A2(n7414), .B1(n6554), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9055 ( .A1(n7747), .A2(n7416), .B1(n6666), .B2(n7745), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9056 ( .A1(n7760), .A2(n7416), .B1(n6425), .B2(n7762), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9057 ( .A(n8889), .ZN(n8890) );
  OAI22_X2 U9058 ( .A1(n7445), .A2(n8890), .B1(n4605), .B2(n1588), .ZN(
        ID_EX_REG_ID_EX_REG_N120) );
  OAI22_X2 U9059 ( .A1(n7626), .A2(n7417), .B1(n6659), .B2(n7624), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9060 ( .A1(n7630), .A2(n7417), .B1(n6498), .B2(n7628), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9061 ( .A1(n7634), .A2(n7417), .B1(n6771), .B2(n7632), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9062 ( .A1(n7639), .A2(n7417), .B1(n7059), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9063 ( .A1(n7643), .A2(n7418), .B1(n6930), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9064 ( .A1(n7647), .A2(n7418), .B1(n7023), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9065 ( .A1(n7651), .A2(n7418), .B1(n7154), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9066 ( .A1(n7654), .A2(n7419), .B1(n6658), .B2(n7652), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9067 ( .A1(n7658), .A2(n7418), .B1(n6418), .B2(n7656), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9068 ( .A1(n7662), .A2(n7419), .B1(n6419), .B2(n7660), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9069 ( .A1(n7666), .A2(n7417), .B1(n6657), .B2(n7664), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9070 ( .A1(n7670), .A2(n7417), .B1(n6470), .B2(n7668), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9071 ( .A1(n7675), .A2(n7419), .B1(n7058), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9072 ( .A1(n7679), .A2(n7419), .B1(n6928), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9073 ( .A1(n7683), .A2(n7418), .B1(n6929), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9074 ( .A1(n7687), .A2(n7419), .B1(n7057), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9075 ( .A1(n7690), .A2(n7418), .B1(n6660), .B2(n7688), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9076 ( .A1(n7694), .A2(n7419), .B1(n6420), .B2(n7692), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9077 ( .A1(n7698), .A2(n7417), .B1(n6163), .B2(n7696), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9078 ( .A1(n7702), .A2(n7417), .B1(n6772), .B2(n7700), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9079 ( .A1(n7706), .A2(n7417), .B1(n6217), .B2(n7704), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9080 ( .A1(n7710), .A2(n7417), .B1(n6069), .B2(n7708), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9081 ( .A1(n7714), .A2(n7418), .B1(n6773), .B2(n7712), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9082 ( .A1(n7718), .A2(n7419), .B1(n6511), .B2(n7716), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9083 ( .A1(n7723), .A2(n7418), .B1(n7155), .B2(n7720), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9084 ( .A1(n7727), .A2(n7418), .B1(n6615), .B2(n7725), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9085 ( .A1(n7732), .A2(n7418), .B1(n6216), .B2(n7730), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9086 ( .A1(n7736), .A2(n7419), .B1(n6120), .B2(n7734), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9087 ( .A1(n7739), .A2(n7417), .B1(n6730), .B2(n7738), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9088 ( .A1(n7744), .A2(n7417), .B1(n6555), .B2(n7742), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9089 ( .A1(n7747), .A2(n7419), .B1(n6661), .B2(n7745), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9090 ( .A1(n7760), .A2(n7419), .B1(n6421), .B2(n7761), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9091 ( .A(n8892), .ZN(n8893) );
  OAI22_X2 U9092 ( .A1(n7445), .A2(n8893), .B1(n4628), .B2(n1588), .ZN(
        ID_EX_REG_ID_EX_REG_N119) );
  OAI22_X2 U9093 ( .A1(n7626), .A2(n7420), .B1(n6654), .B2(n7624), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9094 ( .A1(n7630), .A2(n7421), .B1(n6497), .B2(n7628), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9095 ( .A1(n7634), .A2(n7421), .B1(n6774), .B2(n7632), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9096 ( .A1(n7639), .A2(n7420), .B1(n7056), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9097 ( .A1(n7643), .A2(n7420), .B1(n6384), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9098 ( .A1(n7647), .A2(n7421), .B1(n7022), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9099 ( .A1(n7651), .A2(n7421), .B1(n7156), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9100 ( .A1(n7654), .A2(n7420), .B1(n6653), .B2(n7652), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9101 ( .A1(n6055), .A2(n7657), .B1(n7658), .B2(n7421), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9102 ( .A1(n7662), .A2(n7420), .B1(n6416), .B2(n7660), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9103 ( .A1(n7666), .A2(n7420), .B1(n6652), .B2(n7664), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9104 ( .A1(n6982), .A2(n7669), .B1(n7670), .B2(n7420), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9105 ( .A1(n7675), .A2(n7421), .B1(n7055), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9106 ( .A1(n7679), .A2(n7421), .B1(n6383), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9107 ( .A1(n7683), .A2(n7420), .B1(n6927), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9108 ( .A1(n7687), .A2(n7420), .B1(n7054), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9109 ( .A1(n7690), .A2(n7420), .B1(n6655), .B2(n7688), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9110 ( .A1(n7694), .A2(n7421), .B1(n6417), .B2(n7692), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9111 ( .A1(n7698), .A2(n7421), .B1(n6162), .B2(n7696), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9112 ( .A1(n7702), .A2(n7420), .B1(n6775), .B2(n7700), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9113 ( .A1(n7706), .A2(n7420), .B1(n6215), .B2(n7704), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9114 ( .A1(n7710), .A2(n7421), .B1(n6068), .B2(n7708), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9115 ( .A1(n7714), .A2(n7421), .B1(n6776), .B2(n7712), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9116 ( .A1(n7718), .A2(n7420), .B1(n6510), .B2(n7716), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9117 ( .A1(n7723), .A2(n7420), .B1(n7157), .B2(n7720), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9118 ( .A1(n7727), .A2(n7421), .B1(n6616), .B2(n7725), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9119 ( .A1(n7732), .A2(n7421), .B1(n6214), .B2(n7730), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9120 ( .A1(n7736), .A2(n7421), .B1(n6453), .B2(n7734), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9121 ( .A1(n7739), .A2(n7420), .B1(n6731), .B2(n7738), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9122 ( .A1(n7744), .A2(n7420), .B1(n6556), .B2(n7742), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9123 ( .A1(n7747), .A2(n7421), .B1(n6656), .B2(n7745), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9124 ( .A1(n7760), .A2(n7421), .B1(n6965), .B2(n7762), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9125 ( .A(n7445), .ZN(n8944) );
  NAND2_X2 U9126 ( .A1(n8895), .A2(n8944), .ZN(n8896) );
  NAND2_X2 U9127 ( .A1(n4096), .A2(n8896), .ZN(ID_EX_REG_ID_EX_REG_N129) );
  OAI22_X2 U9128 ( .A1(n7626), .A2(n7422), .B1(n6689), .B2(n7624), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9129 ( .A1(n7630), .A2(n7422), .B1(n5968), .B2(n7629), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9130 ( .A1(n7634), .A2(n7422), .B1(n6777), .B2(n7633), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9131 ( .A1(n7638), .A2(n7423), .B1(n6231), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9132 ( .A1(n7642), .A2(n7423), .B1(n6078), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9133 ( .A1(n7646), .A2(n7423), .B1(n6179), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9134 ( .A1(n7650), .A2(n7422), .B1(n6732), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9135 ( .A1(n7654), .A2(n7423), .B1(n6688), .B2(n7652), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9136 ( .A1(n7658), .A2(n7423), .B1(n6444), .B2(n7656), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9137 ( .A1(n7662), .A2(n7422), .B1(n6106), .B2(n7661), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9138 ( .A1(n7666), .A2(n7422), .B1(n6687), .B2(n7665), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9139 ( .A1(n7670), .A2(n7422), .B1(n6475), .B2(n7668), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9140 ( .A1(n7674), .A2(n7423), .B1(n6229), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9141 ( .A1(n7678), .A2(n7423), .B1(n6076), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9142 ( .A1(n7682), .A2(n7423), .B1(n5941), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9143 ( .A1(n7686), .A2(n7422), .B1(n6228), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9144 ( .A1(n7690), .A2(n7423), .B1(n6690), .B2(n7689), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9145 ( .A1(n7694), .A2(n7423), .B1(n6445), .B2(n7693), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9146 ( .A1(n7698), .A2(n7422), .B1(n5967), .B2(n7697), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9147 ( .A1(n7702), .A2(n7422), .B1(n6778), .B2(n7701), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9148 ( .A1(n7706), .A2(n7422), .B1(n6230), .B2(n7705), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9149 ( .A1(n7710), .A2(n7423), .B1(n6077), .B2(n7709), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9150 ( .A1(n7714), .A2(n7423), .B1(n6779), .B2(n7713), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9151 ( .A1(n7718), .A2(n7423), .B1(n6178), .B2(n7717), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9152 ( .A1(n7723), .A2(n7422), .B1(n7158), .B2(n7721), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9153 ( .A1(n7727), .A2(n7423), .B1(n6617), .B2(n7726), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9154 ( .A1(n3090), .A2(n7423), .B1(n7073), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9155 ( .A1(n7735), .A2(n7422), .B1(n6979), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9156 ( .A1(n7740), .A2(n7422), .B1(n7159), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9157 ( .A1(n7743), .A2(n7422), .B1(n7039), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9158 ( .A1(n7747), .A2(n7423), .B1(n6691), .B2(n7746), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9159 ( .A1(n7760), .A2(n7422), .B1(n6446), .B2(n7762), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9160 ( .A1(n8897), .A2(n8944), .ZN(n8898) );
  NAND2_X2 U9161 ( .A1(n4096), .A2(n8898), .ZN(ID_EX_REG_ID_EX_REG_N128) );
  OAI22_X2 U9162 ( .A1(n7088), .A2(n7625), .B1(n7626), .B2(n7424), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9163 ( .A1(n7630), .A2(n7424), .B1(n5966), .B2(n7629), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9164 ( .A1(n7634), .A2(n7424), .B1(n6780), .B2(n7633), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9165 ( .A1(n7638), .A2(n7425), .B1(n6227), .B2(n7637), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9166 ( .A1(n7642), .A2(n7424), .B1(n6075), .B2(n7641), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9167 ( .A1(n7646), .A2(n7425), .B1(n6177), .B2(n7645), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9168 ( .A1(n7650), .A2(n7425), .B1(n6733), .B2(n7649), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9169 ( .A1(n7087), .A2(n7653), .B1(n3135), .B2(n7425), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9170 ( .A1(n6057), .A2(n7657), .B1(n3133), .B2(n7424), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9171 ( .A1(n7662), .A2(n7425), .B1(n6105), .B2(n7661), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9172 ( .A1(n7666), .A2(n7425), .B1(n6684), .B2(n7665), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9173 ( .A1(n6985), .A2(n7669), .B1(n7670), .B2(n7425), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9174 ( .A1(n7674), .A2(n7424), .B1(n6599), .B2(n7673), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9175 ( .A1(n7678), .A2(n7425), .B1(n6390), .B2(n7677), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9176 ( .A1(n7682), .A2(n7424), .B1(n5940), .B2(n7681), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9177 ( .A1(n7686), .A2(n7425), .B1(n6225), .B2(n7685), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9178 ( .A1(n7690), .A2(n7424), .B1(n6685), .B2(n7689), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9179 ( .A1(n7694), .A2(n7425), .B1(n6442), .B2(n7693), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9180 ( .A1(n7698), .A2(n7425), .B1(n5965), .B2(n7697), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9181 ( .A1(n7702), .A2(n7425), .B1(n6781), .B2(n7701), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9182 ( .A1(n7706), .A2(n7425), .B1(n6226), .B2(n7705), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9183 ( .A1(n7710), .A2(n7424), .B1(n6074), .B2(n7709), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9184 ( .A1(n7714), .A2(n7424), .B1(n6782), .B2(n7713), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9185 ( .A1(n7718), .A2(n7424), .B1(n6176), .B2(n7717), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9186 ( .A1(n7723), .A2(n7425), .B1(n7160), .B2(n7721), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9187 ( .A1(n7727), .A2(n7424), .B1(n6618), .B2(n7726), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9188 ( .A1(n3090), .A2(n7425), .B1(n6600), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9189 ( .A1(n7735), .A2(n7424), .B1(n6457), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9190 ( .A1(n7740), .A2(n7425), .B1(n7161), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9191 ( .A1(n7743), .A2(n7424), .B1(n7040), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9192 ( .A1(n7747), .A2(n7424), .B1(n6686), .B2(n7746), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9193 ( .A1(n7760), .A2(n7424), .B1(n6443), .B2(n7762), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9194 ( .A1(n8899), .A2(n8944), .ZN(n8900) );
  NAND2_X2 U9195 ( .A1(n4096), .A2(n8900), .ZN(ID_EX_REG_ID_EX_REG_N127) );
  OAI22_X2 U9196 ( .A1(n7086), .A2(n7625), .B1(n7626), .B2(n7426), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9197 ( .A1(n7630), .A2(n7426), .B1(n7008), .B2(n7629), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9198 ( .A1(n7634), .A2(n7426), .B1(n7183), .B2(n7633), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9199 ( .A1(n7638), .A2(n7427), .B1(n6598), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9200 ( .A1(n7642), .A2(n7426), .B1(n6389), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9201 ( .A1(n7646), .A2(n7427), .B1(n6175), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9202 ( .A1(n7650), .A2(n7427), .B1(n6734), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9203 ( .A1(n7085), .A2(n7653), .B1(n3135), .B2(n7427), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9204 ( .A1(n6921), .A2(n7657), .B1(n3133), .B2(n7426), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9205 ( .A1(n7662), .A2(n7427), .B1(n6968), .B2(n7661), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9206 ( .A1(n7666), .A2(n7427), .B1(n7124), .B2(n7665), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9207 ( .A1(n6984), .A2(n7669), .B1(n7670), .B2(n7427), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9208 ( .A1(n7674), .A2(n7426), .B1(n6595), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9209 ( .A1(n7678), .A2(n7427), .B1(n6387), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9210 ( .A1(n7682), .A2(n7426), .B1(n6073), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9211 ( .A1(n7686), .A2(n7427), .B1(n6594), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9212 ( .A1(n7690), .A2(n7426), .B1(n7125), .B2(n7689), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9213 ( .A1(n7694), .A2(n7427), .B1(n6969), .B2(n7693), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9214 ( .A1(n7698), .A2(n7427), .B1(n6172), .B2(n7697), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9215 ( .A1(n7702), .A2(n7427), .B1(n7184), .B2(n7701), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9216 ( .A1(n7706), .A2(n7427), .B1(n6597), .B2(n7705), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9217 ( .A1(n7710), .A2(n7426), .B1(n6388), .B2(n7709), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9218 ( .A1(n7714), .A2(n7426), .B1(n7185), .B2(n7713), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9219 ( .A1(n7718), .A2(n7426), .B1(n7030), .B2(n7717), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9220 ( .A1(n7722), .A2(n7427), .B1(n7162), .B2(n7721), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9221 ( .A1(n7727), .A2(n7426), .B1(n7092), .B2(n7726), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9222 ( .A1(n3090), .A2(n7427), .B1(n6596), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9223 ( .A1(n7735), .A2(n7426), .B1(n6456), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9224 ( .A1(n7740), .A2(n7427), .B1(n7163), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9225 ( .A1(n7743), .A2(n7426), .B1(n7041), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9226 ( .A1(n7747), .A2(n7426), .B1(n7126), .B2(n7746), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9227 ( .A1(n7759), .A2(n7426), .B1(n6970), .B2(n7762), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  AND2_X2 U9228 ( .A1(n8901), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N22) );
  OAI22_X2 U9229 ( .A1(n7626), .A2(n7428), .B1(n6651), .B2(n7624), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9230 ( .A1(n7630), .A2(n7428), .B1(n7007), .B2(n7629), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9231 ( .A1(n7634), .A2(n7428), .B1(n7186), .B2(n7633), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9232 ( .A1(n7638), .A2(n7428), .B1(n6585), .B2(n7637), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9233 ( .A1(n7642), .A2(n7429), .B1(n6067), .B2(n7641), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9234 ( .A1(n7646), .A2(n7429), .B1(n6509), .B2(n7645), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9235 ( .A1(n7650), .A2(n7429), .B1(n6735), .B2(n7649), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9236 ( .A1(n7654), .A2(n7430), .B1(n6650), .B2(n7652), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9237 ( .A1(n7658), .A2(n7430), .B1(n6413), .B2(n7656), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9238 ( .A1(n7662), .A2(n7430), .B1(n6964), .B2(n7661), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9239 ( .A1(n7666), .A2(n7428), .B1(n7115), .B2(n7665), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9240 ( .A1(n7670), .A2(n7428), .B1(n6469), .B2(n7668), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9241 ( .A1(n7674), .A2(n7429), .B1(n6213), .B2(n7673), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9242 ( .A1(n7678), .A2(n7430), .B1(n6065), .B2(n7677), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9243 ( .A1(n7682), .A2(n7429), .B1(n6382), .B2(n7681), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9244 ( .A1(n7686), .A2(n7430), .B1(n6583), .B2(n7685), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9245 ( .A1(n7690), .A2(n7429), .B1(n7116), .B2(n7689), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9246 ( .A1(n7694), .A2(n7430), .B1(n6414), .B2(n7693), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9247 ( .A1(n7698), .A2(n7428), .B1(n6496), .B2(n7697), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9248 ( .A1(n7702), .A2(n7428), .B1(n7187), .B2(n7701), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9249 ( .A1(n7706), .A2(n7428), .B1(n6584), .B2(n7705), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9250 ( .A1(n7710), .A2(n7428), .B1(n6066), .B2(n7709), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9251 ( .A1(n7714), .A2(n7429), .B1(n7188), .B2(n7713), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9252 ( .A1(n7718), .A2(n7429), .B1(n7021), .B2(n7717), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9253 ( .A1(n7722), .A2(n7429), .B1(n7164), .B2(n7721), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9254 ( .A1(n7727), .A2(n7429), .B1(n7093), .B2(n7726), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9255 ( .A1(n3090), .A2(n7430), .B1(n7053), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9256 ( .A1(n7735), .A2(n7430), .B1(n6119), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9257 ( .A1(n7740), .A2(n7428), .B1(n7165), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9258 ( .A1(n7743), .A2(n7428), .B1(n7042), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9259 ( .A1(n7747), .A2(n7430), .B1(n7117), .B2(n7746), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9260 ( .A1(n7759), .A2(n7430), .B1(n6415), .B2(n7762), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  AND2_X2 U9261 ( .A1(n8903), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N18) );
  OAI22_X2 U9262 ( .A1(n7078), .A2(n7625), .B1(n7626), .B2(n7431), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9263 ( .A1(n7630), .A2(n7432), .B1(n7006), .B2(n7629), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9264 ( .A1(n7634), .A2(n7431), .B1(n7189), .B2(n7633), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9265 ( .A1(n7638), .A2(n7432), .B1(n6574), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9266 ( .A1(n7642), .A2(n7431), .B1(n5873), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9267 ( .A1(n7646), .A2(n7432), .B1(n6507), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9268 ( .A1(n7650), .A2(n7432), .B1(n6736), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9269 ( .A1(n7077), .A2(n7653), .B1(n7654), .B2(n7432), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9270 ( .A1(n6920), .A2(n7657), .B1(n7658), .B2(n7431), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9271 ( .A1(n7662), .A2(n7432), .B1(n6959), .B2(n7661), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9272 ( .A1(n7666), .A2(n7432), .B1(n7106), .B2(n7665), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9273 ( .A1(n6124), .A2(n7669), .B1(n7670), .B2(n7432), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9274 ( .A1(n7674), .A2(n7431), .B1(n6571), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9275 ( .A1(n7678), .A2(n7431), .B1(n5872), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9276 ( .A1(n7682), .A2(n7431), .B1(n6379), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9277 ( .A1(n7686), .A2(n7432), .B1(n6570), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9278 ( .A1(n7690), .A2(n7431), .B1(n7107), .B2(n7689), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9279 ( .A1(n7694), .A2(n7432), .B1(n6960), .B2(n7693), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9280 ( .A1(n7698), .A2(n7431), .B1(n6493), .B2(n7697), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9281 ( .A1(n7702), .A2(n7432), .B1(n7190), .B2(n7701), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9282 ( .A1(n7706), .A2(n7432), .B1(n6573), .B2(n7705), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9283 ( .A1(n7710), .A2(n7431), .B1(n5934), .B2(n7709), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9284 ( .A1(n7714), .A2(n7431), .B1(n7191), .B2(n7713), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9285 ( .A1(n7718), .A2(n7431), .B1(n7015), .B2(n7717), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9286 ( .A1(n7722), .A2(n7432), .B1(n7166), .B2(n7721), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9287 ( .A1(n7727), .A2(n7431), .B1(n7094), .B2(n7726), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9288 ( .A1(n3090), .A2(n7432), .B1(n6572), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9289 ( .A1(n7735), .A2(n7432), .B1(n5882), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9290 ( .A1(n7740), .A2(n7432), .B1(n7167), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9291 ( .A1(n7743), .A2(n7431), .B1(n7043), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9292 ( .A1(n7747), .A2(n7431), .B1(n7108), .B2(n7746), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9293 ( .A1(n7759), .A2(n7431), .B1(n6961), .B2(n7762), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9294 ( .A(n8905), .ZN(n8906) );
  OAI22_X2 U9295 ( .A1(n7445), .A2(n8906), .B1(n3328), .B2(n1588), .ZN(
        ID_EX_REG_ID_EX_REG_N113) );
  OAI22_X2 U9296 ( .A1(n7076), .A2(n7625), .B1(n7626), .B2(n7433), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9297 ( .A1(n7630), .A2(n7434), .B1(n7005), .B2(n7629), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9298 ( .A1(n7634), .A2(n7433), .B1(n7192), .B2(n7633), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9299 ( .A1(n7638), .A2(n7434), .B1(n6569), .B2(n7637), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9300 ( .A1(n7642), .A2(n7433), .B1(n5871), .B2(n7641), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9301 ( .A1(n7646), .A2(n7434), .B1(n6506), .B2(n7645), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9302 ( .A1(n7650), .A2(n7433), .B1(n6737), .B2(n7649), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9303 ( .A1(n7075), .A2(n7653), .B1(n3135), .B2(n7434), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9304 ( .A1(n6919), .A2(n7657), .B1(n7658), .B2(n7433), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9305 ( .A1(n7662), .A2(n7434), .B1(n6956), .B2(n7661), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9306 ( .A1(n7666), .A2(n7434), .B1(n7103), .B2(n7665), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9307 ( .A1(n6123), .A2(n7669), .B1(n7670), .B2(n7434), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9308 ( .A1(n7674), .A2(n7433), .B1(n6566), .B2(n7673), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9309 ( .A1(n7678), .A2(n7434), .B1(n6376), .B2(n7677), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9310 ( .A1(n7682), .A2(n7433), .B1(n6377), .B2(n7681), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9311 ( .A1(n7686), .A2(n7434), .B1(n6565), .B2(n7685), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9312 ( .A1(n7690), .A2(n7433), .B1(n7104), .B2(n7689), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9313 ( .A1(n7694), .A2(n7434), .B1(n6957), .B2(n7693), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9314 ( .A1(n7698), .A2(n7434), .B1(n6492), .B2(n7697), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9315 ( .A1(n7702), .A2(n7434), .B1(n7193), .B2(n7701), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9316 ( .A1(n7706), .A2(n7434), .B1(n6568), .B2(n7705), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9317 ( .A1(n7710), .A2(n7433), .B1(n6378), .B2(n7709), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9318 ( .A1(n7714), .A2(n7433), .B1(n7194), .B2(n7713), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9319 ( .A1(n7718), .A2(n7433), .B1(n7014), .B2(n7717), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9320 ( .A1(n7722), .A2(n7434), .B1(n7168), .B2(n7721), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9321 ( .A1(n7727), .A2(n7433), .B1(n7095), .B2(n7726), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9322 ( .A1(n3090), .A2(n7434), .B1(n6567), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9323 ( .A1(n7735), .A2(n7433), .B1(n5899), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9324 ( .A1(n7740), .A2(n7434), .B1(n7169), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9325 ( .A1(n7743), .A2(n7433), .B1(n7044), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9326 ( .A1(n7747), .A2(n7433), .B1(n7105), .B2(n7746), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9327 ( .A1(n7759), .A2(n7433), .B1(n6958), .B2(n7762), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  AND2_X2 U9328 ( .A1(n8908), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N16) );
  OAI22_X2 U9329 ( .A1(n7626), .A2(n7435), .B1(n6644), .B2(n7624), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9330 ( .A1(n7630), .A2(n7436), .B1(n7004), .B2(n7629), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9331 ( .A1(n7634), .A2(n8910), .B1(n7195), .B2(n7633), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9332 ( .A1(n7638), .A2(n7435), .B1(n6564), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9333 ( .A1(n7642), .A2(n7436), .B1(n6375), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9334 ( .A1(n7646), .A2(n8910), .B1(n6505), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9335 ( .A1(n7650), .A2(n7435), .B1(n6738), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9336 ( .A1(n7654), .A2(n7436), .B1(n6643), .B2(n7652), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9337 ( .A1(n7658), .A2(n8910), .B1(n6408), .B2(n7656), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9338 ( .A1(n7662), .A2(n7435), .B1(n6953), .B2(n7661), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9339 ( .A1(n7666), .A2(n7436), .B1(n7100), .B2(n7665), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9340 ( .A1(n7670), .A2(n8910), .B1(n6130), .B2(n7668), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9341 ( .A1(n7674), .A2(n7435), .B1(n6209), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9342 ( .A1(n7678), .A2(n7436), .B1(n6062), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9343 ( .A1(n7682), .A2(n8910), .B1(n6373), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9344 ( .A1(n7686), .A2(n7435), .B1(n6562), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9345 ( .A1(n7690), .A2(n7436), .B1(n7101), .B2(n7689), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9346 ( .A1(n7694), .A2(n8910), .B1(n6954), .B2(n7693), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9347 ( .A1(n7698), .A2(n7435), .B1(n6491), .B2(n7697), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9348 ( .A1(n7702), .A2(n7436), .B1(n7196), .B2(n7701), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9349 ( .A1(n7706), .A2(n8910), .B1(n6563), .B2(n7705), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9350 ( .A1(n7710), .A2(n7435), .B1(n6374), .B2(n7709), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9351 ( .A1(n7714), .A2(n7436), .B1(n7197), .B2(n7713), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9352 ( .A1(n7718), .A2(n8910), .B1(n7013), .B2(n7717), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9353 ( .A1(n7722), .A2(n7435), .B1(n7170), .B2(n7721), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9354 ( .A1(n7727), .A2(n7436), .B1(n7096), .B2(n7726), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9355 ( .A1(n3090), .A2(n8910), .B1(n7048), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9356 ( .A1(n7735), .A2(n7435), .B1(n5898), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9357 ( .A1(n7740), .A2(n7436), .B1(n7171), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9358 ( .A1(n7743), .A2(n8910), .B1(n7045), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9359 ( .A1(n7747), .A2(n7435), .B1(n7102), .B2(n7746), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9360 ( .A1(n7759), .A2(n7436), .B1(n6955), .B2(n7762), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9361 ( .A1(n7626), .A2(n7481), .B1(n6640), .B2(n7624), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9362 ( .A1(n7630), .A2(n7481), .B1(n7003), .B2(n7629), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9363 ( .A1(n7634), .A2(n7481), .B1(n7198), .B2(n7633), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9364 ( .A1(n7638), .A2(n7481), .B1(n6208), .B2(n7637), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9365 ( .A1(n7642), .A2(n7481), .B1(n6061), .B2(n7641), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9366 ( .A1(n7646), .A2(n7481), .B1(n6504), .B2(n7645), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9367 ( .A1(n7650), .A2(n7481), .B1(n6739), .B2(n7649), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9368 ( .A1(n7654), .A2(n7481), .B1(n6639), .B2(n7652), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9369 ( .A1(n7658), .A2(n7481), .B1(n6406), .B2(n7656), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9370 ( .A1(n7662), .A2(n7481), .B1(n6951), .B2(n7661), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9371 ( .A1(n7666), .A2(n7481), .B1(n7099), .B2(n7665), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9372 ( .A1(n7670), .A2(n7482), .B1(n6468), .B2(n7668), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9373 ( .A1(n7674), .A2(n7482), .B1(n5906), .B2(n7673), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9374 ( .A1(n7678), .A2(n7482), .B1(n6060), .B2(n7677), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9375 ( .A1(n7682), .A2(n7482), .B1(n6371), .B2(n7681), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9376 ( .A1(n7686), .A2(n7482), .B1(n6561), .B2(n7685), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9377 ( .A1(n7690), .A2(n7482), .B1(n6641), .B2(n7689), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9378 ( .A1(n7694), .A2(n7482), .B1(n6952), .B2(n7693), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9379 ( .A1(n7698), .A2(n7482), .B1(n7002), .B2(n7697), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9380 ( .A1(n7702), .A2(n7482), .B1(n7199), .B2(n7701), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9381 ( .A1(n7706), .A2(n7482), .B1(n6207), .B2(n7705), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9382 ( .A1(n7710), .A2(n7482), .B1(n6372), .B2(n7709), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9383 ( .A1(n7714), .A2(n7482), .B1(n6783), .B2(n7713), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9384 ( .A1(n7718), .A2(n7481), .B1(n6503), .B2(n7717), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9385 ( .A1(n7727), .A2(n7482), .B1(n6619), .B2(n7726), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9386 ( .A1(n3090), .A2(n7481), .B1(n5985), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9387 ( .A1(n7735), .A2(n7482), .B1(n6118), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9388 ( .A1(n7740), .A2(n7481), .B1(n6740), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9389 ( .A1(n7743), .A2(n7482), .B1(n6557), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9390 ( .A1(n7747), .A2(n7481), .B1(n6642), .B2(n7746), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9391 ( .A1(n7759), .A2(n7482), .B1(n6407), .B2(n7762), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9392 ( .A1(n8911), .A2(n8944), .ZN(n8912) );
  NAND2_X2 U9393 ( .A1(n4096), .A2(n8912), .ZN(ID_EX_REG_ID_EX_REG_N133) );
  INV_X4 U9394 ( .A(n8913), .ZN(n9245) );
  INV_X4 U9395 ( .A(n7439), .ZN(n8914) );
  OAI22_X2 U9396 ( .A1(n7626), .A2(n8914), .B1(n6695), .B2(n7624), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9397 ( .A(n7440), .ZN(n8915) );
  OAI22_X2 U9398 ( .A1(n7630), .A2(n8915), .B1(n7010), .B2(n7629), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9399 ( .A(n7441), .ZN(n8916) );
  OAI22_X2 U9400 ( .A1(n7634), .A2(n8916), .B1(n7200), .B2(n7633), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9401 ( .A(n7442), .ZN(n8917) );
  OAI22_X2 U9402 ( .A1(n7638), .A2(n8917), .B1(n6605), .B2(n7636), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9403 ( .A(n7439), .ZN(n8918) );
  OAI22_X2 U9404 ( .A1(n7642), .A2(n8918), .B1(n5877), .B2(n7640), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9405 ( .A(n7440), .ZN(n8919) );
  OAI22_X2 U9406 ( .A1(n7646), .A2(n8919), .B1(n6517), .B2(n7644), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9407 ( .A(n7441), .ZN(n8920) );
  OAI22_X2 U9408 ( .A1(n7650), .A2(n8920), .B1(n6741), .B2(n7648), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9409 ( .A(n7442), .ZN(n8921) );
  OAI22_X2 U9410 ( .A1(n7654), .A2(n8921), .B1(n6694), .B2(n7652), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9411 ( .A(n7439), .ZN(n8922) );
  OAI22_X2 U9412 ( .A1(n7658), .A2(n8922), .B1(n6109), .B2(n7656), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9413 ( .A(n7440), .ZN(n8923) );
  OAI22_X2 U9414 ( .A1(n7662), .A2(n8923), .B1(n6975), .B2(n7661), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9415 ( .A(n7441), .ZN(n8924) );
  OAI22_X2 U9416 ( .A1(n7666), .A2(n8924), .B1(n7130), .B2(n7665), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9417 ( .A1(n7670), .A2(n8917), .B1(n6132), .B2(n7668), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9418 ( .A(n7439), .ZN(n8925) );
  OAI22_X2 U9419 ( .A1(n7674), .A2(n8925), .B1(n6237), .B2(n7672), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9420 ( .A(n7440), .ZN(n8926) );
  OAI22_X2 U9421 ( .A1(n7678), .A2(n8926), .B1(n5876), .B2(n7676), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9422 ( .A1(n7682), .A2(n8920), .B1(n6397), .B2(n7680), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9423 ( .A(n7442), .ZN(n8927) );
  OAI22_X2 U9424 ( .A1(n7686), .A2(n8927), .B1(n6603), .B2(n7684), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9425 ( .A(n7439), .ZN(n8928) );
  OAI22_X2 U9426 ( .A1(n7690), .A2(n8928), .B1(n7131), .B2(n7689), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9427 ( .A(n7440), .ZN(n8929) );
  OAI22_X2 U9428 ( .A1(n7694), .A2(n8929), .B1(n6976), .B2(n7693), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9429 ( .A1(n7698), .A2(n8924), .B1(n6502), .B2(n7697), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9430 ( .A1(n7702), .A2(n8927), .B1(n7201), .B2(n7701), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9431 ( .A(n7439), .ZN(n8930) );
  OAI22_X2 U9432 ( .A1(n7706), .A2(n8930), .B1(n6604), .B2(n7705), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9433 ( .A(n7440), .ZN(n8931) );
  OAI22_X2 U9434 ( .A1(n7710), .A2(n8931), .B1(n6083), .B2(n7709), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9435 ( .A1(n7714), .A2(n8921), .B1(n7202), .B2(n7713), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9436 ( .A(n7442), .ZN(n8932) );
  OAI22_X2 U9437 ( .A1(n7718), .A2(n8932), .B1(n7032), .B2(n7717), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9438 ( .A(n7439), .ZN(n8933) );
  OAI22_X2 U9439 ( .A1(n7722), .A2(n8933), .B1(n7172), .B2(n7721), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U9440 ( .A(n7440), .ZN(n8934) );
  OAI22_X2 U9441 ( .A1(n7727), .A2(n8934), .B1(n7097), .B2(n7726), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9442 ( .A1(n3090), .A2(n8917), .B1(n7074), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9443 ( .A1(n7735), .A2(n8921), .B1(n6980), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9444 ( .A1(n7740), .A2(n8930), .B1(n7173), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9445 ( .A1(n7743), .A2(n8923), .B1(n7046), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9446 ( .A1(n7747), .A2(n8916), .B1(n7132), .B2(n7746), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9447 ( .A1(n7759), .A2(n8932), .B1(n6110), .B2(n7762), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9448 ( .A1(n8935), .A2(n8944), .ZN(n8936) );
  NAND2_X2 U9449 ( .A1(n4096), .A2(n8936), .ZN(ID_EX_REG_ID_EX_REG_N131) );
  OAI22_X2 U9450 ( .A1(n7090), .A2(n7625), .B1(n7626), .B2(n7443), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9451 ( .A1(n7630), .A2(n7443), .B1(n7009), .B2(n7629), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9452 ( .A1(n7634), .A2(n7443), .B1(n7203), .B2(n7633), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9453 ( .A1(n7638), .A2(n7444), .B1(n6235), .B2(n7637), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9454 ( .A1(n7642), .A2(n7443), .B1(n6394), .B2(n7641), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9455 ( .A1(n7646), .A2(n7444), .B1(n6182), .B2(n7645), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9456 ( .A1(n7650), .A2(n7444), .B1(n6742), .B2(n7649), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9457 ( .A1(n7089), .A2(n7653), .B1(n7654), .B2(n7444), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9458 ( .A1(n6922), .A2(n7657), .B1(n7658), .B2(n7443), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9459 ( .A1(n7662), .A2(n7444), .B1(n6971), .B2(n7661), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9460 ( .A1(n7666), .A2(n7444), .B1(n7127), .B2(n7665), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9461 ( .A1(n6986), .A2(n7669), .B1(n7670), .B2(n7444), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9462 ( .A1(n7674), .A2(n7443), .B1(n6233), .B2(n7673), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9463 ( .A1(n7678), .A2(n7444), .B1(n6392), .B2(n7677), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9464 ( .A1(n7682), .A2(n7443), .B1(n6081), .B2(n7681), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9465 ( .A1(n7686), .A2(n7444), .B1(n6602), .B2(n7685), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9466 ( .A1(n7690), .A2(n7443), .B1(n7128), .B2(n7689), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9467 ( .A1(n7694), .A2(n7444), .B1(n6972), .B2(n7693), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9468 ( .A1(n7698), .A2(n7444), .B1(n6173), .B2(n7697), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9469 ( .A1(n7702), .A2(n7444), .B1(n7204), .B2(n7701), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9470 ( .A1(n7706), .A2(n7444), .B1(n6234), .B2(n7705), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9471 ( .A1(n7710), .A2(n7443), .B1(n6393), .B2(n7709), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9472 ( .A1(n7714), .A2(n7443), .B1(n7205), .B2(n7713), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9473 ( .A1(n7718), .A2(n7443), .B1(n7031), .B2(n7717), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9474 ( .A1(n7722), .A2(n7444), .B1(n7174), .B2(n7721), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9475 ( .A1(n7727), .A2(n7443), .B1(n7098), .B2(n7726), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9476 ( .A1(n3090), .A2(n7444), .B1(n5990), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9477 ( .A1(n7735), .A2(n7443), .B1(n6459), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9478 ( .A1(n7740), .A2(n7444), .B1(n7175), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9479 ( .A1(n7743), .A2(n7443), .B1(n7047), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9480 ( .A1(n7747), .A2(n7443), .B1(n7129), .B2(n7746), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9481 ( .A1(n7759), .A2(n7443), .B1(n6973), .B2(n7762), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9482 ( .A1(n8937), .A2(n8944), .ZN(n8938) );
  NAND2_X2 U9483 ( .A1(n4096), .A2(n8938), .ZN(ID_EX_REG_ID_EX_REG_N134) );
  INV_X4 U9484 ( .A(n8939), .ZN(n8940) );
  OAI22_X2 U9485 ( .A1(n7626), .A2(n7455), .B1(n6697), .B2(n7624), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9486 ( .A1(n7630), .A2(n7455), .B1(n7012), .B2(n7629), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9487 ( .A1(n7634), .A2(n7455), .B1(n7206), .B2(n7633), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9488 ( .A1(n7638), .A2(n7455), .B1(n6239), .B2(n7637), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9489 ( .A1(n7642), .A2(n7455), .B1(n5879), .B2(n7641), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9490 ( .A1(n7646), .A2(n7455), .B1(n6519), .B2(n7645), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9491 ( .A1(n7650), .A2(n7455), .B1(n6743), .B2(n7649), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9492 ( .A1(n7654), .A2(n7455), .B1(n6696), .B2(n7652), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9493 ( .A1(n7658), .A2(n7455), .B1(n6111), .B2(n7656), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9494 ( .A1(n7662), .A2(n7455), .B1(n6977), .B2(n7661), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9495 ( .A1(n7666), .A2(n7455), .B1(n7133), .B2(n7665), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9496 ( .A1(n7670), .A2(n7456), .B1(n6133), .B2(n7668), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9497 ( .A1(n7674), .A2(n7456), .B1(n6238), .B2(n7673), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9498 ( .A1(n7678), .A2(n7456), .B1(n5878), .B2(n7677), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9499 ( .A1(n7682), .A2(n7456), .B1(n6398), .B2(n7681), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9500 ( .A1(n7686), .A2(n7456), .B1(n6606), .B2(n7685), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9501 ( .A1(n7690), .A2(n7456), .B1(n7134), .B2(n7689), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9502 ( .A1(n7694), .A2(n7456), .B1(n6978), .B2(n7693), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9503 ( .A1(n7698), .A2(n7456), .B1(n7011), .B2(n7697), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9504 ( .A1(n7702), .A2(n7456), .B1(n7207), .B2(n7701), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9505 ( .A1(n7706), .A2(n7456), .B1(n6607), .B2(n7705), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9506 ( .A1(n7710), .A2(n7456), .B1(n6084), .B2(n7709), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9507 ( .A1(n7714), .A2(n7454), .B1(n6784), .B2(n7713), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9508 ( .A1(n7718), .A2(n7454), .B1(n6518), .B2(n7717), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9509 ( .A1(n7722), .A2(n7454), .B1(n6744), .B2(n7721), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9510 ( .A1(n7727), .A2(n7454), .B1(n6620), .B2(n7726), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9511 ( .A1(n3090), .A2(n7454), .B1(n5995), .B2(n7729), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9512 ( .A1(n7735), .A2(n7454), .B1(n5883), .B2(n7733), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9513 ( .A1(n7740), .A2(n7454), .B1(n6745), .B2(n7737), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9514 ( .A1(n7743), .A2(n7454), .B1(n6558), .B2(n7741), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9515 ( .A1(n7747), .A2(n7455), .B1(n6698), .B2(n7746), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9516 ( .A1(n7759), .A2(n7456), .B1(n6112), .B2(n7761), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9517 ( .A1(n8942), .A2(n8944), .ZN(n8943) );
  NAND2_X2 U9518 ( .A1(n4096), .A2(n8943), .ZN(ID_EX_REG_ID_EX_REG_N132) );
  OAI22_X2 U9519 ( .A1(n6243), .A2(n7624), .B1(n7626), .B2(n5862), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9520 ( .A1(n7630), .A2(n5862), .B1(n5972), .B2(n7628), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9521 ( .A1(n7634), .A2(n5862), .B1(n6785), .B2(n7632), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9522 ( .A1(n7639), .A2(n5862), .B1(n5994), .B2(n7637), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9523 ( .A1(n7643), .A2(n5862), .B1(n6396), .B2(n7641), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9524 ( .A1(n7647), .A2(n5862), .B1(n6184), .B2(n7645), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9525 ( .A1(n7651), .A2(n5862), .B1(n6746), .B2(n7649), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9526 ( .A1(n6242), .A2(n7652), .B1(n7654), .B2(n5862), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9527 ( .A1(n6059), .A2(n7657), .B1(n7658), .B2(n5862), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9528 ( .A1(n7662), .A2(n5862), .B1(n6108), .B2(n7660), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9529 ( .A1(n7666), .A2(n5862), .B1(n6693), .B2(n7664), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9530 ( .A1(n6127), .A2(n7669), .B1(n7670), .B2(n5862), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9531 ( .A1(n7675), .A2(n5862), .B1(n5991), .B2(n7673), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9532 ( .A1(n7679), .A2(n5862), .B1(n6395), .B2(n7677), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9533 ( .A1(n7683), .A2(n5862), .B1(n5943), .B2(n7681), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9534 ( .A1(n7687), .A2(n5862), .B1(n6236), .B2(n7685), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9535 ( .A1(n7690), .A2(n5862), .B1(n6264), .B2(n7688), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9536 ( .A1(n7694), .A2(n5862), .B1(n6449), .B2(n7692), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9537 ( .A1(n7698), .A2(n5862), .B1(n5971), .B2(n7696), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9538 ( .A1(n7702), .A2(n5862), .B1(n6786), .B2(n7700), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9539 ( .A1(n7706), .A2(n5862), .B1(n5993), .B2(n7704), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9540 ( .A1(n7710), .A2(n5862), .B1(n6082), .B2(n7708), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9541 ( .A1(n7714), .A2(n5862), .B1(n6787), .B2(n7712), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9542 ( .A1(n7718), .A2(n5862), .B1(n6183), .B2(n7716), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9543 ( .A1(n7722), .A2(n5862), .B1(n7176), .B2(n7721), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9544 ( .A1(n7727), .A2(n5862), .B1(n6621), .B2(n7725), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9545 ( .A1(n7732), .A2(n5862), .B1(n5992), .B2(n7730), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9546 ( .A1(n7736), .A2(n5862), .B1(n6460), .B2(n7734), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9547 ( .A1(n7739), .A2(n5862), .B1(n6747), .B2(n7738), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9548 ( .A1(n7744), .A2(n5862), .B1(n6559), .B2(n7742), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9549 ( .A1(n7747), .A2(n5862), .B1(n6265), .B2(n7745), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9550 ( .A1(n7759), .A2(n5862), .B1(n6974), .B2(n7761), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9551 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  NAND2_X2 U9552 ( .A1(n4096), .A2(n8946), .ZN(ID_EX_REG_ID_EX_REG_N130) );
  OAI22_X2 U9553 ( .A1(n6241), .A2(n7625), .B1(n7626), .B2(n5863), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9554 ( .A1(n7630), .A2(n5863), .B1(n5970), .B2(n7629), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9555 ( .A1(n7634), .A2(n5863), .B1(n6788), .B2(n7633), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9556 ( .A1(n7638), .A2(n5863), .B1(n5907), .B2(n7637), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9557 ( .A1(n7642), .A2(n5863), .B1(n6080), .B2(n7641), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9558 ( .A1(n7646), .A2(n5863), .B1(n6181), .B2(n7645), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9559 ( .A1(n7650), .A2(n5863), .B1(n6748), .B2(n7649), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9560 ( .A1(n6240), .A2(n7653), .B1(n7654), .B2(n5863), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9561 ( .A1(n6058), .A2(n7656), .B1(n7658), .B2(n5863), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9562 ( .A1(n7662), .A2(n5863), .B1(n6107), .B2(n7661), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9563 ( .A1(n7666), .A2(n5863), .B1(n6692), .B2(n7665), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9564 ( .A1(n6126), .A2(n7668), .B1(n7670), .B2(n5863), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9565 ( .A1(n7674), .A2(n5863), .B1(n6601), .B2(n7673), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9566 ( .A1(n7678), .A2(n5863), .B1(n6391), .B2(n7677), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9567 ( .A1(n7682), .A2(n5863), .B1(n5942), .B2(n7681), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9568 ( .A1(n7686), .A2(n5863), .B1(n6232), .B2(n7685), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9569 ( .A1(n7690), .A2(n5863), .B1(n6262), .B2(n7688), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9570 ( .A1(n7694), .A2(n5863), .B1(n6447), .B2(n7692), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9571 ( .A1(n7698), .A2(n5863), .B1(n5969), .B2(n7697), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9572 ( .A1(n7702), .A2(n5863), .B1(n6789), .B2(n7701), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9573 ( .A1(n7706), .A2(n5863), .B1(n5989), .B2(n7704), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9574 ( .A1(n7710), .A2(n5863), .B1(n6079), .B2(n7708), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9575 ( .A1(n7714), .A2(n5863), .B1(n6790), .B2(n7712), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9576 ( .A1(n7718), .A2(n5863), .B1(n6180), .B2(n7717), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9577 ( .A1(n7722), .A2(n5863), .B1(n7177), .B2(n7721), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9578 ( .A1(n7727), .A2(n5863), .B1(n6622), .B2(n7725), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9579 ( .A1(n3090), .A2(n5863), .B1(n5988), .B2(n7730), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9580 ( .A1(n7735), .A2(n5863), .B1(n6458), .B2(n7734), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9581 ( .A1(n7740), .A2(n5863), .B1(n6749), .B2(n7738), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9582 ( .A1(n7743), .A2(n5863), .B1(n6560), .B2(n7742), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9583 ( .A1(n7747), .A2(n5863), .B1(n6263), .B2(n7745), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U9584 ( .A1(n7759), .A2(n5863), .B1(n6448), .B2(n7761), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U9585 ( .A1(n8948), .A2(n7457), .ZN(n8950) );
  NAND2_X2 U9586 ( .A1(n7458), .A2(n7268), .ZN(n8949) );
  NAND3_X2 U9587 ( .A1(n4817), .A2(n8950), .A3(n8949), .ZN(n10290) );
  AND2_X2 U9588 ( .A1(n10290), .A2(n7774), .ZN(ID_EX_REG_ID_EX_REG_N15) );
  NAND2_X2 U9589 ( .A1(n8952), .A2(n8951), .ZN(n9562) );
  INV_X4 U9590 ( .A(n9886), .ZN(n8963) );
  XNOR2_X2 U9591 ( .A(n9886), .B(n9887), .ZN(n9857) );
  INV_X4 U9592 ( .A(n8966), .ZN(n8970) );
  NAND2_X2 U9593 ( .A1(n6994), .A2(n9843), .ZN(n8969) );
  NAND2_X2 U9594 ( .A1(n8975), .A2(n9544), .ZN(n8968) );
  OAI211_X2 U9595 ( .C1(n9864), .C2(n8970), .A(n8969), .B(n8968), .ZN(n9570)
         );
  INV_X4 U9596 ( .A(n9570), .ZN(n8974) );
  OAI22_X2 U9597 ( .A1(n9877), .A2(n8971), .B1(n9009), .B2(n9182), .ZN(n9549)
         );
  MUX2_X2 U9598 ( .A(n8972), .B(n9549), .S(n9864), .Z(n8973) );
  INV_X4 U9599 ( .A(n8973), .ZN(n8999) );
  OAI22_X2 U9600 ( .A1(n8974), .A2(n10255), .B1(n8999), .B2(n6860), .ZN(n8988)
         );
  INV_X4 U9601 ( .A(n7388), .ZN(n8975) );
  NAND2_X2 U9602 ( .A1(n8975), .A2(n9021), .ZN(n8981) );
  INV_X4 U9603 ( .A(n7386), .ZN(n8976) );
  NAND2_X2 U9604 ( .A1(n8976), .A2(n9537), .ZN(n8980) );
  NAND2_X2 U9605 ( .A1(n7478), .A2(n8977), .ZN(n8979) );
  NAND2_X2 U9606 ( .A1(n10195), .A2(n9120), .ZN(n8978) );
  OAI22_X2 U9607 ( .A1(n7231), .A2(n7392), .B1(n8998), .B2(n7393), .ZN(n8987)
         );
  OAI211_X2 U9608 ( .C1(n10286), .C2(n8991), .A(n8990), .B(n8989), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N90) );
  XNOR2_X2 U9609 ( .A(n8993), .B(n8992), .ZN(n9014) );
  INV_X4 U9610 ( .A(n8994), .ZN(n8997) );
  INV_X4 U9611 ( .A(n8995), .ZN(n8996) );
  OAI22_X2 U9612 ( .A1(n8997), .A2(n6860), .B1(n8996), .B2(n7393), .ZN(n9001)
         );
  OAI22_X2 U9613 ( .A1(n8999), .A2(n10255), .B1(n8998), .B2(n7392), .ZN(n9000)
         );
  INV_X4 U9614 ( .A(n9003), .ZN(n9007) );
  OAI21_X4 U9615 ( .B1(n9007), .B2(n7460), .A(n9005), .ZN(n9008) );
  XNOR2_X2 U9616 ( .A(n9008), .B(n9849), .ZN(n9852) );
  OAI211_X2 U9617 ( .C1(n9014), .C2(n7479), .A(n9013), .B(n9012), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N89) );
  INV_X4 U9618 ( .A(n9964), .ZN(n9015) );
  MUX2_X2 U9619 ( .A(n9018), .B(n9017), .S(n9180), .Z(n9020) );
  NOR2_X4 U9620 ( .A1(n9020), .A2(n9019), .ZN(n9061) );
  NAND2_X2 U9621 ( .A1(n8976), .A2(n9059), .ZN(n9023) );
  NAND2_X2 U9622 ( .A1(n10248), .A2(n9021), .ZN(n9022) );
  INV_X4 U9623 ( .A(n9760), .ZN(n9026) );
  NAND2_X2 U9624 ( .A1(n9753), .A2(n9756), .ZN(n9025) );
  INV_X4 U9625 ( .A(n9182), .ZN(n9027) );
  INV_X4 U9626 ( .A(n7353), .ZN(n10289) );
  NAND2_X2 U9627 ( .A1(n7476), .A2(n9912), .ZN(n9669) );
  INV_X4 U9628 ( .A(n9669), .ZN(n9029) );
  MUX2_X2 U9629 ( .A(n9032), .B(n9031), .S(n9180), .Z(n9033) );
  NAND2_X2 U9630 ( .A1(n9034), .A2(n9033), .ZN(n9808) );
  INV_X4 U9631 ( .A(n9808), .ZN(n9039) );
  NAND2_X2 U9632 ( .A1(n8976), .A2(n9035), .ZN(n9038) );
  NAND2_X2 U9633 ( .A1(n10248), .A2(n9036), .ZN(n9037) );
  OAI211_X2 U9634 ( .C1(n9039), .C2(n7383), .A(n9038), .B(n9037), .ZN(n9040)
         );
  INV_X4 U9635 ( .A(n9040), .ZN(n9065) );
  NAND3_X2 U9636 ( .A1(n7480), .A2(n9047), .A3(n9046), .ZN(n9052) );
  XNOR2_X2 U9637 ( .A(n9871), .B(n9668), .ZN(n9048) );
  INV_X4 U9638 ( .A(n9048), .ZN(n9868) );
  XNOR2_X2 U9639 ( .A(n7366), .B(n7449), .ZN(n9054) );
  XNOR2_X2 U9640 ( .A(n9054), .B(n9786), .ZN(n10085) );
  NAND2_X2 U9641 ( .A1(n7480), .A2(n9058), .ZN(n9074) );
  XNOR2_X2 U9642 ( .A(n9807), .B(n9863), .ZN(n9866) );
  NAND2_X2 U9643 ( .A1(n9143), .A2(n9776), .ZN(n9073) );
  NAND2_X2 U9644 ( .A1(n5852), .A2(n9889), .ZN(n9713) );
  OAI221_X2 U9645 ( .B1(n10105), .B2(n7391), .C1(n9665), .C2(n9804), .A(n9713), 
        .ZN(n9064) );
  AOI211_X4 U9646 ( .C1(n8627), .C2(n9064), .A(n9063), .B(n9062), .ZN(n9818)
         );
  NAND2_X2 U9647 ( .A1(n9618), .A2(n7366), .ZN(n9800) );
  NAND2_X2 U9648 ( .A1(n10257), .A2(n9753), .ZN(n9069) );
  NAND2_X2 U9649 ( .A1(n10264), .A2(n7383), .ZN(n9068) );
  NAND4_X2 U9650 ( .A1(n9074), .A2(n9073), .A3(n9072), .A4(n9071), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N83) );
  INV_X4 U9651 ( .A(n9075), .ZN(n9077) );
  INV_X4 U9652 ( .A(n9500), .ZN(n9076) );
  NAND2_X2 U9653 ( .A1(n9330), .A2(n9499), .ZN(n9084) );
  NAND2_X2 U9654 ( .A1(n7471), .A2(n9079), .ZN(n9080) );
  XNOR2_X2 U9655 ( .A(n9918), .B(n7307), .ZN(n9085) );
  XNOR2_X2 U9656 ( .A(n9085), .B(n9919), .ZN(n9336) );
  INV_X4 U9657 ( .A(n9336), .ZN(n9083) );
  NAND2_X2 U9658 ( .A1(n9084), .A2(n9083), .ZN(n9505) );
  NAND2_X2 U9659 ( .A1(n9085), .A2(n9919), .ZN(n9504) );
  NAND2_X2 U9660 ( .A1(n9505), .A2(n9504), .ZN(n9300) );
  NAND2_X2 U9661 ( .A1(n7471), .A2(n9086), .ZN(n9087) );
  XNOR2_X2 U9662 ( .A(n9929), .B(n7307), .ZN(n9100) );
  XNOR2_X2 U9663 ( .A(n9100), .B(n9930), .ZN(n9495) );
  INV_X4 U9664 ( .A(n9090), .ZN(n9092) );
  NOR2_X4 U9665 ( .A1(n9092), .A2(n9091), .ZN(n9099) );
  INV_X4 U9666 ( .A(n9093), .ZN(n9094) );
  NAND4_X2 U9667 ( .A1(n9095), .A2(n9500), .A3(n9499), .A4(n9504), .ZN(n9096)
         );
  NOR2_X4 U9668 ( .A1(n9097), .A2(n9096), .ZN(n9098) );
  NAND2_X2 U9669 ( .A1(n9100), .A2(n9930), .ZN(n9286) );
  NAND2_X2 U9670 ( .A1(n10223), .A2(n9286), .ZN(n9583) );
  INV_X4 U9671 ( .A(n9583), .ZN(n9105) );
  NAND2_X2 U9672 ( .A1(n7472), .A2(n9101), .ZN(n9137) );
  OAI221_X2 U9673 ( .B1(n7450), .B2(n9137), .C1(n7450), .C2(n9104), .A(n9103), 
        .ZN(n9279) );
  XNOR2_X2 U9674 ( .A(n9105), .B(n9579), .ZN(n9146) );
  NAND2_X2 U9675 ( .A1(n10195), .A2(n10198), .ZN(n9111) );
  NAND2_X2 U9676 ( .A1(n7473), .A2(n9989), .ZN(n9374) );
  NAND2_X2 U9677 ( .A1(n7478), .A2(n10197), .ZN(n9110) );
  NAND2_X2 U9678 ( .A1(n8976), .A2(n10107), .ZN(n9109) );
  NAND2_X2 U9679 ( .A1(n8627), .A2(n9529), .ZN(n9108) );
  NAND2_X2 U9680 ( .A1(n7478), .A2(n9591), .ZN(n9117) );
  NAND2_X2 U9681 ( .A1(n7475), .A2(n9853), .ZN(n9113) );
  NAND2_X2 U9682 ( .A1(n9113), .A2(n9112), .ZN(n10239) );
  NAND2_X2 U9683 ( .A1(n8627), .A2(n10239), .ZN(n9116) );
  NAND2_X2 U9684 ( .A1(n8976), .A2(n10238), .ZN(n9115) );
  NAND2_X2 U9685 ( .A1(n10248), .A2(n9544), .ZN(n9114) );
  NAND4_X2 U9686 ( .A1(n9117), .A2(n9116), .A3(n9115), .A4(n9114), .ZN(n9516)
         );
  NAND2_X2 U9687 ( .A1(n9618), .A2(n9516), .ZN(n9118) );
  NAND2_X2 U9688 ( .A1(n8976), .A2(n9599), .ZN(n9124) );
  NAND2_X2 U9689 ( .A1(n7475), .A2(n7351), .ZN(n9119) );
  NAND2_X2 U9690 ( .A1(n7473), .A2(n10163), .ZN(n9365) );
  NAND2_X2 U9691 ( .A1(n10248), .A2(n10249), .ZN(n9123) );
  NAND2_X2 U9692 ( .A1(n8975), .A2(n9120), .ZN(n9122) );
  NAND2_X2 U9693 ( .A1(n7478), .A2(n10250), .ZN(n9121) );
  NAND4_X2 U9694 ( .A1(n9124), .A2(n9123), .A3(n9122), .A4(n9121), .ZN(n9512)
         );
  INV_X4 U9695 ( .A(n9512), .ZN(n9134) );
  NAND2_X2 U9696 ( .A1(n7475), .A2(n9894), .ZN(n9126) );
  NAND2_X2 U9697 ( .A1(n9126), .A2(n9125), .ZN(n10205) );
  NAND2_X2 U9698 ( .A1(n5864), .A2(n10205), .ZN(n9132) );
  NAND2_X2 U9699 ( .A1(n9128), .A2(n9127), .ZN(n10206) );
  NAND2_X2 U9700 ( .A1(n8975), .A2(n10206), .ZN(n9131) );
  NAND2_X2 U9701 ( .A1(n10248), .A2(n9550), .ZN(n9130) );
  NAND2_X2 U9702 ( .A1(n7478), .A2(n10112), .ZN(n9129) );
  NAND4_X2 U9703 ( .A1(n9132), .A2(n9131), .A3(n9130), .A4(n9129), .ZN(n9604)
         );
  NAND2_X2 U9704 ( .A1(n9753), .A2(n9604), .ZN(n9133) );
  NAND2_X2 U9705 ( .A1(ID_EXEC_OUT[80]), .A2(n5855), .ZN(n9138) );
  XNOR2_X2 U9706 ( .A(n9926), .B(n9927), .ZN(n9139) );
  INV_X4 U9707 ( .A(n9139), .ZN(n9941) );
  OAI211_X2 U9708 ( .C1(n9146), .C2(n7479), .A(n9145), .B(n9144), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N97) );
  INV_X4 U9709 ( .A(n9930), .ZN(n9148) );
  NAND2_X2 U9710 ( .A1(n7473), .A2(n9977), .ZN(n9705) );
  NAND2_X2 U9711 ( .A1(n9189), .A2(n7366), .ZN(n9151) );
  NAND4_X2 U9712 ( .A1(n9153), .A2(n9705), .A3(n9152), .A4(n9151), .ZN(n9667)
         );
  OAI221_X2 U9713 ( .B1(n9156), .B2(n9804), .C1(n9155), .C2(n7391), .A(n9154), 
        .ZN(n9157) );
  MUX2_X2 U9714 ( .A(n9667), .B(n9157), .S(n9180), .Z(n9160) );
  NAND2_X2 U9715 ( .A1(n7390), .A2(n9912), .ZN(n9162) );
  NAND4_X2 U9716 ( .A1(n9163), .A2(n9641), .A3(n9162), .A4(n9161), .ZN(n9436)
         );
  OAI221_X2 U9717 ( .B1(n9168), .B2(n7388), .C1(n9864), .C2(n9438), .A(n9167), 
        .ZN(n9410) );
  NAND2_X2 U9718 ( .A1(ID_EXEC_OUT[64]), .A2(n5855), .ZN(n9171) );
  NAND2_X2 U9719 ( .A1(n7471), .A2(n9169), .ZN(n9170) );
  OAI211_X2 U9720 ( .C1(n5888), .C2(n9293), .A(n9171), .B(n9170), .ZN(n10033)
         );
  XNOR2_X2 U9721 ( .A(n10033), .B(n9318), .ZN(n10051) );
  NAND2_X2 U9722 ( .A1(n9412), .A2(n9173), .ZN(n9206) );
  INV_X4 U9723 ( .A(n10274), .ZN(n9517) );
  NAND2_X2 U9724 ( .A1(n7473), .A2(n9974), .ZN(n9677) );
  NAND2_X2 U9725 ( .A1(n7390), .A2(n9889), .ZN(n9175) );
  NAND4_X2 U9726 ( .A1(n9176), .A2(n9677), .A3(n9175), .A4(n9174), .ZN(n9631)
         );
  INV_X4 U9727 ( .A(n9919), .ZN(n9178) );
  OAI221_X2 U9728 ( .B1(n9179), .B2(n9804), .C1(n9178), .C2(n7391), .A(n9177), 
        .ZN(n9181) );
  MUX2_X2 U9729 ( .A(n9631), .B(n9181), .S(n9180), .Z(n9185) );
  INV_X4 U9730 ( .A(n7351), .ZN(n9183) );
  NAND2_X2 U9731 ( .A1(n9815), .A2(n9318), .ZN(n9194) );
  NAND2_X2 U9732 ( .A1(n7390), .A2(n9909), .ZN(n9188) );
  NAND2_X2 U9733 ( .A1(n7473), .A2(n9964), .ZN(n9353) );
  NAND4_X2 U9734 ( .A1(n9188), .A2(n9187), .A3(n9186), .A4(n9353), .ZN(n9413)
         );
  OAI211_X2 U9735 ( .C1(n9864), .C2(n9414), .A(n9194), .B(n9193), .ZN(n9204)
         );
  NAND2_X2 U9736 ( .A1(n7473), .A2(n9318), .ZN(n9196) );
  NAND2_X2 U9737 ( .A1(n9412), .A2(n9195), .ZN(n9704) );
  INV_X4 U9738 ( .A(n10279), .ZN(n9441) );
  NAND2_X2 U9739 ( .A1(n9441), .A2(n8627), .ZN(n9202) );
  INV_X4 U9740 ( .A(n9197), .ZN(n9199) );
  NAND2_X2 U9741 ( .A1(n6023), .A2(n9318), .ZN(n9198) );
  NAND2_X2 U9742 ( .A1(n9200), .A2(n10033), .ZN(n9201) );
  INV_X4 U9743 ( .A(n9318), .ZN(n10034) );
  NAND2_X2 U9744 ( .A1(ID_EXEC_OUT[66]), .A2(n5855), .ZN(n9219) );
  NAND2_X2 U9745 ( .A1(n7471), .A2(n9215), .ZN(n9218) );
  INV_X4 U9746 ( .A(n7313), .ZN(n9216) );
  NAND2_X2 U9747 ( .A1(n9216), .A2(DMEM_BUS_OUT[2]), .ZN(n9217) );
  NAND3_X4 U9748 ( .A1(n9219), .A2(n9218), .A3(n9217), .ZN(n9445) );
  XNOR2_X2 U9749 ( .A(n9445), .B(n7449), .ZN(n9314) );
  NAND2_X2 U9750 ( .A1(n9314), .A2(n7351), .ZN(n9404) );
  NAND2_X2 U9751 ( .A1(n9221), .A2(n9404), .ZN(n9222) );
  NAND2_X2 U9752 ( .A1(n9400), .A2(n9221), .ZN(n9315) );
  NAND2_X2 U9753 ( .A1(n9222), .A2(n9315), .ZN(n9316) );
  XNOR2_X2 U9754 ( .A(n9477), .B(n7307), .ZN(n9229) );
  NAND2_X2 U9755 ( .A1(ID_EXEC_OUT[68]), .A2(n5855), .ZN(n9232) );
  NAND2_X2 U9756 ( .A1(n7472), .A2(n9230), .ZN(n9231) );
  OAI211_X2 U9757 ( .C1(n5925), .C2(n7313), .A(n9232), .B(n9231), .ZN(n9385)
         );
  XNOR2_X2 U9758 ( .A(n9385), .B(n7307), .ZN(n9233) );
  NAND2_X2 U9759 ( .A1(n9233), .A2(n9964), .ZN(n9489) );
  INV_X4 U9760 ( .A(n9488), .ZN(n9479) );
  XNOR2_X2 U9761 ( .A(n9233), .B(n9964), .ZN(n9482) );
  INV_X4 U9762 ( .A(n9482), .ZN(n9449) );
  NAND2_X2 U9763 ( .A1(n9479), .A2(n9449), .ZN(n9311) );
  NAND2_X2 U9764 ( .A1(ID_EXEC_OUT[69]), .A2(n5855), .ZN(n9236) );
  NAND2_X2 U9765 ( .A1(n7471), .A2(n9234), .ZN(n9235) );
  OAI22_X2 U9766 ( .A1(n9488), .A2(n9489), .B1(n9311), .B2(n9448), .ZN(n9401)
         );
  INV_X4 U9767 ( .A(n9237), .ZN(n9238) );
  AOI22_X2 U9768 ( .A1(n7471), .A2(n9239), .B1(n9238), .B2(n7471), .ZN(n9240)
         );
  XNOR2_X2 U9769 ( .A(n9978), .B(n7307), .ZN(n9258) );
  INV_X4 U9770 ( .A(n9736), .ZN(n9264) );
  OAI211_X2 U9771 ( .C1(n9245), .C2(n7468), .A(n9244), .B(n9243), .ZN(n10134)
         );
  XNOR2_X2 U9772 ( .A(n10134), .B(n7307), .ZN(n9257) );
  NAND2_X2 U9773 ( .A1(n9257), .A2(n10135), .ZN(n9733) );
  INV_X4 U9774 ( .A(n9733), .ZN(n9692) );
  NAND2_X2 U9775 ( .A1(ID_EXEC_OUT[74]), .A2(n5855), .ZN(n9248) );
  NAND2_X2 U9776 ( .A1(n7472), .A2(n9246), .ZN(n9247) );
  XNOR2_X2 U9777 ( .A(n10164), .B(n7307), .ZN(n9254) );
  INV_X4 U9778 ( .A(n9732), .ZN(n10129) );
  NAND2_X2 U9779 ( .A1(ID_EXEC_OUT[75]), .A2(n5855), .ZN(n9251) );
  INV_X4 U9780 ( .A(n10128), .ZN(n10167) );
  XNOR2_X2 U9781 ( .A(n9252), .B(n9989), .ZN(n9253) );
  INV_X4 U9782 ( .A(n9253), .ZN(n10189) );
  XNOR2_X2 U9783 ( .A(n9254), .B(n10163), .ZN(n10168) );
  INV_X4 U9784 ( .A(n10168), .ZN(n9255) );
  OAI21_X4 U9785 ( .B1(n10167), .B2(n10189), .A(n9255), .ZN(n9256) );
  INV_X4 U9786 ( .A(n9694), .ZN(n9259) );
  OAI21_X4 U9787 ( .B1(n9692), .B2(n7326), .A(n9259), .ZN(n9737) );
  INV_X4 U9788 ( .A(n9737), .ZN(n9263) );
  OAI21_X4 U9789 ( .B1(n9264), .B2(n9263), .A(n6989), .ZN(n9653) );
  NAND2_X2 U9790 ( .A1(n9265), .A2(n9977), .ZN(n9304) );
  NAND2_X2 U9791 ( .A1(ID_EXEC_OUT[70]), .A2(n5855), .ZN(n9268) );
  NAND2_X2 U9792 ( .A1(n7472), .A2(n9266), .ZN(n9267) );
  XNOR2_X2 U9793 ( .A(n9310), .B(n9974), .ZN(n9663) );
  INV_X4 U9794 ( .A(n9269), .ZN(n9274) );
  NAND3_X2 U9795 ( .A1(n7380), .A2(DMEM_BUS_OUT[13]), .A3(n7468), .ZN(n9272)
         );
  NAND3_X2 U9796 ( .A1(ID_EXEC_OUT[77]), .A2(n7381), .A3(n7468), .ZN(n9271) );
  OAI211_X2 U9797 ( .C1(n9274), .C2(n7468), .A(n9272), .B(n9271), .ZN(n10263)
         );
  XNOR2_X2 U9798 ( .A(n10263), .B(n7307), .ZN(n9288) );
  XNOR2_X2 U9799 ( .A(n9288), .B(n7353), .ZN(n10269) );
  NAND2_X2 U9800 ( .A1(ID_EXEC_OUT[78]), .A2(n5855), .ZN(n9277) );
  XNOR2_X2 U9801 ( .A(n10104), .B(n7307), .ZN(n9278) );
  INV_X4 U9802 ( .A(n9297), .ZN(n10103) );
  NAND2_X2 U9803 ( .A1(n9579), .A2(n9580), .ZN(n9284) );
  NAND2_X2 U9804 ( .A1(ID_EXEC_OUT[79]), .A2(n5855), .ZN(n9282) );
  OAI211_X2 U9805 ( .C1(n9293), .C2(n6042), .A(n9282), .B(n9281), .ZN(n9924)
         );
  XNOR2_X2 U9806 ( .A(n9924), .B(n7307), .ZN(n9285) );
  XNOR2_X2 U9807 ( .A(n9285), .B(n9925), .ZN(n9584) );
  INV_X4 U9808 ( .A(n9584), .ZN(n9283) );
  NAND2_X2 U9809 ( .A1(n9580), .A2(n9286), .ZN(n10098) );
  INV_X4 U9810 ( .A(n10098), .ZN(n9287) );
  NAND2_X2 U9811 ( .A1(n9287), .A2(n10099), .ZN(n10218) );
  INV_X4 U9812 ( .A(n10269), .ZN(n9295) );
  NAND2_X2 U9813 ( .A1(n10218), .A2(n9295), .ZN(n9289) );
  OAI221_X2 U9814 ( .B1(n10269), .B2(n10219), .C1(n10265), .C2(n9289), .A(
        n10221), .ZN(n9294) );
  NAND2_X2 U9815 ( .A1(ID_EXEC_OUT[76]), .A2(n5855), .ZN(n9292) );
  NAND2_X2 U9816 ( .A1(n7471), .A2(n9290), .ZN(n9291) );
  XNOR2_X2 U9817 ( .A(n10228), .B(n7307), .ZN(n9303) );
  INV_X4 U9818 ( .A(n10226), .ZN(n9296) );
  NAND2_X2 U9819 ( .A1(n9296), .A2(n9295), .ZN(n9298) );
  NAND3_X2 U9820 ( .A1(n10128), .A2(n9656), .A3(n9732), .ZN(n9305) );
  INV_X4 U9821 ( .A(n9304), .ZN(n9660) );
  NAND2_X2 U9822 ( .A1(n9733), .A2(n9736), .ZN(n9654) );
  NOR3_X4 U9823 ( .A1(n9389), .A2(n9626), .A3(n9311), .ZN(n9313) );
  NAND2_X2 U9824 ( .A1(n9310), .A2(n9974), .ZN(n9388) );
  NOR2_X4 U9825 ( .A1(n9313), .A2(n9312), .ZN(n9402) );
  INV_X4 U9826 ( .A(n9324), .ZN(n9327) );
  XNOR2_X2 U9827 ( .A(n9314), .B(n7351), .ZN(n9459) );
  INV_X4 U9828 ( .A(n9459), .ZN(n9447) );
  NAND2_X2 U9829 ( .A1(n9315), .A2(n9447), .ZN(n9317) );
  NAND2_X2 U9830 ( .A1(n9317), .A2(n9316), .ZN(n9320) );
  XNOR2_X2 U9831 ( .A(n9318), .B(n7307), .ZN(n9319) );
  XNOR2_X2 U9832 ( .A(n9319), .B(n10033), .ZN(n9321) );
  INV_X4 U9833 ( .A(n9321), .ZN(n9325) );
  NAND2_X2 U9834 ( .A1(n9320), .A2(n9325), .ZN(n9326) );
  INV_X4 U9835 ( .A(n9320), .ZN(n9322) );
  OAI221_X2 U9836 ( .B1(n9327), .B2(n9326), .C1(n9324), .C2(n9325), .A(n9323), 
        .ZN(n9328) );
  NAND2_X2 U9837 ( .A1(n9329), .A2(n9328), .ZN(n10298) );
  INV_X4 U9838 ( .A(n9330), .ZN(n9335) );
  INV_X4 U9839 ( .A(n9331), .ZN(n9332) );
  INV_X4 U9840 ( .A(n9499), .ZN(n9333) );
  XNOR2_X2 U9841 ( .A(n9337), .B(n9336), .ZN(n9352) );
  INV_X4 U9842 ( .A(n9918), .ZN(n9338) );
  NAND2_X2 U9843 ( .A1(n9339), .A2(n9919), .ZN(n9351) );
  NAND2_X2 U9844 ( .A1(n8976), .A2(n9529), .ZN(n9344) );
  NAND2_X2 U9845 ( .A1(n10248), .A2(n10197), .ZN(n9343) );
  NAND2_X2 U9846 ( .A1(n9813), .A2(n9340), .ZN(n9342) );
  NAND2_X2 U9847 ( .A1(n7478), .A2(n10107), .ZN(n9341) );
  OAI22_X2 U9848 ( .A1(n6807), .A2(n10281), .B1(n6185), .B2(n9646), .ZN(n9349)
         );
  XNOR2_X2 U9849 ( .A(n9918), .B(n9919), .ZN(n9940) );
  AOI22_X2 U9850 ( .A1(n9813), .A2(n10205), .B1(n7478), .B2(n9550), .ZN(n9345)
         );
  NAND2_X2 U9851 ( .A1(n9517), .A2(n9511), .ZN(n9347) );
  OAI221_X2 U9852 ( .B1(n9940), .B2(n9742), .C1(n6805), .C2(n10279), .A(n9347), 
        .ZN(n9348) );
  OAI211_X2 U9853 ( .C1(n7479), .C2(n9352), .A(n9351), .B(n9350), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N95) );
  NAND2_X2 U9854 ( .A1(n10248), .A2(n9412), .ZN(n9639) );
  NAND2_X2 U9855 ( .A1(n9353), .A2(n9704), .ZN(n10172) );
  INV_X4 U9856 ( .A(n10172), .ZN(n9721) );
  INV_X4 U9857 ( .A(n9704), .ZN(n9354) );
  AOI21_X4 U9858 ( .B1(n7473), .B2(n7351), .A(n9354), .ZN(n9722) );
  INV_X4 U9859 ( .A(n9645), .ZN(n9358) );
  NAND2_X2 U9860 ( .A1(n6800), .A2(n9358), .ZN(n9382) );
  NAND2_X2 U9861 ( .A1(n9359), .A2(n9704), .ZN(n9411) );
  INV_X4 U9862 ( .A(n9411), .ZN(n9703) );
  NAND2_X2 U9863 ( .A1(n9360), .A2(n9704), .ZN(n10148) );
  OAI221_X2 U9864 ( .B1(n9703), .B2(n7386), .C1(n9640), .C2(n9806), .A(n9440), 
        .ZN(n9469) );
  NAND2_X2 U9865 ( .A1(n6799), .A2(n9469), .ZN(n9381) );
  NAND2_X2 U9866 ( .A1(n8975), .A2(n9413), .ZN(n9368) );
  NAND2_X2 U9867 ( .A1(n7390), .A2(n9894), .ZN(n9366) );
  AOI22_X2 U9868 ( .A1(n7478), .A2(n9714), .B1(n10195), .B2(n10138), .ZN(n9367) );
  NAND3_X4 U9869 ( .A1(n9369), .A2(n9368), .A3(n9367), .ZN(n9470) );
  NAND2_X2 U9870 ( .A1(n9753), .A2(n9470), .ZN(n9380) );
  NAND2_X2 U9871 ( .A1(n9813), .A2(n9436), .ZN(n9378) );
  NAND2_X2 U9872 ( .A1(n5864), .A2(n9667), .ZN(n9377) );
  NAND2_X2 U9873 ( .A1(n7390), .A2(n9853), .ZN(n9372) );
  NAND2_X2 U9874 ( .A1(n7390), .A2(n9843), .ZN(n9375) );
  AOI22_X2 U9875 ( .A1(n7478), .A2(n9698), .B1(n10248), .B2(n10177), .ZN(n9376) );
  NAND2_X2 U9876 ( .A1(n9618), .A2(n9628), .ZN(n9379) );
  NAND4_X2 U9877 ( .A1(n9382), .A2(n9381), .A3(n9380), .A4(n9379), .ZN(n9383)
         );
  NAND2_X2 U9878 ( .A1(n10257), .A2(n9383), .ZN(n9399) );
  XNOR2_X2 U9879 ( .A(n9385), .B(n9964), .ZN(n10048) );
  INV_X4 U9880 ( .A(n10048), .ZN(n9384) );
  NAND2_X2 U9881 ( .A1(n9143), .A2(n9384), .ZN(n9398) );
  INV_X4 U9882 ( .A(n9385), .ZN(n9965) );
  NAND2_X2 U9883 ( .A1(n9386), .A2(n9964), .ZN(n9397) );
  INV_X4 U9884 ( .A(n9448), .ZN(n9387) );
  NAND2_X2 U9885 ( .A1(n6798), .A2(n9626), .ZN(n9394) );
  INV_X4 U9886 ( .A(n9626), .ZN(n9390) );
  NAND2_X2 U9887 ( .A1(n9389), .A2(n9388), .ZN(n9627) );
  NAND2_X2 U9888 ( .A1(n6798), .A2(n9391), .ZN(n9392) );
  NAND4_X2 U9889 ( .A1(n9395), .A2(n9394), .A3(n9393), .A4(n9392), .ZN(n9396)
         );
  NAND4_X2 U9890 ( .A1(n9396), .A2(n9398), .A3(n9397), .A4(n9399), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N109) );
  INV_X4 U9891 ( .A(n9400), .ZN(n9409) );
  NAND2_X2 U9892 ( .A1(n9459), .A2(n9404), .ZN(n9405) );
  INV_X4 U9893 ( .A(n9401), .ZN(n9403) );
  NAND2_X2 U9894 ( .A1(n9405), .A2(n9409), .ZN(n9406) );
  OAI22_X2 U9895 ( .A1(n9409), .A2(n9408), .B1(n9407), .B2(n9406), .ZN(n9430)
         );
  NAND2_X2 U9896 ( .A1(n9753), .A2(n9410), .ZN(n9423) );
  MUX2_X2 U9897 ( .A(n9412), .B(n9411), .S(n7387), .Z(n9432) );
  NAND2_X2 U9898 ( .A1(n6800), .A2(n9432), .ZN(n9422) );
  NAND2_X2 U9899 ( .A1(n10195), .A2(n9714), .ZN(n9416) );
  NAND2_X2 U9900 ( .A1(n9413), .A2(n10147), .ZN(n9415) );
  INV_X4 U9901 ( .A(n9418), .ZN(n9419) );
  NAND3_X2 U9902 ( .A1(n9423), .A2(n9422), .A3(n9421), .ZN(n9428) );
  XNOR2_X2 U9903 ( .A(n9424), .B(n9970), .ZN(n10050) );
  INV_X4 U9904 ( .A(n9432), .ZN(n9435) );
  NAND2_X2 U9905 ( .A1(n9517), .A2(n9433), .ZN(n9434) );
  XNOR2_X2 U9906 ( .A(n9445), .B(n9968), .ZN(n10052) );
  INV_X4 U9907 ( .A(n9698), .ZN(n9439) );
  NAND2_X2 U9908 ( .A1(n10147), .A2(n9436), .ZN(n9437) );
  OAI221_X2 U9909 ( .B1(n9439), .B2(n10246), .C1(n9438), .C2(n7383), .A(n9437), 
        .ZN(n9466) );
  OAI221_X2 U9910 ( .B1(n9722), .B2(n7388), .C1(n6350), .C2(n7385), .A(n9440), 
        .ZN(n9471) );
  NAND2_X2 U9911 ( .A1(n9441), .A2(n9471), .ZN(n9442) );
  OAI221_X2 U9912 ( .B1(n10052), .B2(n9742), .C1(n9468), .C2(n9646), .A(n9442), 
        .ZN(n9443) );
  INV_X4 U9913 ( .A(n9445), .ZN(n9969) );
  NAND2_X2 U9914 ( .A1(n9446), .A2(n7351), .ZN(n9456) );
  NAND2_X2 U9915 ( .A1(n6916), .A2(n9447), .ZN(n9458) );
  NAND2_X2 U9916 ( .A1(n9488), .A2(n9452), .ZN(n9453) );
  NAND2_X2 U9917 ( .A1(n9626), .A2(n9448), .ZN(n9480) );
  INV_X4 U9918 ( .A(n9462), .ZN(n9451) );
  NAND2_X2 U9919 ( .A1(n9452), .A2(n9489), .ZN(n9454) );
  NAND2_X2 U9920 ( .A1(n9454), .A2(n9453), .ZN(n9460) );
  INV_X4 U9921 ( .A(n9466), .ZN(n9468) );
  XNOR2_X2 U9922 ( .A(n9477), .B(n9966), .ZN(n9788) );
  INV_X4 U9923 ( .A(n9788), .ZN(n9982) );
  NAND2_X2 U9924 ( .A1(n10272), .A2(n9982), .ZN(n9467) );
  INV_X4 U9925 ( .A(n9469), .ZN(n9474) );
  INV_X4 U9926 ( .A(n10281), .ZN(n9513) );
  NAND2_X2 U9927 ( .A1(n9513), .A2(n9471), .ZN(n9472) );
  OAI21_X4 U9928 ( .B1(n9476), .B2(n9475), .A(n10282), .ZN(n9484) );
  INV_X4 U9929 ( .A(n9477), .ZN(n9967) );
  INV_X4 U9930 ( .A(n9480), .ZN(n9481) );
  NOR3_X4 U9931 ( .A1(n7324), .A2(n9482), .A3(n9481), .ZN(n9491) );
  INV_X4 U9932 ( .A(n9495), .ZN(n9508) );
  XNOR2_X2 U9933 ( .A(n9508), .B(n9507), .ZN(n9523) );
  INV_X4 U9934 ( .A(n9929), .ZN(n9509) );
  NAND2_X2 U9935 ( .A1(n9510), .A2(n9930), .ZN(n9522) );
  INV_X4 U9936 ( .A(n9511), .ZN(n9515) );
  NAND2_X2 U9937 ( .A1(n9513), .A2(n9512), .ZN(n9514) );
  XNOR2_X2 U9938 ( .A(n9929), .B(n9930), .ZN(n9943) );
  NAND2_X2 U9939 ( .A1(n9517), .A2(n9516), .ZN(n9518) );
  OAI221_X2 U9940 ( .B1(n9943), .B2(n9742), .C1(n6807), .C2(n10279), .A(n9518), 
        .ZN(n9519) );
  OAI211_X2 U9941 ( .C1(n7479), .C2(n9523), .A(n9522), .B(n9521), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N96) );
  XNOR2_X2 U9942 ( .A(n9911), .B(n9912), .ZN(n9901) );
  INV_X4 U9943 ( .A(n9524), .ZN(n9525) );
  NAND2_X2 U9944 ( .A1(n9526), .A2(n9525), .ZN(n9613) );
  INV_X4 U9945 ( .A(n9613), .ZN(n9528) );
  AOI22_X2 U9946 ( .A1(n9813), .A2(n9530), .B1(n10248), .B2(n9529), .ZN(n9536)
         );
  AOI22_X2 U9947 ( .A1(n8627), .A2(n9537), .B1(n10195), .B2(n9599), .ZN(n9543)
         );
  NAND2_X2 U9948 ( .A1(n7001), .A2(n9843), .ZN(n9548) );
  NAND2_X2 U9949 ( .A1(n6994), .A2(n9853), .ZN(n9547) );
  NAND2_X2 U9950 ( .A1(n10147), .A2(n9544), .ZN(n9546) );
  NAND2_X2 U9951 ( .A1(n9813), .A2(n9591), .ZN(n9545) );
  NAND4_X2 U9952 ( .A1(n9548), .A2(n9547), .A3(n9546), .A4(n9545), .ZN(n9617)
         );
  INV_X4 U9953 ( .A(n9549), .ZN(n9553) );
  NAND2_X2 U9954 ( .A1(n6994), .A2(n9894), .ZN(n9552) );
  NAND2_X2 U9955 ( .A1(n9813), .A2(n9550), .ZN(n9551) );
  OAI211_X2 U9956 ( .C1(n9864), .C2(n9553), .A(n9552), .B(n9551), .ZN(n9571)
         );
  AOI22_X2 U9957 ( .A1(n9753), .A2(n9617), .B1(n9618), .B2(n9571), .ZN(n9554)
         );
  OAI221_X2 U9958 ( .B1(n6806), .B2(n7393), .C1(n6317), .C2(n7392), .A(n9554), 
        .ZN(n9558) );
  NAND2_X2 U9959 ( .A1(n10264), .A2(n9911), .ZN(n9556) );
  INV_X4 U9960 ( .A(n9912), .ZN(n9555) );
  OAI221_X2 U9961 ( .B1(n9901), .B2(n6861), .C1(n9560), .C2(n7479), .A(n9559), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N92) );
  XNOR2_X2 U9962 ( .A(n9888), .B(n9889), .ZN(n9900) );
  INV_X4 U9963 ( .A(n9561), .ZN(n9567) );
  NAND3_X2 U9964 ( .A1(n9563), .A2(n9562), .A3(n7226), .ZN(n9566) );
  INV_X4 U9965 ( .A(n9564), .ZN(n9565) );
  AOI22_X2 U9966 ( .A1(n9753), .A2(n9571), .B1(n9618), .B2(n9570), .ZN(n9572)
         );
  OAI221_X2 U9967 ( .B1(n6806), .B2(n7392), .C1(n7231), .C2(n7393), .A(n9572), 
        .ZN(n9576) );
  NAND2_X2 U9968 ( .A1(n10264), .A2(n9888), .ZN(n9574) );
  INV_X4 U9969 ( .A(n9889), .ZN(n9573) );
  INV_X4 U9970 ( .A(n9579), .ZN(n9582) );
  INV_X4 U9971 ( .A(n9580), .ZN(n9581) );
  NAND2_X2 U9972 ( .A1(n9925), .A2(n9587), .ZN(n9609) );
  NAND2_X2 U9973 ( .A1(n10147), .A2(n10239), .ZN(n9595) );
  NAND2_X2 U9974 ( .A1(n7390), .A2(n7366), .ZN(n9589) );
  NAND2_X2 U9975 ( .A1(n8627), .A2(n10236), .ZN(n9594) );
  NAND2_X2 U9976 ( .A1(n7478), .A2(n10238), .ZN(n9593) );
  NAND2_X2 U9977 ( .A1(n10248), .A2(n9591), .ZN(n9592) );
  NAND2_X2 U9978 ( .A1(n7478), .A2(n10249), .ZN(n9603) );
  NAND2_X2 U9979 ( .A1(n10248), .A2(n10245), .ZN(n9602) );
  NAND2_X2 U9980 ( .A1(n10147), .A2(n10250), .ZN(n9601) );
  NAND2_X2 U9981 ( .A1(n8627), .A2(n9599), .ZN(n9600) );
  NAND2_X2 U9982 ( .A1(n10277), .A2(n9604), .ZN(n9605) );
  OAI221_X2 U9983 ( .B1(n6482), .B2(n10279), .C1(n7138), .C2(n10281), .A(n9605), .ZN(n9606) );
  OAI211_X2 U9984 ( .C1(n7479), .C2(n9610), .A(n9609), .B(n9608), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N98) );
  XNOR2_X2 U9985 ( .A(n9908), .B(n9909), .ZN(n9913) );
  AOI22_X2 U9986 ( .A1(n9618), .A2(n9617), .B1(n9753), .B2(n9616), .ZN(n9619)
         );
  OAI221_X2 U9987 ( .B1(n6317), .B2(n7393), .C1(n7230), .C2(n7392), .A(n9619), 
        .ZN(n9623) );
  INV_X4 U9988 ( .A(n9909), .ZN(n9620) );
  OAI221_X2 U9989 ( .B1(n9913), .B2(n6861), .C1(n9625), .C2(n7479), .A(n9624), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N93) );
  INV_X4 U9990 ( .A(n9628), .ZN(n9630) );
  XNOR2_X2 U9991 ( .A(n9986), .B(n9987), .ZN(n10046) );
  NAND2_X2 U9992 ( .A1(n7478), .A2(n10138), .ZN(n9637) );
  AOI22_X2 U9993 ( .A1(n10195), .A2(n10203), .B1(n8976), .B2(n9714), .ZN(n9636) );
  INV_X4 U9994 ( .A(n10148), .ZN(n9640) );
  NAND2_X2 U9995 ( .A1(n9641), .A2(n9704), .ZN(n10194) );
  INV_X4 U9996 ( .A(n10194), .ZN(n9707) );
  OAI222_X2 U9997 ( .A1(n7035), .A2(n9646), .B1(n9645), .B2(n10281), .C1(n9681), .C2(n10279), .ZN(n9647) );
  OAI221_X2 U9998 ( .B1(n9652), .B2(n9651), .C1(n9650), .C2(n7479), .A(n9649), 
        .ZN(EX_MEM_REGISTER_EX_MEM_REG_N108) );
  XNOR2_X2 U9999 ( .A(n9973), .B(n9974), .ZN(n10013) );
  INV_X4 U10000 ( .A(n9654), .ZN(n9659) );
  NAND2_X2 U10001 ( .A1(n9732), .A2(n10128), .ZN(n9657) );
  XNOR2_X2 U10002 ( .A(n9664), .B(n9663), .ZN(n9689) );
  NAND2_X2 U10003 ( .A1(n8627), .A2(n9667), .ZN(n9674) );
  NAND2_X2 U10004 ( .A1(n7478), .A2(n10177), .ZN(n9673) );
  AOI22_X2 U10005 ( .A1(n10195), .A2(n10237), .B1(n8976), .B2(n9698), .ZN(
        n9672) );
  NAND2_X2 U10006 ( .A1(n9677), .A2(n9704), .ZN(n10247) );
  INV_X4 U10007 ( .A(n10247), .ZN(n9719) );
  NAND2_X2 U10008 ( .A1(n10166), .A2(n10128), .ZN(n9734) );
  INV_X4 U10009 ( .A(n9734), .ZN(n9691) );
  XNOR2_X2 U10010 ( .A(n9695), .B(n9694), .ZN(n9731) );
  XNOR2_X2 U10011 ( .A(n9978), .B(n9979), .ZN(n10012) );
  NAND2_X2 U10012 ( .A1(n10248), .A2(n10236), .ZN(n9702) );
  NAND2_X2 U10013 ( .A1(n10146), .A2(n10237), .ZN(n9701) );
  NAND2_X2 U10014 ( .A1(n10147), .A2(n10177), .ZN(n9700) );
  NAND2_X2 U10015 ( .A1(n9813), .A2(n9698), .ZN(n9699) );
  NAND2_X2 U10016 ( .A1(n9705), .A2(n9704), .ZN(n10196) );
  INV_X4 U10017 ( .A(n10196), .ZN(n9706) );
  OAI22_X2 U10018 ( .A1(n7208), .A2(n6860), .B1(n9746), .B2(n7392), .ZN(n9728)
         );
  NAND2_X2 U10019 ( .A1(n5884), .A2(n10203), .ZN(n9718) );
  NAND2_X2 U10020 ( .A1(n10248), .A2(n10204), .ZN(n9717) );
  NAND2_X2 U10021 ( .A1(n5864), .A2(n10138), .ZN(n9716) );
  NAND2_X2 U10022 ( .A1(n9813), .A2(n9714), .ZN(n9715) );
  NAND4_X2 U10023 ( .A1(n9718), .A2(n9717), .A3(n9716), .A4(n9715), .ZN(n9743)
         );
  INV_X4 U10024 ( .A(n9743), .ZN(n9726) );
  INV_X4 U10025 ( .A(n10245), .ZN(n9720) );
  OAI22_X2 U10026 ( .A1(n7388), .A2(n9720), .B1(n9719), .B2(n7386), .ZN(n9725)
         );
  OAI22_X2 U10027 ( .A1(n10255), .A2(n9726), .B1(n10143), .B2(n7393), .ZN(
        n9727) );
  OAI211_X2 U10028 ( .C1(n9731), .C2(n7479), .A(n9730), .B(n9729), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N105) );
  XNOR2_X2 U10029 ( .A(n6989), .B(n9739), .ZN(n9751) );
  NAND2_X2 U10030 ( .A1(n9741), .A2(n9977), .ZN(n9750) );
  XNOR2_X2 U10031 ( .A(n9976), .B(n9977), .ZN(n10011) );
  NAND2_X2 U10032 ( .A1(n10277), .A2(n9743), .ZN(n9744) );
  OAI221_X2 U10033 ( .B1(n9746), .B2(n10279), .C1(n9745), .C2(n10281), .A(
        n9744), .ZN(n9747) );
  OAI211_X2 U10034 ( .C1(n7479), .C2(n9751), .A(n9750), .B(n9749), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N106) );
  NAND2_X2 U10035 ( .A1(n9753), .A2(n9752), .ZN(n9754) );
  INV_X4 U10036 ( .A(n9756), .ZN(n9757) );
  INV_X4 U10037 ( .A(n9761), .ZN(n9762) );
  XNOR2_X2 U10038 ( .A(n9877), .B(n9764), .ZN(n9879) );
  OAI221_X2 U10039 ( .B1(n9877), .B2(n9769), .C1(n9768), .C2(n10155), .A(n9767), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N85) );
  NAND2_X2 U10040 ( .A1(n9771), .A2(n9770), .ZN(n9787) );
  NAND2_X2 U10041 ( .A1(n6844), .A2(n9787), .ZN(n9796) );
  NAND2_X2 U10042 ( .A1(n9796), .A2(n7378), .ZN(n9834) );
  INV_X4 U10043 ( .A(n9834), .ZN(n10097) );
  INV_X4 U10044 ( .A(n9842), .ZN(n9773) );
  NAND2_X2 U10045 ( .A1(n9943), .A2(n9940), .ZN(n9782) );
  INV_X4 U10046 ( .A(n9781), .ZN(n9951) );
  XNOR2_X2 U10047 ( .A(n10134), .B(n10135), .ZN(n10162) );
  XNOR2_X2 U10048 ( .A(n10164), .B(n10163), .ZN(n10003) );
  XNOR2_X2 U10049 ( .A(n10228), .B(n10234), .ZN(n10232) );
  XNOR2_X2 U10050 ( .A(n10263), .B(n9998), .ZN(n9995) );
  NAND2_X2 U10051 ( .A1(n10127), .A2(n9995), .ZN(n9784) );
  XNOR2_X2 U10052 ( .A(n9787), .B(n9786), .ZN(n9861) );
  INV_X4 U10053 ( .A(n9826), .ZN(n9798) );
  INV_X4 U10054 ( .A(n9796), .ZN(n9797) );
  INV_X4 U10055 ( .A(n9800), .ZN(n9822) );
  NAND2_X2 U10056 ( .A1(n9822), .A2(n7307), .ZN(n9821) );
  INV_X4 U10057 ( .A(n9977), .ZN(n9805) );
  INV_X4 U10058 ( .A(n9925), .ZN(n9803) );
  OAI221_X2 U10059 ( .B1(n9805), .B2(n9804), .C1(n9803), .C2(n7391), .A(n9801), 
        .ZN(n9814) );
  INV_X4 U10060 ( .A(n9806), .ZN(n9813) );
  NAND2_X2 U10061 ( .A1(n9808), .A2(n7383), .ZN(n9809) );
  INV_X4 U10062 ( .A(n9809), .ZN(n9812) );
  NAND2_X2 U10063 ( .A1(n9821), .A2(n9820), .ZN(n9832) );
  NAND2_X2 U10064 ( .A1(n9822), .A2(n7450), .ZN(n9830) );
  INV_X4 U10065 ( .A(n9823), .ZN(n9824) );
  NAND2_X2 U10066 ( .A1(n9824), .A2(n7366), .ZN(n9829) );
  INV_X4 U10067 ( .A(n9861), .ZN(n9825) );
  NAND2_X2 U10068 ( .A1(n9825), .A2(ID_EXEC_OUT[158]), .ZN(n9828) );
  NAND2_X2 U10069 ( .A1(n10084), .A2(n9826), .ZN(n9827) );
  NAND4_X2 U10070 ( .A1(n9830), .A2(n9829), .A3(n9828), .A4(n9827), .ZN(n9831)
         );
  MUX2_X2 U10071 ( .A(n9832), .B(n9831), .S(ID_EXEC_OUT[157]), .Z(n9833) );
  INV_X4 U10072 ( .A(n9833), .ZN(n10095) );
  NAND2_X2 U10073 ( .A1(ID_EXEC_OUT[156]), .A2(n9834), .ZN(n10094) );
  NAND2_X2 U10074 ( .A1(ID_EXEC_OUT[157]), .A2(n9836), .ZN(n9841) );
  NAND2_X2 U10075 ( .A1(n9844), .A2(n9843), .ZN(n9875) );
  INV_X4 U10076 ( .A(n9875), .ZN(n9845) );
  INV_X4 U10077 ( .A(n9913), .ZN(n9904) );
  NAND2_X2 U10078 ( .A1(n9851), .A2(n9850), .ZN(n9854) );
  NAND3_X2 U10079 ( .A1(n9859), .A2(n9858), .A3(n9857), .ZN(n9860) );
  INV_X4 U10080 ( .A(n9869), .ZN(n9865) );
  AOI211_X4 U10081 ( .C1(n9870), .C2(n9869), .A(n9868), .B(n9867), .ZN(n9874)
         );
  NOR2_X4 U10082 ( .A1(n9874), .A2(n9873), .ZN(n9882) );
  NAND3_X2 U10083 ( .A1(n9884), .A2(n9892), .A3(n9883), .ZN(n9885) );
  INV_X4 U10084 ( .A(n9885), .ZN(n9963) );
  INV_X4 U10085 ( .A(n9896), .ZN(n9891) );
  INV_X4 U10086 ( .A(n9888), .ZN(n9890) );
  NAND2_X2 U10087 ( .A1(n9890), .A2(n9889), .ZN(n9897) );
  INV_X4 U10088 ( .A(n9897), .ZN(n9899) );
  NOR3_X4 U10089 ( .A1(n9892), .A2(n9891), .A3(n9899), .ZN(n9936) );
  NAND2_X2 U10090 ( .A1(n9895), .A2(n9894), .ZN(n9898) );
  NAND3_X2 U10091 ( .A1(n9898), .A2(n9897), .A3(n9896), .ZN(n9906) );
  NOR2_X4 U10092 ( .A1(n9900), .A2(n9899), .ZN(n9903) );
  INV_X4 U10093 ( .A(n9901), .ZN(n9902) );
  NAND2_X2 U10094 ( .A1(n9910), .A2(n9909), .ZN(n9923) );
  INV_X4 U10095 ( .A(n9911), .ZN(n9914) );
  NAND3_X2 U10096 ( .A1(n9914), .A2(n9913), .A3(n9912), .ZN(n9922) );
  INV_X4 U10097 ( .A(n9915), .ZN(n9917) );
  INV_X4 U10098 ( .A(n9938), .ZN(n9920) );
  NAND3_X2 U10099 ( .A1(n9923), .A2(n9922), .A3(n9921), .ZN(n9933) );
  NAND2_X2 U10100 ( .A1(n9586), .A2(n9925), .ZN(n9954) );
  INV_X4 U10101 ( .A(n9954), .ZN(n9932) );
  NAND2_X2 U10102 ( .A1(n9509), .A2(n9930), .ZN(n9945) );
  NAND2_X2 U10103 ( .A1(n9946), .A2(n9945), .ZN(n9931) );
  OAI21_X4 U10104 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(n9962) );
  NAND2_X2 U10105 ( .A1(n9938), .A2(n9937), .ZN(n9939) );
  INV_X4 U10106 ( .A(n9943), .ZN(n9944) );
  NAND2_X2 U10107 ( .A1(n9945), .A2(n9944), .ZN(n9948) );
  INV_X4 U10108 ( .A(n9946), .ZN(n9947) );
  NAND2_X2 U10109 ( .A1(n10003), .A2(n10232), .ZN(n9950) );
  INV_X4 U10110 ( .A(n9950), .ZN(n9956) );
  NOR2_X4 U10111 ( .A1(n10191), .A2(n9951), .ZN(n9953) );
  OAI21_X4 U10112 ( .B1(n9959), .B2(n9960), .A(n9958), .ZN(n9961) );
  OAI21_X4 U10113 ( .B1(n9963), .B2(n9962), .A(n9961), .ZN(n10026) );
  NAND2_X2 U10114 ( .A1(n9965), .A2(n9964), .ZN(n10068) );
  NAND2_X2 U10115 ( .A1(n10068), .A2(n10066), .ZN(n10041) );
  NAND2_X2 U10116 ( .A1(n9969), .A2(n9968), .ZN(n10036) );
  NAND2_X2 U10117 ( .A1(n10036), .A2(n10032), .ZN(n9972) );
  NAND2_X2 U10118 ( .A1(n9740), .A2(n9977), .ZN(n10030) );
  INV_X4 U10119 ( .A(n9978), .ZN(n9980) );
  NAND2_X2 U10120 ( .A1(n10066), .A2(n9982), .ZN(n9983) );
  INV_X4 U10121 ( .A(n9983), .ZN(n10054) );
  OAI21_X4 U10122 ( .B1(n10054), .B2(n9985), .A(n10067), .ZN(n10017) );
  INV_X4 U10123 ( .A(n10029), .ZN(n10062) );
  INV_X4 U10124 ( .A(n9989), .ZN(n10217) );
  NAND2_X2 U10125 ( .A1(n9990), .A2(n10163), .ZN(n10005) );
  INV_X4 U10126 ( .A(n10104), .ZN(n9994) );
  INV_X4 U10127 ( .A(n9996), .ZN(n9997) );
  INV_X4 U10128 ( .A(n10003), .ZN(n10170) );
  INV_X4 U10129 ( .A(n10017), .ZN(n10073) );
  INV_X4 U10130 ( .A(n10043), .ZN(n10016) );
  INV_X4 U10131 ( .A(n10013), .ZN(n10014) );
  AOI21_X4 U10132 ( .B1(n10030), .B2(n10015), .A(n10014), .ZN(n10047) );
  XNOR2_X2 U10133 ( .A(n10025), .B(n10051), .ZN(n10081) );
  NAND2_X2 U10134 ( .A1(n7307), .A2(n6828), .ZN(n10080) );
  NAND2_X2 U10135 ( .A1(n10038), .A2(n10051), .ZN(n10039) );
  INV_X4 U10136 ( .A(n10068), .ZN(n10061) );
  NOR2_X4 U10137 ( .A1(n10044), .A2(n10043), .ZN(n10045) );
  AOI211_X4 U10138 ( .C1(n10047), .C2(n10046), .A(n10045), .B(n10062), .ZN(
        n10049) );
  NOR2_X4 U10139 ( .A1(n10049), .A2(n9384), .ZN(n10069) );
  INV_X4 U10140 ( .A(n10052), .ZN(n10053) );
  INV_X4 U10141 ( .A(n10063), .ZN(n10064) );
  AOI211_X4 U10142 ( .C1(n10074), .C2(n10075), .A(n7346), .B(n10072), .ZN(
        n10076) );
  XNOR2_X2 U10143 ( .A(n10077), .B(n10076), .ZN(n10078) );
  XNOR2_X2 U10144 ( .A(n10078), .B(n10081), .ZN(n10088) );
  INV_X4 U10145 ( .A(n10088), .ZN(n10079) );
  INV_X4 U10146 ( .A(n10084), .ZN(n10087) );
  MUX2_X2 U10147 ( .A(n10087), .B(n10086), .S(n10085), .Z(n10090) );
  INV_X4 U10148 ( .A(n10223), .ZN(n10268) );
  XNOR2_X2 U10149 ( .A(n10103), .B(n10102), .ZN(n10126) );
  NAND2_X2 U10150 ( .A1(n10264), .A2(n10104), .ZN(n10106) );
  NAND2_X2 U10151 ( .A1(n5864), .A2(n10197), .ZN(n10111) );
  NAND2_X2 U10152 ( .A1(n10195), .A2(n10196), .ZN(n10110) );
  NAND2_X2 U10153 ( .A1(n8627), .A2(n10107), .ZN(n10109) );
  NAND2_X2 U10154 ( .A1(n7478), .A2(n10198), .ZN(n10108) );
  NAND4_X2 U10155 ( .A1(n10111), .A2(n10110), .A3(n10109), .A4(n10108), .ZN(
        n10275) );
  NAND2_X2 U10156 ( .A1(n5864), .A2(n10206), .ZN(n10116) );
  NAND2_X2 U10157 ( .A1(n9813), .A2(n10204), .ZN(n10115) );
  NAND2_X2 U10158 ( .A1(n10195), .A2(n10112), .ZN(n10114) );
  NAND2_X2 U10159 ( .A1(n10146), .A2(n10205), .ZN(n10113) );
  NAND4_X2 U10160 ( .A1(n10116), .A2(n10115), .A3(n10114), .A4(n10113), .ZN(
        n10276) );
  INV_X4 U10161 ( .A(n10276), .ZN(n10117) );
  OAI221_X2 U10162 ( .B1(n10127), .B2(n6861), .C1(n10126), .C2(n7479), .A(
        n10125), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N99) );
  XNOR2_X2 U10163 ( .A(n10133), .B(n10132), .ZN(n10161) );
  INV_X4 U10164 ( .A(n10135), .ZN(n10136) );
  NAND2_X2 U10165 ( .A1(n8976), .A2(n10203), .ZN(n10142) );
  NAND2_X2 U10166 ( .A1(n10146), .A2(n10204), .ZN(n10141) );
  NAND2_X2 U10167 ( .A1(n10248), .A2(n10206), .ZN(n10140) );
  NAND2_X2 U10168 ( .A1(n8975), .A2(n10138), .ZN(n10139) );
  NAND2_X2 U10169 ( .A1(n10146), .A2(n10194), .ZN(n10152) );
  INV_X4 U10170 ( .A(n7385), .ZN(n10147) );
  NAND2_X2 U10171 ( .A1(n10147), .A2(n10196), .ZN(n10151) );
  NAND2_X2 U10172 ( .A1(n10248), .A2(n10148), .ZN(n10150) );
  NAND2_X2 U10173 ( .A1(n8627), .A2(n10198), .ZN(n10149) );
  OAI221_X2 U10174 ( .B1(n10162), .B2(n6861), .C1(n10161), .C2(n7479), .A(
        n10160), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N104) );
  INV_X4 U10175 ( .A(n10163), .ZN(n10186) );
  NAND2_X2 U10176 ( .A1(n10272), .A2(n10170), .ZN(n10171) );
  NAND2_X2 U10177 ( .A1(n8976), .A2(n10245), .ZN(n10176) );
  NAND2_X2 U10178 ( .A1(n10146), .A2(n10247), .ZN(n10175) );
  NAND2_X2 U10179 ( .A1(n8975), .A2(n10249), .ZN(n10174) );
  NAND2_X2 U10180 ( .A1(n10248), .A2(n10172), .ZN(n10173) );
  AOI22_X2 U10181 ( .A1(n8976), .A2(n10237), .B1(n7478), .B2(n10236), .ZN(
        n10179) );
  AOI22_X2 U10182 ( .A1(n8975), .A2(n10177), .B1(n10195), .B2(n10239), .ZN(
        n10178) );
  NAND2_X2 U10183 ( .A1(n10179), .A2(n10178), .ZN(n10190) );
  NAND2_X2 U10184 ( .A1(n10277), .A2(n10190), .ZN(n10180) );
  OAI221_X2 U10185 ( .B1(n7139), .B2(n10281), .C1(n6804), .C2(n10279), .A(
        n10180), .ZN(n10181) );
  OAI221_X2 U10186 ( .B1(n10186), .B2(n10185), .C1(n10184), .C2(n7479), .A(
        n10183), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N103) );
  XNOR2_X2 U10187 ( .A(n10189), .B(n10188), .ZN(n10215) );
  INV_X4 U10188 ( .A(n10190), .ZN(n10193) );
  NAND2_X2 U10189 ( .A1(n10272), .A2(n10191), .ZN(n10192) );
  INV_X4 U10190 ( .A(n10246), .ZN(n10195) );
  NAND2_X2 U10191 ( .A1(n10195), .A2(n10194), .ZN(n10202) );
  NAND2_X2 U10192 ( .A1(n5884), .A2(n10196), .ZN(n10201) );
  NAND2_X2 U10193 ( .A1(n8975), .A2(n10197), .ZN(n10200) );
  NAND2_X2 U10194 ( .A1(n8976), .A2(n10198), .ZN(n10199) );
  NAND2_X2 U10195 ( .A1(n8975), .A2(n10203), .ZN(n10210) );
  NAND2_X2 U10196 ( .A1(n10147), .A2(n10204), .ZN(n10209) );
  NAND2_X2 U10197 ( .A1(n10248), .A2(n10205), .ZN(n10208) );
  NAND2_X2 U10198 ( .A1(n7478), .A2(n10206), .ZN(n10207) );
  NAND4_X2 U10199 ( .A1(n10210), .A2(n10209), .A3(n10208), .A4(n10207), .ZN(
        n10244) );
  NAND2_X2 U10200 ( .A1(n10277), .A2(n10244), .ZN(n10211) );
  OAI221_X2 U10201 ( .B1(n6804), .B2(n10281), .C1(n7233), .C2(n10279), .A(
        n10211), .ZN(n10212) );
  OAI221_X2 U10202 ( .B1(n10217), .B2(n10216), .C1(n10215), .C2(n7479), .A(
        n10214), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N102) );
  INV_X4 U10203 ( .A(n10218), .ZN(n10220) );
  INV_X4 U10204 ( .A(n10266), .ZN(n10222) );
  XNOR2_X2 U10205 ( .A(n10227), .B(n10226), .ZN(n10262) );
  INV_X4 U10206 ( .A(n10228), .ZN(n10231) );
  NAND2_X2 U10207 ( .A1(n10147), .A2(n10236), .ZN(n10243) );
  NAND2_X2 U10208 ( .A1(n9813), .A2(n10237), .ZN(n10242) );
  NAND2_X2 U10209 ( .A1(n10248), .A2(n10238), .ZN(n10241) );
  NAND2_X2 U10210 ( .A1(n7478), .A2(n10239), .ZN(n10240) );
  OAI22_X2 U10211 ( .A1(n7233), .A2(n7392), .B1(n6188), .B2(n6860), .ZN(n10259) );
  INV_X4 U10212 ( .A(n10244), .ZN(n10256) );
  NAND2_X2 U10213 ( .A1(n10146), .A2(n10245), .ZN(n10254) );
  INV_X4 U10214 ( .A(n10246), .ZN(n10248) );
  NAND2_X2 U10215 ( .A1(n10248), .A2(n10247), .ZN(n10253) );
  NAND2_X2 U10216 ( .A1(n8976), .A2(n10249), .ZN(n10252) );
  NAND2_X2 U10217 ( .A1(n8975), .A2(n10250), .ZN(n10251) );
  OAI22_X2 U10218 ( .A1(n10256), .A2(n10255), .B1(n7232), .B2(n7393), .ZN(
        n10258) );
  OAI211_X2 U10219 ( .C1(n10286), .C2(n10262), .A(n10261), .B(n10260), .ZN(
        EX_MEM_REGISTER_EX_MEM_REG_N101) );
  XNOR2_X2 U10220 ( .A(n10270), .B(n10269), .ZN(n10287) );
  NAND2_X2 U10221 ( .A1(n10272), .A2(n10271), .ZN(n10273) );
  INV_X4 U10222 ( .A(n10275), .ZN(n10280) );
  NAND2_X2 U10223 ( .A1(n10277), .A2(n10276), .ZN(n10278) );
  OAI221_X2 U10224 ( .B1(n7232), .B2(n10281), .C1(n10280), .C2(n10279), .A(
        n10278), .ZN(n10283) );
  OAI221_X2 U10225 ( .B1(n10289), .B2(n10288), .C1(n10287), .C2(n7479), .A(
        n10285), .ZN(EX_MEM_REGISTER_EX_MEM_REG_N100) );
  NAND2_X2 U10226 ( .A1(n6010), .A2(n10290), .ZN(n10292) );
  NAND2_X2 U10227 ( .A1(ID_EX_REG_ID_EX_REG_N95), .A2(n4447), .ZN(n10291) );
  NAND2_X2 U10228 ( .A1(n10292), .A2(n10291), .ZN(n1586) );
  OAI22_X2 U10229 ( .A1(n7722), .A2(n7481), .B1(n6276), .B2(n7720), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_100_ ( .D(DMEM_BUS_IN[31]), .CK(clk), 
        .RN(n7783), .Q(MEM_WB_OUT[100]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_99_ ( .D(DMEM_BUS_IN[30]), .CK(clk), 
        .RN(n7782), .Q(MEM_WB_OUT[99]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_98_ ( .D(DMEM_BUS_IN[29]), .CK(clk), 
        .RN(n7789), .Q(MEM_WB_OUT[98]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_97_ ( .D(DMEM_BUS_IN[28]), .CK(clk), 
        .RN(n7789), .Q(MEM_WB_OUT[97]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_96_ ( .D(DMEM_BUS_IN[27]), .CK(clk), 
        .RN(n7789), .Q(MEM_WB_OUT[96]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_95_ ( .D(DMEM_BUS_IN[26]), .CK(clk), 
        .RN(n7789), .Q(MEM_WB_OUT[95]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_94_ ( .D(DMEM_BUS_IN[25]), .CK(clk), 
        .RN(n7789), .Q(MEM_WB_OUT[94]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_93_ ( .D(DMEM_BUS_IN[24]), .CK(clk), 
        .RN(n7789), .Q(MEM_WB_OUT[93]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_92_ ( .D(DMEM_BUS_IN[23]), .CK(clk), 
        .RN(n7789), .Q(MEM_WB_OUT[92]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_91_ ( .D(DMEM_BUS_IN[22]), .CK(clk), 
        .RN(n7789), .Q(MEM_WB_OUT[91]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_90_ ( .D(DMEM_BUS_IN[21]), .CK(clk), 
        .RN(n7789), .Q(MEM_WB_OUT[90]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_89_ ( .D(DMEM_BUS_IN[20]), .CK(clk), 
        .RN(n7789), .Q(MEM_WB_OUT[89]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_88_ ( .D(DMEM_BUS_IN[19]), .CK(clk), 
        .RN(n7789), .Q(MEM_WB_OUT[88]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_87_ ( .D(DMEM_BUS_IN[18]), .CK(clk), 
        .RN(n7789), .Q(MEM_WB_OUT[87]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_86_ ( .D(DMEM_BUS_IN[17]), .CK(clk), 
        .RN(n7789), .Q(MEM_WB_OUT[86]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_85_ ( .D(DMEM_BUS_IN[16]), .CK(clk), 
        .RN(n7789), .Q(MEM_WB_OUT[85]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_84_ ( .D(DMEM_BUS_IN[15]), .CK(clk), 
        .RN(n7789), .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[31]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_83_ ( .D(DMEM_BUS_IN[14]), .CK(clk), 
        .RN(n7789), .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[30]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_82_ ( .D(DMEM_BUS_IN[13]), .CK(clk), 
        .RN(n7789), .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[29]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_81_ ( .D(DMEM_BUS_IN[12]), .CK(clk), 
        .RN(n7788), .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[28]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_80_ ( .D(DMEM_BUS_IN[11]), .CK(clk), 
        .RN(n7788), .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[27]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_79_ ( .D(DMEM_BUS_IN[10]), .CK(clk), 
        .RN(n7788), .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[26]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_78_ ( .D(DMEM_BUS_IN[9]), .CK(clk), 
        .RN(n7788), .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[25]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_76_ ( .D(DMEM_BUS_IN[7]), .CK(clk), 
        .RN(n7788), .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[23]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_75_ ( .D(DMEM_BUS_IN[6]), .CK(clk), 
        .RN(n7788), .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[22]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_74_ ( .D(DMEM_BUS_IN[5]), .CK(clk), 
        .RN(n7788), .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[21]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_73_ ( .D(DMEM_BUS_IN[4]), .CK(clk), 
        .RN(n7788), .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[20]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_71_ ( .D(DMEM_BUS_IN[2]), .CK(clk), 
        .RN(n7788), .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[18]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_31_ ( .D(IF_ID_REG_IF_ID_REG_N35), .CK(
        clk), .RN(n7776), .Q(IF_ID_OUT[31]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_30_ ( .D(IF_ID_REG_IF_ID_REG_N36), .CK(
        clk), .RN(n7775), .Q(IF_ID_OUT[30]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_20_ ( .D(n1552), .CK(clk), .RN(n7786), 
        .Q(IF_ID_OUT[20]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_19_ ( .D(n1553), .CK(clk), .RN(n7786), 
        .Q(IF_ID_OUT[19]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_18_ ( .D(n1554), .CK(clk), .RN(n7785), 
        .Q(IF_ID_OUT[18]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_17_ ( .D(n1555), .CK(clk), .RN(n7785), 
        .Q(IF_ID_OUT[17]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_16_ ( .D(n1556), .CK(clk), .RN(n7785), 
        .Q(IF_ID_OUT[16]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_15_ ( .D(n1557), .CK(clk), .RN(n7785), 
        .Q(IF_ID_OUT[15]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_14_ ( .D(n1558), .CK(clk), .RN(n7785), 
        .Q(IF_ID_OUT[14]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_13_ ( .D(n1559), .CK(clk), .RN(n7785), 
        .Q(IF_ID_OUT[13]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_12_ ( .D(n1560), .CK(clk), .RN(n7784), 
        .Q(IF_ID_OUT[12]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_11_ ( .D(n1561), .CK(clk), .RN(n7784), 
        .Q(IF_ID_OUT[11]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_10_ ( .D(n1562), .CK(clk), .RN(n7784), 
        .Q(IF_ID_OUT[10]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_9_ ( .D(n1563), .CK(clk), .RN(n7784), 
        .Q(IF_ID_OUT[9]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_8_ ( .D(n1564), .CK(clk), .RN(n7784), 
        .Q(IF_ID_OUT[8]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_7_ ( .D(n1565), .CK(clk), .RN(n7789), 
        .Q(IF_ID_OUT[7]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_6_ ( .D(n1566), .CK(clk), .RN(n7787), 
        .Q(IF_ID_OUT[6]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_5_ ( .D(n1567), .CK(clk), .RN(n7781), 
        .Q(IF_ID_OUT[5]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_4_ ( .D(n1568), .CK(clk), .RN(n7777), 
        .Q(IF_ID_OUT[4]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_3_ ( .D(n1569), .CK(clk), .RN(n7776), 
        .Q(IF_ID_OUT[3]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_2_ ( .D(n1570), .CK(clk), .RN(n7780), 
        .Q(IF_ID_OUT[2]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_1_ ( .D(n1571), .CK(clk), .RN(n7783), 
        .Q(IF_ID_OUT[1]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_0_ ( .D(n1572), .CK(clk), .RN(n7783), 
        .Q(IF_ID_OUT[0]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_29_ ( .D(n1543), .CK(clk), .RN(n7775), 
        .Q(IF_ID_OUT[29]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_45_ ( .D(IF_ID_REG_IF_ID_REG_N21), .CK(
        clk), .RN(n7792), .Q(offset_26_id[7]), .QN(n1641) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_58_ ( .D(IF_ID_REG_IF_ID_REG_N8), .CK(
        clk), .RN(n7790), .Q(ID_STAGE_imm16_aluA[26]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_57_ ( .D(IF_ID_REG_IF_ID_REG_N9), .CK(
        clk), .RN(n7781), .Q(ID_STAGE_imm16_aluA[25]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_55_ ( .D(IF_ID_REG_IF_ID_REG_N11), .CK(
        clk), .RN(n7793), .Q(ID_STAGE_imm16_aluA[23]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_54_ ( .D(IF_ID_REG_IF_ID_REG_N12), .CK(
        clk), .RN(n7786), .Q(ID_STAGE_imm16_aluA[22]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_50_ ( .D(IF_ID_REG_IF_ID_REG_N16), .CK(
        clk), .RN(n7781), .Q(ID_STAGE_imm16_aluA[18]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_28_ ( .D(n1544), .CK(clk), .RN(n7775), 
        .Q(IF_ID_OUT[28]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_27_ ( .D(n1545), .CK(clk), .RN(n7779), 
        .Q(IF_ID_OUT[27]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_26_ ( .D(n1546), .CK(clk), .RN(n7793), 
        .Q(IF_ID_OUT[26]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_25_ ( .D(n1547), .CK(clk), .RN(n7787), 
        .Q(IF_ID_OUT[25]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_24_ ( .D(n1548), .CK(clk), .RN(n7787), 
        .Q(IF_ID_OUT[24]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_23_ ( .D(n1549), .CK(clk), .RN(n7787), 
        .Q(IF_ID_OUT[23]) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[26]), .QN(n2012) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[22]), .QN(n2008) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[10]), .QN(n1996) );
  NAND2_X1 U5669 ( .A1(n7370), .A2(n9964), .ZN(n8274) );
  AOI22_X1 U5670 ( .A1(n7368), .A2(n9230), .B1(n3488), .B2(n3390), .ZN(n3487)
         );
  OAI21_X4 U5673 ( .B1(n8075), .B2(n7922), .A(n7921), .ZN(n9280) );
  OAI21_X4 U5674 ( .B1(n8075), .B2(n7903), .A(n7902), .ZN(n9275) );
  OAI21_X4 U7279 ( .B1(n8075), .B2(n8066), .A(n8065), .ZN(n9249) );
  OAI21_X4 U7280 ( .B1(n8075), .B2(n7968), .A(n7967), .ZN(n9246) );
endmodule

