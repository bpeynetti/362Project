
module and_1_0 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_31 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_30 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_29 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_28 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_27 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_26 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_25 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_24 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_23 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_22 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_21 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_20 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_19 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_18 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_17 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_16 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_15 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_14 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_13 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_12 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_11 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_10 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_9 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_8 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_7 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_6 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_5 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_4 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_3 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_2 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_1_1 ( x, y, z );
  input x, y;
  output z;


  AND2_X2 U1 ( .A1(y), .A2(x), .ZN(z) );
endmodule


module and_32 ( X, Y, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;


  and_1_0 \AND_32BIT[0].AND_1  ( .x(X[0]), .y(Y[0]), .z(Z[0]) );
  and_1_31 \AND_32BIT[1].AND_1  ( .x(X[1]), .y(Y[1]), .z(Z[1]) );
  and_1_30 \AND_32BIT[2].AND_1  ( .x(X[2]), .y(Y[2]), .z(Z[2]) );
  and_1_29 \AND_32BIT[3].AND_1  ( .x(X[3]), .y(Y[3]), .z(Z[3]) );
  and_1_28 \AND_32BIT[4].AND_1  ( .x(X[4]), .y(Y[4]), .z(Z[4]) );
  and_1_27 \AND_32BIT[5].AND_1  ( .x(X[5]), .y(Y[5]), .z(Z[5]) );
  and_1_26 \AND_32BIT[6].AND_1  ( .x(X[6]), .y(Y[6]), .z(Z[6]) );
  and_1_25 \AND_32BIT[7].AND_1  ( .x(X[7]), .y(Y[7]), .z(Z[7]) );
  and_1_24 \AND_32BIT[8].AND_1  ( .x(X[8]), .y(Y[8]), .z(Z[8]) );
  and_1_23 \AND_32BIT[9].AND_1  ( .x(X[9]), .y(Y[9]), .z(Z[9]) );
  and_1_22 \AND_32BIT[10].AND_1  ( .x(X[10]), .y(Y[10]), .z(Z[10]) );
  and_1_21 \AND_32BIT[11].AND_1  ( .x(X[11]), .y(Y[11]), .z(Z[11]) );
  and_1_20 \AND_32BIT[12].AND_1  ( .x(X[12]), .y(Y[12]), .z(Z[12]) );
  and_1_19 \AND_32BIT[13].AND_1  ( .x(X[13]), .y(Y[13]), .z(Z[13]) );
  and_1_18 \AND_32BIT[14].AND_1  ( .x(X[14]), .y(Y[14]), .z(Z[14]) );
  and_1_17 \AND_32BIT[15].AND_1  ( .x(X[15]), .y(Y[15]), .z(Z[15]) );
  and_1_16 \AND_32BIT[16].AND_1  ( .x(X[16]), .y(Y[16]), .z(Z[16]) );
  and_1_15 \AND_32BIT[17].AND_1  ( .x(X[17]), .y(Y[17]), .z(Z[17]) );
  and_1_14 \AND_32BIT[18].AND_1  ( .x(X[18]), .y(Y[18]), .z(Z[18]) );
  and_1_13 \AND_32BIT[19].AND_1  ( .x(X[19]), .y(Y[19]), .z(Z[19]) );
  and_1_12 \AND_32BIT[20].AND_1  ( .x(X[20]), .y(Y[20]), .z(Z[20]) );
  and_1_11 \AND_32BIT[21].AND_1  ( .x(X[21]), .y(Y[21]), .z(Z[21]) );
  and_1_10 \AND_32BIT[22].AND_1  ( .x(X[22]), .y(Y[22]), .z(Z[22]) );
  and_1_9 \AND_32BIT[23].AND_1  ( .x(X[23]), .y(Y[23]), .z(Z[23]) );
  and_1_8 \AND_32BIT[24].AND_1  ( .x(X[24]), .y(Y[24]), .z(Z[24]) );
  and_1_7 \AND_32BIT[25].AND_1  ( .x(X[25]), .y(Y[25]), .z(Z[25]) );
  and_1_6 \AND_32BIT[26].AND_1  ( .x(X[26]), .y(Y[26]), .z(Z[26]) );
  and_1_5 \AND_32BIT[27].AND_1  ( .x(X[27]), .y(Y[27]), .z(Z[27]) );
  and_1_4 \AND_32BIT[28].AND_1  ( .x(X[28]), .y(Y[28]), .z(Z[28]) );
  and_1_3 \AND_32BIT[29].AND_1  ( .x(X[29]), .y(Y[29]), .z(Z[29]) );
  and_1_2 \AND_32BIT[30].AND_1  ( .x(X[30]), .y(Y[30]), .z(Z[30]) );
  and_1_1 \AND_32BIT[31].AND_1  ( .x(X[31]), .y(Y[31]), .z(Z[31]) );
endmodule


module or_1_0 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_31 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_30 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_29 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_28 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_27 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_26 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_25 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_24 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_23 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_22 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_21 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_20 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_19 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_18 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_17 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_16 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_15 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_14 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_13 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_12 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_11 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_10 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_9 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_8 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_7 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_6 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_5 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_4 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_3 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_2 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_1_1 ( x, y, z );
  input x, y;
  output z;


  OR2_X2 U1 ( .A1(x), .A2(y), .ZN(z) );
endmodule


module or_32 ( X, Y, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;


  or_1_0 \OR_32BIT[0].OR_1  ( .x(X[0]), .y(Y[0]), .z(Z[0]) );
  or_1_31 \OR_32BIT[1].OR_1  ( .x(X[1]), .y(Y[1]), .z(Z[1]) );
  or_1_30 \OR_32BIT[2].OR_1  ( .x(X[2]), .y(Y[2]), .z(Z[2]) );
  or_1_29 \OR_32BIT[3].OR_1  ( .x(X[3]), .y(Y[3]), .z(Z[3]) );
  or_1_28 \OR_32BIT[4].OR_1  ( .x(X[4]), .y(Y[4]), .z(Z[4]) );
  or_1_27 \OR_32BIT[5].OR_1  ( .x(X[5]), .y(Y[5]), .z(Z[5]) );
  or_1_26 \OR_32BIT[6].OR_1  ( .x(X[6]), .y(Y[6]), .z(Z[6]) );
  or_1_25 \OR_32BIT[7].OR_1  ( .x(X[7]), .y(Y[7]), .z(Z[7]) );
  or_1_24 \OR_32BIT[8].OR_1  ( .x(X[8]), .y(Y[8]), .z(Z[8]) );
  or_1_23 \OR_32BIT[9].OR_1  ( .x(X[9]), .y(Y[9]), .z(Z[9]) );
  or_1_22 \OR_32BIT[10].OR_1  ( .x(X[10]), .y(Y[10]), .z(Z[10]) );
  or_1_21 \OR_32BIT[11].OR_1  ( .x(X[11]), .y(Y[11]), .z(Z[11]) );
  or_1_20 \OR_32BIT[12].OR_1  ( .x(X[12]), .y(Y[12]), .z(Z[12]) );
  or_1_19 \OR_32BIT[13].OR_1  ( .x(X[13]), .y(Y[13]), .z(Z[13]) );
  or_1_18 \OR_32BIT[14].OR_1  ( .x(X[14]), .y(Y[14]), .z(Z[14]) );
  or_1_17 \OR_32BIT[15].OR_1  ( .x(X[15]), .y(Y[15]), .z(Z[15]) );
  or_1_16 \OR_32BIT[16].OR_1  ( .x(X[16]), .y(Y[16]), .z(Z[16]) );
  or_1_15 \OR_32BIT[17].OR_1  ( .x(X[17]), .y(Y[17]), .z(Z[17]) );
  or_1_14 \OR_32BIT[18].OR_1  ( .x(X[18]), .y(Y[18]), .z(Z[18]) );
  or_1_13 \OR_32BIT[19].OR_1  ( .x(X[19]), .y(Y[19]), .z(Z[19]) );
  or_1_12 \OR_32BIT[20].OR_1  ( .x(X[20]), .y(Y[20]), .z(Z[20]) );
  or_1_11 \OR_32BIT[21].OR_1  ( .x(X[21]), .y(Y[21]), .z(Z[21]) );
  or_1_10 \OR_32BIT[22].OR_1  ( .x(X[22]), .y(Y[22]), .z(Z[22]) );
  or_1_9 \OR_32BIT[23].OR_1  ( .x(X[23]), .y(Y[23]), .z(Z[23]) );
  or_1_8 \OR_32BIT[24].OR_1  ( .x(X[24]), .y(Y[24]), .z(Z[24]) );
  or_1_7 \OR_32BIT[25].OR_1  ( .x(X[25]), .y(Y[25]), .z(Z[25]) );
  or_1_6 \OR_32BIT[26].OR_1  ( .x(X[26]), .y(Y[26]), .z(Z[26]) );
  or_1_5 \OR_32BIT[27].OR_1  ( .x(X[27]), .y(Y[27]), .z(Z[27]) );
  or_1_4 \OR_32BIT[28].OR_1  ( .x(X[28]), .y(Y[28]), .z(Z[28]) );
  or_1_3 \OR_32BIT[29].OR_1  ( .x(X[29]), .y(Y[29]), .z(Z[29]) );
  or_1_2 \OR_32BIT[30].OR_1  ( .x(X[30]), .y(Y[30]), .z(Z[30]) );
  or_1_1 \OR_32BIT[31].OR_1  ( .x(X[31]), .y(Y[31]), .z(Z[31]) );
endmodule


module xor_1_0 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_31 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_30 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_29 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_28 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_27 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_26 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_25 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_24 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_23 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_22 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_21 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_20 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_19 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_18 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_17 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_16 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_15 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_14 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_13 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_12 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_11 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_10 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_9 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_8 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_7 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_6 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_5 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_4 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_3 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_2 ( x, y, z );
  input x, y;
  output z;


  XOR2_X1 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_1_1 ( x, y, z );
  input x, y;
  output z;


  XOR2_X2 U1 ( .A(y), .B(x), .Z(z) );
endmodule


module xor_32 ( X, Y, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;


  xor_1_0 \XOR_32BIT[0].XOR_1  ( .x(X[0]), .y(Y[0]), .z(Z[0]) );
  xor_1_31 \XOR_32BIT[1].XOR_1  ( .x(X[1]), .y(Y[1]), .z(Z[1]) );
  xor_1_30 \XOR_32BIT[2].XOR_1  ( .x(X[2]), .y(Y[2]), .z(Z[2]) );
  xor_1_29 \XOR_32BIT[3].XOR_1  ( .x(X[3]), .y(Y[3]), .z(Z[3]) );
  xor_1_28 \XOR_32BIT[4].XOR_1  ( .x(X[4]), .y(Y[4]), .z(Z[4]) );
  xor_1_27 \XOR_32BIT[5].XOR_1  ( .x(X[5]), .y(Y[5]), .z(Z[5]) );
  xor_1_26 \XOR_32BIT[6].XOR_1  ( .x(X[6]), .y(Y[6]), .z(Z[6]) );
  xor_1_25 \XOR_32BIT[7].XOR_1  ( .x(X[7]), .y(Y[7]), .z(Z[7]) );
  xor_1_24 \XOR_32BIT[8].XOR_1  ( .x(X[8]), .y(Y[8]), .z(Z[8]) );
  xor_1_23 \XOR_32BIT[9].XOR_1  ( .x(X[9]), .y(Y[9]), .z(Z[9]) );
  xor_1_22 \XOR_32BIT[10].XOR_1  ( .x(X[10]), .y(Y[10]), .z(Z[10]) );
  xor_1_21 \XOR_32BIT[11].XOR_1  ( .x(X[11]), .y(Y[11]), .z(Z[11]) );
  xor_1_20 \XOR_32BIT[12].XOR_1  ( .x(X[12]), .y(Y[12]), .z(Z[12]) );
  xor_1_19 \XOR_32BIT[13].XOR_1  ( .x(X[13]), .y(Y[13]), .z(Z[13]) );
  xor_1_18 \XOR_32BIT[14].XOR_1  ( .x(X[14]), .y(Y[14]), .z(Z[14]) );
  xor_1_17 \XOR_32BIT[15].XOR_1  ( .x(X[15]), .y(Y[15]), .z(Z[15]) );
  xor_1_16 \XOR_32BIT[16].XOR_1  ( .x(X[16]), .y(Y[16]), .z(Z[16]) );
  xor_1_15 \XOR_32BIT[17].XOR_1  ( .x(X[17]), .y(Y[17]), .z(Z[17]) );
  xor_1_14 \XOR_32BIT[18].XOR_1  ( .x(X[18]), .y(Y[18]), .z(Z[18]) );
  xor_1_13 \XOR_32BIT[19].XOR_1  ( .x(X[19]), .y(Y[19]), .z(Z[19]) );
  xor_1_12 \XOR_32BIT[20].XOR_1  ( .x(X[20]), .y(Y[20]), .z(Z[20]) );
  xor_1_11 \XOR_32BIT[21].XOR_1  ( .x(X[21]), .y(Y[21]), .z(Z[21]) );
  xor_1_10 \XOR_32BIT[22].XOR_1  ( .x(X[22]), .y(Y[22]), .z(Z[22]) );
  xor_1_9 \XOR_32BIT[23].XOR_1  ( .x(X[23]), .y(Y[23]), .z(Z[23]) );
  xor_1_8 \XOR_32BIT[24].XOR_1  ( .x(X[24]), .y(Y[24]), .z(Z[24]) );
  xor_1_7 \XOR_32BIT[25].XOR_1  ( .x(X[25]), .y(Y[25]), .z(Z[25]) );
  xor_1_6 \XOR_32BIT[26].XOR_1  ( .x(X[26]), .y(Y[26]), .z(Z[26]) );
  xor_1_5 \XOR_32BIT[27].XOR_1  ( .x(X[27]), .y(Y[27]), .z(Z[27]) );
  xor_1_4 \XOR_32BIT[28].XOR_1  ( .x(X[28]), .y(Y[28]), .z(Z[28]) );
  xor_1_3 \XOR_32BIT[29].XOR_1  ( .x(X[29]), .y(Y[29]), .z(Z[29]) );
  xor_1_2 \XOR_32BIT[30].XOR_1  ( .x(X[30]), .y(Y[30]), .z(Z[30]) );
  xor_1_1 \XOR_32BIT[31].XOR_1  ( .x(X[31]), .y(Y[31]), .z(Z[31]) );
endmodule


module not_1_0 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_63 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_62 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_61 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_60 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_59 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_58 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_57 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_56 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_55 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_54 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_53 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_52 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_51 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_50 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_49 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_48 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_47 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_46 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_45 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_44 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_43 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_42 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_41 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_40 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_39 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_38 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_37 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_36 ( x, z );
  input x;
  output z;


  INV_X1 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_35 ( x, z );
  input x;
  output z;


  INV_X1 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_34 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_33 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_32_0 ( X, Z );
  input [0:31] X;
  output [0:31] Z;


  not_1_0 \NOT_32BIT[0].NOT_1  ( .x(X[0]), .z(Z[0]) );
  not_1_63 \NOT_32BIT[1].NOT_1  ( .x(X[1]), .z(Z[1]) );
  not_1_62 \NOT_32BIT[2].NOT_1  ( .x(X[2]), .z(Z[2]) );
  not_1_61 \NOT_32BIT[3].NOT_1  ( .x(X[3]), .z(Z[3]) );
  not_1_60 \NOT_32BIT[4].NOT_1  ( .x(X[4]), .z(Z[4]) );
  not_1_59 \NOT_32BIT[5].NOT_1  ( .x(X[5]), .z(Z[5]) );
  not_1_58 \NOT_32BIT[6].NOT_1  ( .x(X[6]), .z(Z[6]) );
  not_1_57 \NOT_32BIT[7].NOT_1  ( .x(X[7]), .z(Z[7]) );
  not_1_56 \NOT_32BIT[8].NOT_1  ( .x(X[8]), .z(Z[8]) );
  not_1_55 \NOT_32BIT[9].NOT_1  ( .x(X[9]), .z(Z[9]) );
  not_1_54 \NOT_32BIT[10].NOT_1  ( .x(X[10]), .z(Z[10]) );
  not_1_53 \NOT_32BIT[11].NOT_1  ( .x(X[11]), .z(Z[11]) );
  not_1_52 \NOT_32BIT[12].NOT_1  ( .x(X[12]), .z(Z[12]) );
  not_1_51 \NOT_32BIT[13].NOT_1  ( .x(X[13]), .z(Z[13]) );
  not_1_50 \NOT_32BIT[14].NOT_1  ( .x(X[14]), .z(Z[14]) );
  not_1_49 \NOT_32BIT[15].NOT_1  ( .x(X[15]), .z(Z[15]) );
  not_1_48 \NOT_32BIT[16].NOT_1  ( .x(X[16]), .z(Z[16]) );
  not_1_47 \NOT_32BIT[17].NOT_1  ( .x(X[17]), .z(Z[17]) );
  not_1_46 \NOT_32BIT[18].NOT_1  ( .x(X[18]), .z(Z[18]) );
  not_1_45 \NOT_32BIT[19].NOT_1  ( .x(X[19]), .z(Z[19]) );
  not_1_44 \NOT_32BIT[20].NOT_1  ( .x(X[20]), .z(Z[20]) );
  not_1_43 \NOT_32BIT[21].NOT_1  ( .x(X[21]), .z(Z[21]) );
  not_1_42 \NOT_32BIT[22].NOT_1  ( .x(X[22]), .z(Z[22]) );
  not_1_41 \NOT_32BIT[23].NOT_1  ( .x(X[23]), .z(Z[23]) );
  not_1_40 \NOT_32BIT[24].NOT_1  ( .x(X[24]), .z(Z[24]) );
  not_1_39 \NOT_32BIT[25].NOT_1  ( .x(X[25]), .z(Z[25]) );
  not_1_38 \NOT_32BIT[26].NOT_1  ( .x(X[26]), .z(Z[26]) );
  not_1_37 \NOT_32BIT[27].NOT_1  ( .x(X[27]), .z(Z[27]) );
  not_1_36 \NOT_32BIT[28].NOT_1  ( .x(X[28]), .z(Z[28]) );
  not_1_35 \NOT_32BIT[29].NOT_1  ( .x(X[29]), .z(Z[29]) );
  not_1_34 \NOT_32BIT[30].NOT_1  ( .x(X[30]), .z(Z[30]) );
  not_1_33 \NOT_32BIT[31].NOT_1  ( .x(X[31]), .z(Z[31]) );
endmodule


module mux_1_870 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_869 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_868 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_867 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_866 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_865 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_864 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_863 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_862 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_861 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_860 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_859 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_858 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X1 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_857 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_856 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_855 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_854 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_853 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_852 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_851 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_850 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_849 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_848 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_847 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_846 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_845 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_844 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_843 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_842 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_841 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_840 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  NAND2_X2 U1 ( .A1(x), .A2(n1), .ZN(n2) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  NAND2_X2 U3 ( .A1(y), .A2(sel), .ZN(n3) );
  NAND2_X4 U4 ( .A1(n2), .A2(n3), .ZN(z) );
endmodule


module mux_1_839 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2, n3;

  INV_X16 U1 ( .A(x), .ZN(n2) );
  NAND2_X4 U2 ( .A1(n2), .A2(sel), .ZN(n3) );
  OAI21_X4 U3 ( .B1(y), .B2(sel), .A(n3), .ZN(z) );
endmodule


module mux2to1_32bit_27 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(sel), .ZN(n4) );
  INV_X4 U2 ( .A(n4), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(n2) );
  INV_X4 U4 ( .A(n4), .ZN(n3) );
  mux_1_870 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n3), .z(Z[0]) );
  mux_1_869 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n2), .z(Z[1]) );
  mux_1_868 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_867 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n3), .z(Z[3]) );
  mux_1_866 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n2), .z(Z[4]) );
  mux_1_865 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_864 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n3), .z(Z[6]) );
  mux_1_863 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n2), .z(Z[7]) );
  mux_1_862 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_861 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n3), .z(Z[9]) );
  mux_1_860 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n2), .z(Z[10]) );
  mux_1_859 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_858 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n3), .z(Z[12]) );
  mux_1_857 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n3), .z(Z[13]) );
  mux_1_856 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_855 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n1), .z(Z[15]) );
  mux_1_854 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(sel), .z(
        Z[16]) );
  mux_1_853 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(sel), .z(
        Z[17]) );
  mux_1_852 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(sel), .z(
        Z[18]) );
  mux_1_851 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(sel), .z(
        Z[19]) );
  mux_1_850 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(sel), .z(
        Z[20]) );
  mux_1_849 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(sel), .z(
        Z[21]) );
  mux_1_848 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(sel), .z(
        Z[22]) );
  mux_1_847 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(sel), .z(
        Z[23]) );
  mux_1_846 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(sel), .z(
        Z[24]) );
  mux_1_845 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(sel), .z(
        Z[25]) );
  mux_1_844 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(sel), .z(
        Z[26]) );
  mux_1_843 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(sel), .z(
        Z[27]) );
  mux_1_842 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(sel), .z(
        Z[28]) );
  mux_1_841 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(sel), .z(
        Z[29]) );
  mux_1_840 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(sel), .z(
        Z[30]) );
  mux_1_839 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(sel), .z(
        Z[31]) );
endmodule


module fa_0 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1;

  XNOR2_X2 U1 ( .A(b), .B(a), .ZN(n1) );
  XNOR2_X2 U2 ( .A(cin), .B(n1), .ZN(sum) );
endmodule


module fa_63 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4;

  NAND2_X4 U1 ( .A1(n3), .A2(n2), .ZN(cout) );
  XNOR2_X2 U2 ( .A(b), .B(a), .ZN(n4) );
  INV_X4 U3 ( .A(n4), .ZN(n1) );
  NAND2_X2 U4 ( .A1(cin), .A2(n1), .ZN(n3) );
  NAND2_X2 U5 ( .A1(b), .A2(a), .ZN(n2) );
  XNOR2_X2 U6 ( .A(cin), .B(n4), .ZN(sum) );
endmodule


module fa_62 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4;

  NAND2_X4 U1 ( .A1(n3), .A2(n2), .ZN(cout) );
  NAND2_X4 U2 ( .A1(cin), .A2(n1), .ZN(n3) );
  XNOR2_X2 U3 ( .A(b), .B(a), .ZN(n4) );
  INV_X4 U4 ( .A(n4), .ZN(n1) );
  NAND2_X2 U5 ( .A1(b), .A2(a), .ZN(n2) );
  XNOR2_X2 U6 ( .A(cin), .B(n4), .ZN(sum) );
endmodule


module fa_61 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4;

  NAND2_X2 U1 ( .A1(cin), .A2(n1), .ZN(n3) );
  NAND2_X4 U2 ( .A1(n3), .A2(n2), .ZN(cout) );
  XNOR2_X2 U3 ( .A(b), .B(a), .ZN(n4) );
  INV_X4 U4 ( .A(n4), .ZN(n1) );
  NAND2_X2 U5 ( .A1(b), .A2(a), .ZN(n2) );
  XNOR2_X2 U6 ( .A(cin), .B(n4), .ZN(sum) );
endmodule


module fa_60 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(cin), .B(n4), .ZN(sum) );
  NAND2_X4 U2 ( .A1(cin), .A2(n1), .ZN(n3) );
  NAND2_X4 U3 ( .A1(n3), .A2(n2), .ZN(cout) );
  XNOR2_X2 U4 ( .A(b), .B(a), .ZN(n4) );
  INV_X4 U5 ( .A(n4), .ZN(n1) );
  NAND2_X2 U6 ( .A1(b), .A2(a), .ZN(n2) );
endmodule


module fa_59 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5, n6;

  AND2_X4 U1 ( .A1(b), .A2(a), .ZN(n1) );
  AOI21_X4 U5 ( .B1(cin), .B2(n5), .A(n1), .ZN(n4) );
  INV_X8 U6 ( .A(n4), .ZN(cout) );
  XNOR2_X2 U7 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U8 ( .A(n6), .ZN(n5) );
  XNOR2_X1 U2 ( .A(cin), .B(n6), .ZN(sum) );
endmodule


module fa_58 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  INV_X1 U1 ( .A(cin), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(n2) );
  XNOR2_X1 U3 ( .A(n2), .B(n6), .ZN(sum) );
  NAND2_X4 U4 ( .A1(n5), .A2(n4), .ZN(cout) );
  NAND2_X4 U5 ( .A1(cin), .A2(n3), .ZN(n5) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NAND2_X2 U8 ( .A1(b), .A2(a), .ZN(n4) );
endmodule


module fa_57 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6, n8;

  INV_X1 U1 ( .A(n8), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(n2) );
  NAND2_X4 U3 ( .A1(cin), .A2(n3), .ZN(n5) );
  XNOR2_X1 U4 ( .A(n2), .B(n6), .ZN(sum) );
  NAND2_X4 U5 ( .A1(n5), .A2(n4), .ZN(cout) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NAND2_X2 U8 ( .A1(b), .A2(a), .ZN(n4) );
  BUF_X8 U9 ( .A(cin), .Z(n8) );
endmodule


module fa_56 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6, n8;

  INV_X1 U1 ( .A(n8), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(n2) );
  NAND2_X4 U3 ( .A1(cin), .A2(n3), .ZN(n5) );
  XNOR2_X1 U4 ( .A(n2), .B(n6), .ZN(sum) );
  NAND2_X4 U5 ( .A1(n5), .A2(n4), .ZN(cout) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NAND2_X2 U8 ( .A1(b), .A2(a), .ZN(n4) );
  BUF_X16 U9 ( .A(cin), .Z(n8) );
endmodule


module fa_55 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  INV_X1 U1 ( .A(cin), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(n2) );
  NAND2_X4 U3 ( .A1(cin), .A2(n3), .ZN(n5) );
  XNOR2_X1 U4 ( .A(n2), .B(n6), .ZN(sum) );
  NAND2_X4 U5 ( .A1(n5), .A2(n4), .ZN(cout) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NAND2_X2 U8 ( .A1(b), .A2(a), .ZN(n4) );
endmodule


module fa_54 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6, n8;

  INV_X1 U1 ( .A(n8), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(n2) );
  XNOR2_X1 U3 ( .A(n2), .B(n6), .ZN(sum) );
  NAND2_X4 U4 ( .A1(cin), .A2(n3), .ZN(n5) );
  NAND2_X4 U5 ( .A1(n5), .A2(n4), .ZN(cout) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NAND2_X2 U8 ( .A1(b), .A2(a), .ZN(n4) );
  BUF_X32 U9 ( .A(cin), .Z(n8) );
endmodule


module fa_53 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(n5), .ZN(sum) );
  NAND2_X4 U3 ( .A1(n4), .A2(n3), .ZN(cout) );
  NAND2_X4 U4 ( .A1(cin), .A2(n2), .ZN(n4) );
  XNOR2_X2 U5 ( .A(b), .B(a), .ZN(n5) );
  INV_X4 U6 ( .A(n5), .ZN(n2) );
  NAND2_X2 U7 ( .A1(b), .A2(a), .ZN(n3) );
endmodule


module fa_52 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  NAND2_X4 U2 ( .A1(cin), .A2(n2), .ZN(n4) );
  XNOR2_X1 U3 ( .A(n1), .B(n5), .ZN(sum) );
  NAND2_X4 U4 ( .A1(n4), .A2(n3), .ZN(cout) );
  XNOR2_X2 U5 ( .A(b), .B(a), .ZN(n5) );
  INV_X4 U6 ( .A(n5), .ZN(n2) );
  NAND2_X2 U7 ( .A1(b), .A2(a), .ZN(n3) );
endmodule


module fa_51 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  NAND2_X4 U2 ( .A1(n4), .A2(n3), .ZN(cout) );
  NAND2_X4 U3 ( .A1(cin), .A2(n2), .ZN(n4) );
  XNOR2_X1 U4 ( .A(n1), .B(n5), .ZN(sum) );
  XNOR2_X2 U5 ( .A(b), .B(a), .ZN(n5) );
  INV_X4 U6 ( .A(n5), .ZN(n2) );
  NAND2_X2 U7 ( .A1(b), .A2(a), .ZN(n3) );
endmodule


module fa_50 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6, n8;

  INV_X1 U1 ( .A(n8), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(n2) );
  XNOR2_X1 U3 ( .A(n2), .B(n6), .ZN(sum) );
  NAND2_X4 U4 ( .A1(n5), .A2(n4), .ZN(cout) );
  NAND2_X4 U5 ( .A1(cin), .A2(n3), .ZN(n5) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NAND2_X2 U8 ( .A1(b), .A2(a), .ZN(n4) );
  BUF_X32 U9 ( .A(cin), .Z(n8) );
endmodule


module fa_49 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(n5), .ZN(sum) );
  NAND2_X4 U3 ( .A1(n4), .A2(n3), .ZN(cout) );
  NAND2_X4 U4 ( .A1(cin), .A2(n2), .ZN(n4) );
  XNOR2_X2 U5 ( .A(b), .B(a), .ZN(n5) );
  INV_X4 U6 ( .A(n5), .ZN(n2) );
  NAND2_X2 U7 ( .A1(b), .A2(a), .ZN(n3) );
endmodule


module fa_48 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6, n8;

  INV_X1 U1 ( .A(n8), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(n2) );
  XNOR2_X1 U3 ( .A(n2), .B(n6), .ZN(sum) );
  NAND2_X4 U4 ( .A1(n5), .A2(n4), .ZN(cout) );
  NAND2_X4 U5 ( .A1(cin), .A2(n3), .ZN(n5) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NAND2_X2 U8 ( .A1(b), .A2(a), .ZN(n4) );
  BUF_X32 U9 ( .A(cin), .Z(n8) );
endmodule


module fa_47 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6, n8;

  INV_X1 U1 ( .A(n8), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(n2) );
  XNOR2_X1 U3 ( .A(n2), .B(n6), .ZN(sum) );
  NAND2_X4 U4 ( .A1(n5), .A2(n4), .ZN(cout) );
  NAND2_X4 U5 ( .A1(cin), .A2(n3), .ZN(n5) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NAND2_X2 U8 ( .A1(b), .A2(a), .ZN(n4) );
  BUF_X32 U9 ( .A(cin), .Z(n8) );
endmodule


module fa_46 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6, n8;

  INV_X1 U1 ( .A(n8), .ZN(n1) );
  INV_X4 U2 ( .A(n1), .ZN(n2) );
  XNOR2_X1 U3 ( .A(n2), .B(n6), .ZN(sum) );
  NAND2_X4 U4 ( .A1(n5), .A2(n4), .ZN(cout) );
  NAND2_X4 U5 ( .A1(cin), .A2(n3), .ZN(n5) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NAND2_X2 U8 ( .A1(b), .A2(a), .ZN(n4) );
  BUF_X32 U9 ( .A(cin), .Z(n8) );
endmodule


module fa_45 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  NAND2_X4 U2 ( .A1(cin), .A2(n2), .ZN(n4) );
  XNOR2_X1 U3 ( .A(n1), .B(n5), .ZN(sum) );
  NAND2_X4 U4 ( .A1(n4), .A2(n3), .ZN(cout) );
  XNOR2_X2 U5 ( .A(b), .B(a), .ZN(n5) );
  INV_X4 U6 ( .A(n5), .ZN(n2) );
  NAND2_X2 U7 ( .A1(b), .A2(a), .ZN(n3) );
endmodule


module fa_44 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(n5), .ZN(sum) );
  NAND2_X4 U3 ( .A1(cin), .A2(n2), .ZN(n4) );
  NAND2_X4 U4 ( .A1(n4), .A2(n3), .ZN(cout) );
  XNOR2_X2 U5 ( .A(b), .B(a), .ZN(n5) );
  INV_X4 U6 ( .A(n5), .ZN(n2) );
  NAND2_X2 U7 ( .A1(b), .A2(a), .ZN(n3) );
endmodule


module fa_43 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6, n7;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n1), .ZN(n2) );
  INV_X4 U3 ( .A(n2), .ZN(n3) );
  XNOR2_X1 U4 ( .A(n3), .B(n7), .ZN(sum) );
  NAND2_X4 U5 ( .A1(n6), .A2(n5), .ZN(cout) );
  NAND2_X4 U6 ( .A1(cin), .A2(n4), .ZN(n6) );
  XNOR2_X2 U7 ( .A(b), .B(a), .ZN(n7) );
  INV_X4 U8 ( .A(n7), .ZN(n4) );
  NAND2_X2 U9 ( .A1(b), .A2(a), .ZN(n5) );
endmodule


module fa_42 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  NAND2_X4 U2 ( .A1(cin), .A2(n2), .ZN(n4) );
  XNOR2_X1 U3 ( .A(n1), .B(n5), .ZN(sum) );
  NAND2_X4 U4 ( .A1(n4), .A2(n3), .ZN(cout) );
  XNOR2_X2 U5 ( .A(b), .B(a), .ZN(n5) );
  INV_X4 U6 ( .A(n5), .ZN(n2) );
  NAND2_X2 U7 ( .A1(b), .A2(a), .ZN(n3) );
endmodule


module fa_41 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  NAND2_X4 U2 ( .A1(n4), .A2(n3), .ZN(cout) );
  XNOR2_X1 U3 ( .A(n1), .B(n5), .ZN(sum) );
  NAND2_X4 U4 ( .A1(cin), .A2(n2), .ZN(n4) );
  XNOR2_X2 U5 ( .A(b), .B(a), .ZN(n5) );
  INV_X4 U6 ( .A(n5), .ZN(n2) );
  NAND2_X2 U7 ( .A1(b), .A2(a), .ZN(n3) );
endmodule


module fa_40 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  NAND2_X4 U2 ( .A1(cin), .A2(n2), .ZN(n4) );
  XNOR2_X1 U3 ( .A(n1), .B(n5), .ZN(sum) );
  NAND2_X4 U4 ( .A1(n4), .A2(n3), .ZN(cout) );
  XNOR2_X2 U5 ( .A(b), .B(a), .ZN(n5) );
  INV_X4 U6 ( .A(n5), .ZN(n2) );
  NAND2_X2 U7 ( .A1(b), .A2(a), .ZN(n3) );
endmodule


module fa_39 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  NAND2_X4 U2 ( .A1(cin), .A2(n2), .ZN(n4) );
  XNOR2_X1 U3 ( .A(n1), .B(n5), .ZN(sum) );
  NAND2_X4 U4 ( .A1(n4), .A2(n3), .ZN(cout) );
  XNOR2_X2 U5 ( .A(b), .B(a), .ZN(n5) );
  INV_X4 U6 ( .A(n5), .ZN(n2) );
  NAND2_X2 U7 ( .A1(b), .A2(a), .ZN(n3) );
endmodule


module fa_38 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  NAND2_X4 U2 ( .A1(cin), .A2(n2), .ZN(n4) );
  NAND2_X4 U3 ( .A1(n4), .A2(n3), .ZN(cout) );
  XNOR2_X1 U4 ( .A(n1), .B(n5), .ZN(sum) );
  XNOR2_X2 U5 ( .A(b), .B(a), .ZN(n5) );
  INV_X4 U6 ( .A(n5), .ZN(n2) );
  NAND2_X2 U7 ( .A1(b), .A2(a), .ZN(n3) );
endmodule


module fa_37 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  NAND2_X4 U2 ( .A1(cin), .A2(n2), .ZN(n4) );
  NAND2_X4 U3 ( .A1(n4), .A2(n3), .ZN(cout) );
  XNOR2_X1 U4 ( .A(n1), .B(n5), .ZN(sum) );
  XNOR2_X2 U5 ( .A(b), .B(a), .ZN(n5) );
  INV_X4 U6 ( .A(n5), .ZN(n2) );
  NAND2_X2 U7 ( .A1(b), .A2(a), .ZN(n3) );
endmodule


module fa_36 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(n5), .ZN(sum) );
  NAND2_X4 U3 ( .A1(n4), .A2(n3), .ZN(cout) );
  NAND2_X4 U4 ( .A1(cin), .A2(n2), .ZN(n4) );
  XNOR2_X2 U5 ( .A(b), .B(a), .ZN(n5) );
  INV_X4 U6 ( .A(n5), .ZN(n2) );
  NAND2_X2 U7 ( .A1(b), .A2(a), .ZN(n3) );
endmodule


module fa_35 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  BUF_X32 U1 ( .A(n4), .Z(n1) );
  INV_X1 U2 ( .A(n1), .ZN(n2) );
  INV_X8 U3 ( .A(cin), .ZN(n4) );
  NAND2_X1 U4 ( .A1(b), .A2(a), .ZN(n5) );
  BUF_X32 U5 ( .A(n6), .Z(n3) );
  OAI21_X4 U6 ( .B1(n6), .B2(n4), .A(n5), .ZN(cout) );
  XNOR2_X1 U7 ( .A(n2), .B(n3), .ZN(sum) );
  XNOR2_X2 U8 ( .A(b), .B(a), .ZN(n6) );
endmodule


module fa_34 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  INV_X4 U1 ( .A(cin), .ZN(n4) );
  BUF_X32 U2 ( .A(n4), .Z(n1) );
  INV_X1 U3 ( .A(n1), .ZN(n2) );
  NAND2_X2 U4 ( .A1(b), .A2(a), .ZN(n3) );
  OAI21_X4 U5 ( .B1(n4), .B2(n5), .A(n3), .ZN(cout) );
  XNOR2_X1 U6 ( .A(n2), .B(n5), .ZN(sum) );
  XNOR2_X2 U7 ( .A(b), .B(a), .ZN(n5) );
endmodule


module fa_33 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  BUF_X8 U1 ( .A(b), .Z(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(a), .ZN(n2) );
  NAND2_X1 U3 ( .A1(a), .A2(b), .ZN(n4) );
  XOR2_X1 U4 ( .A(n2), .B(n3), .Z(sum) );
  INV_X1 U5 ( .A(cin), .ZN(n3) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n5) );
  OAI21_X4 U7 ( .B1(n5), .B2(n3), .A(n4), .ZN(cout) );
endmodule


module fa_nbit_0 ( A, B, cin, Sum, cout, of );
  input [0:31] A;
  input [0:31] B;
  output [0:31] Sum;
  input cin;
  output cout, of;

  wire   [1:31] carry;

  fa_0 \FA_NBIT[0].FA  ( .a(A[0]), .b(B[0]), .cin(carry[1]), .sum(Sum[0]) );
  fa_63 \FA_NBIT[1].FA  ( .a(A[1]), .b(B[1]), .cin(carry[2]), .sum(Sum[1]), 
        .cout(carry[1]) );
  fa_62 \FA_NBIT[2].FA  ( .a(A[2]), .b(B[2]), .cin(carry[3]), .sum(Sum[2]), 
        .cout(carry[2]) );
  fa_61 \FA_NBIT[3].FA  ( .a(A[3]), .b(B[3]), .cin(carry[4]), .sum(Sum[3]), 
        .cout(carry[3]) );
  fa_60 \FA_NBIT[4].FA  ( .a(A[4]), .b(B[4]), .cin(carry[5]), .sum(Sum[4]), 
        .cout(carry[4]) );
  fa_59 \FA_NBIT[5].FA  ( .a(A[5]), .b(B[5]), .cin(carry[6]), .sum(Sum[5]), 
        .cout(carry[5]) );
  fa_58 \FA_NBIT[6].FA  ( .a(A[6]), .b(B[6]), .cin(carry[7]), .sum(Sum[6]), 
        .cout(carry[6]) );
  fa_57 \FA_NBIT[7].FA  ( .a(A[7]), .b(B[7]), .cin(carry[8]), .sum(Sum[7]), 
        .cout(carry[7]) );
  fa_56 \FA_NBIT[8].FA  ( .a(A[8]), .b(B[8]), .cin(carry[9]), .sum(Sum[8]), 
        .cout(carry[8]) );
  fa_55 \FA_NBIT[9].FA  ( .a(A[9]), .b(B[9]), .cin(carry[10]), .sum(Sum[9]), 
        .cout(carry[9]) );
  fa_54 \FA_NBIT[10].FA  ( .a(A[10]), .b(B[10]), .cin(carry[11]), .sum(Sum[10]), .cout(carry[10]) );
  fa_53 \FA_NBIT[11].FA  ( .a(A[11]), .b(B[11]), .cin(carry[12]), .sum(Sum[11]), .cout(carry[11]) );
  fa_52 \FA_NBIT[12].FA  ( .a(A[12]), .b(B[12]), .cin(carry[13]), .sum(Sum[12]), .cout(carry[12]) );
  fa_51 \FA_NBIT[13].FA  ( .a(A[13]), .b(B[13]), .cin(carry[14]), .sum(Sum[13]), .cout(carry[13]) );
  fa_50 \FA_NBIT[14].FA  ( .a(A[14]), .b(B[14]), .cin(carry[15]), .sum(Sum[14]), .cout(carry[14]) );
  fa_49 \FA_NBIT[15].FA  ( .a(A[15]), .b(B[15]), .cin(carry[16]), .sum(Sum[15]), .cout(carry[15]) );
  fa_48 \FA_NBIT[16].FA  ( .a(A[16]), .b(B[16]), .cin(carry[17]), .sum(Sum[16]), .cout(carry[16]) );
  fa_47 \FA_NBIT[17].FA  ( .a(A[17]), .b(B[17]), .cin(carry[18]), .sum(Sum[17]), .cout(carry[17]) );
  fa_46 \FA_NBIT[18].FA  ( .a(A[18]), .b(B[18]), .cin(carry[19]), .sum(Sum[18]), .cout(carry[18]) );
  fa_45 \FA_NBIT[19].FA  ( .a(A[19]), .b(B[19]), .cin(carry[20]), .sum(Sum[19]), .cout(carry[19]) );
  fa_44 \FA_NBIT[20].FA  ( .a(A[20]), .b(B[20]), .cin(carry[21]), .sum(Sum[20]), .cout(carry[20]) );
  fa_43 \FA_NBIT[21].FA  ( .a(A[21]), .b(B[21]), .cin(carry[22]), .sum(Sum[21]), .cout(carry[21]) );
  fa_42 \FA_NBIT[22].FA  ( .a(A[22]), .b(B[22]), .cin(carry[23]), .sum(Sum[22]), .cout(carry[22]) );
  fa_41 \FA_NBIT[23].FA  ( .a(A[23]), .b(B[23]), .cin(carry[24]), .sum(Sum[23]), .cout(carry[23]) );
  fa_40 \FA_NBIT[24].FA  ( .a(A[24]), .b(B[24]), .cin(carry[25]), .sum(Sum[24]), .cout(carry[24]) );
  fa_39 \FA_NBIT[25].FA  ( .a(A[25]), .b(B[25]), .cin(carry[26]), .sum(Sum[25]), .cout(carry[25]) );
  fa_38 \FA_NBIT[26].FA  ( .a(A[26]), .b(B[26]), .cin(carry[27]), .sum(Sum[26]), .cout(carry[26]) );
  fa_37 \FA_NBIT[27].FA  ( .a(A[27]), .b(B[27]), .cin(carry[28]), .sum(Sum[27]), .cout(carry[27]) );
  fa_36 \FA_NBIT[28].FA  ( .a(A[28]), .b(B[28]), .cin(carry[29]), .sum(Sum[28]), .cout(carry[28]) );
  fa_35 \FA_NBIT[29].FA  ( .a(A[29]), .b(B[29]), .cin(carry[30]), .sum(Sum[29]), .cout(carry[29]) );
  fa_34 \FA_NBIT[30].FA  ( .a(A[30]), .b(B[30]), .cin(carry[31]), .sum(Sum[30]), .cout(carry[30]) );
  fa_33 \FA_NBIT[31].FA  ( .a(A[31]), .b(B[31]), .cin(cin), .sum(Sum[31]), 
        .cout(carry[31]) );
endmodule


module mux_1_832 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_831 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_830 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_829 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_828 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_827 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_826 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_825 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_824 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_823 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_822 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_821 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_820 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_819 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_818 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_817 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_816 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_815 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_814 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_813 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_812 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_811 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_810 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_809 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_808 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_807 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_806 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_805 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_804 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_803 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_802 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_801 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux2to1_32bit_26 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n2) );
  INV_X4 U2 ( .A(n4), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_832 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_831 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_830 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_829 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_828 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_827 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_826 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_825 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_824 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_823 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_822 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10]) );
  mux_1_821 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_820 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12]) );
  mux_1_819 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13]) );
  mux_1_818 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_817 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15]) );
  mux_1_816 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(1'b0), .sel(n2), .z(Z[16])
         );
  mux_1_815 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(1'b0), .sel(n2), .z(Z[17])
         );
  mux_1_814 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(1'b0), .sel(n2), .z(Z[18])
         );
  mux_1_813 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(1'b0), .sel(n2), .z(Z[19])
         );
  mux_1_812 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(1'b0), .sel(n2), .z(Z[20])
         );
  mux_1_811 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(1'b0), .sel(n2), .z(Z[21])
         );
  mux_1_810 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(1'b0), .sel(n2), .z(Z[22])
         );
  mux_1_809 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(1'b0), .sel(n2), .z(Z[23])
         );
  mux_1_808 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(1'b0), .sel(n3), .z(Z[24])
         );
  mux_1_807 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(1'b0), .sel(n3), .z(Z[25])
         );
  mux_1_806 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(1'b0), .sel(n3), .z(Z[26])
         );
  mux_1_805 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(1'b0), .sel(n3), .z(Z[27])
         );
  mux_1_804 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(1'b0), .sel(n3), .z(Z[28])
         );
  mux_1_803 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(1'b0), .sel(n3), .z(Z[29])
         );
  mux_1_802 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(1'b0), .sel(n3), .z(Z[30])
         );
  mux_1_801 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(1'b0), .sel(n3), .z(Z[31])
         );
endmodule


module mux_1_800 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_799 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_798 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_797 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_796 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_795 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_794 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_793 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_792 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_791 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_790 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_789 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_788 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_787 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_786 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_785 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_784 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_783 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_782 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_781 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_780 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_779 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_778 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_777 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_776 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_775 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_774 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_773 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_772 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_771 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_770 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_769 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux2to1_32bit_25 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3;

  INV_X4 U1 ( .A(n3), .ZN(n2) );
  INV_X4 U2 ( .A(n3), .ZN(n1) );
  INV_X4 U3 ( .A(sel), .ZN(n3) );
  mux_1_800 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_799 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_798 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_797 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_796 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_795 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_794 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_793 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_792 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_791 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_790 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10]) );
  mux_1_789 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_788 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12]) );
  mux_1_787 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13]) );
  mux_1_786 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_785 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15]) );
  mux_1_784 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16]) );
  mux_1_783 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17]) );
  mux_1_782 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18]) );
  mux_1_781 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19]) );
  mux_1_780 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_779 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21]) );
  mux_1_778 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_777 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_776 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(1'b0), .sel(sel), .z(Z[24]) );
  mux_1_775 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(1'b0), .sel(n1), .z(Z[25])
         );
  mux_1_774 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(1'b0), .sel(sel), .z(Z[26]) );
  mux_1_773 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(1'b0), .sel(sel), .z(Z[27]) );
  mux_1_772 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(1'b0), .sel(sel), .z(Z[28]) );
  mux_1_771 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(1'b0), .sel(sel), .z(Z[29]) );
  mux_1_770 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(1'b0), .sel(sel), .z(Z[30]) );
  mux_1_769 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(1'b0), .sel(sel), .z(Z[31]) );
endmodule


module mux_1_768 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_767 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_766 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_765 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_764 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_763 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_762 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_761 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_760 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_759 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_758 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_757 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_756 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_755 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_754 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_753 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_752 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_751 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_750 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_749 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_748 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_747 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_746 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_745 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_744 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_743 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_742 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_741 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_740 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_739 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_738 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_737 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux2to1_32bit_24 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3;

  INV_X4 U1 ( .A(n3), .ZN(n2) );
  INV_X4 U2 ( .A(n3), .ZN(n1) );
  INV_X4 U3 ( .A(sel), .ZN(n3) );
  mux_1_768 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_767 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_766 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_765 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_764 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_763 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_762 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_761 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_760 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_759 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_758 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10]) );
  mux_1_757 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_756 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12]) );
  mux_1_755 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13]) );
  mux_1_754 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_753 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15]) );
  mux_1_752 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16]) );
  mux_1_751 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17]) );
  mux_1_750 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18]) );
  mux_1_749 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19]) );
  mux_1_748 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_747 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21]) );
  mux_1_746 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_745 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_744 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(sel), .z(
        Z[24]) );
  mux_1_743 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(sel), .z(
        Z[25]) );
  mux_1_742 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(sel), .z(
        Z[26]) );
  mux_1_741 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(sel), .z(
        Z[27]) );
  mux_1_740 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(1'b0), .sel(sel), .z(Z[28]) );
  mux_1_739 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(1'b0), .sel(sel), .z(Z[29]) );
  mux_1_738 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(1'b0), .sel(sel), .z(Z[30]) );
  mux_1_737 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(1'b0), .sel(sel), .z(Z[31]) );
endmodule


module mux_1_736 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_735 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_734 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_733 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_732 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_731 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_730 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_729 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_728 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_727 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_726 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_725 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_724 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_723 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_722 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_721 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_720 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_719 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_718 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_717 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_716 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_715 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_714 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_713 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_712 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_711 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_710 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_709 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_708 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_707 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_706 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_705 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux2to1_32bit_23 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n2) );
  INV_X4 U2 ( .A(n4), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_736 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_735 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_734 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_733 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_732 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_731 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_730 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_729 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_728 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_727 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_726 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10]) );
  mux_1_725 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_724 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12]) );
  mux_1_723 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13]) );
  mux_1_722 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_721 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15]) );
  mux_1_720 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16]) );
  mux_1_719 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17]) );
  mux_1_718 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18]) );
  mux_1_717 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19]) );
  mux_1_716 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_715 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21]) );
  mux_1_714 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_713 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_712 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n3), .z(Z[24]) );
  mux_1_711 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n3), .z(Z[25]) );
  mux_1_710 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n3), .z(Z[26]) );
  mux_1_709 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n3), .z(Z[27]) );
  mux_1_708 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n3), .z(Z[28]) );
  mux_1_707 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n3), .z(Z[29]) );
  mux_1_706 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(1'b0), .sel(n3), .z(Z[30])
         );
  mux_1_705 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(1'b0), .sel(n3), .z(Z[31])
         );
endmodule


module mux_1_704 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_703 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_702 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_701 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_700 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_699 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_698 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_697 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_696 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_695 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_694 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_693 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_692 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_691 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_690 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_689 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_688 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_687 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_686 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_685 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_684 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_683 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_682 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_681 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_680 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_679 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_678 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_677 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_676 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_675 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_674 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_673 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux2to1_32bit_22 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3;

  INV_X4 U1 ( .A(n3), .ZN(n2) );
  INV_X4 U2 ( .A(n3), .ZN(n1) );
  INV_X4 U3 ( .A(sel), .ZN(n3) );
  mux_1_704 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_703 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_702 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_701 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_700 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_699 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_698 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_697 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_696 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_695 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_694 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10]) );
  mux_1_693 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_692 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12]) );
  mux_1_691 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13]) );
  mux_1_690 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_689 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15]) );
  mux_1_688 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16]) );
  mux_1_687 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17]) );
  mux_1_686 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18]) );
  mux_1_685 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19]) );
  mux_1_684 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_683 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21]) );
  mux_1_682 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_681 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_680 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(sel), .z(
        Z[24]) );
  mux_1_679 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(sel), .z(
        Z[25]) );
  mux_1_678 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(sel), .z(
        Z[26]) );
  mux_1_677 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(sel), .z(
        Z[27]) );
  mux_1_676 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(sel), .z(
        Z[28]) );
  mux_1_675 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(sel), .z(
        Z[29]) );
  mux_1_674 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(sel), .z(
        Z[30]) );
  mux_1_673 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(1'b0), .sel(sel), .z(Z[31]) );
endmodule


module mux_1_672 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_671 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_670 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_669 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_668 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_667 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_666 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_665 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_664 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_663 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_662 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_661 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_660 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_659 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_658 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_657 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_656 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_655 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_654 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_653 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_652 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_651 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_650 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_649 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_648 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_647 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_646 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_645 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_644 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_643 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_642 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_641 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux2to1_32bit_21 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3;

  INV_X4 U1 ( .A(n3), .ZN(n2) );
  INV_X4 U2 ( .A(n3), .ZN(n1) );
  INV_X4 U3 ( .A(sel), .ZN(n3) );
  mux_1_672 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_671 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_670 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_669 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_668 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_667 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_666 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_665 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_664 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_663 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_662 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10]) );
  mux_1_661 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_660 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12]) );
  mux_1_659 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13]) );
  mux_1_658 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_657 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15]) );
  mux_1_656 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16]) );
  mux_1_655 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17]) );
  mux_1_654 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18]) );
  mux_1_653 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19]) );
  mux_1_652 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_651 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21]) );
  mux_1_650 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_649 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_648 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n2), .z(Z[24]) );
  mux_1_647 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(sel), .z(
        Z[25]) );
  mux_1_646 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n2), .z(Z[26]) );
  mux_1_645 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n2), .z(Z[27]) );
  mux_1_644 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(sel), .z(
        Z[28]) );
  mux_1_643 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(sel), .z(
        Z[29]) );
  mux_1_642 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(sel), .z(
        Z[30]) );
  mux_1_641 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(sel), .z(
        Z[31]) );
endmodule


module mux_1_640 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_639 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_638 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_637 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_636 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_635 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_634 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_633 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_632 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_631 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_630 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_629 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_628 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_627 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_626 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_625 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_624 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_623 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_622 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_621 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_620 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_619 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_618 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_617 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_616 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_615 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_614 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_613 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_612 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_611 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_610 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_609 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux2to1_32bit_20 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n2) );
  INV_X4 U2 ( .A(n4), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_640 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_639 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_638 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_637 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_636 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_635 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_634 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_633 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_632 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_631 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_630 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10]) );
  mux_1_629 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_628 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12]) );
  mux_1_627 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13]) );
  mux_1_626 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_625 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15]) );
  mux_1_624 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16]) );
  mux_1_623 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17]) );
  mux_1_622 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18]) );
  mux_1_621 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19]) );
  mux_1_620 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_619 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21]) );
  mux_1_618 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_617 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_616 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n3), .z(Z[24]) );
  mux_1_615 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n3), .z(Z[25]) );
  mux_1_614 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n3), .z(Z[26]) );
  mux_1_613 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n3), .z(Z[27]) );
  mux_1_612 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n3), .z(Z[28]) );
  mux_1_611 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n3), .z(Z[29]) );
  mux_1_610 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(n3), .z(Z[30]) );
  mux_1_609 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n3), .z(Z[31]) );
endmodule


module mux_1_608 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_607 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_606 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_605 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_604 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_603 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_602 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_601 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_600 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_599 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_598 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_597 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_596 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_595 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_594 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_593 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_592 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_591 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_590 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_589 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_588 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_587 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_586 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_585 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_584 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_583 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_582 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_581 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_580 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_579 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_578 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_577 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux2to1_32bit_19 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n2) );
  INV_X4 U2 ( .A(n4), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_608 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_607 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_606 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_605 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_604 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_603 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_602 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_601 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_600 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_599 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_598 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10]) );
  mux_1_597 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_596 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12]) );
  mux_1_595 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13]) );
  mux_1_594 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_593 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15]) );
  mux_1_592 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16]) );
  mux_1_591 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17]) );
  mux_1_590 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18]) );
  mux_1_589 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19]) );
  mux_1_588 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_587 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21]) );
  mux_1_586 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_585 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_584 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n3), .z(Z[24]) );
  mux_1_583 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n3), .z(Z[25]) );
  mux_1_582 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n3), .z(Z[26]) );
  mux_1_581 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n3), .z(Z[27]) );
  mux_1_580 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n3), .z(Z[28]) );
  mux_1_579 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n3), .z(Z[29]) );
  mux_1_578 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(n3), .z(Z[30]) );
  mux_1_577 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n3), .z(Z[31]) );
endmodule


module mux_1_576 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_575 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_574 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_573 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_572 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_571 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_570 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_569 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_568 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_567 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_566 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_565 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_564 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_563 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_562 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_561 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_560 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_559 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_558 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_557 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_556 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_555 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_554 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_553 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_552 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_551 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_550 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_549 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_548 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_547 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_546 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_545 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux2to1_32bit_18 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n2) );
  INV_X4 U2 ( .A(n4), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_576 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_575 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_574 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_573 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_572 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_571 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_570 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_569 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_568 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_567 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_566 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10]) );
  mux_1_565 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_564 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12]) );
  mux_1_563 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13]) );
  mux_1_562 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_561 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15]) );
  mux_1_560 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16]) );
  mux_1_559 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17]) );
  mux_1_558 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18]) );
  mux_1_557 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19]) );
  mux_1_556 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_555 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21]) );
  mux_1_554 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_553 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_552 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n3), .z(Z[24]) );
  mux_1_551 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n3), .z(Z[25]) );
  mux_1_550 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n3), .z(Z[26]) );
  mux_1_549 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n3), .z(Z[27]) );
  mux_1_548 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n3), .z(Z[28]) );
  mux_1_547 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n3), .z(Z[29]) );
  mux_1_546 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(n3), .z(Z[30]) );
  mux_1_545 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n3), .z(Z[31]) );
endmodule


module mux_1_544 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_543 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_542 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_541 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_540 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_539 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_538 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_537 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_536 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_535 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_534 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_533 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_532 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_531 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_530 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_529 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_528 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_527 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_526 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_525 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_524 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_523 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_522 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_521 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_520 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_519 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_518 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_517 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_516 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_515 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_514 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_513 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux2to1_32bit_17 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n2) );
  INV_X4 U2 ( .A(n4), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_544 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_543 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_542 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_541 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_540 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_539 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_538 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_537 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_536 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_535 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_534 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10]) );
  mux_1_533 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_532 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12]) );
  mux_1_531 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13]) );
  mux_1_530 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_529 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15]) );
  mux_1_528 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16]) );
  mux_1_527 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17]) );
  mux_1_526 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18]) );
  mux_1_525 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19]) );
  mux_1_524 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_523 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21]) );
  mux_1_522 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_521 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_520 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n3), .z(Z[24]) );
  mux_1_519 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n3), .z(Z[25]) );
  mux_1_518 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n3), .z(Z[26]) );
  mux_1_517 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n3), .z(Z[27]) );
  mux_1_516 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n3), .z(Z[28]) );
  mux_1_515 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n3), .z(Z[29]) );
  mux_1_514 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(n3), .z(Z[30]) );
  mux_1_513 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n3), .z(Z[31]) );
endmodule


module mux_1_512 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_511 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_510 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_509 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_508 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_507 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_506 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_505 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_504 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_503 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_502 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_501 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_500 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_499 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_498 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_497 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_496 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_495 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_494 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_493 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_492 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_491 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_490 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_489 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_488 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_487 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_486 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_485 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_484 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_483 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_482 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_481 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux2to1_32bit_16 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n2) );
  INV_X4 U2 ( .A(n4), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_512 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_511 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_510 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_509 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_508 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_507 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_506 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_505 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_504 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_503 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_502 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10]) );
  mux_1_501 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_500 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12]) );
  mux_1_499 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13]) );
  mux_1_498 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_497 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15]) );
  mux_1_496 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16]) );
  mux_1_495 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17]) );
  mux_1_494 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18]) );
  mux_1_493 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19]) );
  mux_1_492 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_491 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21]) );
  mux_1_490 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_489 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_488 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n3), .z(Z[24]) );
  mux_1_487 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n3), .z(Z[25]) );
  mux_1_486 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n3), .z(Z[26]) );
  mux_1_485 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n3), .z(Z[27]) );
  mux_1_484 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n3), .z(Z[28]) );
  mux_1_483 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n3), .z(Z[29]) );
  mux_1_482 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(n3), .z(Z[30]) );
  mux_1_481 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n3), .z(Z[31]) );
endmodule


module shift ( X, shamt, arith, right, Z );
  input [0:31] X;
  input [0:4] shamt;
  output [0:31] Z;
  input arith, right;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  wire   [0:31] ltemp0;
  wire   [0:31] ltemp1;
  wire   [0:31] ltemp2;
  wire   [0:31] ltemp3;
  wire   [0:31] ltemp4;
  wire   [0:31] rtemp0;
  wire   [0:31] rtemp1;
  wire   [0:31] rtemp2;
  wire   [0:31] rtemp3;
  wire   [0:31] rtemp4;

  INV_X4 U2 ( .A(n1), .ZN(n2) );
  INV_X4 U3 ( .A(n1), .ZN(n3) );
  INV_X4 U4 ( .A(n12), .ZN(n11) );
  INV_X4 U5 ( .A(shamt[0]), .ZN(n12) );
  INV_X4 U6 ( .A(n10), .ZN(n9) );
  INV_X1 U7 ( .A(shamt[1]), .ZN(n10) );
  INV_X4 U8 ( .A(n8), .ZN(n7) );
  INV_X1 U9 ( .A(shamt[2]), .ZN(n8) );
  INV_X4 U10 ( .A(n1), .ZN(n4) );
  NAND2_X2 U11 ( .A1(arith), .A2(X[0]), .ZN(n1) );
  INV_X4 U12 ( .A(n6), .ZN(n5) );
  INV_X4 U13 ( .A(shamt[4]), .ZN(n6) );
  mux2to1_32bit_26 SHIFTLEFT16 ( .X(X), .Y({X[16:31], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sel(n11), .Z(ltemp0) );
  mux2to1_32bit_25 SHIFTLEFT8 ( .X(ltemp0), .Y({ltemp0[8:31], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sel(n9), .Z(ltemp1) );
  mux2to1_32bit_24 SHIFTLEFT4 ( .X(ltemp1), .Y({ltemp1[4:31], 1'b0, 1'b0, 1'b0, 
        1'b0}), .sel(n7), .Z(ltemp2) );
  mux2to1_32bit_23 SHIFTLEFT2 ( .X(ltemp2), .Y({ltemp2[2:31], 1'b0, 1'b0}), 
        .sel(shamt[3]), .Z(ltemp3) );
  mux2to1_32bit_22 SHIFTLEFT1 ( .X(ltemp3), .Y({ltemp3[1:31], 1'b0}), .sel(n5), 
        .Z(ltemp4) );
  mux2to1_32bit_21 SHIFTRIGHT16 ( .X(X), .Y({n3, n3, n3, n3, n2, n2, n2, n2, 
        n2, n2, n2, n2, n2, n2, n2, n2, X[0:15]}), .sel(n11), .Z(rtemp0) );
  mux2to1_32bit_20 SHIFTRIGHT8 ( .X(rtemp0), .Y({n3, n3, n3, n3, n3, n3, n3, 
        n3, rtemp0[0:23]}), .sel(n9), .Z(rtemp1) );
  mux2to1_32bit_19 SHIFTRIGHT4 ( .X(rtemp1), .Y({n4, n4, n4, n4, rtemp1[0:27]}), .sel(n7), .Z(rtemp2) );
  mux2to1_32bit_18 SHIFTRIGHT2 ( .X(rtemp2), .Y({n4, n4, rtemp2[0:29]}), .sel(
        shamt[3]), .Z(rtemp3) );
  mux2to1_32bit_17 SHIFTRIGHT1 ( .X(rtemp3), .Y({n4, rtemp3[0:30]}), .sel(n5), 
        .Z(rtemp4) );
  mux2to1_32bit_16 LEFTORRIGHT ( .X(ltemp4), .Y(rtemp4), .sel(right), .Z(Z) );
endmodule


module not_1_32 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_31 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_30 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_29 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_28 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_27 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_26 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_25 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_24 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_23 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_22 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_21 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_20 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_19 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_18 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_17 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_16 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_15 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_14 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_13 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_12 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_11 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_10 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_9 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_8 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_7 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_6 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_5 ( x, z );
  input x;
  output z;


  INV_X4 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_4 ( x, z );
  input x;
  output z;


  INV_X32 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_3 ( x, z );
  input x;
  output z;


  INV_X32 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_2 ( x, z );
  input x;
  output z;


  INV_X32 U1 ( .A(x), .ZN(z) );
endmodule


module not_1_1 ( x, z );
  input x;
  output z;


  INV_X32 U1 ( .A(x), .ZN(z) );
endmodule


module not_32_1 ( X, Z );
  input [0:31] X;
  output [0:31] Z;


  not_1_32 \NOT_32BIT[0].NOT_1  ( .x(X[0]), .z(Z[0]) );
  not_1_31 \NOT_32BIT[1].NOT_1  ( .x(X[1]), .z(Z[1]) );
  not_1_30 \NOT_32BIT[2].NOT_1  ( .x(X[2]), .z(Z[2]) );
  not_1_29 \NOT_32BIT[3].NOT_1  ( .x(X[3]), .z(Z[3]) );
  not_1_28 \NOT_32BIT[4].NOT_1  ( .x(X[4]), .z(Z[4]) );
  not_1_27 \NOT_32BIT[5].NOT_1  ( .x(X[5]), .z(Z[5]) );
  not_1_26 \NOT_32BIT[6].NOT_1  ( .x(X[6]), .z(Z[6]) );
  not_1_25 \NOT_32BIT[7].NOT_1  ( .x(X[7]), .z(Z[7]) );
  not_1_24 \NOT_32BIT[8].NOT_1  ( .x(X[8]), .z(Z[8]) );
  not_1_23 \NOT_32BIT[9].NOT_1  ( .x(X[9]), .z(Z[9]) );
  not_1_22 \NOT_32BIT[10].NOT_1  ( .x(X[10]), .z(Z[10]) );
  not_1_21 \NOT_32BIT[11].NOT_1  ( .x(X[11]), .z(Z[11]) );
  not_1_20 \NOT_32BIT[12].NOT_1  ( .x(X[12]), .z(Z[12]) );
  not_1_19 \NOT_32BIT[13].NOT_1  ( .x(X[13]), .z(Z[13]) );
  not_1_18 \NOT_32BIT[14].NOT_1  ( .x(X[14]), .z(Z[14]) );
  not_1_17 \NOT_32BIT[15].NOT_1  ( .x(X[15]), .z(Z[15]) );
  not_1_16 \NOT_32BIT[16].NOT_1  ( .x(X[16]), .z(Z[16]) );
  not_1_15 \NOT_32BIT[17].NOT_1  ( .x(X[17]), .z(Z[17]) );
  not_1_14 \NOT_32BIT[18].NOT_1  ( .x(X[18]), .z(Z[18]) );
  not_1_13 \NOT_32BIT[19].NOT_1  ( .x(X[19]), .z(Z[19]) );
  not_1_12 \NOT_32BIT[20].NOT_1  ( .x(X[20]), .z(Z[20]) );
  not_1_11 \NOT_32BIT[21].NOT_1  ( .x(X[21]), .z(Z[21]) );
  not_1_10 \NOT_32BIT[22].NOT_1  ( .x(X[22]), .z(Z[22]) );
  not_1_9 \NOT_32BIT[23].NOT_1  ( .x(X[23]), .z(Z[23]) );
  not_1_8 \NOT_32BIT[24].NOT_1  ( .x(X[24]), .z(Z[24]) );
  not_1_7 \NOT_32BIT[25].NOT_1  ( .x(X[25]), .z(Z[25]) );
  not_1_6 \NOT_32BIT[26].NOT_1  ( .x(X[26]), .z(Z[26]) );
  not_1_5 \NOT_32BIT[27].NOT_1  ( .x(X[27]), .z(Z[27]) );
  not_1_4 \NOT_32BIT[28].NOT_1  ( .x(X[28]), .z(Z[28]) );
  not_1_3 \NOT_32BIT[29].NOT_1  ( .x(X[29]), .z(Z[29]) );
  not_1_2 \NOT_32BIT[30].NOT_1  ( .x(X[30]), .z(Z[30]) );
  not_1_1 \NOT_32BIT[31].NOT_1  ( .x(X[31]), .z(Z[31]) );
endmodule


module fa_32 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n3, n4, n5, n6, n7, n8, n10, n12, n13, n14, n15;

  NAND2_X4 U7 ( .A1(n3), .A2(n4), .ZN(n6) );
  NAND2_X4 U8 ( .A1(n5), .A2(n6), .ZN(sum) );
  INV_X2 U9 ( .A(n10), .ZN(n4) );
  NAND2_X2 U10 ( .A1(b), .A2(a), .ZN(n8) );
  INV_X4 U11 ( .A(n8), .ZN(n7) );
  XNOR2_X2 U12 ( .A(b), .B(a), .ZN(n10) );
  INV_X8 U1 ( .A(cin), .ZN(n3) );
  INV_X8 U2 ( .A(n13), .ZN(cout) );
  AOI21_X4 U3 ( .B1(cin), .B2(n12), .A(n7), .ZN(n13) );
  INV_X4 U4 ( .A(n10), .ZN(n12) );
  NOR2_X4 U5 ( .A1(n3), .A2(n14), .ZN(n15) );
  INV_X4 U6 ( .A(n10), .ZN(n14) );
  INV_X4 U13 ( .A(n15), .ZN(n5) );
endmodule


module fa_31 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5;

  INV_X4 U1 ( .A(n4), .ZN(n3) );
  NAND2_X2 U2 ( .A1(n5), .A2(n4), .ZN(n1) );
  OAI21_X4 U3 ( .B1(cin), .B2(n3), .A(n1), .ZN(n2) );
  INV_X8 U4 ( .A(n2), .ZN(cout) );
  XNOR2_X1 U5 ( .A(cin), .B(n5), .ZN(sum) );
  NAND2_X2 U6 ( .A1(b), .A2(a), .ZN(n4) );
  XNOR2_X2 U7 ( .A(b), .B(a), .ZN(n5) );
endmodule


module fa_30 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n5, n7, n8;

  AND2_X2 U3 ( .A1(n5), .A2(n3), .ZN(n1) );
  NAND2_X2 U4 ( .A1(b), .A2(a), .ZN(n3) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n5) );
  XNOR2_X2 U1 ( .A(cin), .B(n5), .ZN(sum) );
  OAI21_X4 U2 ( .B1(cin), .B2(n2), .A(n7), .ZN(n8) );
  INV_X4 U5 ( .A(n1), .ZN(n7) );
  INV_X8 U7 ( .A(n8), .ZN(cout) );
  INV_X8 U8 ( .A(n3), .ZN(n2) );
endmodule


module fa_29 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n6, n8, n9;

  XNOR2_X2 U1 ( .A(n1), .B(n6), .ZN(sum) );
  AND2_X2 U3 ( .A1(n6), .A2(n4), .ZN(n2) );
  NAND2_X2 U4 ( .A1(b), .A2(a), .ZN(n4) );
  XNOR2_X2 U7 ( .A(b), .B(a), .ZN(n6) );
  BUF_X4 U2 ( .A(cin), .Z(n1) );
  OAI21_X4 U5 ( .B1(cin), .B2(n3), .A(n8), .ZN(n9) );
  INV_X4 U6 ( .A(n2), .ZN(n8) );
  INV_X8 U8 ( .A(n9), .ZN(cout) );
  INV_X8 U9 ( .A(n4), .ZN(n3) );
endmodule


module fa_28 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR2_X4 U1 ( .A1(cin), .A2(n4), .ZN(n6) );
  INV_X1 U2 ( .A(cin), .ZN(n1) );
  INV_X2 U3 ( .A(n1), .ZN(n2) );
  AND2_X2 U4 ( .A1(n7), .A2(n5), .ZN(n3) );
  XNOR2_X1 U5 ( .A(n2), .B(n7), .ZN(sum) );
  NAND2_X2 U6 ( .A1(b), .A2(a), .ZN(n5) );
  INV_X4 U7 ( .A(n5), .ZN(n4) );
  XNOR2_X2 U8 ( .A(b), .B(a), .ZN(n7) );
  NOR2_X4 U9 ( .A1(n6), .A2(n3), .ZN(cout) );
endmodule


module fa_27 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  BUF_X16 U1 ( .A(cin), .Z(n1) );
  AND2_X2 U2 ( .A1(n6), .A2(n4), .ZN(n2) );
  XNOR2_X1 U3 ( .A(n1), .B(n6), .ZN(sum) );
  NAND2_X2 U4 ( .A1(b), .A2(a), .ZN(n4) );
  INV_X4 U5 ( .A(n4), .ZN(n3) );
  NOR2_X4 U6 ( .A1(cin), .A2(n3), .ZN(n5) );
  XNOR2_X2 U7 ( .A(b), .B(a), .ZN(n6) );
  NOR2_X4 U8 ( .A1(n5), .A2(n2), .ZN(cout) );
endmodule


module fa_26 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  XNOR2_X2 U1 ( .A(n1), .B(n6), .ZN(sum) );
  BUF_X16 U2 ( .A(cin), .Z(n1) );
  AND2_X2 U3 ( .A1(n6), .A2(n4), .ZN(n2) );
  NAND2_X2 U4 ( .A1(b), .A2(a), .ZN(n4) );
  INV_X4 U5 ( .A(n4), .ZN(n3) );
  NOR2_X4 U6 ( .A1(cin), .A2(n3), .ZN(n5) );
  XNOR2_X2 U7 ( .A(b), .B(a), .ZN(n6) );
  NOR2_X4 U8 ( .A1(n5), .A2(n2), .ZN(cout) );
endmodule


module fa_25 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n2, n3, n4, n5, n6, n8, n9, n10;

  AND2_X2 U3 ( .A1(n6), .A2(n4), .ZN(n2) );
  NAND2_X2 U4 ( .A1(b), .A2(a), .ZN(n4) );
  INV_X4 U5 ( .A(n4), .ZN(n3) );
  NOR2_X4 U6 ( .A1(cin), .A2(n3), .ZN(n5) );
  XNOR2_X2 U7 ( .A(b), .B(a), .ZN(n6) );
  NOR2_X4 U8 ( .A1(n5), .A2(n2), .ZN(cout) );
  BUF_X16 U1 ( .A(cin), .Z(n8) );
  INV_X1 U2 ( .A(n8), .ZN(n9) );
  INV_X2 U9 ( .A(n9), .ZN(n10) );
  XNOR2_X1 U10 ( .A(n10), .B(n6), .ZN(sum) );
endmodule


module fa_24 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n3, n4, n6, n8, n9;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  XNOR2_X1 U4 ( .A(n1), .B(n6), .ZN(sum) );
  NAND2_X2 U5 ( .A1(b), .A2(a), .ZN(n4) );
  XNOR2_X2 U7 ( .A(b), .B(a), .ZN(n6) );
  AOI21_X4 U2 ( .B1(cin), .B2(n9), .A(n3), .ZN(n8) );
  INV_X4 U3 ( .A(n8), .ZN(cout) );
  INV_X8 U6 ( .A(n4), .ZN(n3) );
  INV_X4 U8 ( .A(n6), .ZN(n9) );
endmodule


module fa_23 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  NOR2_X4 U2 ( .A1(cin), .A2(n3), .ZN(n5) );
  AND2_X2 U3 ( .A1(n6), .A2(n4), .ZN(n2) );
  XNOR2_X1 U4 ( .A(n1), .B(n6), .ZN(sum) );
  NAND2_X2 U5 ( .A1(b), .A2(a), .ZN(n4) );
  INV_X4 U6 ( .A(n4), .ZN(n3) );
  XNOR2_X2 U7 ( .A(b), .B(a), .ZN(n6) );
  NOR2_X4 U8 ( .A1(n5), .A2(n2), .ZN(cout) );
endmodule


module fa_22 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  BUF_X32 U1 ( .A(cin), .Z(n1) );
  AND2_X2 U2 ( .A1(n6), .A2(n4), .ZN(n2) );
  XNOR2_X1 U3 ( .A(n1), .B(n6), .ZN(sum) );
  NAND2_X2 U4 ( .A1(b), .A2(a), .ZN(n4) );
  INV_X4 U5 ( .A(n4), .ZN(n3) );
  NOR2_X4 U6 ( .A1(cin), .A2(n3), .ZN(n5) );
  XNOR2_X2 U7 ( .A(b), .B(a), .ZN(n6) );
  NOR2_X4 U8 ( .A1(n5), .A2(n2), .ZN(cout) );
endmodule


module fa_21 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X4 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X2 U3 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U4 ( .A(n2), .B(n6), .ZN(sum) );
  NOR2_X4 U5 ( .A1(cin), .A2(n1), .ZN(n5) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NOR2_X4 U8 ( .A1(n5), .A2(n4), .ZN(cout) );
endmodule


module fa_20 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X4 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X2 U3 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U4 ( .A(n2), .B(n6), .ZN(sum) );
  NOR2_X4 U5 ( .A1(cin), .A2(n1), .ZN(n5) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NOR2_X4 U8 ( .A1(n5), .A2(n4), .ZN(cout) );
endmodule


module fa_19 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X4 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X2 U3 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U4 ( .A(n2), .B(n6), .ZN(sum) );
  NOR2_X4 U5 ( .A1(cin), .A2(n1), .ZN(n5) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NOR2_X4 U8 ( .A1(n5), .A2(n4), .ZN(cout) );
endmodule


module fa_18 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X4 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X2 U3 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U4 ( .A(n2), .B(n6), .ZN(sum) );
  NOR2_X4 U5 ( .A1(cin), .A2(n1), .ZN(n5) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NOR2_X4 U8 ( .A1(n5), .A2(n4), .ZN(cout) );
endmodule


module fa_17 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6, n7;

  NOR2_X2 U1 ( .A1(n1), .A2(n4), .ZN(n5) );
  AND2_X4 U2 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U3 ( .A(cin), .Z(n2) );
  XOR2_X1 U4 ( .A(n3), .B(n7), .Z(sum) );
  INV_X1 U5 ( .A(n2), .ZN(n3) );
  NOR2_X4 U6 ( .A1(cin), .A2(n1), .ZN(n6) );
  XNOR2_X2 U7 ( .A(b), .B(a), .ZN(n7) );
  INV_X4 U8 ( .A(n7), .ZN(n4) );
  NOR2_X4 U9 ( .A1(n6), .A2(n5), .ZN(cout) );
endmodule


module fa_16 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X4 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X4 U3 ( .A1(cin), .A2(n1), .ZN(n5) );
  NOR2_X2 U4 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U5 ( .A(n2), .B(n6), .ZN(sum) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NOR2_X4 U8 ( .A1(n5), .A2(n4), .ZN(cout) );
endmodule


module fa_15 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X2 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X4 U3 ( .A1(cin), .A2(n1), .ZN(n5) );
  NOR2_X2 U4 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U5 ( .A(n2), .B(n6), .ZN(sum) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NOR2_X4 U8 ( .A1(n5), .A2(n4), .ZN(cout) );
endmodule


module fa_14 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X2 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X4 U3 ( .A1(cin), .A2(n1), .ZN(n5) );
  NOR2_X2 U4 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U5 ( .A(n2), .B(n6), .ZN(sum) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NOR2_X4 U8 ( .A1(n5), .A2(n4), .ZN(cout) );
endmodule


module fa_13 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X2 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X4 U3 ( .A1(cin), .A2(n1), .ZN(n5) );
  NOR2_X2 U4 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U5 ( .A(n2), .B(n6), .ZN(sum) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NOR2_X4 U8 ( .A1(n5), .A2(n4), .ZN(cout) );
endmodule


module fa_12 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X2 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X4 U3 ( .A1(cin), .A2(n1), .ZN(n5) );
  NOR2_X2 U4 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U5 ( .A(n2), .B(n6), .ZN(sum) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NOR2_X4 U8 ( .A1(n5), .A2(n4), .ZN(cout) );
endmodule


module fa_11 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X4 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X4 U3 ( .A1(cin), .A2(n1), .ZN(n5) );
  NOR2_X4 U4 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U5 ( .A(n2), .B(n6), .ZN(sum) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NOR2_X4 U8 ( .A1(n5), .A2(n4), .ZN(cout) );
endmodule


module fa_10 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X2 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X4 U3 ( .A1(n5), .A2(n4), .ZN(cout) );
  NOR2_X4 U4 ( .A1(cin), .A2(n1), .ZN(n5) );
  NOR2_X2 U5 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U6 ( .A(n2), .B(n6), .ZN(sum) );
  XNOR2_X2 U7 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U8 ( .A(n6), .ZN(n3) );
endmodule


module fa_9 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X2 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X4 U3 ( .A1(cin), .A2(n1), .ZN(n5) );
  NOR2_X2 U4 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U5 ( .A(n2), .B(n6), .ZN(sum) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NOR2_X4 U8 ( .A1(n5), .A2(n4), .ZN(cout) );
endmodule


module fa_8 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X2 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X4 U3 ( .A1(cin), .A2(n1), .ZN(n5) );
  NOR2_X2 U4 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U5 ( .A(n2), .B(n6), .ZN(sum) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NOR2_X4 U8 ( .A1(n5), .A2(n4), .ZN(cout) );
endmodule


module fa_7 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X4 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X4 U3 ( .A1(cin), .A2(n1), .ZN(n5) );
  NOR2_X4 U4 ( .A1(n5), .A2(n4), .ZN(cout) );
  NOR2_X4 U5 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U6 ( .A(n2), .B(n6), .ZN(sum) );
  XNOR2_X2 U7 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U8 ( .A(n6), .ZN(n3) );
endmodule


module fa_6 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X4 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X4 U3 ( .A1(cin), .A2(n1), .ZN(n5) );
  NOR2_X2 U4 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U5 ( .A(n2), .B(n6), .ZN(sum) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NOR2_X4 U8 ( .A1(n5), .A2(n4), .ZN(cout) );
endmodule


module fa_5 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X2 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X4 U3 ( .A1(cin), .A2(n1), .ZN(n5) );
  NOR2_X4 U4 ( .A1(n1), .A2(n3), .ZN(n4) );
  XNOR2_X1 U5 ( .A(n2), .B(n6), .ZN(sum) );
  XNOR2_X2 U6 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U7 ( .A(n6), .ZN(n3) );
  NOR2_X4 U8 ( .A1(n5), .A2(n4), .ZN(cout) );
endmodule


module fa_4 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6;

  AND2_X4 U1 ( .A1(b), .A2(a), .ZN(n1) );
  BUF_X32 U2 ( .A(cin), .Z(n2) );
  NOR2_X4 U3 ( .A1(n5), .A2(n4), .ZN(cout) );
  NOR2_X4 U4 ( .A1(cin), .A2(n1), .ZN(n5) );
  XNOR2_X1 U6 ( .A(n2), .B(n6), .ZN(sum) );
  XNOR2_X2 U7 ( .A(b), .B(a), .ZN(n6) );
  INV_X4 U8 ( .A(n6), .ZN(n3) );
  NOR2_X4 U5 ( .A1(n1), .A2(n3), .ZN(n4) );
endmodule


module fa_3 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  NAND2_X4 U4 ( .A1(n4), .A2(n5), .ZN(n6) );
  BUF_X32 U5 ( .A(cin), .Z(n2) );
  NOR2_X4 U6 ( .A1(n9), .A2(n8), .ZN(cout) );
  NAND2_X2 U7 ( .A1(b), .A2(n7), .ZN(n4) );
  NAND2_X4 U8 ( .A1(n3), .A2(a), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(n10) );
  NOR2_X4 U11 ( .A1(cin), .A2(n1), .ZN(n9) );
  XNOR2_X1 U12 ( .A(n2), .B(n10), .ZN(sum) );
  AND2_X2 U1 ( .A1(b), .A2(a), .ZN(n1) );
  AND2_X4 U2 ( .A1(n3), .A2(n7), .ZN(n8) );
  INV_X2 U3 ( .A(b), .ZN(n3) );
  INV_X4 U9 ( .A(a), .ZN(n7) );
endmodule


module fa_2 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n3, n6, n7, n8, n9, n10, n12, n13, n14;

  NAND2_X4 U3 ( .A1(b), .A2(a), .ZN(n9) );
  BUF_X32 U5 ( .A(n10), .Z(n3) );
  XOR2_X1 U8 ( .A(n14), .B(n7), .Z(sum) );
  INV_X1 U11 ( .A(n3), .ZN(n7) );
  INV_X1 U1 ( .A(n13), .ZN(n6) );
  BUF_X32 U2 ( .A(n8), .Z(n12) );
  NOR2_X4 U4 ( .A1(b), .A2(a), .ZN(n13) );
  NAND2_X1 U6 ( .A1(n6), .A2(n9), .ZN(n10) );
  INV_X1 U7 ( .A(n12), .ZN(n14) );
  INV_X8 U9 ( .A(cin), .ZN(n8) );
  OAI21_X4 U10 ( .B1(n8), .B2(n13), .A(n9), .ZN(cout) );
endmodule


module fa_1 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2, n5;

  INV_X8 U1 ( .A(a), .ZN(n2) );
  INV_X16 U2 ( .A(b), .ZN(n5) );
  INV_X1 U3 ( .A(b), .ZN(n1) );
  XOR2_X1 U4 ( .A(n1), .B(a), .Z(sum) );
  NAND2_X4 U5 ( .A1(n5), .A2(n2), .ZN(cout) );
endmodule


module fa_nbit_1 ( A, B, cin, Sum, cout, of );
  input [0:31] A;
  input [0:31] B;
  output [0:31] Sum;
  input cin;
  output cout, of;
  wire   n3, n1, n4, n5, n6, n7;
  wire   [1:31] carry;

  fa_32 \FA_NBIT[0].FA  ( .a(A[0]), .b(B[0]), .cin(carry[1]), .sum(Sum[0]), 
        .cout(n3) );
  fa_31 \FA_NBIT[1].FA  ( .a(A[1]), .b(B[1]), .cin(carry[2]), .sum(Sum[1]), 
        .cout(carry[1]) );
  fa_30 \FA_NBIT[2].FA  ( .a(A[2]), .b(B[2]), .cin(carry[3]), .sum(Sum[2]), 
        .cout(carry[2]) );
  fa_29 \FA_NBIT[3].FA  ( .a(A[3]), .b(B[3]), .cin(carry[4]), .sum(Sum[3]), 
        .cout(carry[3]) );
  fa_28 \FA_NBIT[4].FA  ( .a(A[4]), .b(B[4]), .cin(carry[5]), .sum(Sum[4]), 
        .cout(carry[4]) );
  fa_27 \FA_NBIT[5].FA  ( .a(A[5]), .b(B[5]), .cin(carry[6]), .sum(Sum[5]), 
        .cout(carry[5]) );
  fa_26 \FA_NBIT[6].FA  ( .a(A[6]), .b(B[6]), .cin(carry[7]), .sum(Sum[6]), 
        .cout(carry[6]) );
  fa_25 \FA_NBIT[7].FA  ( .a(A[7]), .b(B[7]), .cin(carry[8]), .sum(Sum[7]), 
        .cout(carry[7]) );
  fa_24 \FA_NBIT[8].FA  ( .a(A[8]), .b(B[8]), .cin(carry[9]), .sum(Sum[8]), 
        .cout(carry[8]) );
  fa_23 \FA_NBIT[9].FA  ( .a(A[9]), .b(B[9]), .cin(carry[10]), .sum(Sum[9]), 
        .cout(carry[9]) );
  fa_22 \FA_NBIT[10].FA  ( .a(A[10]), .b(B[10]), .cin(carry[11]), .sum(Sum[10]), .cout(carry[10]) );
  fa_21 \FA_NBIT[11].FA  ( .a(A[11]), .b(B[11]), .cin(carry[12]), .sum(Sum[11]), .cout(carry[11]) );
  fa_20 \FA_NBIT[12].FA  ( .a(A[12]), .b(B[12]), .cin(carry[13]), .sum(Sum[12]), .cout(carry[12]) );
  fa_19 \FA_NBIT[13].FA  ( .a(A[13]), .b(B[13]), .cin(carry[14]), .sum(Sum[13]), .cout(carry[13]) );
  fa_18 \FA_NBIT[14].FA  ( .a(A[14]), .b(B[14]), .cin(carry[15]), .sum(Sum[14]), .cout(carry[14]) );
  fa_17 \FA_NBIT[15].FA  ( .a(A[15]), .b(B[15]), .cin(carry[16]), .sum(Sum[15]), .cout(carry[15]) );
  fa_16 \FA_NBIT[16].FA  ( .a(A[16]), .b(B[16]), .cin(carry[17]), .sum(Sum[16]), .cout(carry[16]) );
  fa_15 \FA_NBIT[17].FA  ( .a(A[17]), .b(B[17]), .cin(carry[18]), .sum(Sum[17]), .cout(carry[17]) );
  fa_14 \FA_NBIT[18].FA  ( .a(A[18]), .b(B[18]), .cin(carry[19]), .sum(Sum[18]), .cout(carry[18]) );
  fa_13 \FA_NBIT[19].FA  ( .a(A[19]), .b(B[19]), .cin(carry[20]), .sum(Sum[19]), .cout(carry[19]) );
  fa_12 \FA_NBIT[20].FA  ( .a(A[20]), .b(B[20]), .cin(carry[21]), .sum(Sum[20]), .cout(carry[20]) );
  fa_11 \FA_NBIT[21].FA  ( .a(A[21]), .b(B[21]), .cin(carry[22]), .sum(Sum[21]), .cout(carry[21]) );
  fa_10 \FA_NBIT[22].FA  ( .a(A[22]), .b(B[22]), .cin(carry[23]), .sum(Sum[22]), .cout(carry[22]) );
  fa_9 \FA_NBIT[23].FA  ( .a(A[23]), .b(B[23]), .cin(carry[24]), .sum(Sum[23]), 
        .cout(carry[23]) );
  fa_8 \FA_NBIT[24].FA  ( .a(A[24]), .b(B[24]), .cin(carry[25]), .sum(Sum[24]), 
        .cout(carry[24]) );
  fa_7 \FA_NBIT[25].FA  ( .a(A[25]), .b(B[25]), .cin(carry[26]), .sum(Sum[25]), 
        .cout(carry[25]) );
  fa_6 \FA_NBIT[26].FA  ( .a(A[26]), .b(B[26]), .cin(carry[27]), .sum(Sum[26]), 
        .cout(carry[26]) );
  fa_5 \FA_NBIT[27].FA  ( .a(A[27]), .b(B[27]), .cin(carry[28]), .sum(Sum[27]), 
        .cout(carry[27]) );
  fa_4 \FA_NBIT[28].FA  ( .a(A[28]), .b(B[28]), .cin(carry[29]), .sum(Sum[28]), 
        .cout(carry[28]) );
  fa_3 \FA_NBIT[29].FA  ( .a(A[29]), .b(B[29]), .cin(carry[30]), .sum(Sum[29]), 
        .cout(carry[29]) );
  fa_2 \FA_NBIT[30].FA  ( .a(A[30]), .b(B[30]), .cin(carry[31]), .sum(Sum[30]), 
        .cout(carry[30]) );
  fa_1 \FA_NBIT[31].FA  ( .a(A[31]), .b(B[31]), .cin(1'b1), .sum(Sum[31]), 
        .cout(carry[31]) );
  NAND2_X2 U1 ( .A1(n3), .A2(n1), .ZN(n6) );
  NAND2_X4 U2 ( .A1(n4), .A2(n5), .ZN(n7) );
  NAND2_X4 U4 ( .A1(n6), .A2(n7), .ZN(of) );
  INV_X8 U5 ( .A(n3), .ZN(n4) );
  INV_X4 U6 ( .A(n1), .ZN(n5) );
  INV_X2 U7 ( .A(carry[1]), .ZN(n1) );
endmodule


module zero_1 ( X, z );
  input [0:31] X;
  output z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;

  NOR4_X2 U1 ( .A1(X[5]), .A2(X[6]), .A3(X[7]), .A4(X[8]), .ZN(n7) );
  NAND2_X4 U3 ( .A1(n18), .A2(n17), .ZN(n19) );
  NOR2_X4 U4 ( .A1(n16), .A2(n15), .ZN(n18) );
  NOR2_X4 U5 ( .A1(X[0]), .A2(n19), .ZN(z) );
  NOR2_X2 U6 ( .A1(X[18]), .A2(X[19]), .ZN(n14) );
  OR3_X2 U7 ( .A1(X[14]), .A2(X[13]), .A3(n1), .ZN(n5) );
  OR2_X4 U8 ( .A1(X[15]), .A2(X[16]), .ZN(n1) );
  OR2_X2 U9 ( .A1(X[11]), .A2(X[12]), .ZN(n2) );
  OR3_X2 U10 ( .A1(X[29]), .A2(X[28]), .A3(n3), .ZN(n10) );
  OR2_X4 U11 ( .A1(X[30]), .A2(X[31]), .ZN(n3) );
  OR2_X2 U12 ( .A1(X[26]), .A2(X[27]), .ZN(n4) );
  INV_X2 U13 ( .A(X[1]), .ZN(n17) );
  INV_X2 U14 ( .A(X[2]), .ZN(n8) );
  NOR4_X2 U15 ( .A1(n5), .A2(n2), .A3(X[9]), .A4(X[10]), .ZN(n6) );
  INV_X4 U17 ( .A(X[17]), .ZN(n13) );
  NOR4_X2 U18 ( .A1(X[20]), .A2(X[21]), .A3(X[22]), .A4(X[23]), .ZN(n12) );
  NOR4_X2 U19 ( .A1(n10), .A2(n4), .A3(X[24]), .A4(X[25]), .ZN(n11) );
  NAND4_X2 U20 ( .A1(n14), .A2(n13), .A3(n12), .A4(n11), .ZN(n15) );
  NAND4_X2 U2 ( .A1(n9), .A2(n8), .A3(n7), .A4(n6), .ZN(n16) );
  NOR2_X2 U16 ( .A1(X[3]), .A2(X[4]), .ZN(n9) );
endmodule


module setter ( A, B, seq, sne, sle, slt, sge, sgt );
  input [0:31] A;
  input [0:31] B;
  output seq, sne, sle, slt, sge, sgt;
  wire   sub_of, n12, n1, n2, n3, n4, n5, n6;
  wire   [0:31] b_not;
  wire   [0:31] difference;

  INV_X2 U2 ( .A(difference[0]), .ZN(n4) );
  INV_X1 U4 ( .A(sne), .ZN(n1) );
  INV_X8 U5 ( .A(n12), .ZN(slt) );
  INV_X4 U6 ( .A(sub_of), .ZN(n3) );
  NOR2_X4 U9 ( .A1(slt), .A2(n1), .ZN(sgt) );
  NAND2_X4 U10 ( .A1(n3), .A2(n4), .ZN(n6) );
  NAND2_X4 U12 ( .A1(n5), .A2(n6), .ZN(n12) );
  not_32_1 NEGATE_B ( .X(B), .Z(b_not) );
  fa_nbit_1 FULL_ADDER ( .A(A), .B(b_not), .cin(1'b1), .Sum(difference), .of(
        sub_of) );
  zero_1 CHECK_EQ ( .X(difference), .z(seq) );
  NAND2_X2 U3 ( .A1(difference[0]), .A2(sub_of), .ZN(n5) );
  NAND2_X2 U7 ( .A1(n5), .A2(n6), .ZN(sge) );
  NAND2_X2 U8 ( .A1(n2), .A2(sge), .ZN(sle) );
  BUF_X4 U11 ( .A(sne), .Z(n2) );
  INV_X4 U13 ( .A(seq), .ZN(sne) );
endmodule


module extend_1to32_0 ( x, sign, Z );
  output [0:31] Z;
  input x, sign;
  wire   n1;

  INV_X4 U1 ( .A(n1), .ZN(Z[31]) );
  INV_X8 U2 ( .A(x), .ZN(n1) );
endmodule


module extend_1to32_5 ( x, sign, Z );
  output [0:31] Z;
  input x, sign;
  wire   n1;

  INV_X2 U1 ( .A(x), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(Z[31]) );
endmodule


module extend_1to32_4 ( x, sign, Z );
  output [0:31] Z;
  input x, sign;
  wire   n1;

  INV_X4 U1 ( .A(n1), .ZN(Z[31]) );
  INV_X4 U2 ( .A(x), .ZN(n1) );
endmodule


module extend_1to32_3 ( x, sign, Z );
  output [0:31] Z;
  input x, sign;
  wire   n1;

  INV_X4 U1 ( .A(n1), .ZN(Z[31]) );
  INV_X4 U2 ( .A(x), .ZN(n1) );
endmodule


module extend_1to32_2 ( x, sign, Z );
  output [0:31] Z;
  input x, sign;
  wire   n1;

  INV_X1 U1 ( .A(x), .ZN(n1) );
  INV_X2 U2 ( .A(n1), .ZN(Z[31]) );
endmodule


module extend_1to32_1 ( x, sign, Z );
  output [0:31] Z;
  input x, sign;
  wire   n1;

  INV_X8 U1 ( .A(n1), .ZN(Z[31]) );
  INV_X4 U2 ( .A(x), .ZN(n1) );
endmodule


module mux_1_384 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  NAND2_X2 U2 ( .A1(sel), .A2(y), .ZN(n3) );
  NAND2_X2 U3 ( .A1(x), .A2(n1), .ZN(n2) );
  NAND2_X2 U4 ( .A1(n3), .A2(n2), .ZN(z) );
endmodule


module mux_1_383 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X1 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_382 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  NAND2_X2 U1 ( .A1(y), .A2(sel), .ZN(n3) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  NAND2_X2 U3 ( .A1(x), .A2(n1), .ZN(n2) );
  NAND2_X2 U4 ( .A1(n3), .A2(n2), .ZN(z) );
endmodule


module mux_1_381 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_380 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X1 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_379 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X1 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_378 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_377 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_376 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_375 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_374 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_373 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_372 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_371 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_370 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_369 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_368 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_367 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_366 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_365 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_364 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_363 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_362 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_361 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_360 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_359 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_358 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_357 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_356 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_355 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_354 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_353 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux2to1_32bit_12 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n1) );
  INV_X4 U2 ( .A(n4), .ZN(n2) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_384 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n2), .z(Z[0]) );
  mux_1_383 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n3), .z(Z[1]) );
  mux_1_382 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n2), .z(Z[2]) );
  mux_1_381 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n3), .z(Z[3]) );
  mux_1_380 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n3), .z(Z[4]) );
  mux_1_379 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n3), .z(Z[5]) );
  mux_1_378 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n3), .z(Z[6]) );
  mux_1_377 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n3), .z(Z[7]) );
  mux_1_376 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n3), .z(Z[8]) );
  mux_1_375 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n3), .z(Z[9]) );
  mux_1_374 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n3), .z(Z[10]) );
  mux_1_373 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n3), .z(Z[11]) );
  mux_1_372 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n3), .z(Z[12]) );
  mux_1_371 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n3), .z(Z[13]) );
  mux_1_370 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n3), .z(Z[14]) );
  mux_1_369 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n3), .z(Z[15]) );
  mux_1_368 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n3), .z(Z[16]) );
  mux_1_367 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n3), .z(Z[17]) );
  mux_1_366 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n3), .z(Z[18]) );
  mux_1_365 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n3), .z(Z[19]) );
  mux_1_364 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n3), .z(Z[20]) );
  mux_1_363 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n1), .z(Z[21]) );
  mux_1_362 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n3), .z(Z[22]) );
  mux_1_361 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n1), .z(Z[23]) );
  mux_1_360 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n1), .z(Z[24]) );
  mux_1_359 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n2), .z(Z[25]) );
  mux_1_358 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n1), .z(Z[26]) );
  mux_1_357 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n2), .z(Z[27]) );
  mux_1_356 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n1), .z(Z[28]) );
  mux_1_355 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n1), .z(Z[29]) );
  mux_1_354 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(n2), .z(Z[30]) );
  mux_1_353 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n1), .z(Z[31]) );
endmodule


module mux_1_321 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  INV_X4 U2 ( .A(sel), .ZN(n1) );
  NAND2_X1 U3 ( .A1(x), .A2(n1), .ZN(n2) );
  NAND2_X4 U1 ( .A1(y), .A2(sel), .ZN(n3) );
  NAND2_X4 U4 ( .A1(n3), .A2(n2), .ZN(z) );
endmodule


module mux2to1_32bit_11 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;


  mux_1_321 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(sel), .z(
        Z[31]) );
endmodule


module mux_1_320 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_319 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_318 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_317 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(x), .ZN(n1) );
  NOR2_X2 U2 ( .A1(n1), .A2(sel), .ZN(z) );
endmodule


module mux_1_316 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_315 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_314 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_313 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_312 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_311 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_310 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_309 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_308 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_307 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_306 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_305 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_304 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_303 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_302 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  AND2_X2 U2 ( .A1(x), .A2(n1), .ZN(z) );
endmodule


module mux_1_301 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_300 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_299 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_298 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_297 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_296 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_295 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_294 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_293 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_292 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_291 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_290 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_289 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  NAND2_X4 U2 ( .A1(n3), .A2(n2), .ZN(z) );
  INV_X4 U3 ( .A(sel), .ZN(n1) );
  NAND2_X2 U4 ( .A1(x), .A2(n1), .ZN(n2) );
  NAND2_X4 U1 ( .A1(y), .A2(sel), .ZN(n3) );
endmodule


module mux2to1_32bit_10 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INV_X4 U1 ( .A(n6), .ZN(n1) );
  INV_X4 U2 ( .A(n6), .ZN(n2) );
  INV_X4 U3 ( .A(n6), .ZN(n4) );
  INV_X4 U4 ( .A(n6), .ZN(n3) );
  INV_X4 U5 ( .A(n6), .ZN(n5) );
  INV_X4 U6 ( .A(sel), .ZN(n6) );
  mux_1_320 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(1'b0), .sel(n2), .z(Z[0]) );
  mux_1_319 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(1'b0), .sel(n2), .z(Z[1]) );
  mux_1_318 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(1'b0), .sel(n5), .z(Z[2]) );
  mux_1_317 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(1'b0), .sel(n1), .z(Z[3]) );
  mux_1_316 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(1'b0), .sel(n3), .z(Z[4]) );
  mux_1_315 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(1'b0), .sel(n4), .z(Z[5]) );
  mux_1_314 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(1'b0), .sel(n5), .z(Z[6]) );
  mux_1_313 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(1'b0), .sel(n3), .z(Z[7]) );
  mux_1_312 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(1'b0), .sel(n4), .z(Z[8]) );
  mux_1_311 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(1'b0), .sel(n5), .z(Z[9]) );
  mux_1_310 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(1'b0), .sel(n3), .z(Z[10])
         );
  mux_1_309 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(1'b0), .sel(n4), .z(Z[11])
         );
  mux_1_308 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(1'b0), .sel(n5), .z(Z[12])
         );
  mux_1_307 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(1'b0), .sel(n3), .z(Z[13])
         );
  mux_1_306 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(1'b0), .sel(n4), .z(Z[14])
         );
  mux_1_305 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(1'b0), .sel(n5), .z(Z[15])
         );
  mux_1_304 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(1'b0), .sel(n3), .z(Z[16])
         );
  mux_1_303 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(1'b0), .sel(n4), .z(Z[17])
         );
  mux_1_302 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(1'b0), .sel(sel), .z(Z[18]) );
  mux_1_301 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(1'b0), .sel(n2), .z(Z[19])
         );
  mux_1_300 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(1'b0), .sel(n2), .z(Z[20])
         );
  mux_1_299 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(1'b0), .sel(n2), .z(Z[21])
         );
  mux_1_298 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(1'b0), .sel(n1), .z(Z[22])
         );
  mux_1_297 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(1'b0), .sel(n2), .z(Z[23])
         );
  mux_1_296 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(1'b0), .sel(n1), .z(Z[24])
         );
  mux_1_295 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(1'b0), .sel(n2), .z(Z[25])
         );
  mux_1_294 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(1'b0), .sel(n1), .z(Z[26])
         );
  mux_1_293 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(1'b0), .sel(n2), .z(Z[27])
         );
  mux_1_292 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(1'b0), .sel(n1), .z(Z[28])
         );
  mux_1_291 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(1'b0), .sel(n2), .z(Z[29])
         );
  mux_1_290 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(1'b0), .sel(n1), .z(Z[30])
         );
  mux_1_289 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n2), .z(Z[31]) );
endmodule


module mux4to1_32bit_0 ( in0, in1, in2, in3, sel, Z );
  input [0:31] in0;
  input [0:31] in1;
  input [0:31] in2;
  input [0:31] in3;
  input [0:1] sel;
  output [0:31] Z;
  wire   \bus2[31] ;
  wire   [0:31] bus1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  mux2to1_32bit_12 MUX_BUS1 ( .X(in0), .Y(in1), .sel(sel[1]), .Z(bus1) );
  mux2to1_32bit_11 MUX_BUS2 ( .X({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        in2[31]}), .Y({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, in3[31]}), 
        .sel(sel[1]), .Z({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, \bus2[31] }) );
  mux2to1_32bit_10 MUX_OUT ( .X(bus1), .Y({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \bus2[31] }), .sel(sel[0]), .Z(Z) );
endmodule


module mux_1_257 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  NAND2_X4 U1 ( .A1(x), .A2(n1), .ZN(n3) );
  NAND2_X4 U3 ( .A1(n3), .A2(n2), .ZN(z) );
  INV_X4 U4 ( .A(sel), .ZN(n1) );
  NAND2_X2 U2 ( .A1(y), .A2(sel), .ZN(n2) );
endmodule


module mux2to1_32bit_9 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;


  mux_1_257 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(sel), .z(
        Z[31]) );
endmodule


module mux_1_256 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_255 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_254 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_253 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_252 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_251 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_250 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_249 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_248 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_247 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_246 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_245 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_244 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_243 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_242 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_241 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_240 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_239 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_238 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_237 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_236 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_235 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_234 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_233 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_232 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_231 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_230 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_229 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_228 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_227 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_226 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_225 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux2to1_32bit_8 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n2) );
  INV_X4 U2 ( .A(n4), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_256 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_255 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_254 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_253 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_252 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_251 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_250 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_249 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_248 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_247 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_246 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10]) );
  mux_1_245 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_244 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12]) );
  mux_1_243 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13]) );
  mux_1_242 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_241 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15]) );
  mux_1_240 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16]) );
  mux_1_239 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17]) );
  mux_1_238 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18]) );
  mux_1_237 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19]) );
  mux_1_236 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_235 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21]) );
  mux_1_234 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_233 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_232 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n3), .z(Z[24]) );
  mux_1_231 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n3), .z(Z[25]) );
  mux_1_230 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n3), .z(Z[26]) );
  mux_1_229 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n3), .z(Z[27]) );
  mux_1_228 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n3), .z(Z[28]) );
  mux_1_227 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n3), .z(Z[29]) );
  mux_1_226 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(n3), .z(Z[30]) );
  mux_1_225 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n3), .z(Z[31]) );
endmodule


module mux_1_224 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_223 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_222 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_221 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_220 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_219 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_218 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_217 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_216 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_215 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_214 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_213 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_212 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_211 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_210 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_209 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_208 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_207 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_206 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_205 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_204 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_203 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_202 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_201 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_200 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_199 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_198 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_197 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_196 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_195 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_194 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_193 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  NAND2_X4 U1 ( .A1(n3), .A2(n2), .ZN(z) );
  NAND2_X4 U2 ( .A1(x), .A2(n1), .ZN(n3) );
  INV_X4 U3 ( .A(sel), .ZN(n1) );
  NAND2_X2 U4 ( .A1(y), .A2(sel), .ZN(n2) );
endmodule


module mux2to1_32bit_7 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;


  mux_1_224 \MUX2TO1_32BIT[0].MUX  ( .x(1'b0), .y(Y[0]), .sel(sel), .z(Z[0])
         );
  mux_1_223 \MUX2TO1_32BIT[1].MUX  ( .x(1'b0), .y(Y[1]), .sel(sel), .z(Z[1])
         );
  mux_1_222 \MUX2TO1_32BIT[2].MUX  ( .x(1'b0), .y(Y[2]), .sel(sel), .z(Z[2])
         );
  mux_1_221 \MUX2TO1_32BIT[3].MUX  ( .x(1'b0), .y(Y[3]), .sel(sel), .z(Z[3])
         );
  mux_1_220 \MUX2TO1_32BIT[4].MUX  ( .x(1'b0), .y(Y[4]), .sel(sel), .z(Z[4])
         );
  mux_1_219 \MUX2TO1_32BIT[5].MUX  ( .x(1'b0), .y(Y[5]), .sel(sel), .z(Z[5])
         );
  mux_1_218 \MUX2TO1_32BIT[6].MUX  ( .x(1'b0), .y(Y[6]), .sel(sel), .z(Z[6])
         );
  mux_1_217 \MUX2TO1_32BIT[7].MUX  ( .x(1'b0), .y(Y[7]), .sel(sel), .z(Z[7])
         );
  mux_1_216 \MUX2TO1_32BIT[8].MUX  ( .x(1'b0), .y(Y[8]), .sel(sel), .z(Z[8])
         );
  mux_1_215 \MUX2TO1_32BIT[9].MUX  ( .x(1'b0), .y(Y[9]), .sel(sel), .z(Z[9])
         );
  mux_1_214 \MUX2TO1_32BIT[10].MUX  ( .x(1'b0), .y(Y[10]), .sel(sel), .z(Z[10]) );
  mux_1_213 \MUX2TO1_32BIT[11].MUX  ( .x(1'b0), .y(Y[11]), .sel(sel), .z(Z[11]) );
  mux_1_212 \MUX2TO1_32BIT[12].MUX  ( .x(1'b0), .y(Y[12]), .sel(sel), .z(Z[12]) );
  mux_1_211 \MUX2TO1_32BIT[13].MUX  ( .x(1'b0), .y(Y[13]), .sel(sel), .z(Z[13]) );
  mux_1_210 \MUX2TO1_32BIT[14].MUX  ( .x(1'b0), .y(Y[14]), .sel(sel), .z(Z[14]) );
  mux_1_209 \MUX2TO1_32BIT[15].MUX  ( .x(1'b0), .y(Y[15]), .sel(sel), .z(Z[15]) );
  mux_1_208 \MUX2TO1_32BIT[16].MUX  ( .x(1'b0), .y(Y[16]), .sel(sel), .z(Z[16]) );
  mux_1_207 \MUX2TO1_32BIT[17].MUX  ( .x(1'b0), .y(Y[17]), .sel(sel), .z(Z[17]) );
  mux_1_206 \MUX2TO1_32BIT[18].MUX  ( .x(1'b0), .y(Y[18]), .sel(sel), .z(Z[18]) );
  mux_1_205 \MUX2TO1_32BIT[19].MUX  ( .x(1'b0), .y(Y[19]), .sel(sel), .z(Z[19]) );
  mux_1_204 \MUX2TO1_32BIT[20].MUX  ( .x(1'b0), .y(Y[20]), .sel(sel), .z(Z[20]) );
  mux_1_203 \MUX2TO1_32BIT[21].MUX  ( .x(1'b0), .y(Y[21]), .sel(sel), .z(Z[21]) );
  mux_1_202 \MUX2TO1_32BIT[22].MUX  ( .x(1'b0), .y(Y[22]), .sel(sel), .z(Z[22]) );
  mux_1_201 \MUX2TO1_32BIT[23].MUX  ( .x(1'b0), .y(Y[23]), .sel(sel), .z(Z[23]) );
  mux_1_200 \MUX2TO1_32BIT[24].MUX  ( .x(1'b0), .y(Y[24]), .sel(sel), .z(Z[24]) );
  mux_1_199 \MUX2TO1_32BIT[25].MUX  ( .x(1'b0), .y(Y[25]), .sel(sel), .z(Z[25]) );
  mux_1_198 \MUX2TO1_32BIT[26].MUX  ( .x(1'b0), .y(Y[26]), .sel(sel), .z(Z[26]) );
  mux_1_197 \MUX2TO1_32BIT[27].MUX  ( .x(1'b0), .y(Y[27]), .sel(sel), .z(Z[27]) );
  mux_1_196 \MUX2TO1_32BIT[28].MUX  ( .x(1'b0), .y(Y[28]), .sel(sel), .z(Z[28]) );
  mux_1_195 \MUX2TO1_32BIT[29].MUX  ( .x(1'b0), .y(Y[29]), .sel(sel), .z(Z[29]) );
  mux_1_194 \MUX2TO1_32BIT[30].MUX  ( .x(1'b0), .y(Y[30]), .sel(sel), .z(Z[30]) );
  mux_1_193 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(sel), .z(
        Z[31]) );
endmodule


module mux4to1_32bit_3 ( in0, in1, in2, in3, sel, Z );
  input [0:31] in0;
  input [0:31] in1;
  input [0:31] in2;
  input [0:31] in3;
  input [0:1] sel;
  output [0:31] Z;
  wire   \bus1[31] ;
  wire   [0:31] bus2;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  mux2to1_32bit_9 MUX_BUS1 ( .X({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        in0[31]}), .Y({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, in1[31]}), 
        .sel(sel[1]), .Z({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, \bus1[31] }) );
  mux2to1_32bit_8 MUX_BUS2 ( .X(in2), .Y(in3), .sel(sel[1]), .Z(bus2) );
  mux2to1_32bit_7 MUX_OUT ( .X({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \bus1[31] }), .Y(bus2), .sel(sel[0]), .Z(Z) );
endmodule


module mux_1_448 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2;

  INV_X4 U1 ( .A(x), .ZN(n2) );
  NAND2_X2 U2 ( .A1(sel), .A2(y), .ZN(n1) );
  OAI21_X4 U3 ( .B1(sel), .B2(n2), .A(n1), .ZN(z) );
endmodule


module mux_1_447 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  NAND2_X4 U1 ( .A1(n3), .A2(n2), .ZN(z) );
  NAND2_X4 U2 ( .A1(x), .A2(n1), .ZN(n2) );
  INV_X4 U3 ( .A(sel), .ZN(n1) );
  NAND2_X2 U4 ( .A1(sel), .A2(y), .ZN(n3) );
endmodule


module mux_1_446 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_445 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_444 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_443 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_442 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_441 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_440 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_439 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_438 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_437 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_436 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_435 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_434 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_433 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_432 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_431 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_430 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_429 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_428 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_427 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_426 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_425 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_424 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_423 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_422 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_421 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_420 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_419 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_418 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_417 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  NAND2_X4 U1 ( .A1(x), .A2(n1), .ZN(n3) );
  NAND2_X4 U3 ( .A1(n3), .A2(n2), .ZN(z) );
  INV_X4 U4 ( .A(sel), .ZN(n1) );
  NAND2_X4 U2 ( .A1(y), .A2(sel), .ZN(n2) );
endmodule


module mux2to1_32bit_14 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n1) );
  INV_X4 U2 ( .A(n4), .ZN(n2) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_448 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n3), .z(Z[0]) );
  mux_1_447 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_446 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n3), .z(Z[2]) );
  mux_1_445 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n3), .z(Z[3]) );
  mux_1_444 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n3), .z(Z[4]) );
  mux_1_443 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n3), .z(Z[5]) );
  mux_1_442 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n3), .z(Z[6]) );
  mux_1_441 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n3), .z(Z[7]) );
  mux_1_440 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n3), .z(Z[8]) );
  mux_1_439 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n3), .z(Z[9]) );
  mux_1_438 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n3), .z(Z[10]) );
  mux_1_437 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n3), .z(Z[11]) );
  mux_1_436 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n3), .z(Z[12]) );
  mux_1_435 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n3), .z(Z[13]) );
  mux_1_434 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n3), .z(Z[14]) );
  mux_1_433 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n3), .z(Z[15]) );
  mux_1_432 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n3), .z(Z[16]) );
  mux_1_431 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n3), .z(Z[17]) );
  mux_1_430 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n3), .z(Z[18]) );
  mux_1_429 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n1), .z(Z[19]) );
  mux_1_428 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_427 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n1), .z(Z[21]) );
  mux_1_426 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_425 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n1), .z(Z[23]) );
  mux_1_424 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n2), .z(Z[24]) );
  mux_1_423 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n2), .z(Z[25]) );
  mux_1_422 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n1), .z(Z[26]) );
  mux_1_421 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n2), .z(Z[27]) );
  mux_1_420 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n1), .z(Z[28]) );
  mux_1_419 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n2), .z(Z[29]) );
  mux_1_418 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(n1), .z(Z[30]) );
  mux_1_417 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n2), .z(Z[31]) );
endmodule


module mux8to1_32bit_0 ( in0, in1, in2, in3, in4, in5, in6, in7, sel, Z );
  input [0:31] in0;
  input [0:31] in1;
  input [0:31] in2;
  input [0:31] in3;
  input [0:31] in4;
  input [0:31] in5;
  input [0:31] in6;
  input [0:31] in7;
  input [0:2] sel;
  output [0:31] Z;

  wire   [0:31] bus1;
  wire   [0:31] bus2;

  mux4to1_32bit_0 MUX_BUS1 ( .in0(in0), .in1(in1), .in2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, in2[31]}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, in3[31]}), .sel(sel[1:2]), .Z(bus1) );
  mux4to1_32bit_3 MUX_BUS2 ( .in0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        in4[31]}), .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, in5[31]}), 
        .in2(in6), .in3(in7), .sel(sel[1:2]), .Z(bus2) );
  mux2to1_32bit_14 MUX_OUT ( .X(bus1), .Y(bus2), .sel(sel[0]), .Z(Z) );
endmodule


module mux_1_192 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_191 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_190 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_189 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_188 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_187 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_186 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_185 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_184 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_183 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_182 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_181 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_180 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_179 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_178 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_177 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_176 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_175 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_174 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_173 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_172 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_171 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_170 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_169 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_168 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_167 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_166 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_165 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_164 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_163 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_162 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_161 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux2to1_32bit_6 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n2) );
  INV_X4 U2 ( .A(n4), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_192 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_191 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_190 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_189 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_188 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_187 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_186 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_185 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_184 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_183 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_182 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10]) );
  mux_1_181 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_180 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12]) );
  mux_1_179 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13]) );
  mux_1_178 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_177 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15]) );
  mux_1_176 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16]) );
  mux_1_175 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17]) );
  mux_1_174 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18]) );
  mux_1_173 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19]) );
  mux_1_172 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_171 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21]) );
  mux_1_170 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_169 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_168 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n3), .z(Z[24]) );
  mux_1_167 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n3), .z(Z[25]) );
  mux_1_166 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n3), .z(Z[26]) );
  mux_1_165 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n3), .z(Z[27]) );
  mux_1_164 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n3), .z(Z[28]) );
  mux_1_163 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n3), .z(Z[29]) );
  mux_1_162 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(n3), .z(Z[30]) );
  mux_1_161 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n3), .z(Z[31]) );
endmodule


module mux_1_160 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_159 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_158 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_157 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_156 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_155 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_154 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_153 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_152 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_151 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_150 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_149 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_148 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_147 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_146 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_145 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_144 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_143 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_142 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_141 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_140 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_139 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_138 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_137 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_136 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_135 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_134 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_133 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_132 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_131 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_130 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_129 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  NAND2_X2 U2 ( .A1(x), .A2(n3), .ZN(n2) );
  NAND2_X2 U3 ( .A1(n1), .A2(n2), .ZN(z) );
  INV_X4 U4 ( .A(sel), .ZN(n3) );
  NAND2_X4 U1 ( .A1(y), .A2(sel), .ZN(n1) );
endmodule


module mux2to1_32bit_5 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n2) );
  INV_X4 U2 ( .A(n4), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_160 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(1'b0), .sel(n1), .z(Z[0]) );
  mux_1_159 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(1'b0), .sel(n1), .z(Z[1]) );
  mux_1_158 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(1'b0), .sel(n1), .z(Z[2]) );
  mux_1_157 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(1'b0), .sel(n1), .z(Z[3]) );
  mux_1_156 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(1'b0), .sel(n1), .z(Z[4]) );
  mux_1_155 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(1'b0), .sel(n1), .z(Z[5]) );
  mux_1_154 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(1'b0), .sel(n1), .z(Z[6]) );
  mux_1_153 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(1'b0), .sel(n1), .z(Z[7]) );
  mux_1_152 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(1'b0), .sel(n1), .z(Z[8]) );
  mux_1_151 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(1'b0), .sel(n1), .z(Z[9]) );
  mux_1_150 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(1'b0), .sel(n1), .z(Z[10])
         );
  mux_1_149 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(1'b0), .sel(n1), .z(Z[11])
         );
  mux_1_148 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(1'b0), .sel(n2), .z(Z[12])
         );
  mux_1_147 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(1'b0), .sel(n2), .z(Z[13])
         );
  mux_1_146 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(1'b0), .sel(n2), .z(Z[14])
         );
  mux_1_145 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(1'b0), .sel(n2), .z(Z[15])
         );
  mux_1_144 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(1'b0), .sel(n2), .z(Z[16])
         );
  mux_1_143 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(1'b0), .sel(n2), .z(Z[17])
         );
  mux_1_142 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(1'b0), .sel(n2), .z(Z[18])
         );
  mux_1_141 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(1'b0), .sel(n2), .z(Z[19])
         );
  mux_1_140 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(1'b0), .sel(n2), .z(Z[20])
         );
  mux_1_139 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(1'b0), .sel(n2), .z(Z[21])
         );
  mux_1_138 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(1'b0), .sel(n2), .z(Z[22])
         );
  mux_1_137 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(1'b0), .sel(n2), .z(Z[23])
         );
  mux_1_136 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(1'b0), .sel(n3), .z(Z[24])
         );
  mux_1_135 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(1'b0), .sel(n3), .z(Z[25])
         );
  mux_1_134 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(1'b0), .sel(n3), .z(Z[26])
         );
  mux_1_133 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(1'b0), .sel(n3), .z(Z[27])
         );
  mux_1_132 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(1'b0), .sel(n3), .z(Z[28])
         );
  mux_1_131 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(1'b0), .sel(n3), .z(Z[29])
         );
  mux_1_130 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(1'b0), .sel(n3), .z(Z[30])
         );
  mux_1_129 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n3), .z(Z[31]) );
endmodule


module mux_1_128 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_127 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_126 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_125 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_124 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_123 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_122 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_121 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_120 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_119 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_118 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_117 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_116 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_115 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_114 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_113 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_112 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_111 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_110 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_109 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_108 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_107 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_106 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_105 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_104 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_103 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_102 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_101 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_100 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_99 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_98 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_97 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux2to1_32bit_4 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n2) );
  INV_X4 U2 ( .A(n4), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_128 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_127 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_126 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_125 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_124 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_123 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_122 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_121 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_120 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_119 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_118 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10]) );
  mux_1_117 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_116 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12]) );
  mux_1_115 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13]) );
  mux_1_114 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_113 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15]) );
  mux_1_112 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16]) );
  mux_1_111 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17]) );
  mux_1_110 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18]) );
  mux_1_109 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19]) );
  mux_1_108 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_107 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21]) );
  mux_1_106 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_105 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_104 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n3), .z(Z[24]) );
  mux_1_103 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n3), .z(Z[25]) );
  mux_1_102 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n3), .z(Z[26]) );
  mux_1_101 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n3), .z(Z[27]) );
  mux_1_100 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n3), .z(Z[28]) );
  mux_1_99 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n3), .z(Z[29])
         );
  mux_1_98 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(n3), .z(Z[30])
         );
  mux_1_97 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n3), .z(Z[31])
         );
endmodule


module mux4to1_32bit_2 ( in0, in1, in2, in3, sel, Z );
  input [0:31] in0;
  input [0:31] in1;
  input [0:31] in2;
  input [0:31] in3;
  input [0:1] sel;
  output [0:31] Z;

  wire   [0:31] bus1;
  wire   [0:31] bus2;

  mux2to1_32bit_6 MUX_BUS1 ( .X(in0), .Y(in1), .sel(sel[1]), .Z(bus1) );
  mux2to1_32bit_5 MUX_BUS2 ( .X(in2), .Y({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, in3[31]}), .sel(sel[1]), .Z(bus2) );
  mux2to1_32bit_4 MUX_OUT ( .X(bus1), .Y(bus2), .sel(sel[0]), .Z(Z) );
endmodule


module mux_1_96 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_95 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_94 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_93 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_92 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_91 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_90 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_89 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_88 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_87 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_86 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_85 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_84 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_83 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_82 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_81 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_80 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_79 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_78 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_77 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_76 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_75 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_74 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_73 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_72 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_71 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_70 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_69 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_68 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_67 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_66 ( x, y, sel, z );
  input x, y, sel;
  output z;


  AND2_X4 U1 ( .A1(y), .A2(sel), .ZN(z) );
endmodule


module mux_1_65 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  NAND2_X4 U1 ( .A1(x), .A2(n1), .ZN(n2) );
  NAND2_X2 U2 ( .A1(y), .A2(sel), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n1) );
  NAND2_X4 U3 ( .A1(n2), .A2(n3), .ZN(z) );
endmodule


module mux2to1_32bit_3 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3;

  INV_X4 U1 ( .A(n3), .ZN(n1) );
  INV_X4 U2 ( .A(n3), .ZN(n2) );
  INV_X4 U3 ( .A(sel), .ZN(n3) );
  mux_1_96 \MUX2TO1_32BIT[0].MUX  ( .x(1'b0), .y(Y[0]), .sel(sel), .z(Z[0]) );
  mux_1_95 \MUX2TO1_32BIT[1].MUX  ( .x(1'b0), .y(Y[1]), .sel(n2), .z(Z[1]) );
  mux_1_94 \MUX2TO1_32BIT[2].MUX  ( .x(1'b0), .y(Y[2]), .sel(n2), .z(Z[2]) );
  mux_1_93 \MUX2TO1_32BIT[3].MUX  ( .x(1'b0), .y(Y[3]), .sel(n2), .z(Z[3]) );
  mux_1_92 \MUX2TO1_32BIT[4].MUX  ( .x(1'b0), .y(Y[4]), .sel(n2), .z(Z[4]) );
  mux_1_91 \MUX2TO1_32BIT[5].MUX  ( .x(1'b0), .y(Y[5]), .sel(n2), .z(Z[5]) );
  mux_1_90 \MUX2TO1_32BIT[6].MUX  ( .x(1'b0), .y(Y[6]), .sel(n2), .z(Z[6]) );
  mux_1_89 \MUX2TO1_32BIT[7].MUX  ( .x(1'b0), .y(Y[7]), .sel(n2), .z(Z[7]) );
  mux_1_88 \MUX2TO1_32BIT[8].MUX  ( .x(1'b0), .y(Y[8]), .sel(n2), .z(Z[8]) );
  mux_1_87 \MUX2TO1_32BIT[9].MUX  ( .x(1'b0), .y(Y[9]), .sel(n2), .z(Z[9]) );
  mux_1_86 \MUX2TO1_32BIT[10].MUX  ( .x(1'b0), .y(Y[10]), .sel(n2), .z(Z[10])
         );
  mux_1_85 \MUX2TO1_32BIT[11].MUX  ( .x(1'b0), .y(Y[11]), .sel(n2), .z(Z[11])
         );
  mux_1_84 \MUX2TO1_32BIT[12].MUX  ( .x(1'b0), .y(Y[12]), .sel(n2), .z(Z[12])
         );
  mux_1_83 \MUX2TO1_32BIT[13].MUX  ( .x(1'b0), .y(Y[13]), .sel(n2), .z(Z[13])
         );
  mux_1_82 \MUX2TO1_32BIT[14].MUX  ( .x(1'b0), .y(Y[14]), .sel(n2), .z(Z[14])
         );
  mux_1_81 \MUX2TO1_32BIT[15].MUX  ( .x(1'b0), .y(Y[15]), .sel(n2), .z(Z[15])
         );
  mux_1_80 \MUX2TO1_32BIT[16].MUX  ( .x(1'b0), .y(Y[16]), .sel(n2), .z(Z[16])
         );
  mux_1_79 \MUX2TO1_32BIT[17].MUX  ( .x(1'b0), .y(Y[17]), .sel(n2), .z(Z[17])
         );
  mux_1_78 \MUX2TO1_32BIT[18].MUX  ( .x(1'b0), .y(Y[18]), .sel(n1), .z(Z[18])
         );
  mux_1_77 \MUX2TO1_32BIT[19].MUX  ( .x(1'b0), .y(Y[19]), .sel(n1), .z(Z[19])
         );
  mux_1_76 \MUX2TO1_32BIT[20].MUX  ( .x(1'b0), .y(Y[20]), .sel(n1), .z(Z[20])
         );
  mux_1_75 \MUX2TO1_32BIT[21].MUX  ( .x(1'b0), .y(Y[21]), .sel(n1), .z(Z[21])
         );
  mux_1_74 \MUX2TO1_32BIT[22].MUX  ( .x(1'b0), .y(Y[22]), .sel(n1), .z(Z[22])
         );
  mux_1_73 \MUX2TO1_32BIT[23].MUX  ( .x(1'b0), .y(Y[23]), .sel(n1), .z(Z[23])
         );
  mux_1_72 \MUX2TO1_32BIT[24].MUX  ( .x(1'b0), .y(Y[24]), .sel(n1), .z(Z[24])
         );
  mux_1_71 \MUX2TO1_32BIT[25].MUX  ( .x(1'b0), .y(Y[25]), .sel(n1), .z(Z[25])
         );
  mux_1_70 \MUX2TO1_32BIT[26].MUX  ( .x(1'b0), .y(Y[26]), .sel(n1), .z(Z[26])
         );
  mux_1_69 \MUX2TO1_32BIT[27].MUX  ( .x(1'b0), .y(Y[27]), .sel(n1), .z(Z[27])
         );
  mux_1_68 \MUX2TO1_32BIT[28].MUX  ( .x(1'b0), .y(Y[28]), .sel(n1), .z(Z[28])
         );
  mux_1_67 \MUX2TO1_32BIT[29].MUX  ( .x(1'b0), .y(Y[29]), .sel(n1), .z(Z[29])
         );
  mux_1_66 \MUX2TO1_32BIT[30].MUX  ( .x(1'b0), .y(Y[30]), .sel(n1), .z(Z[30])
         );
  mux_1_65 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n1), .z(Z[31])
         );
endmodule


module mux_1_64 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_63 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_62 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_61 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_60 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_59 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_58 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_57 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_56 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_55 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_54 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_53 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_52 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_51 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_50 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_49 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_48 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_47 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_46 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_45 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_44 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_43 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_42 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_41 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_40 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_39 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_38 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_37 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_36 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_35 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_34 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_33 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux2to1_32bit_2 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n2) );
  INV_X4 U2 ( .A(n4), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_64 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_63 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_62 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_61 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_60 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_59 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_58 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_57 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_56 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_55 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_54 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10])
         );
  mux_1_53 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11])
         );
  mux_1_52 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12])
         );
  mux_1_51 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13])
         );
  mux_1_50 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14])
         );
  mux_1_49 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15])
         );
  mux_1_48 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16])
         );
  mux_1_47 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17])
         );
  mux_1_46 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18])
         );
  mux_1_45 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19])
         );
  mux_1_44 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20])
         );
  mux_1_43 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21])
         );
  mux_1_42 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22])
         );
  mux_1_41 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23])
         );
  mux_1_40 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n3), .z(Z[24])
         );
  mux_1_39 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n3), .z(Z[25])
         );
  mux_1_38 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n3), .z(Z[26])
         );
  mux_1_37 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n3), .z(Z[27])
         );
  mux_1_36 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n3), .z(Z[28])
         );
  mux_1_35 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n3), .z(Z[29])
         );
  mux_1_34 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(n3), .z(Z[30])
         );
  mux_1_33 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n3), .z(Z[31])
         );
endmodule


module mux_1_32 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_31 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_30 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_29 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_28 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_27 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_26 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_25 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_24 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_23 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_22 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_21 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_20 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_19 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_18 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_17 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_16 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_15 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_14 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_13 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_12 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_11 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_10 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_9 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_8 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_7 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_6 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_5 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_4 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_3 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_2 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_1 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux2to1_32bit_1 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n2) );
  INV_X4 U2 ( .A(n4), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_32 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_31 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_30 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_29 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_28 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_27 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_26 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_25 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_24 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_23 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_22 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10])
         );
  mux_1_21 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11])
         );
  mux_1_20 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12])
         );
  mux_1_19 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13])
         );
  mux_1_18 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14])
         );
  mux_1_17 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15])
         );
  mux_1_16 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16])
         );
  mux_1_15 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17])
         );
  mux_1_14 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18])
         );
  mux_1_13 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19])
         );
  mux_1_12 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20])
         );
  mux_1_11 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21])
         );
  mux_1_10 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22])
         );
  mux_1_9 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23])
         );
  mux_1_8 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n3), .z(Z[24])
         );
  mux_1_7 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n3), .z(Z[25])
         );
  mux_1_6 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n3), .z(Z[26])
         );
  mux_1_5 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n3), .z(Z[27])
         );
  mux_1_4 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n3), .z(Z[28])
         );
  mux_1_3 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n3), .z(Z[29])
         );
  mux_1_2 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(n3), .z(Z[30])
         );
  mux_1_1 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n3), .z(Z[31])
         );
endmodule


module mux4to1_32bit_1 ( in0, in1, in2, in3, sel, Z );
  input [0:31] in0;
  input [0:31] in1;
  input [0:31] in2;
  input [0:31] in3;
  input [0:1] sel;
  output [0:31] Z;

  wire   [0:31] bus1;
  wire   [0:31] bus2;

  mux2to1_32bit_3 MUX_BUS1 ( .X({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        in0[31]}), .Y(in1), .sel(sel[1]), .Z(bus1) );
  mux2to1_32bit_2 MUX_BUS2 ( .X(in2), .Y(in3), .sel(sel[1]), .Z(bus2) );
  mux2to1_32bit_1 MUX_OUT ( .X(bus1), .Y(bus2), .sel(sel[0]), .Z(Z) );
endmodule


module mux_1_416 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_415 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_414 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_413 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_412 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_411 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_410 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_409 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_408 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_407 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_406 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_405 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_404 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_403 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_402 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_401 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_400 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_399 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_398 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_397 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_396 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_395 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_394 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_393 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_392 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_391 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_390 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_389 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_388 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_387 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_386 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_385 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  INV_X4 U1 ( .A(sel), .ZN(n1) );
  NAND2_X2 U2 ( .A1(x), .A2(n1), .ZN(n3) );
  NAND2_X2 U3 ( .A1(y), .A2(sel), .ZN(n2) );
  NAND2_X2 U4 ( .A1(n3), .A2(n2), .ZN(z) );
endmodule


module mux2to1_32bit_13 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INV_X4 U1 ( .A(n6), .ZN(n1) );
  INV_X4 U2 ( .A(n6), .ZN(n2) );
  INV_X4 U3 ( .A(n6), .ZN(n4) );
  INV_X4 U4 ( .A(n6), .ZN(n3) );
  INV_X4 U5 ( .A(n6), .ZN(n5) );
  INV_X4 U6 ( .A(sel), .ZN(n6) );
  mux_1_416 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n5), .z(Z[0]) );
  mux_1_415 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n5), .z(Z[1]) );
  mux_1_414 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n5), .z(Z[2]) );
  mux_1_413 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n5), .z(Z[3]) );
  mux_1_412 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n3), .z(Z[4]) );
  mux_1_411 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n4), .z(Z[5]) );
  mux_1_410 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(sel), .z(Z[6])
         );
  mux_1_409 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n3), .z(Z[7]) );
  mux_1_408 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n4), .z(Z[8]) );
  mux_1_407 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(sel), .z(Z[9])
         );
  mux_1_406 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n3), .z(Z[10]) );
  mux_1_405 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n4), .z(Z[11]) );
  mux_1_404 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(sel), .z(
        Z[12]) );
  mux_1_403 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n3), .z(Z[13]) );
  mux_1_402 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n4), .z(Z[14]) );
  mux_1_401 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(sel), .z(
        Z[15]) );
  mux_1_400 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n3), .z(Z[16]) );
  mux_1_399 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n4), .z(Z[17]) );
  mux_1_398 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n5), .z(Z[18]) );
  mux_1_397 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n1), .z(Z[19]) );
  mux_1_396 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_395 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21]) );
  mux_1_394 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n1), .z(Z[22]) );
  mux_1_393 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_392 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n1), .z(Z[24]) );
  mux_1_391 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n2), .z(Z[25]) );
  mux_1_390 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n1), .z(Z[26]) );
  mux_1_389 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n2), .z(Z[27]) );
  mux_1_388 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n1), .z(Z[28]) );
  mux_1_387 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n2), .z(Z[29]) );
  mux_1_386 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(n1), .z(Z[30]) );
  mux_1_385 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n2), .z(Z[31]) );
endmodule


module mux8to1_32bit_1 ( in0, in1, in2, in3, in4, in5, in6, in7, sel, Z );
  input [0:31] in0;
  input [0:31] in1;
  input [0:31] in2;
  input [0:31] in3;
  input [0:31] in4;
  input [0:31] in5;
  input [0:31] in6;
  input [0:31] in7;
  input [0:2] sel;
  output [0:31] Z;

  wire   [0:31] bus1;
  wire   [0:31] bus2;

  mux4to1_32bit_2 MUX_BUS1 ( .in0(in0), .in1(in1), .in2(in2), .in3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, in3[31]}), .sel(sel[1:2]), .Z(bus1) );
  mux4to1_32bit_1 MUX_BUS2 ( .in0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        in4[31]}), .in1(in5), .in2(in6), .in3(in7), .sel(sel[1:2]), .Z(bus2)
         );
  mux2to1_32bit_13 MUX_OUT ( .X(bus1), .Y(bus2), .sel(sel[0]), .Z(Z) );
endmodule


module mux_1_480 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2;

  INV_X4 U1 ( .A(x), .ZN(n2) );
  NAND2_X2 U2 ( .A1(sel), .A2(y), .ZN(n1) );
  OAI21_X4 U3 ( .B1(n2), .B2(sel), .A(n1), .ZN(z) );
endmodule


module mux_1_479 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  NAND2_X4 U1 ( .A1(n2), .A2(n3), .ZN(z) );
  NAND2_X4 U2 ( .A1(x), .A2(n1), .ZN(n2) );
  INV_X4 U3 ( .A(sel), .ZN(n1) );
  NAND2_X2 U4 ( .A1(sel), .A2(y), .ZN(n3) );
endmodule


module mux_1_478 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_477 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_476 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_475 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_474 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_473 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_472 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_471 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_470 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_469 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_468 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_467 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_466 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_465 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_464 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_463 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_462 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_461 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_460 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_459 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_458 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_457 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_456 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_455 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_454 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_453 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_452 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_451 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_450 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_449 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  NAND2_X4 U1 ( .A1(y), .A2(sel), .ZN(n2) );
  NAND2_X4 U2 ( .A1(x), .A2(n1), .ZN(n3) );
  NAND2_X4 U3 ( .A1(n3), .A2(n2), .ZN(z) );
  INV_X4 U4 ( .A(sel), .ZN(n1) );
endmodule


module mux2to1_32bit_15 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3, n4;

  INV_X4 U1 ( .A(n4), .ZN(n1) );
  INV_X4 U2 ( .A(n4), .ZN(n2) );
  INV_X4 U3 ( .A(n4), .ZN(n3) );
  INV_X4 U4 ( .A(sel), .ZN(n4) );
  mux_1_480 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n3), .z(Z[0]) );
  mux_1_479 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_478 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(sel), .z(Z[2])
         );
  mux_1_477 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(sel), .z(Z[3])
         );
  mux_1_476 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(sel), .z(Z[4])
         );
  mux_1_475 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(sel), .z(Z[5])
         );
  mux_1_474 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(sel), .z(Z[6])
         );
  mux_1_473 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(sel), .z(Z[7])
         );
  mux_1_472 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(sel), .z(Z[8])
         );
  mux_1_471 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(sel), .z(Z[9])
         );
  mux_1_470 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(sel), .z(
        Z[10]) );
  mux_1_469 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(sel), .z(
        Z[11]) );
  mux_1_468 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(sel), .z(
        Z[12]) );
  mux_1_467 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(sel), .z(
        Z[13]) );
  mux_1_466 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(sel), .z(
        Z[14]) );
  mux_1_465 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(sel), .z(
        Z[15]) );
  mux_1_464 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(sel), .z(
        Z[16]) );
  mux_1_463 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(sel), .z(
        Z[17]) );
  mux_1_462 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(sel), .z(
        Z[18]) );
  mux_1_461 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n3), .z(Z[19]) );
  mux_1_460 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_459 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n1), .z(Z[21]) );
  mux_1_458 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_457 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n1), .z(Z[23]) );
  mux_1_456 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n2), .z(Z[24]) );
  mux_1_455 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n2), .z(Z[25]) );
  mux_1_454 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n1), .z(Z[26]) );
  mux_1_453 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n2), .z(Z[27]) );
  mux_1_452 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n1), .z(Z[28]) );
  mux_1_451 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n2), .z(Z[29]) );
  mux_1_450 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(n1), .z(Z[30]) );
  mux_1_449 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n3), .z(Z[31]) );
endmodule


module mux16to1_32bit ( in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, 
        in11, in12, in13, in14, in15, sel, Z );
  input [0:31] in0;
  input [0:31] in1;
  input [0:31] in2;
  input [0:31] in3;
  input [0:31] in4;
  input [0:31] in5;
  input [0:31] in6;
  input [0:31] in7;
  input [0:31] in8;
  input [0:31] in9;
  input [0:31] in10;
  input [0:31] in11;
  input [0:31] in12;
  input [0:31] in13;
  input [0:31] in14;
  input [0:31] in15;
  input [0:3] sel;
  output [0:31] Z;
  wire   n1, n2;
  wire   [0:31] bus1;
  wire   [0:31] bus2;

  INV_X4 U1 ( .A(n2), .ZN(n1) );
  INV_X1 U2 ( .A(sel[3]), .ZN(n2) );
  mux8to1_32bit_0 MUX_BUS1 ( .in0(in0), .in1(in1), .in2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, in2[31]}), .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, in3[31]}), .in4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        in4[31]}), .in5({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, in5[31]}), 
        .in6(in6), .in7(in7), .sel({sel[1:2], n1}), .Z(bus1) );
  mux8to1_32bit_1 MUX_BUS2 ( .in0(in8), .in1(in9), .in2(in10), .in3({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, in11[31]}), .in4({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, in12[31]}), .in5(in13), .in6(in14), .in7(in15), 
        .sel({sel[1:2], n1}), .Z(bus2) );
  mux2to1_32bit_15 MUX_OUT ( .X(bus1), .Y(bus2), .sel(sel[0]), .Z(Z) );
endmodule


module alu ( A, B, ctrl, ALUout, zero, of );
  input [0:31] A;
  input [0:31] B;
  input [0:3] ctrl;
  output [0:31] ALUout;
  output zero, of;
  wire   n3, sne_1bit, sle_1bit, slt_1bit, sge_1bit, sgt_1bit, \seq_out[31] ,
         \sne_out[31] , \sle_out[31] , \slt_out[31] , \sge_out[31] ,
         \sgt_out[31] , n1, n4;
  wire   [0:31] and_out;
  wire   [0:31] or_out;
  wire   [0:31] xor_out;
  wire   [0:31] b_not;
  wire   [0:31] add_sub_in;
  wire   [0:31] add_sub_out;
  wire   [0:31] shift_out;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185;

  BUF_X4 U2 ( .A(B[30]), .Z(n1) );
  and_32 AND_32 ( .X(A), .Y({B[0:29], n1, n4}), .Z(and_out) );
  or_32 OR_32 ( .X(A), .Y({B[0:29], n1, n4}), .Z(or_out) );
  xor_32 XOR_32 ( .X(A), .Y({B[0:29], n1, n4}), .Z(xor_out) );
  not_32_0 NEGATE_B ( .X(B), .Z(b_not) );
  mux2to1_32bit_27 ADD_OR_SUB ( .X(B), .Y(b_not), .sel(ctrl[3]), .Z(add_sub_in) );
  fa_nbit_0 FULL_ADDER ( .A(A), .B(add_sub_in), .cin(ctrl[3]), .Sum(
        add_sub_out) );
  shift SHIFTER ( .X(A), .shamt(B[27:31]), .arith(ctrl[1]), .right(ctrl[2]), 
        .Z(shift_out) );
  setter SET_FLAGS ( .A(A), .B(B), .seq(n3), .sne(sne_1bit), .sle(sle_1bit), 
        .slt(slt_1bit), .sge(sge_1bit), .sgt(sgt_1bit) );
  extend_1to32_0 EXTEND_SEQ ( .x(n3), .sign(1'b0), .Z({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, \seq_out[31] }) );
  extend_1to32_5 EXTEND_SNE ( .x(sne_1bit), .sign(1'b0), .Z({
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, \sne_out[31] }) );
  extend_1to32_4 EXTEND_SLE ( .x(sle_1bit), .sign(1'b0), .Z({
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, \sle_out[31] }) );
  extend_1to32_3 EXTEND_SLT ( .x(slt_1bit), .sign(1'b0), .Z({
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, 
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, 
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, 
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, 
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, 
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, 
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, 
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, 
        SYNOPSYS_UNCONNECTED__123, \slt_out[31] }) );
  extend_1to32_2 EXTEND_SGE ( .x(sge_1bit), .sign(1'b0), .Z({
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, \sge_out[31] }) );
  extend_1to32_1 EXTEND_SGT ( .x(sgt_1bit), .sign(1'b0), .Z({
        SYNOPSYS_UNCONNECTED__155, SYNOPSYS_UNCONNECTED__156, 
        SYNOPSYS_UNCONNECTED__157, SYNOPSYS_UNCONNECTED__158, 
        SYNOPSYS_UNCONNECTED__159, SYNOPSYS_UNCONNECTED__160, 
        SYNOPSYS_UNCONNECTED__161, SYNOPSYS_UNCONNECTED__162, 
        SYNOPSYS_UNCONNECTED__163, SYNOPSYS_UNCONNECTED__164, 
        SYNOPSYS_UNCONNECTED__165, SYNOPSYS_UNCONNECTED__166, 
        SYNOPSYS_UNCONNECTED__167, SYNOPSYS_UNCONNECTED__168, 
        SYNOPSYS_UNCONNECTED__169, SYNOPSYS_UNCONNECTED__170, 
        SYNOPSYS_UNCONNECTED__171, SYNOPSYS_UNCONNECTED__172, 
        SYNOPSYS_UNCONNECTED__173, SYNOPSYS_UNCONNECTED__174, 
        SYNOPSYS_UNCONNECTED__175, SYNOPSYS_UNCONNECTED__176, 
        SYNOPSYS_UNCONNECTED__177, SYNOPSYS_UNCONNECTED__178, 
        SYNOPSYS_UNCONNECTED__179, SYNOPSYS_UNCONNECTED__180, 
        SYNOPSYS_UNCONNECTED__181, SYNOPSYS_UNCONNECTED__182, 
        SYNOPSYS_UNCONNECTED__183, SYNOPSYS_UNCONNECTED__184, 
        SYNOPSYS_UNCONNECTED__185, \sgt_out[31] }) );
  mux16to1_32bit FINAL_MUX ( .in0(add_sub_out), .in1(add_sub_out), .in2({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \slt_out[31] }), .in3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \sle_out[31] }), .in4({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, \sgt_out[31] }), .in5({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, \sge_out[31] }), .in6(and_out), .in7(shift_out), 
        .in8(and_out), .in9(shift_out), .in10(shift_out), .in11({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \seq_out[31] }), .in12({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, \sne_out[31] }), .in13(and_out), .in14(or_out), 
        .in15(xor_out), .sel(ctrl), .Z(ALUout) );
  BUF_X4 U4 ( .A(B[31]), .Z(n4) );
endmodule


module mux_1_0 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  AND2_X4 U1 ( .A1(sel), .A2(y), .ZN(n1) );
  INV_X2 U2 ( .A(n3), .ZN(z) );
  INV_X4 U3 ( .A(sel), .ZN(n2) );
  AOI21_X2 U4 ( .B1(x), .B2(n2), .A(n1), .ZN(n3) );
endmodule


module mux_1_999 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X1 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_998 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X1 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_997 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X1 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_996 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X1 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_995 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X1 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_994 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_993 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_992 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_991 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_990 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_989 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_988 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_987 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_986 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_985 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_984 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_983 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_982 ( x, y, sel, z );
  input x, y, sel;
  output z;


  MUX2_X2 U1 ( .A(x), .B(y), .S(sel), .Z(z) );
endmodule


module mux_1_981 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_980 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_979 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_978 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_977 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_976 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_975 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_974 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_973 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_972 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_971 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_970 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_969 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n3;

  NAND2_X4 U1 ( .A1(x), .A2(n1), .ZN(n3) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  NAND2_X2 U3 ( .A1(y), .A2(sel), .ZN(n2) );
  NAND2_X2 U4 ( .A1(n3), .A2(n2), .ZN(z) );
endmodule


module mux2to1_32bit_0 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3;

  INV_X4 U1 ( .A(n3), .ZN(n1) );
  INV_X4 U2 ( .A(n3), .ZN(n2) );
  INV_X4 U3 ( .A(sel), .ZN(n3) );
  mux_1_0 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n2), .z(Z[0]) );
  mux_1_999 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(sel), .z(Z[1])
         );
  mux_1_998 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(sel), .z(Z[2])
         );
  mux_1_997 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(sel), .z(Z[3])
         );
  mux_1_996 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(sel), .z(Z[4])
         );
  mux_1_995 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(sel), .z(Z[5])
         );
  mux_1_994 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(sel), .z(Z[6])
         );
  mux_1_993 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(sel), .z(Z[7])
         );
  mux_1_992 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(sel), .z(Z[8])
         );
  mux_1_991 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(sel), .z(Z[9])
         );
  mux_1_990 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(sel), .z(
        Z[10]) );
  mux_1_989 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(sel), .z(
        Z[11]) );
  mux_1_988 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(sel), .z(
        Z[12]) );
  mux_1_987 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(sel), .z(
        Z[13]) );
  mux_1_986 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(sel), .z(
        Z[14]) );
  mux_1_985 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(sel), .z(
        Z[15]) );
  mux_1_984 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(sel), .z(
        Z[16]) );
  mux_1_983 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(sel), .z(
        Z[17]) );
  mux_1_982 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(sel), .z(
        Z[18]) );
  mux_1_981 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19]) );
  mux_1_980 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n1), .z(Z[20]) );
  mux_1_979 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n1), .z(Z[21]) );
  mux_1_978 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n1), .z(Z[22]) );
  mux_1_977 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_976 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(n1), .z(Z[24]) );
  mux_1_975 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(n2), .z(Z[25]) );
  mux_1_974 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(n1), .z(Z[26]) );
  mux_1_973 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(n2), .z(Z[27]) );
  mux_1_972 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(n1), .z(Z[28]) );
  mux_1_971 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(n2), .z(Z[29]) );
  mux_1_970 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(n1), .z(Z[30]) );
  mux_1_969 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(n1), .z(Z[31]) );
endmodule


module multiplier_DW01_add_0 ( A, B, CI, SUM, CO );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [15:2] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(SUM[16]), .S(SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X2 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X4 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module multiplier_DW01_add_1 ( A, B, CI, SUM, CO );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [15:2] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(SUM[16]), .S(SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X2 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X4 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module multiplier_DW01_add_3 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16, n17,
         n33;
  wire   [32:18] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(n33), .CO(carry[18]), .S(SUM[17]) );
  XOR2_X2 U1 ( .A(B[33]), .B(n17), .Z(SUM[33]) );
  AND2_X4 U2 ( .A1(B[45]), .A2(n11), .ZN(n2) );
  AND2_X4 U3 ( .A1(B[43]), .A2(n12), .ZN(n3) );
  AND2_X4 U4 ( .A1(B[41]), .A2(n13), .ZN(n4) );
  AND2_X4 U5 ( .A1(B[39]), .A2(n14), .ZN(n5) );
  AND2_X4 U6 ( .A1(B[37]), .A2(n15), .ZN(n6) );
  AND2_X4 U7 ( .A1(B[35]), .A2(n16), .ZN(n7) );
  AND2_X4 U8 ( .A1(B[33]), .A2(n17), .ZN(n8) );
  XOR2_X2 U9 ( .A(B[32]), .B(carry[32]), .Z(SUM[32]) );
  AND2_X4 U10 ( .A1(B[46]), .A2(n2), .ZN(n10) );
  AND2_X4 U11 ( .A1(B[44]), .A2(n3), .ZN(n11) );
  AND2_X4 U12 ( .A1(B[42]), .A2(n4), .ZN(n12) );
  AND2_X4 U13 ( .A1(B[40]), .A2(n5), .ZN(n13) );
  AND2_X4 U14 ( .A1(B[38]), .A2(n6), .ZN(n14) );
  AND2_X4 U15 ( .A1(B[36]), .A2(n7), .ZN(n15) );
  AND2_X4 U16 ( .A1(B[34]), .A2(n8), .ZN(n16) );
  AND2_X4 U17 ( .A1(B[32]), .A2(carry[32]), .ZN(n17) );
  XOR2_X2 U18 ( .A(B[34]), .B(n8), .Z(SUM[34]) );
  XOR2_X2 U19 ( .A(B[35]), .B(n16), .Z(SUM[35]) );
  XOR2_X2 U20 ( .A(B[36]), .B(n7), .Z(SUM[36]) );
  XOR2_X2 U21 ( .A(B[37]), .B(n15), .Z(SUM[37]) );
  XOR2_X2 U22 ( .A(B[38]), .B(n6), .Z(SUM[38]) );
  XOR2_X2 U23 ( .A(B[39]), .B(n14), .Z(SUM[39]) );
  XOR2_X2 U24 ( .A(B[40]), .B(n5), .Z(SUM[40]) );
  XOR2_X2 U25 ( .A(B[41]), .B(n13), .Z(SUM[41]) );
  XOR2_X2 U26 ( .A(B[42]), .B(n4), .Z(SUM[42]) );
  XOR2_X2 U27 ( .A(B[43]), .B(n12), .Z(SUM[43]) );
  XOR2_X2 U28 ( .A(B[44]), .B(n3), .Z(SUM[44]) );
  XOR2_X2 U29 ( .A(B[45]), .B(n11), .Z(SUM[45]) );
  XOR2_X2 U30 ( .A(B[46]), .B(n2), .Z(SUM[46]) );
  XOR2_X2 U31 ( .A(B[47]), .B(n10), .Z(SUM[47]) );
  AND2_X4 U32 ( .A1(B[47]), .A2(n10), .ZN(SUM[48]) );
  AND2_X4 U33 ( .A1(B[16]), .A2(A[16]), .ZN(n33) );
  XOR2_X2 U34 ( .A(B[16]), .B(A[16]), .Z(SUM[16]) );
  BUF_X32 U35 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X32 U36 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X32 U37 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X32 U38 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X32 U39 ( .A(A[4]), .Z(SUM[4]) );
  BUF_X32 U40 ( .A(A[5]), .Z(SUM[5]) );
  BUF_X32 U41 ( .A(A[6]), .Z(SUM[6]) );
  BUF_X32 U42 ( .A(A[7]), .Z(SUM[7]) );
  BUF_X32 U43 ( .A(A[8]), .Z(SUM[8]) );
  BUF_X32 U44 ( .A(A[9]), .Z(SUM[9]) );
  BUF_X32 U45 ( .A(A[10]), .Z(SUM[10]) );
  BUF_X32 U46 ( .A(A[11]), .Z(SUM[11]) );
  BUF_X32 U47 ( .A(A[12]), .Z(SUM[12]) );
  BUF_X32 U48 ( .A(A[13]), .Z(SUM[13]) );
  BUF_X32 U49 ( .A(A[14]), .Z(SUM[14]) );
  BUF_X32 U50 ( .A(A[15]), .Z(SUM[15]) );
endmodule


module multiplier_DW01_add_2 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;
  wire   [49:34] carry;

  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(n14), .CO(carry[34]), .S(SUM[33]) );
  AND2_X4 U1 ( .A1(A[60]), .A2(n8), .ZN(n1) );
  AND2_X4 U2 ( .A1(A[58]), .A2(n9), .ZN(n2) );
  AND2_X4 U3 ( .A1(A[56]), .A2(n10), .ZN(n3) );
  AND2_X4 U4 ( .A1(A[54]), .A2(n11), .ZN(n4) );
  AND2_X4 U5 ( .A1(A[52]), .A2(n12), .ZN(n5) );
  AND2_X4 U6 ( .A1(A[50]), .A2(n13), .ZN(n6) );
  AND2_X4 U7 ( .A1(A[61]), .A2(n1), .ZN(n7) );
  AND2_X4 U8 ( .A1(A[59]), .A2(n2), .ZN(n8) );
  AND2_X4 U9 ( .A1(A[57]), .A2(n3), .ZN(n9) );
  AND2_X4 U10 ( .A1(A[55]), .A2(n4), .ZN(n10) );
  AND2_X4 U11 ( .A1(A[53]), .A2(n5), .ZN(n11) );
  AND2_X4 U12 ( .A1(A[51]), .A2(n6), .ZN(n12) );
  AND2_X4 U13 ( .A1(A[49]), .A2(carry[49]), .ZN(n13) );
  AND2_X4 U14 ( .A1(B[32]), .A2(A[32]), .ZN(n14) );
  AND2_X4 U15 ( .A1(A[62]), .A2(n7), .ZN(n15) );
  XOR2_X2 U16 ( .A(A[49]), .B(carry[49]), .Z(SUM[49]) );
  XOR2_X2 U17 ( .A(B[32]), .B(A[32]), .Z(SUM[32]) );
  XOR2_X2 U18 ( .A(A[50]), .B(n13), .Z(SUM[50]) );
  XOR2_X2 U19 ( .A(A[51]), .B(n6), .Z(SUM[51]) );
  XOR2_X2 U20 ( .A(A[52]), .B(n12), .Z(SUM[52]) );
  XOR2_X2 U21 ( .A(A[53]), .B(n5), .Z(SUM[53]) );
  XOR2_X2 U22 ( .A(A[54]), .B(n11), .Z(SUM[54]) );
  XOR2_X2 U23 ( .A(A[55]), .B(n4), .Z(SUM[55]) );
  XOR2_X2 U24 ( .A(A[56]), .B(n10), .Z(SUM[56]) );
  XOR2_X2 U25 ( .A(A[57]), .B(n3), .Z(SUM[57]) );
  XOR2_X2 U26 ( .A(A[58]), .B(n9), .Z(SUM[58]) );
  XOR2_X2 U27 ( .A(A[59]), .B(n2), .Z(SUM[59]) );
  XOR2_X2 U28 ( .A(A[60]), .B(n8), .Z(SUM[60]) );
  XOR2_X2 U29 ( .A(A[61]), .B(n1), .Z(SUM[61]) );
  XOR2_X2 U30 ( .A(A[62]), .B(n7), .Z(SUM[62]) );
  XOR2_X2 U31 ( .A(A[63]), .B(n15), .Z(SUM[63]) );
  BUF_X32 U32 ( .A(B[0]), .Z(SUM[0]) );
  BUF_X32 U33 ( .A(B[1]), .Z(SUM[1]) );
  BUF_X32 U34 ( .A(B[2]), .Z(SUM[2]) );
  BUF_X32 U35 ( .A(B[3]), .Z(SUM[3]) );
  BUF_X32 U36 ( .A(B[4]), .Z(SUM[4]) );
  BUF_X32 U37 ( .A(B[5]), .Z(SUM[5]) );
  BUF_X32 U38 ( .A(B[6]), .Z(SUM[6]) );
  BUF_X32 U39 ( .A(B[7]), .Z(SUM[7]) );
  BUF_X32 U40 ( .A(B[8]), .Z(SUM[8]) );
  BUF_X32 U41 ( .A(B[9]), .Z(SUM[9]) );
  BUF_X32 U42 ( .A(B[10]), .Z(SUM[10]) );
  BUF_X32 U43 ( .A(B[11]), .Z(SUM[11]) );
  BUF_X32 U44 ( .A(B[12]), .Z(SUM[12]) );
  BUF_X32 U45 ( .A(B[13]), .Z(SUM[13]) );
  BUF_X32 U46 ( .A(B[14]), .Z(SUM[14]) );
  BUF_X32 U47 ( .A(B[15]), .Z(SUM[15]) );
  BUF_X32 U48 ( .A(B[16]), .Z(SUM[16]) );
  BUF_X32 U49 ( .A(B[17]), .Z(SUM[17]) );
  BUF_X32 U50 ( .A(B[18]), .Z(SUM[18]) );
  BUF_X32 U51 ( .A(B[19]), .Z(SUM[19]) );
  BUF_X32 U52 ( .A(B[20]), .Z(SUM[20]) );
  BUF_X32 U53 ( .A(B[21]), .Z(SUM[21]) );
  BUF_X32 U54 ( .A(B[22]), .Z(SUM[22]) );
  BUF_X32 U55 ( .A(B[23]), .Z(SUM[23]) );
  BUF_X32 U56 ( .A(B[24]), .Z(SUM[24]) );
  BUF_X32 U57 ( .A(B[25]), .Z(SUM[25]) );
  BUF_X32 U58 ( .A(B[26]), .Z(SUM[26]) );
  BUF_X32 U59 ( .A(B[27]), .Z(SUM[27]) );
  BUF_X32 U60 ( .A(B[28]), .Z(SUM[28]) );
  BUF_X32 U61 ( .A(B[29]), .Z(SUM[29]) );
  BUF_X32 U62 ( .A(B[30]), .Z(SUM[30]) );
  BUF_X32 U63 ( .A(B[31]), .Z(SUM[31]) );
endmodule


module multiplier_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [31:1] carry;

  FA_X1 U2_31 ( .A(A[31]), .B(n2), .CI(carry[31]), .S(DIFF[31]) );
  FA_X1 U2_30 ( .A(A[30]), .B(n3), .CI(carry[30]), .CO(carry[31]), .S(DIFF[30]) );
  FA_X1 U2_29 ( .A(A[29]), .B(n4), .CI(carry[29]), .CO(carry[30]), .S(DIFF[29]) );
  FA_X1 U2_28 ( .A(A[28]), .B(n5), .CI(carry[28]), .CO(carry[29]), .S(DIFF[28]) );
  FA_X1 U2_27 ( .A(A[27]), .B(n6), .CI(carry[27]), .CO(carry[28]), .S(DIFF[27]) );
  FA_X1 U2_26 ( .A(A[26]), .B(n7), .CI(carry[26]), .CO(carry[27]), .S(DIFF[26]) );
  FA_X1 U2_25 ( .A(A[25]), .B(n8), .CI(carry[25]), .CO(carry[26]), .S(DIFF[25]) );
  FA_X1 U2_24 ( .A(A[24]), .B(n9), .CI(carry[24]), .CO(carry[25]), .S(DIFF[24]) );
  FA_X1 U2_23 ( .A(A[23]), .B(n10), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FA_X1 U2_22 ( .A(A[22]), .B(n11), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FA_X1 U2_21 ( .A(A[21]), .B(n12), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FA_X1 U2_20 ( .A(A[20]), .B(n13), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FA_X1 U2_19 ( .A(A[19]), .B(n14), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FA_X1 U2_18 ( .A(A[18]), .B(n15), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FA_X1 U2_17 ( .A(A[17]), .B(n16), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FA_X1 U2_16 ( .A(A[16]), .B(n17), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FA_X1 U2_15 ( .A(A[15]), .B(n18), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FA_X1 U2_14 ( .A(A[14]), .B(n19), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(n20), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(n21), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(n22), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FA_X1 U2_10 ( .A(A[10]), .B(n23), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n24), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FA_X1 U2_8 ( .A(A[8]), .B(n25), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FA_X1 U2_7 ( .A(A[7]), .B(n26), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n27), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n28), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n29), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n30), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n31), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n32), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  NAND2_X2 U1 ( .A1(B[0]), .A2(n1), .ZN(carry[1]) );
  XNOR2_X2 U2 ( .A(n33), .B(A[0]), .ZN(DIFF[0]) );
  INV_X4 U3 ( .A(A[0]), .ZN(n1) );
  INV_X4 U4 ( .A(B[31]), .ZN(n2) );
  INV_X4 U5 ( .A(B[30]), .ZN(n3) );
  INV_X4 U6 ( .A(B[29]), .ZN(n4) );
  INV_X4 U7 ( .A(B[28]), .ZN(n5) );
  INV_X4 U8 ( .A(B[27]), .ZN(n6) );
  INV_X4 U9 ( .A(B[26]), .ZN(n7) );
  INV_X4 U10 ( .A(B[25]), .ZN(n8) );
  INV_X4 U11 ( .A(B[24]), .ZN(n9) );
  INV_X4 U12 ( .A(B[23]), .ZN(n10) );
  INV_X4 U13 ( .A(B[22]), .ZN(n11) );
  INV_X4 U14 ( .A(B[21]), .ZN(n12) );
  INV_X4 U15 ( .A(B[20]), .ZN(n13) );
  INV_X4 U16 ( .A(B[19]), .ZN(n14) );
  INV_X4 U17 ( .A(B[18]), .ZN(n15) );
  INV_X4 U18 ( .A(B[17]), .ZN(n16) );
  INV_X4 U19 ( .A(B[16]), .ZN(n17) );
  INV_X4 U20 ( .A(B[15]), .ZN(n18) );
  INV_X4 U21 ( .A(B[14]), .ZN(n19) );
  INV_X4 U22 ( .A(B[13]), .ZN(n20) );
  INV_X4 U23 ( .A(B[12]), .ZN(n21) );
  INV_X4 U24 ( .A(B[11]), .ZN(n22) );
  INV_X4 U25 ( .A(B[10]), .ZN(n23) );
  INV_X4 U26 ( .A(B[9]), .ZN(n24) );
  INV_X4 U27 ( .A(B[8]), .ZN(n25) );
  INV_X4 U28 ( .A(B[7]), .ZN(n26) );
  INV_X4 U29 ( .A(B[6]), .ZN(n27) );
  INV_X4 U30 ( .A(B[5]), .ZN(n28) );
  INV_X4 U31 ( .A(B[4]), .ZN(n29) );
  INV_X4 U32 ( .A(B[3]), .ZN(n30) );
  INV_X4 U33 ( .A(B[2]), .ZN(n31) );
  INV_X4 U34 ( .A(B[1]), .ZN(n32) );
  INV_X4 U35 ( .A(B[0]), .ZN(n33) );
endmodule


module multiplier_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [31:1] carry;

  FA_X1 U2_31 ( .A(A[31]), .B(n2), .CI(carry[31]), .S(DIFF[31]) );
  FA_X1 U2_30 ( .A(A[30]), .B(n3), .CI(carry[30]), .CO(carry[31]), .S(DIFF[30]) );
  FA_X1 U2_29 ( .A(A[29]), .B(n4), .CI(carry[29]), .CO(carry[30]), .S(DIFF[29]) );
  FA_X1 U2_28 ( .A(A[28]), .B(n5), .CI(carry[28]), .CO(carry[29]), .S(DIFF[28]) );
  FA_X1 U2_27 ( .A(A[27]), .B(n6), .CI(carry[27]), .CO(carry[28]), .S(DIFF[27]) );
  FA_X1 U2_26 ( .A(A[26]), .B(n7), .CI(carry[26]), .CO(carry[27]), .S(DIFF[26]) );
  FA_X1 U2_25 ( .A(A[25]), .B(n8), .CI(carry[25]), .CO(carry[26]), .S(DIFF[25]) );
  FA_X1 U2_24 ( .A(A[24]), .B(n9), .CI(carry[24]), .CO(carry[25]), .S(DIFF[24]) );
  FA_X1 U2_23 ( .A(A[23]), .B(n10), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FA_X1 U2_22 ( .A(A[22]), .B(n11), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FA_X1 U2_21 ( .A(A[21]), .B(n12), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FA_X1 U2_20 ( .A(A[20]), .B(n13), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FA_X1 U2_19 ( .A(A[19]), .B(n14), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FA_X1 U2_18 ( .A(A[18]), .B(n15), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FA_X1 U2_17 ( .A(A[17]), .B(n16), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FA_X1 U2_16 ( .A(A[16]), .B(n17), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FA_X1 U2_15 ( .A(A[15]), .B(n18), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FA_X1 U2_14 ( .A(A[14]), .B(n19), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(n20), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(n21), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(n22), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FA_X1 U2_10 ( .A(A[10]), .B(n23), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n24), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FA_X1 U2_8 ( .A(A[8]), .B(n25), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FA_X1 U2_7 ( .A(A[7]), .B(n26), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n27), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n28), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n29), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n30), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n31), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n32), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  NAND2_X2 U1 ( .A1(B[0]), .A2(n1), .ZN(carry[1]) );
  XNOR2_X2 U2 ( .A(n33), .B(A[0]), .ZN(DIFF[0]) );
  INV_X4 U3 ( .A(A[0]), .ZN(n1) );
  INV_X4 U4 ( .A(B[31]), .ZN(n2) );
  INV_X4 U5 ( .A(B[30]), .ZN(n3) );
  INV_X4 U6 ( .A(B[29]), .ZN(n4) );
  INV_X4 U7 ( .A(B[28]), .ZN(n5) );
  INV_X4 U8 ( .A(B[27]), .ZN(n6) );
  INV_X4 U9 ( .A(B[26]), .ZN(n7) );
  INV_X4 U10 ( .A(B[25]), .ZN(n8) );
  INV_X4 U11 ( .A(B[24]), .ZN(n9) );
  INV_X4 U12 ( .A(B[23]), .ZN(n10) );
  INV_X4 U13 ( .A(B[22]), .ZN(n11) );
  INV_X4 U14 ( .A(B[21]), .ZN(n12) );
  INV_X4 U15 ( .A(B[20]), .ZN(n13) );
  INV_X4 U16 ( .A(B[19]), .ZN(n14) );
  INV_X4 U17 ( .A(B[18]), .ZN(n15) );
  INV_X4 U18 ( .A(B[17]), .ZN(n16) );
  INV_X4 U19 ( .A(B[16]), .ZN(n17) );
  INV_X4 U20 ( .A(B[15]), .ZN(n18) );
  INV_X4 U21 ( .A(B[14]), .ZN(n19) );
  INV_X4 U22 ( .A(B[13]), .ZN(n20) );
  INV_X4 U23 ( .A(B[12]), .ZN(n21) );
  INV_X4 U24 ( .A(B[11]), .ZN(n22) );
  INV_X4 U25 ( .A(B[10]), .ZN(n23) );
  INV_X4 U26 ( .A(B[9]), .ZN(n24) );
  INV_X4 U27 ( .A(B[8]), .ZN(n25) );
  INV_X4 U28 ( .A(B[7]), .ZN(n26) );
  INV_X4 U29 ( .A(B[6]), .ZN(n27) );
  INV_X4 U30 ( .A(B[5]), .ZN(n28) );
  INV_X4 U31 ( .A(B[4]), .ZN(n29) );
  INV_X4 U32 ( .A(B[3]), .ZN(n30) );
  INV_X4 U33 ( .A(B[2]), .ZN(n31) );
  INV_X4 U34 ( .A(B[1]), .ZN(n32) );
  INV_X4 U35 ( .A(B[0]), .ZN(n33) );
endmodule


module multiplier_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   \ab[16][15] , \ab[16][14] , \ab[16][13] , \ab[16][12] , \ab[16][11] ,
         \ab[16][10] , \ab[16][9] , \ab[16][8] , \ab[16][7] , \ab[16][6] ,
         \ab[16][5] , \ab[16][4] , \ab[16][3] , \ab[16][2] , \ab[16][1] ,
         \ab[16][0] , \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] ,
         \ab[15][11] , \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] ,
         \ab[15][6] , \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] ,
         \ab[15][1] , \ab[15][0] , \ab[14][15] , \ab[14][14] , \ab[14][13] ,
         \ab[14][12] , \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] ,
         \ab[14][7] , \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] ,
         \ab[14][2] , \ab[14][1] , \ab[14][0] , \ab[13][15] , \ab[13][14] ,
         \ab[13][13] , \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] ,
         \ab[13][8] , \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] ,
         \ab[13][3] , \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][15] ,
         \ab[12][14] , \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] ,
         \ab[12][9] , \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] ,
         \ab[12][4] , \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] ,
         \ab[11][15] , \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] ,
         \ab[11][10] , \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] ,
         \ab[11][5] , \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] ,
         \ab[11][0] , \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] ,
         \ab[10][11] , \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] ,
         \ab[10][6] , \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] ,
         \ab[10][1] , \ab[10][0] , \ab[9][15] , \ab[9][14] , \ab[9][13] ,
         \ab[9][12] , \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] ,
         \ab[9][7] , \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] ,
         \ab[9][2] , \ab[9][1] , \ab[9][0] , \ab[8][15] , \ab[8][14] ,
         \ab[8][13] , \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] ,
         \ab[8][8] , \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] ,
         \ab[8][3] , \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][15] ,
         \ab[7][14] , \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] ,
         \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] ,
         \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] ,
         \ab[6][15] , \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] ,
         \ab[6][10] , \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] ,
         \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] ,
         \ab[6][0] , \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] ,
         \ab[5][11] , \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] ,
         \ab[5][6] , \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] ,
         \ab[5][1] , \ab[5][0] , \ab[4][15] , \ab[4][14] , \ab[4][13] ,
         \ab[4][12] , \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] ,
         \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] ,
         \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][15] , \ab[3][14] ,
         \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] ,
         \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] ,
         \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][15] ,
         \ab[2][14] , \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] ,
         \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] ,
         \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] ,
         \ab[1][16] , \ab[1][15] , \ab[1][14] , \ab[1][13] , \ab[1][12] ,
         \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][8] , \ab[1][7] ,
         \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] ,
         \ab[1][1] , \ab[1][0] , \ab[0][16] , \ab[0][15] , \ab[0][14] ,
         \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] ,
         \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] ,
         \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[15][15] ,
         \CARRYB[15][14] , \CARRYB[15][13] , \CARRYB[15][12] ,
         \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] ,
         \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] ,
         \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] ,
         \CARRYB[14][15] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \CARRYB[13][15] , \CARRYB[13][14] , \CARRYB[13][13] ,
         \CARRYB[13][12] , \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] ,
         \CARRYB[13][8] , \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] ,
         \CARRYB[13][0] , \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][15] , \CARRYB[10][14] , \CARRYB[10][13] ,
         \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] ,
         \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] ,
         \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] ,
         \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] ,
         \CARRYB[9][0] , \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] ,
         \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] ,
         \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] ,
         \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] ,
         \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] ,
         \CARRYB[5][0] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][13] ,
         \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] ,
         \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[15][16] , \SUMB[15][15] , \SUMB[15][14] ,
         \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] , \SUMB[15][10] ,
         \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] , \SUMB[15][6] ,
         \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] , \SUMB[15][2] ,
         \SUMB[15][1] , \SUMB[14][16] , \SUMB[14][15] , \SUMB[14][14] ,
         \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] ,
         \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] ,
         \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] ,
         \SUMB[14][1] , \SUMB[13][16] , \SUMB[13][15] , \SUMB[13][14] ,
         \SUMB[13][13] , \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] ,
         \SUMB[13][9] , \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][6] ,
         \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] ,
         \SUMB[13][1] , \SUMB[12][16] , \SUMB[12][15] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][16] , \SUMB[11][15] , \SUMB[11][14] ,
         \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] , \SUMB[11][10] ,
         \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] , \SUMB[11][6] ,
         \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] , \SUMB[11][2] ,
         \SUMB[11][1] , \SUMB[10][16] , \SUMB[10][15] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][16] , \SUMB[9][15] , \SUMB[9][14] ,
         \SUMB[9][13] , \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] ,
         \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] ,
         \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][16] ,
         \SUMB[8][15] , \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] ,
         \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] ,
         \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] ,
         \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][16] , \SUMB[7][15] ,
         \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] , \SUMB[6][13] ,
         \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] , \SUMB[6][9] ,
         \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] ,
         \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][16] ,
         \SUMB[5][15] , \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] ,
         \SUMB[5][11] , \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] ,
         \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] ,
         \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][16] , \SUMB[4][15] ,
         \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] ,
         \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] , \SUMB[3][13] ,
         \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] , \SUMB[3][9] ,
         \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] ,
         \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][16] ,
         \SUMB[2][15] , \SUMB[2][14] , \SUMB[2][13] , \SUMB[2][12] ,
         \SUMB[2][11] , \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] ,
         \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , \CARRYB[30][0] , \CARRYB[29][1] ,
         \CARRYB[29][0] , \CARRYB[28][2] , \CARRYB[28][1] , \CARRYB[28][0] ,
         \CARRYB[27][3] , \CARRYB[27][2] , \CARRYB[27][1] , \CARRYB[27][0] ,
         \CARRYB[26][4] , \CARRYB[26][3] , \CARRYB[26][2] , \CARRYB[26][1] ,
         \CARRYB[26][0] , \CARRYB[25][5] , \CARRYB[25][4] , \CARRYB[25][3] ,
         \CARRYB[25][2] , \CARRYB[25][1] , \CARRYB[25][0] , \CARRYB[24][6] ,
         \CARRYB[24][5] , \CARRYB[24][4] , \CARRYB[24][3] , \CARRYB[24][2] ,
         \CARRYB[24][1] , \CARRYB[24][0] , \CARRYB[23][7] , \CARRYB[23][6] ,
         \CARRYB[23][5] , \CARRYB[23][4] , \CARRYB[23][3] , \CARRYB[23][2] ,
         \CARRYB[23][1] , \CARRYB[23][0] , \CARRYB[22][8] , \CARRYB[22][7] ,
         \CARRYB[22][6] , \CARRYB[22][5] , \CARRYB[22][4] , \CARRYB[22][3] ,
         \CARRYB[22][2] , \CARRYB[22][1] , \CARRYB[22][0] , \CARRYB[21][9] ,
         \CARRYB[21][8] , \CARRYB[21][7] , \CARRYB[21][6] , \CARRYB[21][5] ,
         \CARRYB[21][4] , \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] ,
         \CARRYB[21][0] , \CARRYB[20][10] , \CARRYB[20][9] , \CARRYB[20][8] ,
         \CARRYB[20][7] , \CARRYB[20][6] , \CARRYB[20][5] , \CARRYB[20][4] ,
         \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] , \CARRYB[20][0] ,
         \CARRYB[19][11] , \CARRYB[19][10] , \CARRYB[19][9] , \CARRYB[19][8] ,
         \CARRYB[19][7] , \CARRYB[19][6] , \CARRYB[19][5] , \CARRYB[19][4] ,
         \CARRYB[19][3] , \CARRYB[19][2] , \CARRYB[19][1] , \CARRYB[19][0] ,
         \CARRYB[18][12] , \CARRYB[18][11] , \CARRYB[18][10] , \CARRYB[18][9] ,
         \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][6] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] ,
         \CARRYB[18][0] , \CARRYB[17][13] , \CARRYB[17][12] , \CARRYB[17][11] ,
         \CARRYB[17][10] , \CARRYB[17][9] , \CARRYB[17][8] , \CARRYB[17][7] ,
         \CARRYB[17][6] , \CARRYB[17][5] , \CARRYB[17][4] , \CARRYB[17][3] ,
         \CARRYB[17][2] , \CARRYB[17][1] , \CARRYB[17][0] , \CARRYB[16][14] ,
         \CARRYB[16][13] , \CARRYB[16][12] , \CARRYB[16][11] ,
         \CARRYB[16][10] , \CARRYB[16][9] , \CARRYB[16][8] , \CARRYB[16][7] ,
         \CARRYB[16][6] , \CARRYB[16][5] , \CARRYB[16][4] , \CARRYB[16][3] ,
         \CARRYB[16][2] , \CARRYB[16][1] , \CARRYB[16][0] , \SUMB[30][1] ,
         \SUMB[29][2] , \SUMB[29][1] , \SUMB[28][3] , \SUMB[28][2] ,
         \SUMB[28][1] , \SUMB[27][4] , \SUMB[27][3] , \SUMB[27][2] ,
         \SUMB[27][1] , \SUMB[26][5] , \SUMB[26][4] , \SUMB[26][3] ,
         \SUMB[26][2] , \SUMB[26][1] , \SUMB[25][6] , \SUMB[25][5] ,
         \SUMB[25][4] , \SUMB[25][3] , \SUMB[25][2] , \SUMB[25][1] ,
         \SUMB[24][7] , \SUMB[24][6] , \SUMB[24][5] , \SUMB[24][4] ,
         \SUMB[24][3] , \SUMB[24][2] , \SUMB[24][1] , \SUMB[23][8] ,
         \SUMB[23][7] , \SUMB[23][6] , \SUMB[23][5] , \SUMB[23][4] ,
         \SUMB[23][3] , \SUMB[23][2] , \SUMB[23][1] , \SUMB[22][9] ,
         \SUMB[22][8] , \SUMB[22][7] , \SUMB[22][6] , \SUMB[22][5] ,
         \SUMB[22][4] , \SUMB[22][3] , \SUMB[22][2] , \SUMB[22][1] ,
         \SUMB[21][10] , \SUMB[21][9] , \SUMB[21][8] , \SUMB[21][7] ,
         \SUMB[21][6] , \SUMB[21][5] , \SUMB[21][4] , \SUMB[21][3] ,
         \SUMB[21][2] , \SUMB[21][1] , \SUMB[20][11] , \SUMB[20][10] ,
         \SUMB[20][9] , \SUMB[20][8] , \SUMB[20][7] , \SUMB[20][6] ,
         \SUMB[20][5] , \SUMB[20][4] , \SUMB[20][3] , \SUMB[20][2] ,
         \SUMB[20][1] , \SUMB[19][12] , \SUMB[19][11] , \SUMB[19][10] ,
         \SUMB[19][9] , \SUMB[19][8] , \SUMB[19][7] , \SUMB[19][6] ,
         \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] , \SUMB[19][2] ,
         \SUMB[19][1] , \SUMB[18][13] , \SUMB[18][12] , \SUMB[18][11] ,
         \SUMB[18][10] , \SUMB[18][9] , \SUMB[18][8] , \SUMB[18][7] ,
         \SUMB[18][6] , \SUMB[18][5] , \SUMB[18][4] , \SUMB[18][3] ,
         \SUMB[18][2] , \SUMB[18][1] , \SUMB[17][14] , \SUMB[17][13] ,
         \SUMB[17][12] , \SUMB[17][11] , \SUMB[17][10] , \SUMB[17][9] ,
         \SUMB[17][8] , \SUMB[17][7] , \SUMB[17][6] , \SUMB[17][5] ,
         \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] , \SUMB[17][1] ,
         \SUMB[16][15] , \SUMB[16][14] , \SUMB[16][13] , \SUMB[16][12] ,
         \SUMB[16][11] , \SUMB[16][10] , \SUMB[16][9] , \SUMB[16][8] ,
         \SUMB[16][7] , \SUMB[16][6] , \SUMB[16][5] , \SUMB[16][4] ,
         \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] , n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299;

  FA_X1 S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(PRODUCT[16]) );
  FA_X1 S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA_X1 S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), 
        .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA_X1 S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), 
        .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA_X1 S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA_X1 S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), 
        .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA_X1 S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), 
        .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA_X1 S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA_X1 S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA_X1 S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA_X1 S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), 
        .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA_X1 S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(\SUMB[15][12] ), 
        .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FA_X1 S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), 
        .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FA_X1 S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(\SUMB[15][14] ), 
        .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FA_X1 S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(\SUMB[15][15] ), 
        .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FA_X1 S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), 
        .S(\SUMB[16][15] ) );
  FA_X1 S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), 
        .CO(\CARRYB[15][0] ), .S(PRODUCT[15]) );
  FA_X1 S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), 
        .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA_X1 S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), 
        .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA_X1 S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), 
        .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA_X1 S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA_X1 S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA_X1 S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), 
        .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA_X1 S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), 
        .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA_X1 S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), 
        .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA_X1 S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA_X1 S2_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA_X1 S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA_X1 S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA_X1 S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA_X1 S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA_X1 S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), 
        .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FA_X1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(PRODUCT[14]) );
  FA_X1 S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA_X1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA_X1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA_X1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA_X1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA_X1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA_X1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA_X1 S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA_X1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA_X1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA_X1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA_X1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA_X1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA_X1 S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA_X1 S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\SUMB[13][16] ), 
        .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA_X1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(PRODUCT[13]) );
  FA_X1 S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA_X1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA_X1 S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA_X1 S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA_X1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA_X1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA_X1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA_X1 S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA_X1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA_X1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA_X1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA_X1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA_X1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA_X1 S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA_X1 S2_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\SUMB[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA_X1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(PRODUCT[12]) );
  FA_X1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA_X1 S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA_X1 S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA_X1 S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA_X1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA_X1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA_X1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA_X1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA_X1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA_X1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA_X1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA_X1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA_X1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA_X1 S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA_X1 S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\SUMB[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA_X1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(PRODUCT[11]) );
  FA_X1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA_X1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA_X1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA_X1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA_X1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA_X1 S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA_X1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA_X1 S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA_X1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA_X1 S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA_X1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA_X1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA_X1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA_X1 S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA_X1 S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA_X1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(PRODUCT[10]) );
  FA_X1 S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA_X1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA_X1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA_X1 S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA_X1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA_X1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA_X1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA_X1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA_X1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA_X1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA_X1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA_X1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA_X1 S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA_X1 S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA_X1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(PRODUCT[9]) );
  FA_X1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA_X1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA_X1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA_X1 S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA_X1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA_X1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA_X1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA_X1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA_X1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA_X1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA_X1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA_X1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA_X1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA_X1 S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA_X1 S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), 
        .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA_X1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(PRODUCT[8]) );
  FA_X1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA_X1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA_X1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA_X1 S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA_X1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA_X1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA_X1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA_X1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA_X1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA_X1 S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA_X1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA_X1 S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA_X1 S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA_X1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(PRODUCT[7]) );
  FA_X1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA_X1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA_X1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA_X1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA_X1 S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA_X1 S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA_X1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA_X1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA_X1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA_X1 S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA_X1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA_X1 S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA_X1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA_X1 S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA_X1 S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA_X1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(PRODUCT[6]) );
  FA_X1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA_X1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA_X1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA_X1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA_X1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA_X1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA_X1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA_X1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA_X1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA_X1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA_X1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA_X1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA_X1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA_X1 S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA_X1 S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA_X1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(PRODUCT[5]) );
  FA_X1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA_X1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA_X1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA_X1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA_X1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA_X1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA_X1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA_X1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA_X1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA_X1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA_X1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA_X1 S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA_X1 S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA_X1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(PRODUCT[4]) );
  FA_X1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA_X1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA_X1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA_X1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA_X1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA_X1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA_X1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA_X1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA_X1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA_X1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA_X1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA_X1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA_X1 S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA_X1 S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA_X1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(PRODUCT[3]) );
  FA_X1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA_X1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA_X1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA_X1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA_X1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA_X1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA_X1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA_X1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA_X1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA_X1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA_X1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA_X1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA_X1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA_X1 S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA_X1 S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), 
        .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(n33), .CI(n48), .CO(\CARRYB[2][0] ), .S(
        PRODUCT[2]) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(n32), .CI(n47), .CO(\CARRYB[2][1] ), .S(
        \SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(n31), .CI(n46), .CO(\CARRYB[2][2] ), .S(
        \SUMB[2][2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2][3] ), .B(n30), .CI(n45), .CO(\CARRYB[2][3] ), .S(
        \SUMB[2][3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2][4] ), .B(n29), .CI(n44), .CO(\CARRYB[2][4] ), .S(
        \SUMB[2][4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2][5] ), .B(n28), .CI(n43), .CO(\CARRYB[2][5] ), .S(
        \SUMB[2][5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2][6] ), .B(n27), .CI(n42), .CO(\CARRYB[2][6] ), .S(
        \SUMB[2][6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(n26), .CI(n41), .CO(\CARRYB[2][7] ), .S(
        \SUMB[2][7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(n25), .CI(n40), .CO(\CARRYB[2][8] ), .S(
        \SUMB[2][8] ) );
  FA_X1 S2_2_9 ( .A(\ab[2][9] ), .B(n24), .CI(n39), .CO(\CARRYB[2][9] ), .S(
        \SUMB[2][9] ) );
  FA_X1 S2_2_10 ( .A(\ab[2][10] ), .B(n23), .CI(n38), .CO(\CARRYB[2][10] ), 
        .S(\SUMB[2][10] ) );
  FA_X1 S2_2_11 ( .A(\ab[2][11] ), .B(n22), .CI(n37), .CO(\CARRYB[2][11] ), 
        .S(\SUMB[2][11] ) );
  FA_X1 S2_2_12 ( .A(\ab[2][12] ), .B(n21), .CI(n36), .CO(\CARRYB[2][12] ), 
        .S(\SUMB[2][12] ) );
  FA_X1 S2_2_13 ( .A(\ab[2][13] ), .B(n20), .CI(n35), .CO(\CARRYB[2][13] ), 
        .S(\SUMB[2][13] ) );
  FA_X1 S2_2_14 ( .A(\ab[2][14] ), .B(n19), .CI(n34), .CO(\CARRYB[2][14] ), 
        .S(\SUMB[2][14] ) );
  FA_X1 S2_2_15 ( .A(\ab[2][15] ), .B(n18), .CI(\ab[1][16] ), .CO(
        \CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  XNOR2_X2 U2 ( .A(\CARRYB[30][0] ), .B(\SUMB[30][1] ), .ZN(n3) );
  INV_X4 U3 ( .A(n3), .ZN(PRODUCT[31]) );
  XNOR2_X2 U4 ( .A(\CARRYB[20][10] ), .B(\SUMB[20][11] ), .ZN(n4) );
  INV_X4 U5 ( .A(n4), .ZN(\SUMB[21][10] ) );
  XNOR2_X2 U6 ( .A(\CARRYB[19][11] ), .B(\SUMB[19][12] ), .ZN(n5) );
  INV_X4 U7 ( .A(n5), .ZN(\SUMB[20][11] ) );
  XNOR2_X2 U8 ( .A(\CARRYB[18][12] ), .B(\SUMB[18][13] ), .ZN(n6) );
  INV_X4 U9 ( .A(n6), .ZN(\SUMB[19][12] ) );
  XNOR2_X2 U10 ( .A(\CARRYB[17][13] ), .B(\SUMB[17][14] ), .ZN(n7) );
  INV_X4 U11 ( .A(n7), .ZN(\SUMB[18][13] ) );
  XNOR2_X2 U12 ( .A(\CARRYB[16][14] ), .B(\SUMB[16][15] ), .ZN(n8) );
  INV_X4 U13 ( .A(n8), .ZN(\SUMB[17][14] ) );
  XNOR2_X2 U14 ( .A(\CARRYB[29][1] ), .B(\SUMB[29][2] ), .ZN(n9) );
  INV_X4 U15 ( .A(n9), .ZN(\SUMB[30][1] ) );
  XNOR2_X2 U16 ( .A(\CARRYB[28][2] ), .B(\SUMB[28][3] ), .ZN(n10) );
  INV_X4 U17 ( .A(n10), .ZN(\SUMB[29][2] ) );
  XNOR2_X2 U18 ( .A(\CARRYB[27][3] ), .B(\SUMB[27][4] ), .ZN(n11) );
  INV_X4 U19 ( .A(n11), .ZN(\SUMB[28][3] ) );
  XNOR2_X2 U20 ( .A(\CARRYB[26][4] ), .B(\SUMB[26][5] ), .ZN(n12) );
  INV_X4 U21 ( .A(n12), .ZN(\SUMB[27][4] ) );
  XNOR2_X2 U22 ( .A(\CARRYB[25][5] ), .B(\SUMB[25][6] ), .ZN(n13) );
  INV_X4 U23 ( .A(n13), .ZN(\SUMB[26][5] ) );
  XNOR2_X2 U24 ( .A(\CARRYB[24][6] ), .B(\SUMB[24][7] ), .ZN(n14) );
  INV_X4 U25 ( .A(n14), .ZN(\SUMB[25][6] ) );
  XNOR2_X2 U26 ( .A(\CARRYB[23][7] ), .B(\SUMB[23][8] ), .ZN(n15) );
  INV_X4 U27 ( .A(n15), .ZN(\SUMB[24][7] ) );
  XNOR2_X2 U28 ( .A(\CARRYB[22][8] ), .B(\SUMB[22][9] ), .ZN(n16) );
  INV_X4 U29 ( .A(n16), .ZN(\SUMB[23][8] ) );
  XNOR2_X2 U30 ( .A(\CARRYB[21][9] ), .B(\SUMB[21][10] ), .ZN(n17) );
  INV_X4 U31 ( .A(n17), .ZN(\SUMB[22][9] ) );
  AND2_X4 U32 ( .A1(\ab[0][16] ), .A2(\ab[1][15] ), .ZN(n18) );
  AND2_X4 U33 ( .A1(\ab[0][15] ), .A2(\ab[1][14] ), .ZN(n19) );
  AND2_X4 U34 ( .A1(\ab[0][14] ), .A2(\ab[1][13] ), .ZN(n20) );
  AND2_X4 U35 ( .A1(\ab[0][13] ), .A2(\ab[1][12] ), .ZN(n21) );
  AND2_X4 U36 ( .A1(\ab[0][12] ), .A2(\ab[1][11] ), .ZN(n22) );
  AND2_X4 U37 ( .A1(\ab[0][11] ), .A2(\ab[1][10] ), .ZN(n23) );
  AND2_X4 U38 ( .A1(\ab[0][10] ), .A2(\ab[1][9] ), .ZN(n24) );
  AND2_X4 U39 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .ZN(n25) );
  AND2_X4 U40 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .ZN(n26) );
  AND2_X4 U41 ( .A1(\ab[0][7] ), .A2(\ab[1][6] ), .ZN(n27) );
  AND2_X4 U42 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .ZN(n28) );
  AND2_X4 U43 ( .A1(\ab[0][5] ), .A2(\ab[1][4] ), .ZN(n29) );
  AND2_X4 U44 ( .A1(\ab[0][4] ), .A2(\ab[1][3] ), .ZN(n30) );
  AND2_X4 U45 ( .A1(\ab[0][3] ), .A2(\ab[1][2] ), .ZN(n31) );
  AND2_X4 U46 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .ZN(n32) );
  AND2_X4 U47 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .ZN(n33) );
  XOR2_X2 U48 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(n34) );
  XOR2_X2 U49 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(n35) );
  XOR2_X2 U50 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(n36) );
  XOR2_X2 U51 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(n37) );
  XOR2_X2 U52 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(n38) );
  XOR2_X2 U53 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(n39) );
  XOR2_X2 U54 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(n40) );
  XOR2_X2 U55 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(n41) );
  XOR2_X2 U56 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(n42) );
  XOR2_X2 U57 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(n43) );
  XOR2_X2 U58 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(n44) );
  XOR2_X2 U59 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(n45) );
  XOR2_X2 U60 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(n46) );
  XOR2_X2 U61 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(n47) );
  XOR2_X2 U62 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(n48) );
  XOR2_X2 U63 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  AND2_X2 U64 ( .A1(B[1]), .A2(A[1]), .ZN(\ab[1][1] ) );
  INV_X4 U65 ( .A(B[3]), .ZN(n50) );
  INV_X4 U66 ( .A(B[0]), .ZN(n54) );
  INV_X4 U67 ( .A(B[1]), .ZN(n53) );
  INV_X4 U68 ( .A(B[2]), .ZN(n52) );
  INV_X4 U69 ( .A(A[0]), .ZN(n59) );
  INV_X4 U70 ( .A(A[1]), .ZN(n58) );
  INV_X4 U71 ( .A(A[2]), .ZN(n57) );
  INV_X4 U72 ( .A(A[3]), .ZN(n55) );
  INV_X4 U73 ( .A(B[3]), .ZN(n51) );
  INV_X4 U74 ( .A(A[3]), .ZN(n56) );
  INV_X4 U75 ( .A(B[11]), .ZN(n65) );
  INV_X4 U76 ( .A(B[12]), .ZN(n64) );
  INV_X4 U77 ( .A(B[13]), .ZN(n63) );
  INV_X4 U78 ( .A(B[14]), .ZN(n62) );
  INV_X4 U79 ( .A(B[15]), .ZN(n61) );
  INV_X4 U80 ( .A(A[10]), .ZN(n81) );
  INV_X4 U81 ( .A(A[11]), .ZN(n80) );
  INV_X4 U82 ( .A(A[12]), .ZN(n79) );
  INV_X4 U83 ( .A(A[13]), .ZN(n78) );
  INV_X4 U84 ( .A(A[14]), .ZN(n77) );
  INV_X4 U85 ( .A(A[15]), .ZN(n76) );
  INV_X4 U86 ( .A(B[16]), .ZN(n60) );
  INV_X4 U87 ( .A(A[16]), .ZN(n75) );
  INV_X4 U88 ( .A(A[9]), .ZN(n82) );
  INV_X4 U89 ( .A(B[4]), .ZN(n72) );
  INV_X4 U90 ( .A(B[5]), .ZN(n71) );
  INV_X4 U91 ( .A(B[6]), .ZN(n70) );
  INV_X4 U92 ( .A(B[7]), .ZN(n69) );
  INV_X4 U93 ( .A(B[8]), .ZN(n68) );
  INV_X4 U94 ( .A(B[9]), .ZN(n67) );
  INV_X4 U95 ( .A(B[10]), .ZN(n66) );
  INV_X4 U96 ( .A(A[4]), .ZN(n87) );
  INV_X4 U97 ( .A(A[5]), .ZN(n86) );
  INV_X4 U98 ( .A(A[6]), .ZN(n85) );
  INV_X4 U99 ( .A(A[7]), .ZN(n84) );
  INV_X4 U100 ( .A(A[8]), .ZN(n83) );
  INV_X4 U206 ( .A(B[2]), .ZN(n73) );
  INV_X4 U207 ( .A(B[0]), .ZN(n74) );
  INV_X4 U208 ( .A(A[2]), .ZN(n88) );
  INV_X4 U209 ( .A(A[0]), .ZN(n89) );
  NOR2_X1 U210 ( .A1(n82), .A2(n67), .ZN(\ab[9][9] ) );
  NOR2_X1 U211 ( .A1(n82), .A2(n68), .ZN(\ab[9][8] ) );
  NOR2_X1 U212 ( .A1(n82), .A2(n69), .ZN(\ab[9][7] ) );
  NOR2_X1 U213 ( .A1(n82), .A2(n70), .ZN(\ab[9][6] ) );
  NOR2_X1 U214 ( .A1(n82), .A2(n71), .ZN(\ab[9][5] ) );
  NOR2_X1 U215 ( .A1(n82), .A2(n72), .ZN(\ab[9][4] ) );
  NOR2_X1 U216 ( .A1(n82), .A2(n51), .ZN(\ab[9][3] ) );
  NOR2_X1 U217 ( .A1(n82), .A2(n52), .ZN(\ab[9][2] ) );
  NOR2_X1 U218 ( .A1(n82), .A2(n53), .ZN(\ab[9][1] ) );
  NOR2_X1 U219 ( .A1(n82), .A2(n60), .ZN(\SUMB[9][16] ) );
  NOR2_X1 U220 ( .A1(n82), .A2(n61), .ZN(\ab[9][15] ) );
  NOR2_X1 U221 ( .A1(n82), .A2(n62), .ZN(\ab[9][14] ) );
  NOR2_X1 U222 ( .A1(n82), .A2(n63), .ZN(\ab[9][13] ) );
  NOR2_X1 U223 ( .A1(n82), .A2(n64), .ZN(\ab[9][12] ) );
  NOR2_X1 U224 ( .A1(n82), .A2(n65), .ZN(\ab[9][11] ) );
  NOR2_X1 U225 ( .A1(n82), .A2(n66), .ZN(\ab[9][10] ) );
  NOR2_X1 U226 ( .A1(n82), .A2(n54), .ZN(\ab[9][0] ) );
  NOR2_X1 U227 ( .A1(n67), .A2(n83), .ZN(\ab[8][9] ) );
  NOR2_X1 U228 ( .A1(n68), .A2(n83), .ZN(\ab[8][8] ) );
  NOR2_X1 U229 ( .A1(n69), .A2(n83), .ZN(\ab[8][7] ) );
  NOR2_X1 U230 ( .A1(n70), .A2(n83), .ZN(\ab[8][6] ) );
  NOR2_X1 U231 ( .A1(n71), .A2(n83), .ZN(\ab[8][5] ) );
  NOR2_X1 U232 ( .A1(n72), .A2(n83), .ZN(\ab[8][4] ) );
  NOR2_X1 U233 ( .A1(n51), .A2(n83), .ZN(\ab[8][3] ) );
  NOR2_X1 U234 ( .A1(n52), .A2(n83), .ZN(\ab[8][2] ) );
  NOR2_X1 U235 ( .A1(n53), .A2(n83), .ZN(\ab[8][1] ) );
  NOR2_X1 U236 ( .A1(n60), .A2(n83), .ZN(\SUMB[8][16] ) );
  NOR2_X1 U237 ( .A1(n61), .A2(n83), .ZN(\ab[8][15] ) );
  NOR2_X1 U238 ( .A1(n62), .A2(n83), .ZN(\ab[8][14] ) );
  NOR2_X1 U239 ( .A1(n63), .A2(n83), .ZN(\ab[8][13] ) );
  NOR2_X1 U240 ( .A1(n64), .A2(n83), .ZN(\ab[8][12] ) );
  NOR2_X1 U241 ( .A1(n65), .A2(n83), .ZN(\ab[8][11] ) );
  NOR2_X1 U242 ( .A1(n66), .A2(n83), .ZN(\ab[8][10] ) );
  NOR2_X1 U243 ( .A1(n74), .A2(n83), .ZN(\ab[8][0] ) );
  NOR2_X1 U244 ( .A1(n67), .A2(n84), .ZN(\ab[7][9] ) );
  NOR2_X1 U245 ( .A1(n68), .A2(n84), .ZN(\ab[7][8] ) );
  NOR2_X1 U246 ( .A1(n69), .A2(n84), .ZN(\ab[7][7] ) );
  NOR2_X1 U247 ( .A1(n70), .A2(n84), .ZN(\ab[7][6] ) );
  NOR2_X1 U248 ( .A1(n71), .A2(n84), .ZN(\ab[7][5] ) );
  NOR2_X1 U249 ( .A1(n72), .A2(n84), .ZN(\ab[7][4] ) );
  NOR2_X1 U250 ( .A1(n51), .A2(n84), .ZN(\ab[7][3] ) );
  NOR2_X1 U251 ( .A1(n52), .A2(n84), .ZN(\ab[7][2] ) );
  NOR2_X1 U252 ( .A1(n53), .A2(n84), .ZN(\ab[7][1] ) );
  NOR2_X1 U253 ( .A1(n60), .A2(n84), .ZN(\SUMB[7][16] ) );
  NOR2_X1 U254 ( .A1(n61), .A2(n84), .ZN(\ab[7][15] ) );
  NOR2_X1 U255 ( .A1(n62), .A2(n84), .ZN(\ab[7][14] ) );
  NOR2_X1 U256 ( .A1(n63), .A2(n84), .ZN(\ab[7][13] ) );
  NOR2_X1 U257 ( .A1(n64), .A2(n84), .ZN(\ab[7][12] ) );
  NOR2_X1 U258 ( .A1(n65), .A2(n84), .ZN(\ab[7][11] ) );
  NOR2_X1 U259 ( .A1(n66), .A2(n84), .ZN(\ab[7][10] ) );
  NOR2_X1 U260 ( .A1(n74), .A2(n84), .ZN(\ab[7][0] ) );
  NOR2_X1 U261 ( .A1(n67), .A2(n85), .ZN(\ab[6][9] ) );
  NOR2_X1 U262 ( .A1(n68), .A2(n85), .ZN(\ab[6][8] ) );
  NOR2_X1 U263 ( .A1(n69), .A2(n85), .ZN(\ab[6][7] ) );
  NOR2_X1 U264 ( .A1(n70), .A2(n85), .ZN(\ab[6][6] ) );
  NOR2_X1 U265 ( .A1(n71), .A2(n85), .ZN(\ab[6][5] ) );
  NOR2_X1 U266 ( .A1(n72), .A2(n85), .ZN(\ab[6][4] ) );
  NOR2_X1 U267 ( .A1(n51), .A2(n85), .ZN(\ab[6][3] ) );
  NOR2_X1 U268 ( .A1(n52), .A2(n85), .ZN(\ab[6][2] ) );
  NOR2_X1 U269 ( .A1(n53), .A2(n85), .ZN(\ab[6][1] ) );
  NOR2_X1 U270 ( .A1(n60), .A2(n85), .ZN(\SUMB[6][16] ) );
  NOR2_X1 U271 ( .A1(n61), .A2(n85), .ZN(\ab[6][15] ) );
  NOR2_X1 U272 ( .A1(n62), .A2(n85), .ZN(\ab[6][14] ) );
  NOR2_X1 U273 ( .A1(n63), .A2(n85), .ZN(\ab[6][13] ) );
  NOR2_X1 U274 ( .A1(n64), .A2(n85), .ZN(\ab[6][12] ) );
  NOR2_X1 U275 ( .A1(n65), .A2(n85), .ZN(\ab[6][11] ) );
  NOR2_X1 U276 ( .A1(n66), .A2(n85), .ZN(\ab[6][10] ) );
  NOR2_X1 U277 ( .A1(n74), .A2(n85), .ZN(\ab[6][0] ) );
  NOR2_X1 U278 ( .A1(n67), .A2(n86), .ZN(\ab[5][9] ) );
  NOR2_X1 U279 ( .A1(n68), .A2(n86), .ZN(\ab[5][8] ) );
  NOR2_X1 U280 ( .A1(n69), .A2(n86), .ZN(\ab[5][7] ) );
  NOR2_X1 U281 ( .A1(n70), .A2(n86), .ZN(\ab[5][6] ) );
  NOR2_X1 U282 ( .A1(n71), .A2(n86), .ZN(\ab[5][5] ) );
  NOR2_X1 U283 ( .A1(n72), .A2(n86), .ZN(\ab[5][4] ) );
  NOR2_X1 U284 ( .A1(n51), .A2(n86), .ZN(\ab[5][3] ) );
  NOR2_X1 U285 ( .A1(n52), .A2(n86), .ZN(\ab[5][2] ) );
  NOR2_X1 U286 ( .A1(n53), .A2(n86), .ZN(\ab[5][1] ) );
  NOR2_X1 U287 ( .A1(n60), .A2(n86), .ZN(\SUMB[5][16] ) );
  NOR2_X1 U288 ( .A1(n61), .A2(n86), .ZN(\ab[5][15] ) );
  NOR2_X1 U289 ( .A1(n62), .A2(n86), .ZN(\ab[5][14] ) );
  NOR2_X1 U290 ( .A1(n63), .A2(n86), .ZN(\ab[5][13] ) );
  NOR2_X1 U291 ( .A1(n64), .A2(n86), .ZN(\ab[5][12] ) );
  NOR2_X1 U292 ( .A1(n65), .A2(n86), .ZN(\ab[5][11] ) );
  NOR2_X1 U293 ( .A1(n66), .A2(n86), .ZN(\ab[5][10] ) );
  NOR2_X1 U294 ( .A1(n74), .A2(n86), .ZN(\ab[5][0] ) );
  NOR2_X1 U295 ( .A1(n67), .A2(n87), .ZN(\ab[4][9] ) );
  NOR2_X1 U296 ( .A1(n68), .A2(n87), .ZN(\ab[4][8] ) );
  NOR2_X1 U297 ( .A1(n69), .A2(n87), .ZN(\ab[4][7] ) );
  NOR2_X1 U298 ( .A1(n70), .A2(n87), .ZN(\ab[4][6] ) );
  NOR2_X1 U299 ( .A1(n71), .A2(n87), .ZN(\ab[4][5] ) );
  NOR2_X1 U300 ( .A1(n72), .A2(n87), .ZN(\ab[4][4] ) );
  NOR2_X1 U301 ( .A1(n51), .A2(n87), .ZN(\ab[4][3] ) );
  NOR2_X1 U302 ( .A1(n52), .A2(n87), .ZN(\ab[4][2] ) );
  NOR2_X1 U303 ( .A1(n53), .A2(n87), .ZN(\ab[4][1] ) );
  NOR2_X1 U304 ( .A1(n60), .A2(n87), .ZN(\SUMB[4][16] ) );
  NOR2_X1 U305 ( .A1(n61), .A2(n87), .ZN(\ab[4][15] ) );
  NOR2_X1 U306 ( .A1(n62), .A2(n87), .ZN(\ab[4][14] ) );
  NOR2_X1 U307 ( .A1(n63), .A2(n87), .ZN(\ab[4][13] ) );
  NOR2_X1 U308 ( .A1(n64), .A2(n87), .ZN(\ab[4][12] ) );
  NOR2_X1 U309 ( .A1(n65), .A2(n87), .ZN(\ab[4][11] ) );
  NOR2_X1 U310 ( .A1(n66), .A2(n87), .ZN(\ab[4][10] ) );
  NOR2_X1 U311 ( .A1(n74), .A2(n87), .ZN(\ab[4][0] ) );
  NOR2_X1 U312 ( .A1(n67), .A2(n56), .ZN(\ab[3][9] ) );
  NOR2_X1 U313 ( .A1(n68), .A2(n56), .ZN(\ab[3][8] ) );
  NOR2_X1 U314 ( .A1(n69), .A2(n56), .ZN(\ab[3][7] ) );
  NOR2_X1 U315 ( .A1(n70), .A2(n56), .ZN(\ab[3][6] ) );
  NOR2_X1 U316 ( .A1(n71), .A2(n56), .ZN(\ab[3][5] ) );
  NOR2_X1 U317 ( .A1(n72), .A2(n56), .ZN(\ab[3][4] ) );
  NOR2_X1 U318 ( .A1(n51), .A2(n56), .ZN(\ab[3][3] ) );
  NOR2_X1 U319 ( .A1(n52), .A2(n56), .ZN(\ab[3][2] ) );
  NOR2_X1 U320 ( .A1(n53), .A2(n55), .ZN(\ab[3][1] ) );
  NOR2_X1 U321 ( .A1(n60), .A2(n55), .ZN(\SUMB[3][16] ) );
  NOR2_X1 U322 ( .A1(n61), .A2(n55), .ZN(\ab[3][15] ) );
  NOR2_X1 U323 ( .A1(n62), .A2(n55), .ZN(\ab[3][14] ) );
  NOR2_X1 U324 ( .A1(n63), .A2(n55), .ZN(\ab[3][13] ) );
  NOR2_X1 U325 ( .A1(n64), .A2(n55), .ZN(\ab[3][12] ) );
  NOR2_X1 U326 ( .A1(n65), .A2(n55), .ZN(\ab[3][11] ) );
  NOR2_X1 U327 ( .A1(n66), .A2(n55), .ZN(\ab[3][10] ) );
  NOR2_X1 U328 ( .A1(n74), .A2(n55), .ZN(\ab[3][0] ) );
  NOR2_X1 U329 ( .A1(n67), .A2(n57), .ZN(\ab[2][9] ) );
  NOR2_X1 U330 ( .A1(n68), .A2(n57), .ZN(\ab[2][8] ) );
  NOR2_X1 U331 ( .A1(n69), .A2(n57), .ZN(\ab[2][7] ) );
  NOR2_X1 U332 ( .A1(n70), .A2(n57), .ZN(\ab[2][6] ) );
  NOR2_X1 U333 ( .A1(n71), .A2(n57), .ZN(\ab[2][5] ) );
  NOR2_X1 U334 ( .A1(n72), .A2(n57), .ZN(\ab[2][4] ) );
  NOR2_X1 U335 ( .A1(n51), .A2(n57), .ZN(\ab[2][3] ) );
  NOR2_X1 U336 ( .A1(n52), .A2(n57), .ZN(\ab[2][2] ) );
  NOR2_X1 U337 ( .A1(n53), .A2(n88), .ZN(\ab[2][1] ) );
  NOR2_X1 U338 ( .A1(n60), .A2(n88), .ZN(\SUMB[2][16] ) );
  NOR2_X1 U339 ( .A1(n61), .A2(n88), .ZN(\ab[2][15] ) );
  NOR2_X1 U340 ( .A1(n62), .A2(n88), .ZN(\ab[2][14] ) );
  NOR2_X1 U341 ( .A1(n63), .A2(n88), .ZN(\ab[2][13] ) );
  NOR2_X1 U342 ( .A1(n64), .A2(n88), .ZN(\ab[2][12] ) );
  NOR2_X1 U343 ( .A1(n65), .A2(n88), .ZN(\ab[2][11] ) );
  NOR2_X1 U344 ( .A1(n66), .A2(n88), .ZN(\ab[2][10] ) );
  NOR2_X1 U345 ( .A1(n74), .A2(n57), .ZN(\ab[2][0] ) );
  NOR2_X1 U346 ( .A1(n67), .A2(n58), .ZN(\ab[1][9] ) );
  NOR2_X1 U347 ( .A1(n68), .A2(n58), .ZN(\ab[1][8] ) );
  NOR2_X1 U348 ( .A1(n69), .A2(n58), .ZN(\ab[1][7] ) );
  NOR2_X1 U349 ( .A1(n70), .A2(n58), .ZN(\ab[1][6] ) );
  NOR2_X1 U350 ( .A1(n71), .A2(n58), .ZN(\ab[1][5] ) );
  NOR2_X1 U351 ( .A1(n72), .A2(n58), .ZN(\ab[1][4] ) );
  NOR2_X1 U352 ( .A1(n51), .A2(n58), .ZN(\ab[1][3] ) );
  NOR2_X1 U353 ( .A1(n73), .A2(n58), .ZN(\ab[1][2] ) );
  NOR2_X1 U354 ( .A1(n60), .A2(n58), .ZN(\ab[1][16] ) );
  NOR2_X1 U355 ( .A1(n61), .A2(n58), .ZN(\ab[1][15] ) );
  NOR2_X1 U356 ( .A1(n62), .A2(n58), .ZN(\ab[1][14] ) );
  NOR2_X1 U357 ( .A1(n63), .A2(n58), .ZN(\ab[1][13] ) );
  NOR2_X1 U358 ( .A1(n64), .A2(n58), .ZN(\ab[1][12] ) );
  NOR2_X1 U359 ( .A1(n65), .A2(n58), .ZN(\ab[1][11] ) );
  NOR2_X1 U360 ( .A1(n66), .A2(n58), .ZN(\ab[1][10] ) );
  NOR2_X1 U361 ( .A1(n74), .A2(n58), .ZN(\ab[1][0] ) );
  NOR2_X1 U362 ( .A1(n67), .A2(n75), .ZN(\ab[16][9] ) );
  NOR2_X1 U363 ( .A1(n68), .A2(n75), .ZN(\ab[16][8] ) );
  NOR2_X1 U364 ( .A1(n69), .A2(n75), .ZN(\ab[16][7] ) );
  NOR2_X1 U365 ( .A1(n70), .A2(n75), .ZN(\ab[16][6] ) );
  NOR2_X1 U366 ( .A1(n71), .A2(n75), .ZN(\ab[16][5] ) );
  NOR2_X1 U367 ( .A1(n72), .A2(n75), .ZN(\ab[16][4] ) );
  NOR2_X1 U368 ( .A1(n50), .A2(n75), .ZN(\ab[16][3] ) );
  NOR2_X1 U369 ( .A1(n73), .A2(n75), .ZN(\ab[16][2] ) );
  NOR2_X1 U370 ( .A1(n53), .A2(n75), .ZN(\ab[16][1] ) );
  NOR2_X1 U371 ( .A1(n61), .A2(n75), .ZN(\ab[16][15] ) );
  NOR2_X1 U372 ( .A1(n62), .A2(n75), .ZN(\ab[16][14] ) );
  NOR2_X1 U373 ( .A1(n63), .A2(n75), .ZN(\ab[16][13] ) );
  NOR2_X1 U374 ( .A1(n64), .A2(n75), .ZN(\ab[16][12] ) );
  NOR2_X1 U375 ( .A1(n65), .A2(n75), .ZN(\ab[16][11] ) );
  NOR2_X1 U376 ( .A1(n66), .A2(n75), .ZN(\ab[16][10] ) );
  NOR2_X1 U377 ( .A1(n54), .A2(n75), .ZN(\ab[16][0] ) );
  NOR2_X1 U378 ( .A1(n67), .A2(n76), .ZN(\ab[15][9] ) );
  NOR2_X1 U379 ( .A1(n68), .A2(n76), .ZN(\ab[15][8] ) );
  NOR2_X1 U380 ( .A1(n69), .A2(n76), .ZN(\ab[15][7] ) );
  NOR2_X1 U381 ( .A1(n70), .A2(n76), .ZN(\ab[15][6] ) );
  NOR2_X1 U382 ( .A1(n71), .A2(n76), .ZN(\ab[15][5] ) );
  NOR2_X1 U383 ( .A1(n72), .A2(n76), .ZN(\ab[15][4] ) );
  NOR2_X1 U384 ( .A1(n50), .A2(n76), .ZN(\ab[15][3] ) );
  NOR2_X1 U385 ( .A1(n73), .A2(n76), .ZN(\ab[15][2] ) );
  NOR2_X1 U386 ( .A1(n53), .A2(n76), .ZN(\ab[15][1] ) );
  NOR2_X1 U387 ( .A1(n60), .A2(n76), .ZN(\SUMB[15][16] ) );
  NOR2_X1 U388 ( .A1(n61), .A2(n76), .ZN(\ab[15][15] ) );
  NOR2_X1 U389 ( .A1(n62), .A2(n76), .ZN(\ab[15][14] ) );
  NOR2_X1 U390 ( .A1(n63), .A2(n76), .ZN(\ab[15][13] ) );
  NOR2_X1 U391 ( .A1(n64), .A2(n76), .ZN(\ab[15][12] ) );
  NOR2_X1 U392 ( .A1(n65), .A2(n76), .ZN(\ab[15][11] ) );
  NOR2_X1 U393 ( .A1(n66), .A2(n76), .ZN(\ab[15][10] ) );
  NOR2_X1 U394 ( .A1(n54), .A2(n76), .ZN(\ab[15][0] ) );
  NOR2_X1 U395 ( .A1(n67), .A2(n77), .ZN(\ab[14][9] ) );
  NOR2_X1 U396 ( .A1(n68), .A2(n77), .ZN(\ab[14][8] ) );
  NOR2_X1 U397 ( .A1(n69), .A2(n77), .ZN(\ab[14][7] ) );
  NOR2_X1 U398 ( .A1(n70), .A2(n77), .ZN(\ab[14][6] ) );
  NOR2_X1 U399 ( .A1(n71), .A2(n77), .ZN(\ab[14][5] ) );
  NOR2_X1 U400 ( .A1(n72), .A2(n77), .ZN(\ab[14][4] ) );
  NOR2_X1 U401 ( .A1(n50), .A2(n77), .ZN(\ab[14][3] ) );
  NOR2_X1 U402 ( .A1(n73), .A2(n77), .ZN(\ab[14][2] ) );
  NOR2_X1 U403 ( .A1(n53), .A2(n77), .ZN(\ab[14][1] ) );
  NOR2_X1 U404 ( .A1(n60), .A2(n77), .ZN(\SUMB[14][16] ) );
  NOR2_X1 U405 ( .A1(n61), .A2(n77), .ZN(\ab[14][15] ) );
  NOR2_X1 U406 ( .A1(n62), .A2(n77), .ZN(\ab[14][14] ) );
  NOR2_X1 U407 ( .A1(n63), .A2(n77), .ZN(\ab[14][13] ) );
  NOR2_X1 U408 ( .A1(n64), .A2(n77), .ZN(\ab[14][12] ) );
  NOR2_X1 U409 ( .A1(n65), .A2(n77), .ZN(\ab[14][11] ) );
  NOR2_X1 U410 ( .A1(n66), .A2(n77), .ZN(\ab[14][10] ) );
  NOR2_X1 U411 ( .A1(n54), .A2(n77), .ZN(\ab[14][0] ) );
  NOR2_X1 U412 ( .A1(n67), .A2(n78), .ZN(\ab[13][9] ) );
  NOR2_X1 U413 ( .A1(n68), .A2(n78), .ZN(\ab[13][8] ) );
  NOR2_X1 U414 ( .A1(n69), .A2(n78), .ZN(\ab[13][7] ) );
  NOR2_X1 U415 ( .A1(n70), .A2(n78), .ZN(\ab[13][6] ) );
  NOR2_X1 U416 ( .A1(n71), .A2(n78), .ZN(\ab[13][5] ) );
  NOR2_X1 U417 ( .A1(n72), .A2(n78), .ZN(\ab[13][4] ) );
  NOR2_X1 U418 ( .A1(n50), .A2(n78), .ZN(\ab[13][3] ) );
  NOR2_X1 U419 ( .A1(n73), .A2(n78), .ZN(\ab[13][2] ) );
  NOR2_X1 U420 ( .A1(n53), .A2(n78), .ZN(\ab[13][1] ) );
  NOR2_X1 U421 ( .A1(n60), .A2(n78), .ZN(\SUMB[13][16] ) );
  NOR2_X1 U422 ( .A1(n61), .A2(n78), .ZN(\ab[13][15] ) );
  NOR2_X1 U423 ( .A1(n62), .A2(n78), .ZN(\ab[13][14] ) );
  NOR2_X1 U424 ( .A1(n63), .A2(n78), .ZN(\ab[13][13] ) );
  NOR2_X1 U425 ( .A1(n64), .A2(n78), .ZN(\ab[13][12] ) );
  NOR2_X1 U426 ( .A1(n65), .A2(n78), .ZN(\ab[13][11] ) );
  NOR2_X1 U427 ( .A1(n66), .A2(n78), .ZN(\ab[13][10] ) );
  NOR2_X1 U428 ( .A1(n54), .A2(n78), .ZN(\ab[13][0] ) );
  NOR2_X1 U429 ( .A1(n67), .A2(n79), .ZN(\ab[12][9] ) );
  NOR2_X1 U430 ( .A1(n68), .A2(n79), .ZN(\ab[12][8] ) );
  NOR2_X1 U431 ( .A1(n69), .A2(n79), .ZN(\ab[12][7] ) );
  NOR2_X1 U432 ( .A1(n70), .A2(n79), .ZN(\ab[12][6] ) );
  NOR2_X1 U433 ( .A1(n71), .A2(n79), .ZN(\ab[12][5] ) );
  NOR2_X1 U434 ( .A1(n72), .A2(n79), .ZN(\ab[12][4] ) );
  NOR2_X1 U435 ( .A1(n50), .A2(n79), .ZN(\ab[12][3] ) );
  NOR2_X1 U436 ( .A1(n73), .A2(n79), .ZN(\ab[12][2] ) );
  NOR2_X1 U437 ( .A1(n53), .A2(n79), .ZN(\ab[12][1] ) );
  NOR2_X1 U438 ( .A1(n60), .A2(n79), .ZN(\SUMB[12][16] ) );
  NOR2_X1 U439 ( .A1(n61), .A2(n79), .ZN(\ab[12][15] ) );
  NOR2_X1 U440 ( .A1(n62), .A2(n79), .ZN(\ab[12][14] ) );
  NOR2_X1 U441 ( .A1(n63), .A2(n79), .ZN(\ab[12][13] ) );
  NOR2_X1 U442 ( .A1(n64), .A2(n79), .ZN(\ab[12][12] ) );
  NOR2_X1 U443 ( .A1(n65), .A2(n79), .ZN(\ab[12][11] ) );
  NOR2_X1 U444 ( .A1(n66), .A2(n79), .ZN(\ab[12][10] ) );
  NOR2_X1 U445 ( .A1(n54), .A2(n79), .ZN(\ab[12][0] ) );
  NOR2_X1 U446 ( .A1(n67), .A2(n80), .ZN(\ab[11][9] ) );
  NOR2_X1 U447 ( .A1(n68), .A2(n80), .ZN(\ab[11][8] ) );
  NOR2_X1 U448 ( .A1(n69), .A2(n80), .ZN(\ab[11][7] ) );
  NOR2_X1 U449 ( .A1(n70), .A2(n80), .ZN(\ab[11][6] ) );
  NOR2_X1 U450 ( .A1(n71), .A2(n80), .ZN(\ab[11][5] ) );
  NOR2_X1 U451 ( .A1(n72), .A2(n80), .ZN(\ab[11][4] ) );
  NOR2_X1 U452 ( .A1(n50), .A2(n80), .ZN(\ab[11][3] ) );
  NOR2_X1 U453 ( .A1(n73), .A2(n80), .ZN(\ab[11][2] ) );
  NOR2_X1 U454 ( .A1(n53), .A2(n80), .ZN(\ab[11][1] ) );
  NOR2_X1 U455 ( .A1(n60), .A2(n80), .ZN(\SUMB[11][16] ) );
  NOR2_X1 U456 ( .A1(n61), .A2(n80), .ZN(\ab[11][15] ) );
  NOR2_X1 U457 ( .A1(n62), .A2(n80), .ZN(\ab[11][14] ) );
  NOR2_X1 U458 ( .A1(n63), .A2(n80), .ZN(\ab[11][13] ) );
  NOR2_X1 U459 ( .A1(n64), .A2(n80), .ZN(\ab[11][12] ) );
  NOR2_X1 U460 ( .A1(n65), .A2(n80), .ZN(\ab[11][11] ) );
  NOR2_X1 U461 ( .A1(n66), .A2(n80), .ZN(\ab[11][10] ) );
  NOR2_X1 U462 ( .A1(n54), .A2(n80), .ZN(\ab[11][0] ) );
  NOR2_X1 U463 ( .A1(n67), .A2(n81), .ZN(\ab[10][9] ) );
  NOR2_X1 U464 ( .A1(n68), .A2(n81), .ZN(\ab[10][8] ) );
  NOR2_X1 U465 ( .A1(n69), .A2(n81), .ZN(\ab[10][7] ) );
  NOR2_X1 U466 ( .A1(n70), .A2(n81), .ZN(\ab[10][6] ) );
  NOR2_X1 U467 ( .A1(n71), .A2(n81), .ZN(\ab[10][5] ) );
  NOR2_X1 U468 ( .A1(n72), .A2(n81), .ZN(\ab[10][4] ) );
  NOR2_X1 U469 ( .A1(n50), .A2(n81), .ZN(\ab[10][3] ) );
  NOR2_X1 U470 ( .A1(n73), .A2(n81), .ZN(\ab[10][2] ) );
  NOR2_X1 U471 ( .A1(n53), .A2(n81), .ZN(\ab[10][1] ) );
  NOR2_X1 U472 ( .A1(n60), .A2(n81), .ZN(\SUMB[10][16] ) );
  NOR2_X1 U473 ( .A1(n61), .A2(n81), .ZN(\ab[10][15] ) );
  NOR2_X1 U474 ( .A1(n62), .A2(n81), .ZN(\ab[10][14] ) );
  NOR2_X1 U475 ( .A1(n63), .A2(n81), .ZN(\ab[10][13] ) );
  NOR2_X1 U476 ( .A1(n64), .A2(n81), .ZN(\ab[10][12] ) );
  NOR2_X1 U477 ( .A1(n65), .A2(n81), .ZN(\ab[10][11] ) );
  NOR2_X1 U478 ( .A1(n66), .A2(n81), .ZN(\ab[10][10] ) );
  NOR2_X1 U479 ( .A1(n54), .A2(n81), .ZN(\ab[10][0] ) );
  NOR2_X1 U480 ( .A1(n67), .A2(n59), .ZN(\ab[0][9] ) );
  NOR2_X1 U481 ( .A1(n68), .A2(n59), .ZN(\ab[0][8] ) );
  NOR2_X1 U482 ( .A1(n69), .A2(n59), .ZN(\ab[0][7] ) );
  NOR2_X1 U483 ( .A1(n70), .A2(n59), .ZN(\ab[0][6] ) );
  NOR2_X1 U484 ( .A1(n71), .A2(n59), .ZN(\ab[0][5] ) );
  NOR2_X1 U485 ( .A1(n72), .A2(n59), .ZN(\ab[0][4] ) );
  NOR2_X1 U486 ( .A1(n50), .A2(n59), .ZN(\ab[0][3] ) );
  NOR2_X1 U487 ( .A1(n52), .A2(n59), .ZN(\ab[0][2] ) );
  NOR2_X1 U488 ( .A1(n53), .A2(n89), .ZN(\ab[0][1] ) );
  NOR2_X1 U489 ( .A1(n60), .A2(n89), .ZN(\ab[0][16] ) );
  NOR2_X1 U490 ( .A1(n61), .A2(n89), .ZN(\ab[0][15] ) );
  NOR2_X1 U491 ( .A1(n62), .A2(n89), .ZN(\ab[0][14] ) );
  NOR2_X1 U492 ( .A1(n63), .A2(n89), .ZN(\ab[0][13] ) );
  NOR2_X1 U493 ( .A1(n64), .A2(n89), .ZN(\ab[0][12] ) );
  NOR2_X1 U494 ( .A1(n65), .A2(n89), .ZN(\ab[0][11] ) );
  NOR2_X1 U495 ( .A1(n66), .A2(n89), .ZN(\ab[0][10] ) );
  NOR2_X1 U496 ( .A1(n54), .A2(n59), .ZN(PRODUCT[0]) );
  NAND2_X2 U101 ( .A1(\SUMB[21][9] ), .A2(\CARRYB[21][8] ), .ZN(n90) );
  INV_X4 U102 ( .A(n90), .ZN(\CARRYB[22][8] ) );
  XNOR2_X2 U103 ( .A(\CARRYB[21][8] ), .B(\SUMB[21][9] ), .ZN(n91) );
  INV_X4 U104 ( .A(n91), .ZN(\SUMB[22][8] ) );
  NAND2_X2 U105 ( .A1(\SUMB[21][8] ), .A2(\CARRYB[21][7] ), .ZN(n92) );
  INV_X4 U106 ( .A(n92), .ZN(\CARRYB[22][7] ) );
  XNOR2_X2 U107 ( .A(\CARRYB[21][7] ), .B(\SUMB[21][8] ), .ZN(n93) );
  INV_X4 U108 ( .A(n93), .ZN(\SUMB[22][7] ) );
  NAND2_X2 U109 ( .A1(\SUMB[21][7] ), .A2(\CARRYB[21][6] ), .ZN(n94) );
  INV_X4 U110 ( .A(n94), .ZN(\CARRYB[22][6] ) );
  XNOR2_X2 U111 ( .A(\CARRYB[21][6] ), .B(\SUMB[21][7] ), .ZN(n95) );
  INV_X4 U112 ( .A(n95), .ZN(\SUMB[22][6] ) );
  NAND2_X2 U113 ( .A1(\SUMB[21][6] ), .A2(\CARRYB[21][5] ), .ZN(n96) );
  INV_X4 U114 ( .A(n96), .ZN(\CARRYB[22][5] ) );
  XNOR2_X2 U115 ( .A(\CARRYB[21][5] ), .B(\SUMB[21][6] ), .ZN(n97) );
  INV_X4 U116 ( .A(n97), .ZN(\SUMB[22][5] ) );
  NAND2_X2 U117 ( .A1(\SUMB[21][5] ), .A2(\CARRYB[21][4] ), .ZN(n98) );
  INV_X4 U118 ( .A(n98), .ZN(\CARRYB[22][4] ) );
  XNOR2_X2 U119 ( .A(\CARRYB[21][4] ), .B(\SUMB[21][5] ), .ZN(n99) );
  INV_X4 U120 ( .A(n99), .ZN(\SUMB[22][4] ) );
  NAND2_X2 U121 ( .A1(\SUMB[21][4] ), .A2(\CARRYB[21][3] ), .ZN(n100) );
  INV_X4 U122 ( .A(n100), .ZN(\CARRYB[22][3] ) );
  XNOR2_X2 U123 ( .A(\CARRYB[21][3] ), .B(\SUMB[21][4] ), .ZN(n101) );
  INV_X4 U124 ( .A(n101), .ZN(\SUMB[22][3] ) );
  NAND2_X2 U125 ( .A1(\SUMB[21][3] ), .A2(\CARRYB[21][2] ), .ZN(n102) );
  INV_X4 U126 ( .A(n102), .ZN(\CARRYB[22][2] ) );
  XNOR2_X2 U127 ( .A(\CARRYB[21][2] ), .B(\SUMB[21][3] ), .ZN(n103) );
  INV_X4 U128 ( .A(n103), .ZN(\SUMB[22][2] ) );
  NAND2_X2 U129 ( .A1(\SUMB[21][2] ), .A2(\CARRYB[21][1] ), .ZN(n104) );
  INV_X4 U130 ( .A(n104), .ZN(\CARRYB[22][1] ) );
  XNOR2_X2 U131 ( .A(\CARRYB[21][1] ), .B(\SUMB[21][2] ), .ZN(n105) );
  INV_X4 U132 ( .A(n105), .ZN(\SUMB[22][1] ) );
  NAND2_X2 U133 ( .A1(\SUMB[21][1] ), .A2(\CARRYB[21][0] ), .ZN(n106) );
  INV_X4 U134 ( .A(n106), .ZN(\CARRYB[22][0] ) );
  XNOR2_X2 U135 ( .A(\CARRYB[21][0] ), .B(\SUMB[21][1] ), .ZN(n107) );
  INV_X4 U136 ( .A(n107), .ZN(PRODUCT[22]) );
  NAND2_X2 U137 ( .A1(\SUMB[22][8] ), .A2(\CARRYB[22][7] ), .ZN(n108) );
  INV_X4 U138 ( .A(n108), .ZN(\CARRYB[23][7] ) );
  XNOR2_X2 U139 ( .A(\CARRYB[22][7] ), .B(\SUMB[22][8] ), .ZN(n109) );
  INV_X4 U140 ( .A(n109), .ZN(\SUMB[23][7] ) );
  NAND2_X2 U141 ( .A1(\SUMB[22][7] ), .A2(\CARRYB[22][6] ), .ZN(n110) );
  INV_X4 U142 ( .A(n110), .ZN(\CARRYB[23][6] ) );
  XNOR2_X2 U143 ( .A(\CARRYB[22][6] ), .B(\SUMB[22][7] ), .ZN(n111) );
  INV_X4 U144 ( .A(n111), .ZN(\SUMB[23][6] ) );
  NAND2_X2 U145 ( .A1(\SUMB[22][6] ), .A2(\CARRYB[22][5] ), .ZN(n112) );
  INV_X4 U146 ( .A(n112), .ZN(\CARRYB[23][5] ) );
  XNOR2_X2 U147 ( .A(\CARRYB[22][5] ), .B(\SUMB[22][6] ), .ZN(n113) );
  INV_X4 U148 ( .A(n113), .ZN(\SUMB[23][5] ) );
  NAND2_X2 U149 ( .A1(\SUMB[22][5] ), .A2(\CARRYB[22][4] ), .ZN(n114) );
  INV_X4 U150 ( .A(n114), .ZN(\CARRYB[23][4] ) );
  XNOR2_X2 U151 ( .A(\CARRYB[22][4] ), .B(\SUMB[22][5] ), .ZN(n115) );
  INV_X4 U152 ( .A(n115), .ZN(\SUMB[23][4] ) );
  NAND2_X2 U153 ( .A1(\SUMB[22][4] ), .A2(\CARRYB[22][3] ), .ZN(n116) );
  INV_X4 U154 ( .A(n116), .ZN(\CARRYB[23][3] ) );
  XNOR2_X2 U155 ( .A(\CARRYB[22][3] ), .B(\SUMB[22][4] ), .ZN(n117) );
  INV_X4 U156 ( .A(n117), .ZN(\SUMB[23][3] ) );
  NAND2_X2 U157 ( .A1(\SUMB[22][3] ), .A2(\CARRYB[22][2] ), .ZN(n118) );
  INV_X4 U158 ( .A(n118), .ZN(\CARRYB[23][2] ) );
  XNOR2_X2 U159 ( .A(\CARRYB[22][2] ), .B(\SUMB[22][3] ), .ZN(n119) );
  INV_X4 U160 ( .A(n119), .ZN(\SUMB[23][2] ) );
  NAND2_X2 U161 ( .A1(\SUMB[22][2] ), .A2(\CARRYB[22][1] ), .ZN(n120) );
  INV_X4 U162 ( .A(n120), .ZN(\CARRYB[23][1] ) );
  XNOR2_X2 U163 ( .A(\CARRYB[22][1] ), .B(\SUMB[22][2] ), .ZN(n121) );
  INV_X4 U164 ( .A(n121), .ZN(\SUMB[23][1] ) );
  NAND2_X2 U165 ( .A1(\SUMB[22][1] ), .A2(\CARRYB[22][0] ), .ZN(n122) );
  INV_X4 U166 ( .A(n122), .ZN(\CARRYB[23][0] ) );
  XNOR2_X2 U167 ( .A(\CARRYB[22][0] ), .B(\SUMB[22][1] ), .ZN(n123) );
  INV_X4 U168 ( .A(n123), .ZN(PRODUCT[23]) );
  NAND2_X2 U169 ( .A1(\SUMB[23][7] ), .A2(\CARRYB[23][6] ), .ZN(n124) );
  INV_X4 U170 ( .A(n124), .ZN(\CARRYB[24][6] ) );
  XNOR2_X2 U171 ( .A(\CARRYB[23][6] ), .B(\SUMB[23][7] ), .ZN(n125) );
  INV_X4 U172 ( .A(n125), .ZN(\SUMB[24][6] ) );
  NAND2_X2 U173 ( .A1(\SUMB[23][6] ), .A2(\CARRYB[23][5] ), .ZN(n126) );
  INV_X4 U174 ( .A(n126), .ZN(\CARRYB[24][5] ) );
  XNOR2_X2 U175 ( .A(\CARRYB[23][5] ), .B(\SUMB[23][6] ), .ZN(n127) );
  INV_X4 U176 ( .A(n127), .ZN(\SUMB[24][5] ) );
  NAND2_X2 U177 ( .A1(\SUMB[23][5] ), .A2(\CARRYB[23][4] ), .ZN(n128) );
  INV_X4 U178 ( .A(n128), .ZN(\CARRYB[24][4] ) );
  XNOR2_X2 U179 ( .A(\CARRYB[23][4] ), .B(\SUMB[23][5] ), .ZN(n129) );
  INV_X4 U180 ( .A(n129), .ZN(\SUMB[24][4] ) );
  NAND2_X2 U181 ( .A1(\SUMB[23][4] ), .A2(\CARRYB[23][3] ), .ZN(n130) );
  INV_X4 U182 ( .A(n130), .ZN(\CARRYB[24][3] ) );
  XNOR2_X2 U183 ( .A(\CARRYB[23][3] ), .B(\SUMB[23][4] ), .ZN(n131) );
  INV_X4 U184 ( .A(n131), .ZN(\SUMB[24][3] ) );
  NAND2_X2 U185 ( .A1(\SUMB[23][3] ), .A2(\CARRYB[23][2] ), .ZN(n132) );
  INV_X4 U186 ( .A(n132), .ZN(\CARRYB[24][2] ) );
  XNOR2_X2 U187 ( .A(\CARRYB[23][2] ), .B(\SUMB[23][3] ), .ZN(n133) );
  INV_X4 U188 ( .A(n133), .ZN(\SUMB[24][2] ) );
  NAND2_X2 U189 ( .A1(\SUMB[23][2] ), .A2(\CARRYB[23][1] ), .ZN(n134) );
  INV_X4 U190 ( .A(n134), .ZN(\CARRYB[24][1] ) );
  XNOR2_X2 U191 ( .A(\CARRYB[23][1] ), .B(\SUMB[23][2] ), .ZN(n135) );
  INV_X4 U192 ( .A(n135), .ZN(\SUMB[24][1] ) );
  NAND2_X2 U193 ( .A1(\SUMB[23][1] ), .A2(\CARRYB[23][0] ), .ZN(n136) );
  INV_X4 U194 ( .A(n136), .ZN(\CARRYB[24][0] ) );
  XNOR2_X2 U195 ( .A(\CARRYB[23][0] ), .B(\SUMB[23][1] ), .ZN(n137) );
  INV_X4 U196 ( .A(n137), .ZN(PRODUCT[24]) );
  NAND2_X2 U197 ( .A1(\SUMB[24][6] ), .A2(\CARRYB[24][5] ), .ZN(n138) );
  INV_X4 U198 ( .A(n138), .ZN(\CARRYB[25][5] ) );
  XNOR2_X2 U199 ( .A(\CARRYB[24][5] ), .B(\SUMB[24][6] ), .ZN(n139) );
  INV_X4 U200 ( .A(n139), .ZN(\SUMB[25][5] ) );
  NAND2_X2 U201 ( .A1(\SUMB[24][5] ), .A2(\CARRYB[24][4] ), .ZN(n140) );
  INV_X4 U202 ( .A(n140), .ZN(\CARRYB[25][4] ) );
  XNOR2_X2 U203 ( .A(\CARRYB[24][4] ), .B(\SUMB[24][5] ), .ZN(n141) );
  INV_X4 U204 ( .A(n141), .ZN(\SUMB[25][4] ) );
  NAND2_X2 U205 ( .A1(\SUMB[24][4] ), .A2(\CARRYB[24][3] ), .ZN(n142) );
  INV_X4 U497 ( .A(n142), .ZN(\CARRYB[25][3] ) );
  XNOR2_X2 U498 ( .A(\CARRYB[24][3] ), .B(\SUMB[24][4] ), .ZN(n143) );
  INV_X4 U499 ( .A(n143), .ZN(\SUMB[25][3] ) );
  NAND2_X2 U500 ( .A1(\SUMB[24][3] ), .A2(\CARRYB[24][2] ), .ZN(n144) );
  INV_X4 U501 ( .A(n144), .ZN(\CARRYB[25][2] ) );
  XNOR2_X2 U502 ( .A(\CARRYB[24][2] ), .B(\SUMB[24][3] ), .ZN(n145) );
  INV_X4 U503 ( .A(n145), .ZN(\SUMB[25][2] ) );
  NAND2_X2 U504 ( .A1(\SUMB[24][2] ), .A2(\CARRYB[24][1] ), .ZN(n146) );
  INV_X4 U505 ( .A(n146), .ZN(\CARRYB[25][1] ) );
  XNOR2_X2 U506 ( .A(\CARRYB[24][1] ), .B(\SUMB[24][2] ), .ZN(n147) );
  INV_X4 U507 ( .A(n147), .ZN(\SUMB[25][1] ) );
  NAND2_X2 U508 ( .A1(\SUMB[24][1] ), .A2(\CARRYB[24][0] ), .ZN(n148) );
  INV_X4 U509 ( .A(n148), .ZN(\CARRYB[25][0] ) );
  XNOR2_X2 U510 ( .A(\CARRYB[24][0] ), .B(\SUMB[24][1] ), .ZN(n149) );
  INV_X4 U511 ( .A(n149), .ZN(PRODUCT[25]) );
  NAND2_X2 U512 ( .A1(\SUMB[25][5] ), .A2(\CARRYB[25][4] ), .ZN(n150) );
  INV_X4 U513 ( .A(n150), .ZN(\CARRYB[26][4] ) );
  XNOR2_X2 U514 ( .A(\CARRYB[25][4] ), .B(\SUMB[25][5] ), .ZN(n151) );
  INV_X4 U515 ( .A(n151), .ZN(\SUMB[26][4] ) );
  NAND2_X2 U516 ( .A1(\SUMB[25][4] ), .A2(\CARRYB[25][3] ), .ZN(n152) );
  INV_X4 U517 ( .A(n152), .ZN(\CARRYB[26][3] ) );
  XNOR2_X2 U518 ( .A(\CARRYB[25][3] ), .B(\SUMB[25][4] ), .ZN(n153) );
  INV_X4 U519 ( .A(n153), .ZN(\SUMB[26][3] ) );
  NAND2_X2 U520 ( .A1(\SUMB[25][3] ), .A2(\CARRYB[25][2] ), .ZN(n154) );
  INV_X4 U521 ( .A(n154), .ZN(\CARRYB[26][2] ) );
  XNOR2_X2 U522 ( .A(\CARRYB[25][2] ), .B(\SUMB[25][3] ), .ZN(n155) );
  INV_X4 U523 ( .A(n155), .ZN(\SUMB[26][2] ) );
  NAND2_X2 U524 ( .A1(\SUMB[25][2] ), .A2(\CARRYB[25][1] ), .ZN(n156) );
  INV_X4 U525 ( .A(n156), .ZN(\CARRYB[26][1] ) );
  XNOR2_X2 U526 ( .A(\CARRYB[25][1] ), .B(\SUMB[25][2] ), .ZN(n157) );
  INV_X4 U527 ( .A(n157), .ZN(\SUMB[26][1] ) );
  NAND2_X2 U528 ( .A1(\SUMB[25][1] ), .A2(\CARRYB[25][0] ), .ZN(n158) );
  INV_X4 U529 ( .A(n158), .ZN(\CARRYB[26][0] ) );
  XNOR2_X2 U530 ( .A(\CARRYB[25][0] ), .B(\SUMB[25][1] ), .ZN(n159) );
  INV_X4 U531 ( .A(n159), .ZN(PRODUCT[26]) );
  NAND2_X2 U532 ( .A1(\SUMB[26][4] ), .A2(\CARRYB[26][3] ), .ZN(n160) );
  INV_X4 U533 ( .A(n160), .ZN(\CARRYB[27][3] ) );
  XNOR2_X2 U534 ( .A(\CARRYB[26][3] ), .B(\SUMB[26][4] ), .ZN(n161) );
  INV_X4 U535 ( .A(n161), .ZN(\SUMB[27][3] ) );
  NAND2_X2 U536 ( .A1(\SUMB[26][3] ), .A2(\CARRYB[26][2] ), .ZN(n162) );
  INV_X4 U537 ( .A(n162), .ZN(\CARRYB[27][2] ) );
  XNOR2_X2 U538 ( .A(\CARRYB[26][2] ), .B(\SUMB[26][3] ), .ZN(n163) );
  INV_X4 U539 ( .A(n163), .ZN(\SUMB[27][2] ) );
  NAND2_X2 U540 ( .A1(\SUMB[26][2] ), .A2(\CARRYB[26][1] ), .ZN(n164) );
  INV_X4 U541 ( .A(n164), .ZN(\CARRYB[27][1] ) );
  XNOR2_X2 U542 ( .A(\CARRYB[26][1] ), .B(\SUMB[26][2] ), .ZN(n165) );
  INV_X4 U543 ( .A(n165), .ZN(\SUMB[27][1] ) );
  NAND2_X2 U544 ( .A1(\SUMB[26][1] ), .A2(\CARRYB[26][0] ), .ZN(n166) );
  INV_X4 U545 ( .A(n166), .ZN(\CARRYB[27][0] ) );
  XNOR2_X2 U546 ( .A(\CARRYB[26][0] ), .B(\SUMB[26][1] ), .ZN(n167) );
  INV_X4 U547 ( .A(n167), .ZN(PRODUCT[27]) );
  NAND2_X2 U548 ( .A1(\SUMB[27][3] ), .A2(\CARRYB[27][2] ), .ZN(n168) );
  INV_X4 U549 ( .A(n168), .ZN(\CARRYB[28][2] ) );
  XNOR2_X2 U550 ( .A(\CARRYB[27][2] ), .B(\SUMB[27][3] ), .ZN(n169) );
  INV_X4 U551 ( .A(n169), .ZN(\SUMB[28][2] ) );
  NAND2_X2 U552 ( .A1(\SUMB[27][2] ), .A2(\CARRYB[27][1] ), .ZN(n170) );
  INV_X4 U553 ( .A(n170), .ZN(\CARRYB[28][1] ) );
  XNOR2_X2 U554 ( .A(\CARRYB[27][1] ), .B(\SUMB[27][2] ), .ZN(n171) );
  INV_X4 U555 ( .A(n171), .ZN(\SUMB[28][1] ) );
  NAND2_X2 U556 ( .A1(\SUMB[27][1] ), .A2(\CARRYB[27][0] ), .ZN(n172) );
  INV_X4 U557 ( .A(n172), .ZN(\CARRYB[28][0] ) );
  XNOR2_X2 U558 ( .A(\CARRYB[27][0] ), .B(\SUMB[27][1] ), .ZN(n173) );
  INV_X4 U559 ( .A(n173), .ZN(PRODUCT[28]) );
  NAND2_X2 U560 ( .A1(\SUMB[28][2] ), .A2(\CARRYB[28][1] ), .ZN(n174) );
  INV_X4 U561 ( .A(n174), .ZN(\CARRYB[29][1] ) );
  XNOR2_X2 U562 ( .A(\CARRYB[28][1] ), .B(\SUMB[28][2] ), .ZN(n175) );
  INV_X4 U563 ( .A(n175), .ZN(\SUMB[29][1] ) );
  NAND2_X2 U564 ( .A1(\SUMB[28][1] ), .A2(\CARRYB[28][0] ), .ZN(n176) );
  INV_X4 U565 ( .A(n176), .ZN(\CARRYB[29][0] ) );
  XNOR2_X2 U566 ( .A(\CARRYB[28][0] ), .B(\SUMB[28][1] ), .ZN(n177) );
  INV_X4 U567 ( .A(n177), .ZN(PRODUCT[29]) );
  NAND2_X2 U568 ( .A1(\SUMB[29][1] ), .A2(\CARRYB[29][0] ), .ZN(n178) );
  INV_X4 U569 ( .A(n178), .ZN(\CARRYB[30][0] ) );
  XNOR2_X2 U570 ( .A(\CARRYB[29][0] ), .B(\SUMB[29][1] ), .ZN(n179) );
  INV_X4 U571 ( .A(n179), .ZN(PRODUCT[30]) );
  NAND2_X2 U572 ( .A1(\SUMB[16][9] ), .A2(\CARRYB[16][8] ), .ZN(n180) );
  INV_X4 U573 ( .A(n180), .ZN(\CARRYB[17][8] ) );
  XNOR2_X2 U574 ( .A(\CARRYB[16][8] ), .B(\SUMB[16][9] ), .ZN(n181) );
  INV_X4 U575 ( .A(n181), .ZN(\SUMB[17][8] ) );
  NAND2_X2 U576 ( .A1(\SUMB[16][8] ), .A2(\CARRYB[16][7] ), .ZN(n182) );
  INV_X4 U577 ( .A(n182), .ZN(\CARRYB[17][7] ) );
  XNOR2_X2 U578 ( .A(\CARRYB[16][7] ), .B(\SUMB[16][8] ), .ZN(n183) );
  INV_X4 U579 ( .A(n183), .ZN(\SUMB[17][7] ) );
  NAND2_X2 U580 ( .A1(\SUMB[16][7] ), .A2(\CARRYB[16][6] ), .ZN(n184) );
  INV_X4 U581 ( .A(n184), .ZN(\CARRYB[17][6] ) );
  XNOR2_X2 U582 ( .A(\CARRYB[16][6] ), .B(\SUMB[16][7] ), .ZN(n185) );
  INV_X4 U583 ( .A(n185), .ZN(\SUMB[17][6] ) );
  NAND2_X2 U584 ( .A1(\SUMB[16][6] ), .A2(\CARRYB[16][5] ), .ZN(n186) );
  INV_X4 U585 ( .A(n186), .ZN(\CARRYB[17][5] ) );
  XNOR2_X2 U586 ( .A(\CARRYB[16][5] ), .B(\SUMB[16][6] ), .ZN(n187) );
  INV_X4 U587 ( .A(n187), .ZN(\SUMB[17][5] ) );
  NAND2_X2 U588 ( .A1(\SUMB[16][5] ), .A2(\CARRYB[16][4] ), .ZN(n188) );
  INV_X4 U589 ( .A(n188), .ZN(\CARRYB[17][4] ) );
  XNOR2_X2 U590 ( .A(\CARRYB[16][4] ), .B(\SUMB[16][5] ), .ZN(n189) );
  INV_X4 U591 ( .A(n189), .ZN(\SUMB[17][4] ) );
  NAND2_X2 U592 ( .A1(\SUMB[16][4] ), .A2(\CARRYB[16][3] ), .ZN(n190) );
  INV_X4 U593 ( .A(n190), .ZN(\CARRYB[17][3] ) );
  XNOR2_X2 U594 ( .A(\CARRYB[16][3] ), .B(\SUMB[16][4] ), .ZN(n191) );
  INV_X4 U595 ( .A(n191), .ZN(\SUMB[17][3] ) );
  NAND2_X2 U596 ( .A1(\SUMB[16][3] ), .A2(\CARRYB[16][2] ), .ZN(n192) );
  INV_X4 U597 ( .A(n192), .ZN(\CARRYB[17][2] ) );
  XNOR2_X2 U598 ( .A(\CARRYB[16][2] ), .B(\SUMB[16][3] ), .ZN(n193) );
  INV_X4 U599 ( .A(n193), .ZN(\SUMB[17][2] ) );
  NAND2_X2 U600 ( .A1(\SUMB[16][2] ), .A2(\CARRYB[16][1] ), .ZN(n194) );
  INV_X4 U601 ( .A(n194), .ZN(\CARRYB[17][1] ) );
  XNOR2_X2 U602 ( .A(\CARRYB[16][1] ), .B(\SUMB[16][2] ), .ZN(n195) );
  INV_X4 U603 ( .A(n195), .ZN(\SUMB[17][1] ) );
  NAND2_X2 U604 ( .A1(\SUMB[16][14] ), .A2(\CARRYB[16][13] ), .ZN(n196) );
  INV_X4 U605 ( .A(n196), .ZN(\CARRYB[17][13] ) );
  XNOR2_X2 U606 ( .A(\CARRYB[16][13] ), .B(\SUMB[16][14] ), .ZN(n197) );
  INV_X4 U607 ( .A(n197), .ZN(\SUMB[17][13] ) );
  NAND2_X2 U608 ( .A1(\SUMB[16][13] ), .A2(\CARRYB[16][12] ), .ZN(n198) );
  INV_X4 U609 ( .A(n198), .ZN(\CARRYB[17][12] ) );
  XNOR2_X2 U610 ( .A(\CARRYB[16][12] ), .B(\SUMB[16][13] ), .ZN(n199) );
  INV_X4 U611 ( .A(n199), .ZN(\SUMB[17][12] ) );
  NAND2_X2 U612 ( .A1(\SUMB[16][12] ), .A2(\CARRYB[16][11] ), .ZN(n200) );
  INV_X4 U613 ( .A(n200), .ZN(\CARRYB[17][11] ) );
  XNOR2_X2 U614 ( .A(\CARRYB[16][11] ), .B(\SUMB[16][12] ), .ZN(n201) );
  INV_X4 U615 ( .A(n201), .ZN(\SUMB[17][11] ) );
  NAND2_X2 U616 ( .A1(\SUMB[16][11] ), .A2(\CARRYB[16][10] ), .ZN(n202) );
  INV_X4 U617 ( .A(n202), .ZN(\CARRYB[17][10] ) );
  XNOR2_X2 U618 ( .A(\CARRYB[16][10] ), .B(\SUMB[16][11] ), .ZN(n203) );
  INV_X4 U619 ( .A(n203), .ZN(\SUMB[17][10] ) );
  NAND2_X2 U620 ( .A1(\SUMB[16][1] ), .A2(\CARRYB[16][0] ), .ZN(n204) );
  INV_X4 U621 ( .A(n204), .ZN(\CARRYB[17][0] ) );
  XNOR2_X2 U622 ( .A(\CARRYB[16][0] ), .B(\SUMB[16][1] ), .ZN(n205) );
  INV_X4 U623 ( .A(n205), .ZN(PRODUCT[17]) );
  NAND2_X2 U624 ( .A1(\SUMB[16][10] ), .A2(\CARRYB[16][9] ), .ZN(n206) );
  INV_X4 U625 ( .A(n206), .ZN(\CARRYB[17][9] ) );
  XNOR2_X2 U626 ( .A(\CARRYB[16][9] ), .B(\SUMB[16][10] ), .ZN(n207) );
  INV_X4 U627 ( .A(n207), .ZN(\SUMB[17][9] ) );
  NAND2_X2 U628 ( .A1(\SUMB[17][9] ), .A2(\CARRYB[17][8] ), .ZN(n208) );
  INV_X4 U629 ( .A(n208), .ZN(\CARRYB[18][8] ) );
  XNOR2_X2 U630 ( .A(\CARRYB[17][8] ), .B(\SUMB[17][9] ), .ZN(n209) );
  INV_X4 U631 ( .A(n209), .ZN(\SUMB[18][8] ) );
  NAND2_X2 U632 ( .A1(\SUMB[17][8] ), .A2(\CARRYB[17][7] ), .ZN(n210) );
  INV_X4 U633 ( .A(n210), .ZN(\CARRYB[18][7] ) );
  XNOR2_X2 U634 ( .A(\CARRYB[17][7] ), .B(\SUMB[17][8] ), .ZN(n211) );
  INV_X4 U635 ( .A(n211), .ZN(\SUMB[18][7] ) );
  NAND2_X2 U636 ( .A1(\SUMB[17][7] ), .A2(\CARRYB[17][6] ), .ZN(n212) );
  INV_X4 U637 ( .A(n212), .ZN(\CARRYB[18][6] ) );
  XNOR2_X2 U638 ( .A(\CARRYB[17][6] ), .B(\SUMB[17][7] ), .ZN(n213) );
  INV_X4 U639 ( .A(n213), .ZN(\SUMB[18][6] ) );
  NAND2_X2 U640 ( .A1(\SUMB[17][6] ), .A2(\CARRYB[17][5] ), .ZN(n214) );
  INV_X4 U641 ( .A(n214), .ZN(\CARRYB[18][5] ) );
  XNOR2_X2 U642 ( .A(\CARRYB[17][5] ), .B(\SUMB[17][6] ), .ZN(n215) );
  INV_X4 U643 ( .A(n215), .ZN(\SUMB[18][5] ) );
  NAND2_X2 U644 ( .A1(\SUMB[17][5] ), .A2(\CARRYB[17][4] ), .ZN(n216) );
  INV_X4 U645 ( .A(n216), .ZN(\CARRYB[18][4] ) );
  XNOR2_X2 U646 ( .A(\CARRYB[17][4] ), .B(\SUMB[17][5] ), .ZN(n217) );
  INV_X4 U647 ( .A(n217), .ZN(\SUMB[18][4] ) );
  NAND2_X2 U648 ( .A1(\SUMB[17][4] ), .A2(\CARRYB[17][3] ), .ZN(n218) );
  INV_X4 U649 ( .A(n218), .ZN(\CARRYB[18][3] ) );
  XNOR2_X2 U650 ( .A(\CARRYB[17][3] ), .B(\SUMB[17][4] ), .ZN(n219) );
  INV_X4 U651 ( .A(n219), .ZN(\SUMB[18][3] ) );
  NAND2_X2 U652 ( .A1(\SUMB[17][3] ), .A2(\CARRYB[17][2] ), .ZN(n220) );
  INV_X4 U653 ( .A(n220), .ZN(\CARRYB[18][2] ) );
  XNOR2_X2 U654 ( .A(\CARRYB[17][2] ), .B(\SUMB[17][3] ), .ZN(n221) );
  INV_X4 U655 ( .A(n221), .ZN(\SUMB[18][2] ) );
  NAND2_X2 U656 ( .A1(\SUMB[17][2] ), .A2(\CARRYB[17][1] ), .ZN(n222) );
  INV_X4 U657 ( .A(n222), .ZN(\CARRYB[18][1] ) );
  XNOR2_X2 U658 ( .A(\CARRYB[17][1] ), .B(\SUMB[17][2] ), .ZN(n223) );
  INV_X4 U659 ( .A(n223), .ZN(\SUMB[18][1] ) );
  NAND2_X2 U660 ( .A1(\SUMB[17][13] ), .A2(\CARRYB[17][12] ), .ZN(n224) );
  INV_X4 U661 ( .A(n224), .ZN(\CARRYB[18][12] ) );
  XNOR2_X2 U662 ( .A(\CARRYB[17][12] ), .B(\SUMB[17][13] ), .ZN(n225) );
  INV_X4 U663 ( .A(n225), .ZN(\SUMB[18][12] ) );
  NAND2_X2 U664 ( .A1(\SUMB[17][12] ), .A2(\CARRYB[17][11] ), .ZN(n226) );
  INV_X4 U665 ( .A(n226), .ZN(\CARRYB[18][11] ) );
  XNOR2_X2 U666 ( .A(\CARRYB[17][11] ), .B(\SUMB[17][12] ), .ZN(n227) );
  INV_X4 U667 ( .A(n227), .ZN(\SUMB[18][11] ) );
  NAND2_X2 U668 ( .A1(\SUMB[17][11] ), .A2(\CARRYB[17][10] ), .ZN(n228) );
  INV_X4 U669 ( .A(n228), .ZN(\CARRYB[18][10] ) );
  XNOR2_X2 U670 ( .A(\CARRYB[17][10] ), .B(\SUMB[17][11] ), .ZN(n229) );
  INV_X4 U671 ( .A(n229), .ZN(\SUMB[18][10] ) );
  NAND2_X2 U672 ( .A1(\SUMB[17][1] ), .A2(\CARRYB[17][0] ), .ZN(n230) );
  INV_X4 U673 ( .A(n230), .ZN(\CARRYB[18][0] ) );
  XNOR2_X2 U674 ( .A(\CARRYB[17][0] ), .B(\SUMB[17][1] ), .ZN(n231) );
  INV_X4 U675 ( .A(n231), .ZN(PRODUCT[18]) );
  NAND2_X2 U676 ( .A1(\SUMB[17][10] ), .A2(\CARRYB[17][9] ), .ZN(n232) );
  INV_X4 U677 ( .A(n232), .ZN(\CARRYB[18][9] ) );
  XNOR2_X2 U678 ( .A(\CARRYB[17][9] ), .B(\SUMB[17][10] ), .ZN(n233) );
  INV_X4 U679 ( .A(n233), .ZN(\SUMB[18][9] ) );
  NAND2_X2 U680 ( .A1(\SUMB[18][9] ), .A2(\CARRYB[18][8] ), .ZN(n234) );
  INV_X4 U681 ( .A(n234), .ZN(\CARRYB[19][8] ) );
  XNOR2_X2 U682 ( .A(\CARRYB[18][8] ), .B(\SUMB[18][9] ), .ZN(n235) );
  INV_X4 U683 ( .A(n235), .ZN(\SUMB[19][8] ) );
  NAND2_X2 U684 ( .A1(\SUMB[18][8] ), .A2(\CARRYB[18][7] ), .ZN(n236) );
  INV_X4 U685 ( .A(n236), .ZN(\CARRYB[19][7] ) );
  XNOR2_X2 U686 ( .A(\CARRYB[18][7] ), .B(\SUMB[18][8] ), .ZN(n237) );
  INV_X4 U687 ( .A(n237), .ZN(\SUMB[19][7] ) );
  NAND2_X2 U688 ( .A1(\SUMB[18][7] ), .A2(\CARRYB[18][6] ), .ZN(n238) );
  INV_X4 U689 ( .A(n238), .ZN(\CARRYB[19][6] ) );
  XNOR2_X2 U690 ( .A(\CARRYB[18][6] ), .B(\SUMB[18][7] ), .ZN(n239) );
  INV_X4 U691 ( .A(n239), .ZN(\SUMB[19][6] ) );
  NAND2_X2 U692 ( .A1(\SUMB[18][6] ), .A2(\CARRYB[18][5] ), .ZN(n240) );
  INV_X4 U693 ( .A(n240), .ZN(\CARRYB[19][5] ) );
  XNOR2_X2 U694 ( .A(\CARRYB[18][5] ), .B(\SUMB[18][6] ), .ZN(n241) );
  INV_X4 U695 ( .A(n241), .ZN(\SUMB[19][5] ) );
  NAND2_X2 U696 ( .A1(\SUMB[18][5] ), .A2(\CARRYB[18][4] ), .ZN(n242) );
  INV_X4 U697 ( .A(n242), .ZN(\CARRYB[19][4] ) );
  XNOR2_X2 U698 ( .A(\CARRYB[18][4] ), .B(\SUMB[18][5] ), .ZN(n243) );
  INV_X4 U699 ( .A(n243), .ZN(\SUMB[19][4] ) );
  NAND2_X2 U700 ( .A1(\SUMB[18][4] ), .A2(\CARRYB[18][3] ), .ZN(n244) );
  INV_X4 U701 ( .A(n244), .ZN(\CARRYB[19][3] ) );
  XNOR2_X2 U702 ( .A(\CARRYB[18][3] ), .B(\SUMB[18][4] ), .ZN(n245) );
  INV_X4 U703 ( .A(n245), .ZN(\SUMB[19][3] ) );
  NAND2_X2 U704 ( .A1(\SUMB[18][3] ), .A2(\CARRYB[18][2] ), .ZN(n246) );
  INV_X4 U705 ( .A(n246), .ZN(\CARRYB[19][2] ) );
  XNOR2_X2 U706 ( .A(\CARRYB[18][2] ), .B(\SUMB[18][3] ), .ZN(n247) );
  INV_X4 U707 ( .A(n247), .ZN(\SUMB[19][2] ) );
  NAND2_X2 U708 ( .A1(\SUMB[18][2] ), .A2(\CARRYB[18][1] ), .ZN(n248) );
  INV_X4 U709 ( .A(n248), .ZN(\CARRYB[19][1] ) );
  XNOR2_X2 U710 ( .A(\CARRYB[18][1] ), .B(\SUMB[18][2] ), .ZN(n249) );
  INV_X4 U711 ( .A(n249), .ZN(\SUMB[19][1] ) );
  NAND2_X2 U712 ( .A1(\SUMB[18][12] ), .A2(\CARRYB[18][11] ), .ZN(n250) );
  INV_X4 U713 ( .A(n250), .ZN(\CARRYB[19][11] ) );
  XNOR2_X2 U714 ( .A(\CARRYB[18][11] ), .B(\SUMB[18][12] ), .ZN(n251) );
  INV_X4 U715 ( .A(n251), .ZN(\SUMB[19][11] ) );
  NAND2_X2 U716 ( .A1(\SUMB[18][11] ), .A2(\CARRYB[18][10] ), .ZN(n252) );
  INV_X4 U717 ( .A(n252), .ZN(\CARRYB[19][10] ) );
  XNOR2_X2 U718 ( .A(\CARRYB[18][10] ), .B(\SUMB[18][11] ), .ZN(n253) );
  INV_X4 U719 ( .A(n253), .ZN(\SUMB[19][10] ) );
  NAND2_X2 U720 ( .A1(\SUMB[18][1] ), .A2(\CARRYB[18][0] ), .ZN(n254) );
  INV_X4 U721 ( .A(n254), .ZN(\CARRYB[19][0] ) );
  XNOR2_X2 U722 ( .A(\CARRYB[18][0] ), .B(\SUMB[18][1] ), .ZN(n255) );
  INV_X4 U723 ( .A(n255), .ZN(PRODUCT[19]) );
  NAND2_X2 U724 ( .A1(\SUMB[18][10] ), .A2(\CARRYB[18][9] ), .ZN(n256) );
  INV_X4 U725 ( .A(n256), .ZN(\CARRYB[19][9] ) );
  XNOR2_X2 U726 ( .A(\CARRYB[18][9] ), .B(\SUMB[18][10] ), .ZN(n257) );
  INV_X4 U727 ( .A(n257), .ZN(\SUMB[19][9] ) );
  NAND2_X2 U728 ( .A1(\SUMB[19][9] ), .A2(\CARRYB[19][8] ), .ZN(n258) );
  INV_X4 U729 ( .A(n258), .ZN(\CARRYB[20][8] ) );
  XNOR2_X2 U730 ( .A(\CARRYB[19][8] ), .B(\SUMB[19][9] ), .ZN(n259) );
  INV_X4 U731 ( .A(n259), .ZN(\SUMB[20][8] ) );
  NAND2_X2 U732 ( .A1(\SUMB[19][8] ), .A2(\CARRYB[19][7] ), .ZN(n260) );
  INV_X4 U733 ( .A(n260), .ZN(\CARRYB[20][7] ) );
  XNOR2_X2 U734 ( .A(\CARRYB[19][7] ), .B(\SUMB[19][8] ), .ZN(n261) );
  INV_X4 U735 ( .A(n261), .ZN(\SUMB[20][7] ) );
  NAND2_X2 U736 ( .A1(\SUMB[19][7] ), .A2(\CARRYB[19][6] ), .ZN(n262) );
  INV_X4 U737 ( .A(n262), .ZN(\CARRYB[20][6] ) );
  XNOR2_X2 U738 ( .A(\CARRYB[19][6] ), .B(\SUMB[19][7] ), .ZN(n263) );
  INV_X4 U739 ( .A(n263), .ZN(\SUMB[20][6] ) );
  NAND2_X2 U740 ( .A1(\SUMB[19][6] ), .A2(\CARRYB[19][5] ), .ZN(n264) );
  INV_X4 U741 ( .A(n264), .ZN(\CARRYB[20][5] ) );
  XNOR2_X2 U742 ( .A(\CARRYB[19][5] ), .B(\SUMB[19][6] ), .ZN(n265) );
  INV_X4 U743 ( .A(n265), .ZN(\SUMB[20][5] ) );
  NAND2_X2 U744 ( .A1(\SUMB[19][5] ), .A2(\CARRYB[19][4] ), .ZN(n266) );
  INV_X4 U745 ( .A(n266), .ZN(\CARRYB[20][4] ) );
  XNOR2_X2 U746 ( .A(\CARRYB[19][4] ), .B(\SUMB[19][5] ), .ZN(n267) );
  INV_X4 U747 ( .A(n267), .ZN(\SUMB[20][4] ) );
  NAND2_X2 U748 ( .A1(\SUMB[19][4] ), .A2(\CARRYB[19][3] ), .ZN(n268) );
  INV_X4 U749 ( .A(n268), .ZN(\CARRYB[20][3] ) );
  XNOR2_X2 U750 ( .A(\CARRYB[19][3] ), .B(\SUMB[19][4] ), .ZN(n269) );
  INV_X4 U751 ( .A(n269), .ZN(\SUMB[20][3] ) );
  NAND2_X2 U752 ( .A1(\SUMB[19][3] ), .A2(\CARRYB[19][2] ), .ZN(n270) );
  INV_X4 U753 ( .A(n270), .ZN(\CARRYB[20][2] ) );
  XNOR2_X2 U754 ( .A(\CARRYB[19][2] ), .B(\SUMB[19][3] ), .ZN(n271) );
  INV_X4 U755 ( .A(n271), .ZN(\SUMB[20][2] ) );
  NAND2_X2 U756 ( .A1(\SUMB[19][2] ), .A2(\CARRYB[19][1] ), .ZN(n272) );
  INV_X4 U757 ( .A(n272), .ZN(\CARRYB[20][1] ) );
  XNOR2_X2 U758 ( .A(\CARRYB[19][1] ), .B(\SUMB[19][2] ), .ZN(n273) );
  INV_X4 U759 ( .A(n273), .ZN(\SUMB[20][1] ) );
  NAND2_X2 U760 ( .A1(\SUMB[19][11] ), .A2(\CARRYB[19][10] ), .ZN(n274) );
  INV_X4 U761 ( .A(n274), .ZN(\CARRYB[20][10] ) );
  XNOR2_X2 U762 ( .A(\CARRYB[19][10] ), .B(\SUMB[19][11] ), .ZN(n275) );
  INV_X4 U763 ( .A(n275), .ZN(\SUMB[20][10] ) );
  NAND2_X2 U764 ( .A1(\SUMB[19][1] ), .A2(\CARRYB[19][0] ), .ZN(n276) );
  INV_X4 U765 ( .A(n276), .ZN(\CARRYB[20][0] ) );
  XNOR2_X2 U766 ( .A(\CARRYB[19][0] ), .B(\SUMB[19][1] ), .ZN(n277) );
  INV_X4 U767 ( .A(n277), .ZN(PRODUCT[20]) );
  NAND2_X2 U768 ( .A1(\SUMB[19][10] ), .A2(\CARRYB[19][9] ), .ZN(n278) );
  INV_X4 U769 ( .A(n278), .ZN(\CARRYB[20][9] ) );
  XNOR2_X2 U770 ( .A(\CARRYB[19][9] ), .B(\SUMB[19][10] ), .ZN(n279) );
  INV_X4 U771 ( .A(n279), .ZN(\SUMB[20][9] ) );
  NAND2_X2 U772 ( .A1(\SUMB[20][9] ), .A2(\CARRYB[20][8] ), .ZN(n280) );
  INV_X4 U773 ( .A(n280), .ZN(\CARRYB[21][8] ) );
  XNOR2_X2 U774 ( .A(\CARRYB[20][8] ), .B(\SUMB[20][9] ), .ZN(n281) );
  INV_X4 U775 ( .A(n281), .ZN(\SUMB[21][8] ) );
  NAND2_X2 U776 ( .A1(\SUMB[20][8] ), .A2(\CARRYB[20][7] ), .ZN(n282) );
  INV_X4 U777 ( .A(n282), .ZN(\CARRYB[21][7] ) );
  XNOR2_X2 U778 ( .A(\CARRYB[20][7] ), .B(\SUMB[20][8] ), .ZN(n283) );
  INV_X4 U779 ( .A(n283), .ZN(\SUMB[21][7] ) );
  NAND2_X2 U780 ( .A1(\SUMB[20][7] ), .A2(\CARRYB[20][6] ), .ZN(n284) );
  INV_X4 U781 ( .A(n284), .ZN(\CARRYB[21][6] ) );
  XNOR2_X2 U782 ( .A(\CARRYB[20][6] ), .B(\SUMB[20][7] ), .ZN(n285) );
  INV_X4 U783 ( .A(n285), .ZN(\SUMB[21][6] ) );
  NAND2_X2 U784 ( .A1(\SUMB[20][6] ), .A2(\CARRYB[20][5] ), .ZN(n286) );
  INV_X4 U785 ( .A(n286), .ZN(\CARRYB[21][5] ) );
  XNOR2_X2 U786 ( .A(\CARRYB[20][5] ), .B(\SUMB[20][6] ), .ZN(n287) );
  INV_X4 U787 ( .A(n287), .ZN(\SUMB[21][5] ) );
  NAND2_X2 U788 ( .A1(\SUMB[20][5] ), .A2(\CARRYB[20][4] ), .ZN(n288) );
  INV_X4 U789 ( .A(n288), .ZN(\CARRYB[21][4] ) );
  XNOR2_X2 U790 ( .A(\CARRYB[20][4] ), .B(\SUMB[20][5] ), .ZN(n289) );
  INV_X4 U791 ( .A(n289), .ZN(\SUMB[21][4] ) );
  NAND2_X2 U792 ( .A1(\SUMB[20][4] ), .A2(\CARRYB[20][3] ), .ZN(n290) );
  INV_X4 U793 ( .A(n290), .ZN(\CARRYB[21][3] ) );
  XNOR2_X2 U794 ( .A(\CARRYB[20][3] ), .B(\SUMB[20][4] ), .ZN(n291) );
  INV_X4 U795 ( .A(n291), .ZN(\SUMB[21][3] ) );
  NAND2_X2 U796 ( .A1(\SUMB[20][3] ), .A2(\CARRYB[20][2] ), .ZN(n292) );
  INV_X4 U797 ( .A(n292), .ZN(\CARRYB[21][2] ) );
  XNOR2_X2 U798 ( .A(\CARRYB[20][2] ), .B(\SUMB[20][3] ), .ZN(n293) );
  INV_X4 U799 ( .A(n293), .ZN(\SUMB[21][2] ) );
  NAND2_X2 U800 ( .A1(\SUMB[20][2] ), .A2(\CARRYB[20][1] ), .ZN(n294) );
  INV_X4 U801 ( .A(n294), .ZN(\CARRYB[21][1] ) );
  XNOR2_X2 U802 ( .A(\CARRYB[20][1] ), .B(\SUMB[20][2] ), .ZN(n295) );
  INV_X4 U803 ( .A(n295), .ZN(\SUMB[21][1] ) );
  NAND2_X2 U804 ( .A1(\SUMB[20][1] ), .A2(\CARRYB[20][0] ), .ZN(n296) );
  INV_X4 U805 ( .A(n296), .ZN(\CARRYB[21][0] ) );
  XNOR2_X2 U806 ( .A(\CARRYB[20][0] ), .B(\SUMB[20][1] ), .ZN(n297) );
  INV_X4 U807 ( .A(n297), .ZN(PRODUCT[21]) );
  NAND2_X2 U808 ( .A1(\SUMB[20][10] ), .A2(\CARRYB[20][9] ), .ZN(n298) );
  INV_X4 U809 ( .A(n298), .ZN(\CARRYB[21][9] ) );
  XNOR2_X2 U810 ( .A(\CARRYB[20][9] ), .B(\SUMB[20][10] ), .ZN(n299) );
  INV_X4 U811 ( .A(n299), .ZN(\SUMB[21][9] ) );
endmodule


module multiplier_DW01_add_5 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70;

  OR2_X4 U2 ( .A1(B[15]), .A2(A[15]), .ZN(n1) );
  AND2_X4 U3 ( .A1(n1), .A2(n70), .ZN(SUM[15]) );
  INV_X4 U4 ( .A(B[29]), .ZN(n3) );
  INV_X4 U5 ( .A(n21), .ZN(n4) );
  INV_X4 U6 ( .A(n23), .ZN(n5) );
  INV_X4 U7 ( .A(n29), .ZN(n6) );
  INV_X4 U8 ( .A(n31), .ZN(n7) );
  INV_X4 U9 ( .A(n37), .ZN(n8) );
  INV_X4 U10 ( .A(n39), .ZN(n9) );
  INV_X4 U11 ( .A(n45), .ZN(n10) );
  INV_X4 U12 ( .A(n47), .ZN(n11) );
  INV_X4 U13 ( .A(n53), .ZN(n12) );
  INV_X4 U14 ( .A(n55), .ZN(n13) );
  INV_X4 U15 ( .A(n61), .ZN(n14) );
  INV_X4 U16 ( .A(n63), .ZN(n15) );
  INV_X4 U17 ( .A(n68), .ZN(n16) );
  INV_X4 U18 ( .A(n70), .ZN(n17) );
  XOR2_X1 U19 ( .A(n3), .B(n18), .Z(SUM[29]) );
  AOI21_X1 U20 ( .B1(n19), .B2(n4), .A(n20), .ZN(n18) );
  XOR2_X1 U21 ( .A(n19), .B(n22), .Z(SUM[28]) );
  NOR2_X1 U22 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U23 ( .A1(B[28]), .A2(A[28]), .ZN(n21) );
  AND2_X1 U24 ( .A1(B[28]), .A2(A[28]), .ZN(n20) );
  OAI21_X1 U25 ( .B1(n23), .B2(n24), .A(n25), .ZN(n19) );
  XOR2_X1 U26 ( .A(n26), .B(n24), .Z(SUM[27]) );
  AOI21_X1 U27 ( .B1(n6), .B2(n27), .A(n28), .ZN(n24) );
  NAND2_X1 U28 ( .A1(n5), .A2(n25), .ZN(n26) );
  NAND2_X1 U29 ( .A1(B[27]), .A2(A[27]), .ZN(n25) );
  NOR2_X1 U30 ( .A1(B[27]), .A2(A[27]), .ZN(n23) );
  XOR2_X1 U31 ( .A(n27), .B(n30), .Z(SUM[26]) );
  NOR2_X1 U32 ( .A1(n28), .A2(n29), .ZN(n30) );
  NOR2_X1 U33 ( .A1(B[26]), .A2(A[26]), .ZN(n29) );
  AND2_X1 U34 ( .A1(B[26]), .A2(A[26]), .ZN(n28) );
  OAI21_X1 U35 ( .B1(n31), .B2(n32), .A(n33), .ZN(n27) );
  XOR2_X1 U36 ( .A(n34), .B(n32), .Z(SUM[25]) );
  AOI21_X1 U37 ( .B1(n8), .B2(n35), .A(n36), .ZN(n32) );
  NAND2_X1 U38 ( .A1(n7), .A2(n33), .ZN(n34) );
  NAND2_X1 U39 ( .A1(B[25]), .A2(A[25]), .ZN(n33) );
  NOR2_X1 U40 ( .A1(B[25]), .A2(A[25]), .ZN(n31) );
  XOR2_X1 U41 ( .A(n35), .B(n38), .Z(SUM[24]) );
  NOR2_X1 U42 ( .A1(n36), .A2(n37), .ZN(n38) );
  NOR2_X1 U43 ( .A1(B[24]), .A2(A[24]), .ZN(n37) );
  AND2_X1 U44 ( .A1(B[24]), .A2(A[24]), .ZN(n36) );
  OAI21_X1 U45 ( .B1(n39), .B2(n40), .A(n41), .ZN(n35) );
  XOR2_X1 U46 ( .A(n42), .B(n40), .Z(SUM[23]) );
  AOI21_X1 U47 ( .B1(n10), .B2(n43), .A(n44), .ZN(n40) );
  NAND2_X1 U48 ( .A1(n9), .A2(n41), .ZN(n42) );
  NAND2_X1 U49 ( .A1(B[23]), .A2(A[23]), .ZN(n41) );
  NOR2_X1 U50 ( .A1(B[23]), .A2(A[23]), .ZN(n39) );
  XOR2_X1 U51 ( .A(n43), .B(n46), .Z(SUM[22]) );
  NOR2_X1 U52 ( .A1(n44), .A2(n45), .ZN(n46) );
  NOR2_X1 U53 ( .A1(B[22]), .A2(A[22]), .ZN(n45) );
  AND2_X1 U54 ( .A1(B[22]), .A2(A[22]), .ZN(n44) );
  OAI21_X1 U55 ( .B1(n47), .B2(n48), .A(n49), .ZN(n43) );
  XOR2_X1 U56 ( .A(n50), .B(n48), .Z(SUM[21]) );
  AOI21_X1 U57 ( .B1(n12), .B2(n51), .A(n52), .ZN(n48) );
  NAND2_X1 U58 ( .A1(n11), .A2(n49), .ZN(n50) );
  NAND2_X1 U59 ( .A1(B[21]), .A2(A[21]), .ZN(n49) );
  NOR2_X1 U60 ( .A1(B[21]), .A2(A[21]), .ZN(n47) );
  XOR2_X1 U61 ( .A(n51), .B(n54), .Z(SUM[20]) );
  NOR2_X1 U62 ( .A1(n52), .A2(n53), .ZN(n54) );
  NOR2_X1 U63 ( .A1(B[20]), .A2(A[20]), .ZN(n53) );
  AND2_X1 U64 ( .A1(B[20]), .A2(A[20]), .ZN(n52) );
  OAI21_X1 U65 ( .B1(n55), .B2(n56), .A(n57), .ZN(n51) );
  XOR2_X1 U66 ( .A(n58), .B(n56), .Z(SUM[19]) );
  AOI21_X1 U67 ( .B1(n14), .B2(n59), .A(n60), .ZN(n56) );
  NAND2_X1 U68 ( .A1(n13), .A2(n57), .ZN(n58) );
  NAND2_X1 U69 ( .A1(B[19]), .A2(A[19]), .ZN(n57) );
  NOR2_X1 U70 ( .A1(B[19]), .A2(A[19]), .ZN(n55) );
  XOR2_X1 U71 ( .A(n59), .B(n62), .Z(SUM[18]) );
  NOR2_X1 U72 ( .A1(n60), .A2(n61), .ZN(n62) );
  NOR2_X1 U73 ( .A1(B[18]), .A2(A[18]), .ZN(n61) );
  AND2_X1 U74 ( .A1(B[18]), .A2(A[18]), .ZN(n60) );
  OAI21_X1 U75 ( .B1(n63), .B2(n64), .A(n65), .ZN(n59) );
  XOR2_X1 U76 ( .A(n66), .B(n64), .Z(SUM[17]) );
  AOI21_X1 U77 ( .B1(n16), .B2(n17), .A(n67), .ZN(n64) );
  NAND2_X1 U78 ( .A1(n15), .A2(n65), .ZN(n66) );
  NAND2_X1 U79 ( .A1(B[17]), .A2(A[17]), .ZN(n65) );
  NOR2_X1 U80 ( .A1(B[17]), .A2(A[17]), .ZN(n63) );
  XOR2_X1 U81 ( .A(n17), .B(n69), .Z(SUM[16]) );
  NOR2_X1 U82 ( .A1(n67), .A2(n68), .ZN(n69) );
  NOR2_X1 U83 ( .A1(B[16]), .A2(A[16]), .ZN(n68) );
  AND2_X1 U84 ( .A1(B[16]), .A2(A[16]), .ZN(n67) );
  NAND2_X1 U85 ( .A1(B[15]), .A2(A[15]), .ZN(n70) );
  BUF_X32 U86 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X32 U87 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X32 U88 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X32 U89 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X32 U90 ( .A(A[4]), .Z(SUM[4]) );
  BUF_X32 U91 ( .A(A[5]), .Z(SUM[5]) );
  BUF_X32 U92 ( .A(A[6]), .Z(SUM[6]) );
  BUF_X32 U93 ( .A(A[7]), .Z(SUM[7]) );
  BUF_X32 U94 ( .A(A[8]), .Z(SUM[8]) );
  BUF_X32 U95 ( .A(A[9]), .Z(SUM[9]) );
  BUF_X32 U96 ( .A(A[10]), .Z(SUM[10]) );
  BUF_X32 U97 ( .A(A[11]), .Z(SUM[11]) );
  BUF_X32 U98 ( .A(A[12]), .Z(SUM[12]) );
  BUF_X32 U99 ( .A(A[13]), .Z(SUM[13]) );
  BUF_X32 U100 ( .A(A[14]), .Z(SUM[14]) );
endmodule


module multiplier_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [15:0] A;
  input [15:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] ,
         \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] ,
         \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] ,
         \ab[15][0] , \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] ,
         \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] ,
         \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][15] , \ab[13][14] , \ab[13][13] ,
         \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] ,
         \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] ,
         \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][15] , \ab[12][14] ,
         \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] ,
         \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] ,
         \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][15] ,
         \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] ,
         \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] ,
         \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] ,
         \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] ,
         \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][15] , \ab[8][14] , \ab[8][13] ,
         \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][15] , \ab[7][14] ,
         \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] , \ab[7][9] ,
         \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] ,
         \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][15] ,
         \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] ,
         \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] ,
         \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][15] , \ab[3][14] , \ab[3][13] ,
         \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][15] , \ab[2][14] ,
         \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] , \ab[2][9] ,
         \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] ,
         \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][15] ,
         \ab[1][14] , \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] ,
         \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] ,
         \ab[0][15] , \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] ,
         \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] ,
         \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] ,
         \CARRYB[15][14] , \CARRYB[15][13] , \CARRYB[15][12] ,
         \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] ,
         \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] ,
         \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] ,
         \CARRYB[14][14] , \CARRYB[14][13] , \CARRYB[14][12] ,
         \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] ,
         \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] ,
         \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][14] , \CARRYB[12][13] , \CARRYB[12][12] ,
         \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] ,
         \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] ,
         \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] ,
         \CARRYB[11][14] , \CARRYB[11][13] , \CARRYB[11][12] ,
         \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] ,
         \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] ,
         \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] ,
         \CARRYB[10][14] , \CARRYB[10][13] , \CARRYB[10][12] ,
         \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] ,
         \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] ,
         \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] ,
         \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] ,
         \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] ,
         \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][14] ,
         \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] ,
         \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] ,
         \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] ,
         \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] ,
         \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] ,
         \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] ,
         \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] ,
         \CARRYB[5][14] , \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] ,
         \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] ,
         \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] ,
         \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][14] ,
         \CARRYB[4][13] , \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] ,
         \CARRYB[4][9] , \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] ,
         \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] ,
         \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][14] , \CARRYB[3][13] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] ,
         \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] ,
         \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] ,
         \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[15][0] , \SUMB[14][14] ,
         \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] ,
         \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] ,
         \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] ,
         \SUMB[14][1] , \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] ,
         \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] ,
         \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] ,
         \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] ,
         \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] ,
         \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] ,
         \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][14] , \SUMB[8][13] ,
         \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] ,
         \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] ,
         \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \A1[12] ,
         \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] ,
         \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] , n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94;

  FA_X1 S4_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), .CO(
        \CARRYB[15][0] ), .S(\SUMB[15][0] ) );
  FA_X1 S4_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), .CO(
        \CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA_X1 S4_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), .CO(
        \CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA_X1 S4_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), .CO(
        \CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA_X1 S4_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), .CO(
        \CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA_X1 S4_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), .CO(
        \CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA_X1 S4_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), .CO(
        \CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA_X1 S4_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), .CO(
        \CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA_X1 S4_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), .CO(
        \CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA_X1 S4_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), .CO(
        \CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA_X1 S4_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA_X1 S4_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA_X1 S4_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA_X1 S4_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA_X1 S5_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\ab[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA_X1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FA_X1 S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA_X1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA_X1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA_X1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA_X1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA_X1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA_X1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA_X1 S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA_X1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA_X1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA_X1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA_X1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA_X1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA_X1 S3_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\ab[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA_X1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA_X1 S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA_X1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA_X1 S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA_X1 S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA_X1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA_X1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA_X1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA_X1 S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA_X1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA_X1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA_X1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA_X1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA_X1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA_X1 S3_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\ab[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA_X1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA_X1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA_X1 S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA_X1 S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA_X1 S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA_X1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA_X1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA_X1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA_X1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA_X1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA_X1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA_X1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA_X1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA_X1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA_X1 S3_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\ab[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA_X1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA_X1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA_X1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA_X1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA_X1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA_X1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA_X1 S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA_X1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA_X1 S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA_X1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA_X1 S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA_X1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA_X1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA_X1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA_X1 S3_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\ab[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA_X1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA_X1 S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA_X1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA_X1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA_X1 S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA_X1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA_X1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA_X1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA_X1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA_X1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA_X1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA_X1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA_X1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA_X1 S3_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\ab[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA_X1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA_X1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA_X1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA_X1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA_X1 S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA_X1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA_X1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA_X1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA_X1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA_X1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA_X1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA_X1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA_X1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA_X1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA_X1 S3_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\ab[8][15] ), .CO(
        \CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA_X1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA_X1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA_X1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA_X1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA_X1 S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA_X1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA_X1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA_X1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA_X1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA_X1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA_X1 S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA_X1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA_X1 S3_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\ab[7][15] ), .CO(
        \CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA_X1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA_X1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA_X1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA_X1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA_X1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA_X1 S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA_X1 S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA_X1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA_X1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA_X1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA_X1 S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA_X1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA_X1 S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA_X1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA_X1 S3_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\ab[6][15] ), .CO(
        \CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA_X1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA_X1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA_X1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA_X1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA_X1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA_X1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA_X1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA_X1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA_X1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA_X1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA_X1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA_X1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA_X1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA_X1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA_X1 S3_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\ab[5][15] ), .CO(
        \CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA_X1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA_X1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA_X1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA_X1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA_X1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA_X1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA_X1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA_X1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA_X1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA_X1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA_X1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA_X1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA_X1 S3_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\ab[4][15] ), .CO(
        \CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA_X1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA_X1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA_X1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA_X1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA_X1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA_X1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA_X1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA_X1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA_X1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA_X1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA_X1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA_X1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA_X1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA_X1 S3_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\ab[3][15] ), .CO(
        \CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA_X1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA_X1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA_X1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA_X1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA_X1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA_X1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA_X1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA_X1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA_X1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA_X1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA_X1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA_X1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA_X1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA_X1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA_X1 S3_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\ab[2][15] ), .CO(
        \CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(n16), .CI(n45), .CO(\CARRYB[2][0] ), .S(
        \A1[0] ) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(n15), .CI(n44), .CO(\CARRYB[2][1] ), .S(
        \SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(n14), .CI(n43), .CO(\CARRYB[2][2] ), .S(
        \SUMB[2][2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2][3] ), .B(n13), .CI(n42), .CO(\CARRYB[2][3] ), .S(
        \SUMB[2][3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2][4] ), .B(n12), .CI(n41), .CO(\CARRYB[2][4] ), .S(
        \SUMB[2][4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2][5] ), .B(n11), .CI(n40), .CO(\CARRYB[2][5] ), .S(
        \SUMB[2][5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2][6] ), .B(n10), .CI(n39), .CO(\CARRYB[2][6] ), .S(
        \SUMB[2][6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(n9), .CI(n38), .CO(\CARRYB[2][7] ), .S(
        \SUMB[2][7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(n8), .CI(n37), .CO(\CARRYB[2][8] ), .S(
        \SUMB[2][8] ) );
  FA_X1 S2_2_9 ( .A(\ab[2][9] ), .B(n7), .CI(n36), .CO(\CARRYB[2][9] ), .S(
        \SUMB[2][9] ) );
  FA_X1 S2_2_10 ( .A(\ab[2][10] ), .B(n6), .CI(n35), .CO(\CARRYB[2][10] ), .S(
        \SUMB[2][10] ) );
  FA_X1 S2_2_11 ( .A(\ab[2][11] ), .B(n5), .CI(n34), .CO(\CARRYB[2][11] ), .S(
        \SUMB[2][11] ) );
  FA_X1 S2_2_12 ( .A(\ab[2][12] ), .B(n4), .CI(n33), .CO(\CARRYB[2][12] ), .S(
        \SUMB[2][12] ) );
  FA_X1 S2_2_13 ( .A(\ab[2][13] ), .B(n3), .CI(n32), .CO(\CARRYB[2][13] ), .S(
        \SUMB[2][13] ) );
  FA_X1 S3_2_14 ( .A(\ab[2][14] ), .B(n31), .CI(\ab[1][15] ), .CO(
        \CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  AND2_X4 U2 ( .A1(\ab[0][14] ), .A2(\ab[1][13] ), .ZN(n3) );
  AND2_X4 U3 ( .A1(\ab[0][13] ), .A2(\ab[1][12] ), .ZN(n4) );
  AND2_X4 U4 ( .A1(\ab[0][12] ), .A2(\ab[1][11] ), .ZN(n5) );
  AND2_X4 U5 ( .A1(\ab[0][11] ), .A2(\ab[1][10] ), .ZN(n6) );
  AND2_X4 U6 ( .A1(\ab[0][10] ), .A2(\ab[1][9] ), .ZN(n7) );
  AND2_X4 U7 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .ZN(n8) );
  AND2_X4 U8 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .ZN(n9) );
  AND2_X4 U9 ( .A1(\ab[0][7] ), .A2(\ab[1][6] ), .ZN(n10) );
  AND2_X4 U10 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .ZN(n11) );
  AND2_X4 U11 ( .A1(\ab[0][5] ), .A2(\ab[1][4] ), .ZN(n12) );
  AND2_X4 U12 ( .A1(\ab[0][4] ), .A2(\ab[1][3] ), .ZN(n13) );
  AND2_X4 U13 ( .A1(\ab[0][3] ), .A2(\ab[1][2] ), .ZN(n14) );
  AND2_X4 U14 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .ZN(n15) );
  AND2_X4 U15 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .ZN(n16) );
  XOR2_X2 U16 ( .A(\CARRYB[15][14] ), .B(\ab[15][15] ), .Z(n17) );
  XOR2_X2 U17 ( .A(\CARRYB[15][12] ), .B(\SUMB[15][13] ), .Z(n18) );
  XOR2_X2 U18 ( .A(\CARRYB[15][10] ), .B(\SUMB[15][11] ), .Z(n19) );
  XOR2_X2 U19 ( .A(\CARRYB[15][8] ), .B(\SUMB[15][9] ), .Z(n20) );
  XOR2_X2 U20 ( .A(\CARRYB[15][6] ), .B(\SUMB[15][7] ), .Z(n21) );
  XOR2_X2 U21 ( .A(\CARRYB[15][4] ), .B(\SUMB[15][5] ), .Z(n22) );
  XOR2_X2 U22 ( .A(\CARRYB[15][2] ), .B(\SUMB[15][3] ), .Z(n23) );
  XOR2_X2 U23 ( .A(\CARRYB[15][1] ), .B(\SUMB[15][2] ), .Z(n24) );
  XOR2_X2 U24 ( .A(\CARRYB[15][13] ), .B(\SUMB[15][14] ), .Z(n25) );
  XOR2_X2 U25 ( .A(\CARRYB[15][11] ), .B(\SUMB[15][12] ), .Z(n26) );
  XOR2_X2 U26 ( .A(\CARRYB[15][9] ), .B(\SUMB[15][10] ), .Z(n27) );
  XOR2_X2 U27 ( .A(\CARRYB[15][7] ), .B(\SUMB[15][8] ), .Z(n28) );
  XOR2_X2 U28 ( .A(\CARRYB[15][5] ), .B(\SUMB[15][6] ), .Z(n29) );
  XOR2_X2 U29 ( .A(\CARRYB[15][3] ), .B(\SUMB[15][4] ), .Z(n30) );
  AND2_X4 U30 ( .A1(\ab[0][15] ), .A2(\ab[1][14] ), .ZN(n31) );
  XOR2_X2 U31 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(n32) );
  XOR2_X2 U32 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(n33) );
  XOR2_X2 U33 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(n34) );
  XOR2_X2 U34 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(n35) );
  XOR2_X2 U35 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(n36) );
  XOR2_X2 U36 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(n37) );
  XOR2_X2 U37 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(n38) );
  XOR2_X2 U38 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(n39) );
  XOR2_X2 U39 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(n40) );
  XOR2_X2 U40 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(n41) );
  XOR2_X2 U41 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(n42) );
  XOR2_X2 U42 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(n43) );
  XOR2_X2 U43 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(n44) );
  XOR2_X2 U44 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(n45) );
  XOR2_X2 U45 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  AND2_X4 U46 ( .A1(\CARRYB[15][13] ), .A2(\SUMB[15][14] ), .ZN(n47) );
  AND2_X4 U47 ( .A1(\CARRYB[15][11] ), .A2(\SUMB[15][12] ), .ZN(n48) );
  AND2_X4 U48 ( .A1(\CARRYB[15][9] ), .A2(\SUMB[15][10] ), .ZN(n49) );
  AND2_X4 U49 ( .A1(\CARRYB[15][7] ), .A2(\SUMB[15][8] ), .ZN(n50) );
  AND2_X4 U50 ( .A1(\CARRYB[15][5] ), .A2(\SUMB[15][6] ), .ZN(n51) );
  AND2_X4 U51 ( .A1(\CARRYB[15][3] ), .A2(\SUMB[15][4] ), .ZN(n52) );
  AND2_X4 U52 ( .A1(\CARRYB[15][1] ), .A2(\SUMB[15][2] ), .ZN(n53) );
  AND2_X4 U53 ( .A1(\CARRYB[15][12] ), .A2(\SUMB[15][13] ), .ZN(n54) );
  AND2_X4 U54 ( .A1(\CARRYB[15][10] ), .A2(\SUMB[15][11] ), .ZN(n55) );
  AND2_X4 U55 ( .A1(\CARRYB[15][8] ), .A2(\SUMB[15][9] ), .ZN(n56) );
  AND2_X4 U56 ( .A1(\CARRYB[15][6] ), .A2(\SUMB[15][7] ), .ZN(n57) );
  AND2_X4 U57 ( .A1(\CARRYB[15][4] ), .A2(\SUMB[15][5] ), .ZN(n58) );
  AND2_X4 U58 ( .A1(\CARRYB[15][2] ), .A2(\SUMB[15][3] ), .ZN(n59) );
  AND2_X4 U59 ( .A1(\CARRYB[15][0] ), .A2(\SUMB[15][1] ), .ZN(n60) );
  XOR2_X2 U60 ( .A(\CARRYB[15][0] ), .B(\SUMB[15][1] ), .Z(n61) );
  AND2_X4 U61 ( .A1(\CARRYB[15][14] ), .A2(\ab[15][15] ), .ZN(n62) );
  INV_X4 U62 ( .A(A[9]), .ZN(n69) );
  INV_X4 U63 ( .A(B[8]), .ZN(n86) );
  INV_X4 U64 ( .A(B[7]), .ZN(n87) );
  INV_X4 U65 ( .A(B[1]), .ZN(n93) );
  INV_X4 U66 ( .A(B[2]), .ZN(n92) );
  INV_X4 U67 ( .A(B[3]), .ZN(n91) );
  INV_X4 U68 ( .A(B[4]), .ZN(n90) );
  INV_X4 U69 ( .A(B[5]), .ZN(n89) );
  INV_X4 U70 ( .A(B[6]), .ZN(n88) );
  INV_X4 U71 ( .A(B[10]), .ZN(n84) );
  INV_X4 U72 ( .A(B[9]), .ZN(n85) );
  INV_X4 U73 ( .A(B[12]), .ZN(n82) );
  INV_X4 U74 ( .A(B[11]), .ZN(n83) );
  INV_X4 U75 ( .A(B[14]), .ZN(n80) );
  INV_X4 U76 ( .A(B[13]), .ZN(n81) );
  INV_X4 U77 ( .A(B[15]), .ZN(n79) );
  INV_X4 U78 ( .A(B[0]), .ZN(n94) );
  INV_X4 U79 ( .A(A[0]), .ZN(n78) );
  INV_X4 U80 ( .A(A[1]), .ZN(n77) );
  INV_X4 U81 ( .A(A[3]), .ZN(n75) );
  INV_X4 U82 ( .A(A[4]), .ZN(n74) );
  INV_X4 U83 ( .A(A[5]), .ZN(n73) );
  INV_X4 U84 ( .A(A[6]), .ZN(n72) );
  INV_X4 U85 ( .A(A[7]), .ZN(n71) );
  INV_X4 U86 ( .A(A[8]), .ZN(n70) );
  INV_X4 U87 ( .A(A[10]), .ZN(n68) );
  INV_X4 U88 ( .A(A[11]), .ZN(n67) );
  INV_X4 U89 ( .A(A[12]), .ZN(n66) );
  INV_X4 U90 ( .A(A[13]), .ZN(n65) );
  INV_X4 U91 ( .A(A[14]), .ZN(n64) );
  INV_X4 U92 ( .A(A[15]), .ZN(n63) );
  INV_X4 U93 ( .A(A[2]), .ZN(n76) );
  NOR2_X1 U95 ( .A1(n69), .A2(n85), .ZN(\ab[9][9] ) );
  NOR2_X1 U96 ( .A1(n69), .A2(n86), .ZN(\ab[9][8] ) );
  NOR2_X1 U97 ( .A1(n69), .A2(n87), .ZN(\ab[9][7] ) );
  NOR2_X1 U98 ( .A1(n69), .A2(n88), .ZN(\ab[9][6] ) );
  NOR2_X1 U99 ( .A1(n69), .A2(n89), .ZN(\ab[9][5] ) );
  NOR2_X1 U100 ( .A1(n69), .A2(n90), .ZN(\ab[9][4] ) );
  NOR2_X1 U101 ( .A1(n69), .A2(n91), .ZN(\ab[9][3] ) );
  NOR2_X1 U102 ( .A1(n69), .A2(n92), .ZN(\ab[9][2] ) );
  NOR2_X1 U103 ( .A1(n69), .A2(n93), .ZN(\ab[9][1] ) );
  NOR2_X1 U104 ( .A1(n69), .A2(n79), .ZN(\ab[9][15] ) );
  NOR2_X1 U105 ( .A1(n69), .A2(n80), .ZN(\ab[9][14] ) );
  NOR2_X1 U106 ( .A1(n69), .A2(n81), .ZN(\ab[9][13] ) );
  NOR2_X1 U107 ( .A1(n69), .A2(n82), .ZN(\ab[9][12] ) );
  NOR2_X1 U108 ( .A1(n69), .A2(n83), .ZN(\ab[9][11] ) );
  NOR2_X1 U109 ( .A1(n69), .A2(n84), .ZN(\ab[9][10] ) );
  NOR2_X1 U110 ( .A1(n69), .A2(n94), .ZN(\ab[9][0] ) );
  NOR2_X1 U111 ( .A1(n85), .A2(n70), .ZN(\ab[8][9] ) );
  NOR2_X1 U112 ( .A1(n86), .A2(n70), .ZN(\ab[8][8] ) );
  NOR2_X1 U113 ( .A1(n87), .A2(n70), .ZN(\ab[8][7] ) );
  NOR2_X1 U114 ( .A1(n88), .A2(n70), .ZN(\ab[8][6] ) );
  NOR2_X1 U115 ( .A1(n89), .A2(n70), .ZN(\ab[8][5] ) );
  NOR2_X1 U116 ( .A1(n90), .A2(n70), .ZN(\ab[8][4] ) );
  NOR2_X1 U117 ( .A1(n91), .A2(n70), .ZN(\ab[8][3] ) );
  NOR2_X1 U118 ( .A1(n92), .A2(n70), .ZN(\ab[8][2] ) );
  NOR2_X1 U119 ( .A1(n93), .A2(n70), .ZN(\ab[8][1] ) );
  NOR2_X1 U120 ( .A1(n79), .A2(n70), .ZN(\ab[8][15] ) );
  NOR2_X1 U121 ( .A1(n80), .A2(n70), .ZN(\ab[8][14] ) );
  NOR2_X1 U122 ( .A1(n81), .A2(n70), .ZN(\ab[8][13] ) );
  NOR2_X1 U123 ( .A1(n82), .A2(n70), .ZN(\ab[8][12] ) );
  NOR2_X1 U124 ( .A1(n83), .A2(n70), .ZN(\ab[8][11] ) );
  NOR2_X1 U125 ( .A1(n84), .A2(n70), .ZN(\ab[8][10] ) );
  NOR2_X1 U126 ( .A1(n94), .A2(n70), .ZN(\ab[8][0] ) );
  NOR2_X1 U127 ( .A1(n85), .A2(n71), .ZN(\ab[7][9] ) );
  NOR2_X1 U128 ( .A1(n86), .A2(n71), .ZN(\ab[7][8] ) );
  NOR2_X1 U129 ( .A1(n87), .A2(n71), .ZN(\ab[7][7] ) );
  NOR2_X1 U130 ( .A1(n88), .A2(n71), .ZN(\ab[7][6] ) );
  NOR2_X1 U131 ( .A1(n89), .A2(n71), .ZN(\ab[7][5] ) );
  NOR2_X1 U132 ( .A1(n90), .A2(n71), .ZN(\ab[7][4] ) );
  NOR2_X1 U133 ( .A1(n91), .A2(n71), .ZN(\ab[7][3] ) );
  NOR2_X1 U134 ( .A1(n92), .A2(n71), .ZN(\ab[7][2] ) );
  NOR2_X1 U135 ( .A1(n93), .A2(n71), .ZN(\ab[7][1] ) );
  NOR2_X1 U136 ( .A1(n79), .A2(n71), .ZN(\ab[7][15] ) );
  NOR2_X1 U137 ( .A1(n80), .A2(n71), .ZN(\ab[7][14] ) );
  NOR2_X1 U138 ( .A1(n81), .A2(n71), .ZN(\ab[7][13] ) );
  NOR2_X1 U139 ( .A1(n82), .A2(n71), .ZN(\ab[7][12] ) );
  NOR2_X1 U140 ( .A1(n83), .A2(n71), .ZN(\ab[7][11] ) );
  NOR2_X1 U141 ( .A1(n84), .A2(n71), .ZN(\ab[7][10] ) );
  NOR2_X1 U142 ( .A1(n94), .A2(n71), .ZN(\ab[7][0] ) );
  NOR2_X1 U143 ( .A1(n85), .A2(n72), .ZN(\ab[6][9] ) );
  NOR2_X1 U144 ( .A1(n86), .A2(n72), .ZN(\ab[6][8] ) );
  NOR2_X1 U145 ( .A1(n87), .A2(n72), .ZN(\ab[6][7] ) );
  NOR2_X1 U146 ( .A1(n88), .A2(n72), .ZN(\ab[6][6] ) );
  NOR2_X1 U147 ( .A1(n89), .A2(n72), .ZN(\ab[6][5] ) );
  NOR2_X1 U148 ( .A1(n90), .A2(n72), .ZN(\ab[6][4] ) );
  NOR2_X1 U149 ( .A1(n91), .A2(n72), .ZN(\ab[6][3] ) );
  NOR2_X1 U150 ( .A1(n92), .A2(n72), .ZN(\ab[6][2] ) );
  NOR2_X1 U151 ( .A1(n93), .A2(n72), .ZN(\ab[6][1] ) );
  NOR2_X1 U152 ( .A1(n79), .A2(n72), .ZN(\ab[6][15] ) );
  NOR2_X1 U153 ( .A1(n80), .A2(n72), .ZN(\ab[6][14] ) );
  NOR2_X1 U154 ( .A1(n81), .A2(n72), .ZN(\ab[6][13] ) );
  NOR2_X1 U155 ( .A1(n82), .A2(n72), .ZN(\ab[6][12] ) );
  NOR2_X1 U156 ( .A1(n83), .A2(n72), .ZN(\ab[6][11] ) );
  NOR2_X1 U157 ( .A1(n84), .A2(n72), .ZN(\ab[6][10] ) );
  NOR2_X1 U158 ( .A1(n94), .A2(n72), .ZN(\ab[6][0] ) );
  NOR2_X1 U159 ( .A1(n85), .A2(n73), .ZN(\ab[5][9] ) );
  NOR2_X1 U160 ( .A1(n86), .A2(n73), .ZN(\ab[5][8] ) );
  NOR2_X1 U161 ( .A1(n87), .A2(n73), .ZN(\ab[5][7] ) );
  NOR2_X1 U162 ( .A1(n88), .A2(n73), .ZN(\ab[5][6] ) );
  NOR2_X1 U163 ( .A1(n89), .A2(n73), .ZN(\ab[5][5] ) );
  NOR2_X1 U164 ( .A1(n90), .A2(n73), .ZN(\ab[5][4] ) );
  NOR2_X1 U165 ( .A1(n91), .A2(n73), .ZN(\ab[5][3] ) );
  NOR2_X1 U166 ( .A1(n92), .A2(n73), .ZN(\ab[5][2] ) );
  NOR2_X1 U167 ( .A1(n93), .A2(n73), .ZN(\ab[5][1] ) );
  NOR2_X1 U168 ( .A1(n79), .A2(n73), .ZN(\ab[5][15] ) );
  NOR2_X1 U169 ( .A1(n80), .A2(n73), .ZN(\ab[5][14] ) );
  NOR2_X1 U170 ( .A1(n81), .A2(n73), .ZN(\ab[5][13] ) );
  NOR2_X1 U171 ( .A1(n82), .A2(n73), .ZN(\ab[5][12] ) );
  NOR2_X1 U172 ( .A1(n83), .A2(n73), .ZN(\ab[5][11] ) );
  NOR2_X1 U173 ( .A1(n84), .A2(n73), .ZN(\ab[5][10] ) );
  NOR2_X1 U174 ( .A1(n94), .A2(n73), .ZN(\ab[5][0] ) );
  NOR2_X1 U175 ( .A1(n85), .A2(n74), .ZN(\ab[4][9] ) );
  NOR2_X1 U176 ( .A1(n86), .A2(n74), .ZN(\ab[4][8] ) );
  NOR2_X1 U177 ( .A1(n87), .A2(n74), .ZN(\ab[4][7] ) );
  NOR2_X1 U178 ( .A1(n88), .A2(n74), .ZN(\ab[4][6] ) );
  NOR2_X1 U179 ( .A1(n89), .A2(n74), .ZN(\ab[4][5] ) );
  NOR2_X1 U180 ( .A1(n90), .A2(n74), .ZN(\ab[4][4] ) );
  NOR2_X1 U181 ( .A1(n91), .A2(n74), .ZN(\ab[4][3] ) );
  NOR2_X1 U182 ( .A1(n92), .A2(n74), .ZN(\ab[4][2] ) );
  NOR2_X1 U183 ( .A1(n93), .A2(n74), .ZN(\ab[4][1] ) );
  NOR2_X1 U184 ( .A1(n79), .A2(n74), .ZN(\ab[4][15] ) );
  NOR2_X1 U185 ( .A1(n80), .A2(n74), .ZN(\ab[4][14] ) );
  NOR2_X1 U186 ( .A1(n81), .A2(n74), .ZN(\ab[4][13] ) );
  NOR2_X1 U187 ( .A1(n82), .A2(n74), .ZN(\ab[4][12] ) );
  NOR2_X1 U188 ( .A1(n83), .A2(n74), .ZN(\ab[4][11] ) );
  NOR2_X1 U189 ( .A1(n84), .A2(n74), .ZN(\ab[4][10] ) );
  NOR2_X1 U190 ( .A1(n94), .A2(n74), .ZN(\ab[4][0] ) );
  NOR2_X1 U191 ( .A1(n85), .A2(n75), .ZN(\ab[3][9] ) );
  NOR2_X1 U192 ( .A1(n86), .A2(n75), .ZN(\ab[3][8] ) );
  NOR2_X1 U193 ( .A1(n87), .A2(n75), .ZN(\ab[3][7] ) );
  NOR2_X1 U194 ( .A1(n88), .A2(n75), .ZN(\ab[3][6] ) );
  NOR2_X1 U195 ( .A1(n89), .A2(n75), .ZN(\ab[3][5] ) );
  NOR2_X1 U196 ( .A1(n90), .A2(n75), .ZN(\ab[3][4] ) );
  NOR2_X1 U197 ( .A1(n91), .A2(n75), .ZN(\ab[3][3] ) );
  NOR2_X1 U198 ( .A1(n92), .A2(n75), .ZN(\ab[3][2] ) );
  NOR2_X1 U199 ( .A1(n93), .A2(n75), .ZN(\ab[3][1] ) );
  NOR2_X1 U200 ( .A1(n79), .A2(n75), .ZN(\ab[3][15] ) );
  NOR2_X1 U201 ( .A1(n80), .A2(n75), .ZN(\ab[3][14] ) );
  NOR2_X1 U202 ( .A1(n81), .A2(n75), .ZN(\ab[3][13] ) );
  NOR2_X1 U203 ( .A1(n82), .A2(n75), .ZN(\ab[3][12] ) );
  NOR2_X1 U204 ( .A1(n83), .A2(n75), .ZN(\ab[3][11] ) );
  NOR2_X1 U205 ( .A1(n84), .A2(n75), .ZN(\ab[3][10] ) );
  NOR2_X1 U206 ( .A1(n94), .A2(n75), .ZN(\ab[3][0] ) );
  NOR2_X1 U207 ( .A1(n85), .A2(n76), .ZN(\ab[2][9] ) );
  NOR2_X1 U208 ( .A1(n86), .A2(n76), .ZN(\ab[2][8] ) );
  NOR2_X1 U209 ( .A1(n87), .A2(n76), .ZN(\ab[2][7] ) );
  NOR2_X1 U210 ( .A1(n88), .A2(n76), .ZN(\ab[2][6] ) );
  NOR2_X1 U211 ( .A1(n89), .A2(n76), .ZN(\ab[2][5] ) );
  NOR2_X1 U212 ( .A1(n90), .A2(n76), .ZN(\ab[2][4] ) );
  NOR2_X1 U213 ( .A1(n91), .A2(n76), .ZN(\ab[2][3] ) );
  NOR2_X1 U214 ( .A1(n92), .A2(n76), .ZN(\ab[2][2] ) );
  NOR2_X1 U215 ( .A1(n93), .A2(n76), .ZN(\ab[2][1] ) );
  NOR2_X1 U216 ( .A1(n79), .A2(n76), .ZN(\ab[2][15] ) );
  NOR2_X1 U217 ( .A1(n80), .A2(n76), .ZN(\ab[2][14] ) );
  NOR2_X1 U218 ( .A1(n81), .A2(n76), .ZN(\ab[2][13] ) );
  NOR2_X1 U219 ( .A1(n82), .A2(n76), .ZN(\ab[2][12] ) );
  NOR2_X1 U220 ( .A1(n83), .A2(n76), .ZN(\ab[2][11] ) );
  NOR2_X1 U221 ( .A1(n84), .A2(n76), .ZN(\ab[2][10] ) );
  NOR2_X1 U222 ( .A1(n94), .A2(n76), .ZN(\ab[2][0] ) );
  NOR2_X1 U223 ( .A1(n85), .A2(n77), .ZN(\ab[1][9] ) );
  NOR2_X1 U224 ( .A1(n86), .A2(n77), .ZN(\ab[1][8] ) );
  NOR2_X1 U225 ( .A1(n87), .A2(n77), .ZN(\ab[1][7] ) );
  NOR2_X1 U226 ( .A1(n88), .A2(n77), .ZN(\ab[1][6] ) );
  NOR2_X1 U227 ( .A1(n89), .A2(n77), .ZN(\ab[1][5] ) );
  NOR2_X1 U228 ( .A1(n90), .A2(n77), .ZN(\ab[1][4] ) );
  NOR2_X1 U229 ( .A1(n91), .A2(n77), .ZN(\ab[1][3] ) );
  NOR2_X1 U230 ( .A1(n92), .A2(n77), .ZN(\ab[1][2] ) );
  NOR2_X1 U231 ( .A1(n93), .A2(n77), .ZN(\ab[1][1] ) );
  NOR2_X1 U232 ( .A1(n79), .A2(n77), .ZN(\ab[1][15] ) );
  NOR2_X1 U233 ( .A1(n80), .A2(n77), .ZN(\ab[1][14] ) );
  NOR2_X1 U234 ( .A1(n81), .A2(n77), .ZN(\ab[1][13] ) );
  NOR2_X1 U235 ( .A1(n82), .A2(n77), .ZN(\ab[1][12] ) );
  NOR2_X1 U236 ( .A1(n83), .A2(n77), .ZN(\ab[1][11] ) );
  NOR2_X1 U237 ( .A1(n84), .A2(n77), .ZN(\ab[1][10] ) );
  NOR2_X1 U238 ( .A1(n94), .A2(n77), .ZN(\ab[1][0] ) );
  NOR2_X1 U239 ( .A1(n85), .A2(n63), .ZN(\ab[15][9] ) );
  NOR2_X1 U240 ( .A1(n86), .A2(n63), .ZN(\ab[15][8] ) );
  NOR2_X1 U241 ( .A1(n87), .A2(n63), .ZN(\ab[15][7] ) );
  NOR2_X1 U242 ( .A1(n88), .A2(n63), .ZN(\ab[15][6] ) );
  NOR2_X1 U243 ( .A1(n89), .A2(n63), .ZN(\ab[15][5] ) );
  NOR2_X1 U244 ( .A1(n90), .A2(n63), .ZN(\ab[15][4] ) );
  NOR2_X1 U245 ( .A1(n91), .A2(n63), .ZN(\ab[15][3] ) );
  NOR2_X1 U246 ( .A1(n92), .A2(n63), .ZN(\ab[15][2] ) );
  NOR2_X1 U247 ( .A1(n93), .A2(n63), .ZN(\ab[15][1] ) );
  NOR2_X1 U248 ( .A1(n79), .A2(n63), .ZN(\ab[15][15] ) );
  NOR2_X1 U249 ( .A1(n80), .A2(n63), .ZN(\ab[15][14] ) );
  NOR2_X1 U250 ( .A1(n81), .A2(n63), .ZN(\ab[15][13] ) );
  NOR2_X1 U251 ( .A1(n82), .A2(n63), .ZN(\ab[15][12] ) );
  NOR2_X1 U252 ( .A1(n83), .A2(n63), .ZN(\ab[15][11] ) );
  NOR2_X1 U253 ( .A1(n84), .A2(n63), .ZN(\ab[15][10] ) );
  NOR2_X1 U254 ( .A1(n94), .A2(n63), .ZN(\ab[15][0] ) );
  NOR2_X1 U255 ( .A1(n85), .A2(n64), .ZN(\ab[14][9] ) );
  NOR2_X1 U256 ( .A1(n86), .A2(n64), .ZN(\ab[14][8] ) );
  NOR2_X1 U257 ( .A1(n87), .A2(n64), .ZN(\ab[14][7] ) );
  NOR2_X1 U258 ( .A1(n88), .A2(n64), .ZN(\ab[14][6] ) );
  NOR2_X1 U259 ( .A1(n89), .A2(n64), .ZN(\ab[14][5] ) );
  NOR2_X1 U260 ( .A1(n90), .A2(n64), .ZN(\ab[14][4] ) );
  NOR2_X1 U261 ( .A1(n91), .A2(n64), .ZN(\ab[14][3] ) );
  NOR2_X1 U262 ( .A1(n92), .A2(n64), .ZN(\ab[14][2] ) );
  NOR2_X1 U263 ( .A1(n93), .A2(n64), .ZN(\ab[14][1] ) );
  NOR2_X1 U264 ( .A1(n79), .A2(n64), .ZN(\ab[14][15] ) );
  NOR2_X1 U265 ( .A1(n80), .A2(n64), .ZN(\ab[14][14] ) );
  NOR2_X1 U266 ( .A1(n81), .A2(n64), .ZN(\ab[14][13] ) );
  NOR2_X1 U267 ( .A1(n82), .A2(n64), .ZN(\ab[14][12] ) );
  NOR2_X1 U268 ( .A1(n83), .A2(n64), .ZN(\ab[14][11] ) );
  NOR2_X1 U269 ( .A1(n84), .A2(n64), .ZN(\ab[14][10] ) );
  NOR2_X1 U270 ( .A1(n94), .A2(n64), .ZN(\ab[14][0] ) );
  NOR2_X1 U271 ( .A1(n85), .A2(n65), .ZN(\ab[13][9] ) );
  NOR2_X1 U272 ( .A1(n86), .A2(n65), .ZN(\ab[13][8] ) );
  NOR2_X1 U273 ( .A1(n87), .A2(n65), .ZN(\ab[13][7] ) );
  NOR2_X1 U274 ( .A1(n88), .A2(n65), .ZN(\ab[13][6] ) );
  NOR2_X1 U275 ( .A1(n89), .A2(n65), .ZN(\ab[13][5] ) );
  NOR2_X1 U276 ( .A1(n90), .A2(n65), .ZN(\ab[13][4] ) );
  NOR2_X1 U277 ( .A1(n91), .A2(n65), .ZN(\ab[13][3] ) );
  NOR2_X1 U278 ( .A1(n92), .A2(n65), .ZN(\ab[13][2] ) );
  NOR2_X1 U279 ( .A1(n93), .A2(n65), .ZN(\ab[13][1] ) );
  NOR2_X1 U280 ( .A1(n79), .A2(n65), .ZN(\ab[13][15] ) );
  NOR2_X1 U281 ( .A1(n80), .A2(n65), .ZN(\ab[13][14] ) );
  NOR2_X1 U282 ( .A1(n81), .A2(n65), .ZN(\ab[13][13] ) );
  NOR2_X1 U283 ( .A1(n82), .A2(n65), .ZN(\ab[13][12] ) );
  NOR2_X1 U284 ( .A1(n83), .A2(n65), .ZN(\ab[13][11] ) );
  NOR2_X1 U285 ( .A1(n84), .A2(n65), .ZN(\ab[13][10] ) );
  NOR2_X1 U286 ( .A1(n94), .A2(n65), .ZN(\ab[13][0] ) );
  NOR2_X1 U287 ( .A1(n85), .A2(n66), .ZN(\ab[12][9] ) );
  NOR2_X1 U288 ( .A1(n86), .A2(n66), .ZN(\ab[12][8] ) );
  NOR2_X1 U289 ( .A1(n87), .A2(n66), .ZN(\ab[12][7] ) );
  NOR2_X1 U290 ( .A1(n88), .A2(n66), .ZN(\ab[12][6] ) );
  NOR2_X1 U291 ( .A1(n89), .A2(n66), .ZN(\ab[12][5] ) );
  NOR2_X1 U292 ( .A1(n90), .A2(n66), .ZN(\ab[12][4] ) );
  NOR2_X1 U293 ( .A1(n91), .A2(n66), .ZN(\ab[12][3] ) );
  NOR2_X1 U294 ( .A1(n92), .A2(n66), .ZN(\ab[12][2] ) );
  NOR2_X1 U295 ( .A1(n93), .A2(n66), .ZN(\ab[12][1] ) );
  NOR2_X1 U296 ( .A1(n79), .A2(n66), .ZN(\ab[12][15] ) );
  NOR2_X1 U297 ( .A1(n80), .A2(n66), .ZN(\ab[12][14] ) );
  NOR2_X1 U298 ( .A1(n81), .A2(n66), .ZN(\ab[12][13] ) );
  NOR2_X1 U299 ( .A1(n82), .A2(n66), .ZN(\ab[12][12] ) );
  NOR2_X1 U300 ( .A1(n83), .A2(n66), .ZN(\ab[12][11] ) );
  NOR2_X1 U301 ( .A1(n84), .A2(n66), .ZN(\ab[12][10] ) );
  NOR2_X1 U302 ( .A1(n94), .A2(n66), .ZN(\ab[12][0] ) );
  NOR2_X1 U303 ( .A1(n85), .A2(n67), .ZN(\ab[11][9] ) );
  NOR2_X1 U304 ( .A1(n86), .A2(n67), .ZN(\ab[11][8] ) );
  NOR2_X1 U305 ( .A1(n87), .A2(n67), .ZN(\ab[11][7] ) );
  NOR2_X1 U306 ( .A1(n88), .A2(n67), .ZN(\ab[11][6] ) );
  NOR2_X1 U307 ( .A1(n89), .A2(n67), .ZN(\ab[11][5] ) );
  NOR2_X1 U308 ( .A1(n90), .A2(n67), .ZN(\ab[11][4] ) );
  NOR2_X1 U309 ( .A1(n91), .A2(n67), .ZN(\ab[11][3] ) );
  NOR2_X1 U310 ( .A1(n92), .A2(n67), .ZN(\ab[11][2] ) );
  NOR2_X1 U311 ( .A1(n93), .A2(n67), .ZN(\ab[11][1] ) );
  NOR2_X1 U312 ( .A1(n79), .A2(n67), .ZN(\ab[11][15] ) );
  NOR2_X1 U313 ( .A1(n80), .A2(n67), .ZN(\ab[11][14] ) );
  NOR2_X1 U314 ( .A1(n81), .A2(n67), .ZN(\ab[11][13] ) );
  NOR2_X1 U315 ( .A1(n82), .A2(n67), .ZN(\ab[11][12] ) );
  NOR2_X1 U316 ( .A1(n83), .A2(n67), .ZN(\ab[11][11] ) );
  NOR2_X1 U317 ( .A1(n84), .A2(n67), .ZN(\ab[11][10] ) );
  NOR2_X1 U318 ( .A1(n94), .A2(n67), .ZN(\ab[11][0] ) );
  NOR2_X1 U319 ( .A1(n85), .A2(n68), .ZN(\ab[10][9] ) );
  NOR2_X1 U320 ( .A1(n86), .A2(n68), .ZN(\ab[10][8] ) );
  NOR2_X1 U321 ( .A1(n87), .A2(n68), .ZN(\ab[10][7] ) );
  NOR2_X1 U322 ( .A1(n88), .A2(n68), .ZN(\ab[10][6] ) );
  NOR2_X1 U323 ( .A1(n89), .A2(n68), .ZN(\ab[10][5] ) );
  NOR2_X1 U324 ( .A1(n90), .A2(n68), .ZN(\ab[10][4] ) );
  NOR2_X1 U325 ( .A1(n91), .A2(n68), .ZN(\ab[10][3] ) );
  NOR2_X1 U326 ( .A1(n92), .A2(n68), .ZN(\ab[10][2] ) );
  NOR2_X1 U327 ( .A1(n93), .A2(n68), .ZN(\ab[10][1] ) );
  NOR2_X1 U328 ( .A1(n79), .A2(n68), .ZN(\ab[10][15] ) );
  NOR2_X1 U329 ( .A1(n80), .A2(n68), .ZN(\ab[10][14] ) );
  NOR2_X1 U330 ( .A1(n81), .A2(n68), .ZN(\ab[10][13] ) );
  NOR2_X1 U331 ( .A1(n82), .A2(n68), .ZN(\ab[10][12] ) );
  NOR2_X1 U332 ( .A1(n83), .A2(n68), .ZN(\ab[10][11] ) );
  NOR2_X1 U333 ( .A1(n84), .A2(n68), .ZN(\ab[10][10] ) );
  NOR2_X1 U334 ( .A1(n94), .A2(n68), .ZN(\ab[10][0] ) );
  NOR2_X1 U335 ( .A1(n85), .A2(n78), .ZN(\ab[0][9] ) );
  NOR2_X1 U336 ( .A1(n86), .A2(n78), .ZN(\ab[0][8] ) );
  NOR2_X1 U337 ( .A1(n87), .A2(n78), .ZN(\ab[0][7] ) );
  NOR2_X1 U338 ( .A1(n88), .A2(n78), .ZN(\ab[0][6] ) );
  NOR2_X1 U339 ( .A1(n89), .A2(n78), .ZN(\ab[0][5] ) );
  NOR2_X1 U340 ( .A1(n90), .A2(n78), .ZN(\ab[0][4] ) );
  NOR2_X1 U341 ( .A1(n91), .A2(n78), .ZN(\ab[0][3] ) );
  NOR2_X1 U342 ( .A1(n92), .A2(n78), .ZN(\ab[0][2] ) );
  NOR2_X1 U343 ( .A1(n93), .A2(n78), .ZN(\ab[0][1] ) );
  NOR2_X1 U344 ( .A1(n79), .A2(n78), .ZN(\ab[0][15] ) );
  NOR2_X1 U345 ( .A1(n80), .A2(n78), .ZN(\ab[0][14] ) );
  NOR2_X1 U346 ( .A1(n81), .A2(n78), .ZN(\ab[0][13] ) );
  NOR2_X1 U347 ( .A1(n82), .A2(n78), .ZN(\ab[0][12] ) );
  NOR2_X1 U348 ( .A1(n83), .A2(n78), .ZN(\ab[0][11] ) );
  NOR2_X1 U349 ( .A1(n84), .A2(n78), .ZN(\ab[0][10] ) );
  NOR2_X1 U350 ( .A1(n94), .A2(n78), .ZN(PRODUCT[0]) );
  multiplier_DW01_add_5 FS_1 ( .A({1'b0, n17, n25, n18, n26, n19, n27, n20, 
        n28, n21, n29, n22, n30, n23, n24, n61, \SUMB[15][0] , \A1[12] , 
        \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , 
        \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({n62, n47, n54, n48, 
        n55, n49, n56, n50, n57, n51, n58, n52, n59, n53, n60, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .CI(1'b0), .SUM(PRODUCT[31:2]) );
endmodule


module multiplier_DW01_add_6 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70;

  OR2_X4 U2 ( .A1(B[15]), .A2(A[15]), .ZN(n1) );
  AND2_X4 U3 ( .A1(n1), .A2(n70), .ZN(SUM[15]) );
  INV_X4 U4 ( .A(B[29]), .ZN(n3) );
  INV_X4 U5 ( .A(n21), .ZN(n4) );
  INV_X4 U6 ( .A(n23), .ZN(n5) );
  INV_X4 U7 ( .A(n29), .ZN(n6) );
  INV_X4 U8 ( .A(n31), .ZN(n7) );
  INV_X4 U9 ( .A(n37), .ZN(n8) );
  INV_X4 U10 ( .A(n39), .ZN(n9) );
  INV_X4 U11 ( .A(n45), .ZN(n10) );
  INV_X4 U12 ( .A(n47), .ZN(n11) );
  INV_X4 U13 ( .A(n53), .ZN(n12) );
  INV_X4 U14 ( .A(n55), .ZN(n13) );
  INV_X4 U15 ( .A(n61), .ZN(n14) );
  INV_X4 U16 ( .A(n63), .ZN(n15) );
  INV_X4 U17 ( .A(n68), .ZN(n16) );
  INV_X4 U18 ( .A(n70), .ZN(n17) );
  XOR2_X1 U19 ( .A(n3), .B(n18), .Z(SUM[29]) );
  AOI21_X1 U20 ( .B1(n19), .B2(n4), .A(n20), .ZN(n18) );
  XOR2_X1 U21 ( .A(n19), .B(n22), .Z(SUM[28]) );
  NOR2_X1 U22 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U23 ( .A1(B[28]), .A2(A[28]), .ZN(n21) );
  AND2_X1 U24 ( .A1(B[28]), .A2(A[28]), .ZN(n20) );
  OAI21_X1 U25 ( .B1(n23), .B2(n24), .A(n25), .ZN(n19) );
  XOR2_X1 U26 ( .A(n26), .B(n24), .Z(SUM[27]) );
  AOI21_X1 U27 ( .B1(n6), .B2(n27), .A(n28), .ZN(n24) );
  NAND2_X1 U28 ( .A1(n5), .A2(n25), .ZN(n26) );
  NAND2_X1 U29 ( .A1(B[27]), .A2(A[27]), .ZN(n25) );
  NOR2_X1 U30 ( .A1(B[27]), .A2(A[27]), .ZN(n23) );
  XOR2_X1 U31 ( .A(n27), .B(n30), .Z(SUM[26]) );
  NOR2_X1 U32 ( .A1(n28), .A2(n29), .ZN(n30) );
  NOR2_X1 U33 ( .A1(B[26]), .A2(A[26]), .ZN(n29) );
  AND2_X1 U34 ( .A1(B[26]), .A2(A[26]), .ZN(n28) );
  OAI21_X1 U35 ( .B1(n31), .B2(n32), .A(n33), .ZN(n27) );
  XOR2_X1 U36 ( .A(n34), .B(n32), .Z(SUM[25]) );
  AOI21_X1 U37 ( .B1(n8), .B2(n35), .A(n36), .ZN(n32) );
  NAND2_X1 U38 ( .A1(n7), .A2(n33), .ZN(n34) );
  NAND2_X1 U39 ( .A1(B[25]), .A2(A[25]), .ZN(n33) );
  NOR2_X1 U40 ( .A1(B[25]), .A2(A[25]), .ZN(n31) );
  XOR2_X1 U41 ( .A(n35), .B(n38), .Z(SUM[24]) );
  NOR2_X1 U42 ( .A1(n36), .A2(n37), .ZN(n38) );
  NOR2_X1 U43 ( .A1(B[24]), .A2(A[24]), .ZN(n37) );
  AND2_X1 U44 ( .A1(B[24]), .A2(A[24]), .ZN(n36) );
  OAI21_X1 U45 ( .B1(n39), .B2(n40), .A(n41), .ZN(n35) );
  XOR2_X1 U46 ( .A(n42), .B(n40), .Z(SUM[23]) );
  AOI21_X1 U47 ( .B1(n10), .B2(n43), .A(n44), .ZN(n40) );
  NAND2_X1 U48 ( .A1(n9), .A2(n41), .ZN(n42) );
  NAND2_X1 U49 ( .A1(B[23]), .A2(A[23]), .ZN(n41) );
  NOR2_X1 U50 ( .A1(B[23]), .A2(A[23]), .ZN(n39) );
  XOR2_X1 U51 ( .A(n43), .B(n46), .Z(SUM[22]) );
  NOR2_X1 U52 ( .A1(n44), .A2(n45), .ZN(n46) );
  NOR2_X1 U53 ( .A1(B[22]), .A2(A[22]), .ZN(n45) );
  AND2_X1 U54 ( .A1(B[22]), .A2(A[22]), .ZN(n44) );
  OAI21_X1 U55 ( .B1(n47), .B2(n48), .A(n49), .ZN(n43) );
  XOR2_X1 U56 ( .A(n50), .B(n48), .Z(SUM[21]) );
  AOI21_X1 U57 ( .B1(n12), .B2(n51), .A(n52), .ZN(n48) );
  NAND2_X1 U58 ( .A1(n11), .A2(n49), .ZN(n50) );
  NAND2_X1 U59 ( .A1(B[21]), .A2(A[21]), .ZN(n49) );
  NOR2_X1 U60 ( .A1(B[21]), .A2(A[21]), .ZN(n47) );
  XOR2_X1 U61 ( .A(n51), .B(n54), .Z(SUM[20]) );
  NOR2_X1 U62 ( .A1(n52), .A2(n53), .ZN(n54) );
  NOR2_X1 U63 ( .A1(B[20]), .A2(A[20]), .ZN(n53) );
  AND2_X1 U64 ( .A1(B[20]), .A2(A[20]), .ZN(n52) );
  OAI21_X1 U65 ( .B1(n55), .B2(n56), .A(n57), .ZN(n51) );
  XOR2_X1 U66 ( .A(n58), .B(n56), .Z(SUM[19]) );
  AOI21_X1 U67 ( .B1(n14), .B2(n59), .A(n60), .ZN(n56) );
  NAND2_X1 U68 ( .A1(n13), .A2(n57), .ZN(n58) );
  NAND2_X1 U69 ( .A1(B[19]), .A2(A[19]), .ZN(n57) );
  NOR2_X1 U70 ( .A1(B[19]), .A2(A[19]), .ZN(n55) );
  XOR2_X1 U71 ( .A(n59), .B(n62), .Z(SUM[18]) );
  NOR2_X1 U72 ( .A1(n60), .A2(n61), .ZN(n62) );
  NOR2_X1 U73 ( .A1(B[18]), .A2(A[18]), .ZN(n61) );
  AND2_X1 U74 ( .A1(B[18]), .A2(A[18]), .ZN(n60) );
  OAI21_X1 U75 ( .B1(n63), .B2(n64), .A(n65), .ZN(n59) );
  XOR2_X1 U76 ( .A(n66), .B(n64), .Z(SUM[17]) );
  AOI21_X1 U77 ( .B1(n16), .B2(n17), .A(n67), .ZN(n64) );
  NAND2_X1 U78 ( .A1(n15), .A2(n65), .ZN(n66) );
  NAND2_X1 U79 ( .A1(B[17]), .A2(A[17]), .ZN(n65) );
  NOR2_X1 U80 ( .A1(B[17]), .A2(A[17]), .ZN(n63) );
  XOR2_X1 U81 ( .A(n17), .B(n69), .Z(SUM[16]) );
  NOR2_X1 U82 ( .A1(n67), .A2(n68), .ZN(n69) );
  NOR2_X1 U83 ( .A1(B[16]), .A2(A[16]), .ZN(n68) );
  AND2_X1 U84 ( .A1(B[16]), .A2(A[16]), .ZN(n67) );
  NAND2_X1 U85 ( .A1(B[15]), .A2(A[15]), .ZN(n70) );
  BUF_X4 U86 ( .A(A[9]), .Z(SUM[9]) );
  BUF_X4 U87 ( .A(A[8]), .Z(SUM[8]) );
  BUF_X4 U88 ( .A(A[7]), .Z(SUM[7]) );
  BUF_X4 U89 ( .A(A[6]), .Z(SUM[6]) );
  BUF_X4 U90 ( .A(A[5]), .Z(SUM[5]) );
  BUF_X4 U91 ( .A(A[4]), .Z(SUM[4]) );
  BUF_X4 U92 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X4 U93 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X4 U94 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X4 U95 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X32 U96 ( .A(A[10]), .Z(SUM[10]) );
  BUF_X32 U97 ( .A(A[11]), .Z(SUM[11]) );
  BUF_X32 U98 ( .A(A[12]), .Z(SUM[12]) );
  BUF_X32 U99 ( .A(A[13]), .Z(SUM[13]) );
  BUF_X32 U100 ( .A(A[14]), .Z(SUM[14]) );
endmodule


module multiplier_DW02_mult_2 ( A, B, TC, PRODUCT );
  input [15:0] A;
  input [15:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] ,
         \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] ,
         \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] ,
         \ab[15][0] , \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] ,
         \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] ,
         \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][15] , \ab[13][14] , \ab[13][13] ,
         \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] ,
         \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] ,
         \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][15] , \ab[12][14] ,
         \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] ,
         \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] ,
         \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][15] ,
         \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] ,
         \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] ,
         \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] ,
         \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] ,
         \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][15] , \ab[8][14] , \ab[8][13] ,
         \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][15] , \ab[7][14] ,
         \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] , \ab[7][9] ,
         \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] ,
         \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][15] ,
         \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] ,
         \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] ,
         \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][15] , \ab[3][14] , \ab[3][13] ,
         \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][15] , \ab[2][14] ,
         \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] , \ab[2][9] ,
         \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] ,
         \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][15] ,
         \ab[1][14] , \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] ,
         \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] ,
         \ab[0][15] , \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] ,
         \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] ,
         \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] ,
         \CARRYB[15][14] , \CARRYB[15][13] , \CARRYB[15][12] ,
         \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] ,
         \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] ,
         \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] ,
         \CARRYB[14][14] , \CARRYB[14][13] , \CARRYB[14][12] ,
         \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] ,
         \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] ,
         \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][14] , \CARRYB[12][13] , \CARRYB[12][12] ,
         \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] ,
         \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] ,
         \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] ,
         \CARRYB[11][14] , \CARRYB[11][13] , \CARRYB[11][12] ,
         \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] ,
         \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] ,
         \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] ,
         \CARRYB[10][14] , \CARRYB[10][13] , \CARRYB[10][12] ,
         \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] ,
         \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] ,
         \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] ,
         \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] ,
         \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] ,
         \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][14] ,
         \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] ,
         \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] ,
         \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] ,
         \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] ,
         \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] ,
         \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] ,
         \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] ,
         \CARRYB[5][14] , \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] ,
         \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] ,
         \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] ,
         \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][14] ,
         \CARRYB[4][13] , \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] ,
         \CARRYB[4][9] , \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] ,
         \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] ,
         \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][14] , \CARRYB[3][13] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] ,
         \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] ,
         \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] ,
         \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[15][0] , \SUMB[14][14] ,
         \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] ,
         \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] ,
         \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] ,
         \SUMB[14][1] , \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] ,
         \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] ,
         \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] ,
         \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] ,
         \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] ,
         \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] ,
         \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][14] , \SUMB[8][13] ,
         \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] ,
         \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] ,
         \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \A1[12] ,
         \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] ,
         \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] , n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94;

  FA_X1 S4_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), .CO(
        \CARRYB[15][0] ), .S(\SUMB[15][0] ) );
  FA_X1 S4_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), .CO(
        \CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA_X1 S4_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), .CO(
        \CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA_X1 S4_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), .CO(
        \CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA_X1 S4_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), .CO(
        \CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA_X1 S4_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), .CO(
        \CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA_X1 S4_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), .CO(
        \CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA_X1 S4_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), .CO(
        \CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA_X1 S4_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), .CO(
        \CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA_X1 S4_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), .CO(
        \CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA_X1 S4_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA_X1 S4_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA_X1 S4_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA_X1 S4_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA_X1 S5_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\ab[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA_X1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FA_X1 S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA_X1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA_X1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA_X1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA_X1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA_X1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA_X1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA_X1 S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA_X1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA_X1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA_X1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA_X1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA_X1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA_X1 S3_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\ab[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA_X1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA_X1 S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA_X1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA_X1 S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA_X1 S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA_X1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA_X1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA_X1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA_X1 S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA_X1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA_X1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA_X1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA_X1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA_X1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA_X1 S3_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\ab[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA_X1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA_X1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA_X1 S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA_X1 S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA_X1 S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA_X1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA_X1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA_X1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA_X1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA_X1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA_X1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA_X1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA_X1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA_X1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA_X1 S3_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\ab[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA_X1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA_X1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA_X1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA_X1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA_X1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA_X1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA_X1 S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA_X1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA_X1 S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA_X1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA_X1 S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA_X1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA_X1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA_X1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA_X1 S3_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\ab[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA_X1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA_X1 S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA_X1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA_X1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA_X1 S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA_X1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA_X1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA_X1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA_X1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA_X1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA_X1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA_X1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA_X1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA_X1 S3_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\ab[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA_X1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA_X1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA_X1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA_X1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA_X1 S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA_X1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA_X1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA_X1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA_X1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA_X1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA_X1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA_X1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA_X1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA_X1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA_X1 S3_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\ab[8][15] ), .CO(
        \CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA_X1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA_X1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA_X1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA_X1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA_X1 S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA_X1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA_X1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA_X1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA_X1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA_X1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA_X1 S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA_X1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA_X1 S3_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\ab[7][15] ), .CO(
        \CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA_X1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA_X1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA_X1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA_X1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA_X1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA_X1 S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA_X1 S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA_X1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA_X1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA_X1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA_X1 S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA_X1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA_X1 S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA_X1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA_X1 S3_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\ab[6][15] ), .CO(
        \CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA_X1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA_X1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA_X1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA_X1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA_X1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA_X1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA_X1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA_X1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA_X1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA_X1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA_X1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA_X1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA_X1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA_X1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA_X1 S3_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\ab[5][15] ), .CO(
        \CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA_X1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA_X1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA_X1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA_X1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA_X1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA_X1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA_X1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA_X1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA_X1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA_X1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA_X1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA_X1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA_X1 S3_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\ab[4][15] ), .CO(
        \CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA_X1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA_X1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA_X1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA_X1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA_X1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA_X1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA_X1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA_X1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA_X1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA_X1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA_X1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA_X1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA_X1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA_X1 S3_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\ab[3][15] ), .CO(
        \CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA_X1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA_X1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA_X1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA_X1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA_X1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA_X1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA_X1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA_X1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA_X1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA_X1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA_X1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA_X1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA_X1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA_X1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA_X1 S3_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\ab[2][15] ), .CO(
        \CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(n16), .CI(n45), .CO(\CARRYB[2][0] ), .S(
        \A1[0] ) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(n15), .CI(n44), .CO(\CARRYB[2][1] ), .S(
        \SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(n14), .CI(n43), .CO(\CARRYB[2][2] ), .S(
        \SUMB[2][2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2][3] ), .B(n13), .CI(n42), .CO(\CARRYB[2][3] ), .S(
        \SUMB[2][3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2][4] ), .B(n12), .CI(n41), .CO(\CARRYB[2][4] ), .S(
        \SUMB[2][4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2][5] ), .B(n11), .CI(n40), .CO(\CARRYB[2][5] ), .S(
        \SUMB[2][5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2][6] ), .B(n10), .CI(n39), .CO(\CARRYB[2][6] ), .S(
        \SUMB[2][6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(n9), .CI(n38), .CO(\CARRYB[2][7] ), .S(
        \SUMB[2][7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(n8), .CI(n37), .CO(\CARRYB[2][8] ), .S(
        \SUMB[2][8] ) );
  FA_X1 S2_2_9 ( .A(\ab[2][9] ), .B(n7), .CI(n36), .CO(\CARRYB[2][9] ), .S(
        \SUMB[2][9] ) );
  FA_X1 S2_2_10 ( .A(\ab[2][10] ), .B(n6), .CI(n35), .CO(\CARRYB[2][10] ), .S(
        \SUMB[2][10] ) );
  FA_X1 S2_2_11 ( .A(\ab[2][11] ), .B(n5), .CI(n34), .CO(\CARRYB[2][11] ), .S(
        \SUMB[2][11] ) );
  FA_X1 S2_2_12 ( .A(\ab[2][12] ), .B(n4), .CI(n33), .CO(\CARRYB[2][12] ), .S(
        \SUMB[2][12] ) );
  FA_X1 S2_2_13 ( .A(\ab[2][13] ), .B(n3), .CI(n32), .CO(\CARRYB[2][13] ), .S(
        \SUMB[2][13] ) );
  FA_X1 S3_2_14 ( .A(\ab[2][14] ), .B(n31), .CI(\ab[1][15] ), .CO(
        \CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  AND2_X4 U2 ( .A1(\ab[0][14] ), .A2(\ab[1][13] ), .ZN(n3) );
  AND2_X4 U3 ( .A1(\ab[0][13] ), .A2(\ab[1][12] ), .ZN(n4) );
  AND2_X4 U4 ( .A1(\ab[0][12] ), .A2(\ab[1][11] ), .ZN(n5) );
  AND2_X4 U5 ( .A1(\ab[0][11] ), .A2(\ab[1][10] ), .ZN(n6) );
  AND2_X4 U6 ( .A1(\ab[0][10] ), .A2(\ab[1][9] ), .ZN(n7) );
  AND2_X4 U7 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .ZN(n8) );
  AND2_X4 U8 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .ZN(n9) );
  AND2_X4 U9 ( .A1(\ab[0][7] ), .A2(\ab[1][6] ), .ZN(n10) );
  AND2_X4 U10 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .ZN(n11) );
  AND2_X4 U11 ( .A1(\ab[0][5] ), .A2(\ab[1][4] ), .ZN(n12) );
  AND2_X4 U12 ( .A1(\ab[0][4] ), .A2(\ab[1][3] ), .ZN(n13) );
  AND2_X4 U13 ( .A1(\ab[0][3] ), .A2(\ab[1][2] ), .ZN(n14) );
  AND2_X4 U14 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .ZN(n15) );
  AND2_X4 U15 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .ZN(n16) );
  XOR2_X2 U16 ( .A(\CARRYB[15][14] ), .B(\ab[15][15] ), .Z(n17) );
  XOR2_X2 U17 ( .A(\CARRYB[15][12] ), .B(\SUMB[15][13] ), .Z(n18) );
  XOR2_X2 U18 ( .A(\CARRYB[15][10] ), .B(\SUMB[15][11] ), .Z(n19) );
  XOR2_X2 U19 ( .A(\CARRYB[15][8] ), .B(\SUMB[15][9] ), .Z(n20) );
  XOR2_X2 U20 ( .A(\CARRYB[15][6] ), .B(\SUMB[15][7] ), .Z(n21) );
  XOR2_X2 U21 ( .A(\CARRYB[15][4] ), .B(\SUMB[15][5] ), .Z(n22) );
  XOR2_X2 U22 ( .A(\CARRYB[15][2] ), .B(\SUMB[15][3] ), .Z(n23) );
  XOR2_X2 U23 ( .A(\CARRYB[15][1] ), .B(\SUMB[15][2] ), .Z(n24) );
  XOR2_X2 U24 ( .A(\CARRYB[15][13] ), .B(\SUMB[15][14] ), .Z(n25) );
  XOR2_X2 U25 ( .A(\CARRYB[15][11] ), .B(\SUMB[15][12] ), .Z(n26) );
  XOR2_X2 U26 ( .A(\CARRYB[15][9] ), .B(\SUMB[15][10] ), .Z(n27) );
  XOR2_X2 U27 ( .A(\CARRYB[15][7] ), .B(\SUMB[15][8] ), .Z(n28) );
  XOR2_X2 U28 ( .A(\CARRYB[15][5] ), .B(\SUMB[15][6] ), .Z(n29) );
  XOR2_X2 U29 ( .A(\CARRYB[15][3] ), .B(\SUMB[15][4] ), .Z(n30) );
  AND2_X4 U30 ( .A1(\ab[0][15] ), .A2(\ab[1][14] ), .ZN(n31) );
  XOR2_X2 U31 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(n32) );
  XOR2_X2 U32 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(n33) );
  XOR2_X2 U33 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(n34) );
  XOR2_X2 U34 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(n35) );
  XOR2_X2 U35 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(n36) );
  XOR2_X2 U36 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(n37) );
  XOR2_X2 U37 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(n38) );
  XOR2_X2 U38 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(n39) );
  XOR2_X2 U39 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(n40) );
  XOR2_X2 U40 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(n41) );
  XOR2_X2 U41 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(n42) );
  XOR2_X2 U42 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(n43) );
  XOR2_X2 U43 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(n44) );
  XOR2_X2 U44 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(n45) );
  AND2_X4 U45 ( .A1(\CARRYB[15][13] ), .A2(\SUMB[15][14] ), .ZN(n46) );
  AND2_X4 U46 ( .A1(\CARRYB[15][11] ), .A2(\SUMB[15][12] ), .ZN(n47) );
  AND2_X4 U47 ( .A1(\CARRYB[15][9] ), .A2(\SUMB[15][10] ), .ZN(n48) );
  AND2_X4 U48 ( .A1(\CARRYB[15][7] ), .A2(\SUMB[15][8] ), .ZN(n49) );
  AND2_X4 U49 ( .A1(\CARRYB[15][5] ), .A2(\SUMB[15][6] ), .ZN(n50) );
  AND2_X4 U50 ( .A1(\CARRYB[15][3] ), .A2(\SUMB[15][4] ), .ZN(n51) );
  AND2_X4 U51 ( .A1(\CARRYB[15][1] ), .A2(\SUMB[15][2] ), .ZN(n52) );
  AND2_X4 U52 ( .A1(\CARRYB[15][12] ), .A2(\SUMB[15][13] ), .ZN(n53) );
  AND2_X4 U53 ( .A1(\CARRYB[15][10] ), .A2(\SUMB[15][11] ), .ZN(n54) );
  AND2_X4 U54 ( .A1(\CARRYB[15][8] ), .A2(\SUMB[15][9] ), .ZN(n55) );
  AND2_X4 U55 ( .A1(\CARRYB[15][6] ), .A2(\SUMB[15][7] ), .ZN(n56) );
  AND2_X4 U56 ( .A1(\CARRYB[15][4] ), .A2(\SUMB[15][5] ), .ZN(n57) );
  AND2_X4 U57 ( .A1(\CARRYB[15][2] ), .A2(\SUMB[15][3] ), .ZN(n58) );
  AND2_X4 U58 ( .A1(\CARRYB[15][0] ), .A2(\SUMB[15][1] ), .ZN(n59) );
  XOR2_X2 U59 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  XOR2_X2 U60 ( .A(\CARRYB[15][0] ), .B(\SUMB[15][1] ), .Z(n61) );
  AND2_X4 U61 ( .A1(\CARRYB[15][14] ), .A2(\ab[15][15] ), .ZN(n62) );
  INV_X4 U62 ( .A(A[9]), .ZN(n69) );
  INV_X4 U63 ( .A(B[7]), .ZN(n87) );
  INV_X4 U64 ( .A(B[1]), .ZN(n93) );
  INV_X4 U65 ( .A(B[2]), .ZN(n92) );
  INV_X4 U66 ( .A(B[3]), .ZN(n91) );
  INV_X4 U67 ( .A(B[4]), .ZN(n90) );
  INV_X4 U68 ( .A(B[5]), .ZN(n89) );
  INV_X4 U69 ( .A(B[6]), .ZN(n88) );
  INV_X4 U70 ( .A(B[9]), .ZN(n85) );
  INV_X4 U71 ( .A(B[8]), .ZN(n86) );
  INV_X4 U72 ( .A(B[11]), .ZN(n83) );
  INV_X4 U73 ( .A(B[10]), .ZN(n84) );
  INV_X4 U74 ( .A(B[13]), .ZN(n81) );
  INV_X4 U75 ( .A(B[12]), .ZN(n82) );
  INV_X4 U76 ( .A(B[14]), .ZN(n80) );
  INV_X4 U77 ( .A(B[15]), .ZN(n79) );
  INV_X4 U78 ( .A(B[0]), .ZN(n94) );
  INV_X4 U79 ( .A(A[0]), .ZN(n78) );
  INV_X4 U80 ( .A(A[1]), .ZN(n77) );
  INV_X4 U81 ( .A(A[3]), .ZN(n75) );
  INV_X4 U82 ( .A(A[4]), .ZN(n74) );
  INV_X4 U83 ( .A(A[5]), .ZN(n73) );
  INV_X4 U84 ( .A(A[6]), .ZN(n72) );
  INV_X4 U85 ( .A(A[7]), .ZN(n71) );
  INV_X4 U86 ( .A(A[8]), .ZN(n70) );
  INV_X4 U87 ( .A(A[2]), .ZN(n76) );
  INV_X4 U88 ( .A(A[10]), .ZN(n68) );
  INV_X4 U89 ( .A(A[11]), .ZN(n67) );
  INV_X4 U90 ( .A(A[12]), .ZN(n66) );
  INV_X4 U91 ( .A(A[13]), .ZN(n65) );
  INV_X4 U92 ( .A(A[14]), .ZN(n64) );
  INV_X4 U93 ( .A(A[15]), .ZN(n63) );
  NOR2_X1 U95 ( .A1(n69), .A2(n85), .ZN(\ab[9][9] ) );
  NOR2_X1 U96 ( .A1(n69), .A2(n86), .ZN(\ab[9][8] ) );
  NOR2_X1 U97 ( .A1(n69), .A2(n87), .ZN(\ab[9][7] ) );
  NOR2_X1 U98 ( .A1(n69), .A2(n88), .ZN(\ab[9][6] ) );
  NOR2_X1 U99 ( .A1(n69), .A2(n89), .ZN(\ab[9][5] ) );
  NOR2_X1 U100 ( .A1(n69), .A2(n90), .ZN(\ab[9][4] ) );
  NOR2_X1 U101 ( .A1(n69), .A2(n91), .ZN(\ab[9][3] ) );
  NOR2_X1 U102 ( .A1(n69), .A2(n92), .ZN(\ab[9][2] ) );
  NOR2_X1 U103 ( .A1(n69), .A2(n93), .ZN(\ab[9][1] ) );
  NOR2_X1 U104 ( .A1(n69), .A2(n79), .ZN(\ab[9][15] ) );
  NOR2_X1 U105 ( .A1(n69), .A2(n80), .ZN(\ab[9][14] ) );
  NOR2_X1 U106 ( .A1(n69), .A2(n81), .ZN(\ab[9][13] ) );
  NOR2_X1 U107 ( .A1(n69), .A2(n82), .ZN(\ab[9][12] ) );
  NOR2_X1 U108 ( .A1(n69), .A2(n83), .ZN(\ab[9][11] ) );
  NOR2_X1 U109 ( .A1(n69), .A2(n84), .ZN(\ab[9][10] ) );
  NOR2_X1 U110 ( .A1(n69), .A2(n94), .ZN(\ab[9][0] ) );
  NOR2_X1 U111 ( .A1(n85), .A2(n70), .ZN(\ab[8][9] ) );
  NOR2_X1 U112 ( .A1(n86), .A2(n70), .ZN(\ab[8][8] ) );
  NOR2_X1 U113 ( .A1(n87), .A2(n70), .ZN(\ab[8][7] ) );
  NOR2_X1 U114 ( .A1(n88), .A2(n70), .ZN(\ab[8][6] ) );
  NOR2_X1 U115 ( .A1(n89), .A2(n70), .ZN(\ab[8][5] ) );
  NOR2_X1 U116 ( .A1(n90), .A2(n70), .ZN(\ab[8][4] ) );
  NOR2_X1 U117 ( .A1(n91), .A2(n70), .ZN(\ab[8][3] ) );
  NOR2_X1 U118 ( .A1(n92), .A2(n70), .ZN(\ab[8][2] ) );
  NOR2_X1 U119 ( .A1(n93), .A2(n70), .ZN(\ab[8][1] ) );
  NOR2_X1 U120 ( .A1(n79), .A2(n70), .ZN(\ab[8][15] ) );
  NOR2_X1 U121 ( .A1(n80), .A2(n70), .ZN(\ab[8][14] ) );
  NOR2_X1 U122 ( .A1(n81), .A2(n70), .ZN(\ab[8][13] ) );
  NOR2_X1 U123 ( .A1(n82), .A2(n70), .ZN(\ab[8][12] ) );
  NOR2_X1 U124 ( .A1(n83), .A2(n70), .ZN(\ab[8][11] ) );
  NOR2_X1 U125 ( .A1(n84), .A2(n70), .ZN(\ab[8][10] ) );
  NOR2_X1 U126 ( .A1(n94), .A2(n70), .ZN(\ab[8][0] ) );
  NOR2_X1 U127 ( .A1(n85), .A2(n71), .ZN(\ab[7][9] ) );
  NOR2_X1 U128 ( .A1(n86), .A2(n71), .ZN(\ab[7][8] ) );
  NOR2_X1 U129 ( .A1(n87), .A2(n71), .ZN(\ab[7][7] ) );
  NOR2_X1 U130 ( .A1(n88), .A2(n71), .ZN(\ab[7][6] ) );
  NOR2_X1 U131 ( .A1(n89), .A2(n71), .ZN(\ab[7][5] ) );
  NOR2_X1 U132 ( .A1(n90), .A2(n71), .ZN(\ab[7][4] ) );
  NOR2_X1 U133 ( .A1(n91), .A2(n71), .ZN(\ab[7][3] ) );
  NOR2_X1 U134 ( .A1(n92), .A2(n71), .ZN(\ab[7][2] ) );
  NOR2_X1 U135 ( .A1(n93), .A2(n71), .ZN(\ab[7][1] ) );
  NOR2_X1 U136 ( .A1(n79), .A2(n71), .ZN(\ab[7][15] ) );
  NOR2_X1 U137 ( .A1(n80), .A2(n71), .ZN(\ab[7][14] ) );
  NOR2_X1 U138 ( .A1(n81), .A2(n71), .ZN(\ab[7][13] ) );
  NOR2_X1 U139 ( .A1(n82), .A2(n71), .ZN(\ab[7][12] ) );
  NOR2_X1 U140 ( .A1(n83), .A2(n71), .ZN(\ab[7][11] ) );
  NOR2_X1 U141 ( .A1(n84), .A2(n71), .ZN(\ab[7][10] ) );
  NOR2_X1 U142 ( .A1(n94), .A2(n71), .ZN(\ab[7][0] ) );
  NOR2_X1 U143 ( .A1(n85), .A2(n72), .ZN(\ab[6][9] ) );
  NOR2_X1 U144 ( .A1(n86), .A2(n72), .ZN(\ab[6][8] ) );
  NOR2_X1 U145 ( .A1(n87), .A2(n72), .ZN(\ab[6][7] ) );
  NOR2_X1 U146 ( .A1(n88), .A2(n72), .ZN(\ab[6][6] ) );
  NOR2_X1 U147 ( .A1(n89), .A2(n72), .ZN(\ab[6][5] ) );
  NOR2_X1 U148 ( .A1(n90), .A2(n72), .ZN(\ab[6][4] ) );
  NOR2_X1 U149 ( .A1(n91), .A2(n72), .ZN(\ab[6][3] ) );
  NOR2_X1 U150 ( .A1(n92), .A2(n72), .ZN(\ab[6][2] ) );
  NOR2_X1 U151 ( .A1(n93), .A2(n72), .ZN(\ab[6][1] ) );
  NOR2_X1 U152 ( .A1(n79), .A2(n72), .ZN(\ab[6][15] ) );
  NOR2_X1 U153 ( .A1(n80), .A2(n72), .ZN(\ab[6][14] ) );
  NOR2_X1 U154 ( .A1(n81), .A2(n72), .ZN(\ab[6][13] ) );
  NOR2_X1 U155 ( .A1(n82), .A2(n72), .ZN(\ab[6][12] ) );
  NOR2_X1 U156 ( .A1(n83), .A2(n72), .ZN(\ab[6][11] ) );
  NOR2_X1 U157 ( .A1(n84), .A2(n72), .ZN(\ab[6][10] ) );
  NOR2_X1 U158 ( .A1(n94), .A2(n72), .ZN(\ab[6][0] ) );
  NOR2_X1 U159 ( .A1(n85), .A2(n73), .ZN(\ab[5][9] ) );
  NOR2_X1 U160 ( .A1(n86), .A2(n73), .ZN(\ab[5][8] ) );
  NOR2_X1 U161 ( .A1(n87), .A2(n73), .ZN(\ab[5][7] ) );
  NOR2_X1 U162 ( .A1(n88), .A2(n73), .ZN(\ab[5][6] ) );
  NOR2_X1 U163 ( .A1(n89), .A2(n73), .ZN(\ab[5][5] ) );
  NOR2_X1 U164 ( .A1(n90), .A2(n73), .ZN(\ab[5][4] ) );
  NOR2_X1 U165 ( .A1(n91), .A2(n73), .ZN(\ab[5][3] ) );
  NOR2_X1 U166 ( .A1(n92), .A2(n73), .ZN(\ab[5][2] ) );
  NOR2_X1 U167 ( .A1(n93), .A2(n73), .ZN(\ab[5][1] ) );
  NOR2_X1 U168 ( .A1(n79), .A2(n73), .ZN(\ab[5][15] ) );
  NOR2_X1 U169 ( .A1(n80), .A2(n73), .ZN(\ab[5][14] ) );
  NOR2_X1 U170 ( .A1(n81), .A2(n73), .ZN(\ab[5][13] ) );
  NOR2_X1 U171 ( .A1(n82), .A2(n73), .ZN(\ab[5][12] ) );
  NOR2_X1 U172 ( .A1(n83), .A2(n73), .ZN(\ab[5][11] ) );
  NOR2_X1 U173 ( .A1(n84), .A2(n73), .ZN(\ab[5][10] ) );
  NOR2_X1 U174 ( .A1(n94), .A2(n73), .ZN(\ab[5][0] ) );
  NOR2_X1 U175 ( .A1(n85), .A2(n74), .ZN(\ab[4][9] ) );
  NOR2_X1 U176 ( .A1(n86), .A2(n74), .ZN(\ab[4][8] ) );
  NOR2_X1 U177 ( .A1(n87), .A2(n74), .ZN(\ab[4][7] ) );
  NOR2_X1 U178 ( .A1(n88), .A2(n74), .ZN(\ab[4][6] ) );
  NOR2_X1 U179 ( .A1(n89), .A2(n74), .ZN(\ab[4][5] ) );
  NOR2_X1 U180 ( .A1(n90), .A2(n74), .ZN(\ab[4][4] ) );
  NOR2_X1 U181 ( .A1(n91), .A2(n74), .ZN(\ab[4][3] ) );
  NOR2_X1 U182 ( .A1(n92), .A2(n74), .ZN(\ab[4][2] ) );
  NOR2_X1 U183 ( .A1(n93), .A2(n74), .ZN(\ab[4][1] ) );
  NOR2_X1 U184 ( .A1(n79), .A2(n74), .ZN(\ab[4][15] ) );
  NOR2_X1 U185 ( .A1(n80), .A2(n74), .ZN(\ab[4][14] ) );
  NOR2_X1 U186 ( .A1(n81), .A2(n74), .ZN(\ab[4][13] ) );
  NOR2_X1 U187 ( .A1(n82), .A2(n74), .ZN(\ab[4][12] ) );
  NOR2_X1 U188 ( .A1(n83), .A2(n74), .ZN(\ab[4][11] ) );
  NOR2_X1 U189 ( .A1(n84), .A2(n74), .ZN(\ab[4][10] ) );
  NOR2_X1 U190 ( .A1(n94), .A2(n74), .ZN(\ab[4][0] ) );
  NOR2_X1 U191 ( .A1(n85), .A2(n75), .ZN(\ab[3][9] ) );
  NOR2_X1 U192 ( .A1(n86), .A2(n75), .ZN(\ab[3][8] ) );
  NOR2_X1 U193 ( .A1(n87), .A2(n75), .ZN(\ab[3][7] ) );
  NOR2_X1 U194 ( .A1(n88), .A2(n75), .ZN(\ab[3][6] ) );
  NOR2_X1 U195 ( .A1(n89), .A2(n75), .ZN(\ab[3][5] ) );
  NOR2_X1 U196 ( .A1(n90), .A2(n75), .ZN(\ab[3][4] ) );
  NOR2_X1 U197 ( .A1(n91), .A2(n75), .ZN(\ab[3][3] ) );
  NOR2_X1 U198 ( .A1(n92), .A2(n75), .ZN(\ab[3][2] ) );
  NOR2_X1 U199 ( .A1(n93), .A2(n75), .ZN(\ab[3][1] ) );
  NOR2_X1 U200 ( .A1(n79), .A2(n75), .ZN(\ab[3][15] ) );
  NOR2_X1 U201 ( .A1(n80), .A2(n75), .ZN(\ab[3][14] ) );
  NOR2_X1 U202 ( .A1(n81), .A2(n75), .ZN(\ab[3][13] ) );
  NOR2_X1 U203 ( .A1(n82), .A2(n75), .ZN(\ab[3][12] ) );
  NOR2_X1 U204 ( .A1(n83), .A2(n75), .ZN(\ab[3][11] ) );
  NOR2_X1 U205 ( .A1(n84), .A2(n75), .ZN(\ab[3][10] ) );
  NOR2_X1 U206 ( .A1(n94), .A2(n75), .ZN(\ab[3][0] ) );
  NOR2_X1 U207 ( .A1(n85), .A2(n76), .ZN(\ab[2][9] ) );
  NOR2_X1 U208 ( .A1(n86), .A2(n76), .ZN(\ab[2][8] ) );
  NOR2_X1 U209 ( .A1(n87), .A2(n76), .ZN(\ab[2][7] ) );
  NOR2_X1 U210 ( .A1(n88), .A2(n76), .ZN(\ab[2][6] ) );
  NOR2_X1 U211 ( .A1(n89), .A2(n76), .ZN(\ab[2][5] ) );
  NOR2_X1 U212 ( .A1(n90), .A2(n76), .ZN(\ab[2][4] ) );
  NOR2_X1 U213 ( .A1(n91), .A2(n76), .ZN(\ab[2][3] ) );
  NOR2_X1 U214 ( .A1(n92), .A2(n76), .ZN(\ab[2][2] ) );
  NOR2_X1 U215 ( .A1(n93), .A2(n76), .ZN(\ab[2][1] ) );
  NOR2_X1 U216 ( .A1(n79), .A2(n76), .ZN(\ab[2][15] ) );
  NOR2_X1 U217 ( .A1(n80), .A2(n76), .ZN(\ab[2][14] ) );
  NOR2_X1 U218 ( .A1(n81), .A2(n76), .ZN(\ab[2][13] ) );
  NOR2_X1 U219 ( .A1(n82), .A2(n76), .ZN(\ab[2][12] ) );
  NOR2_X1 U220 ( .A1(n83), .A2(n76), .ZN(\ab[2][11] ) );
  NOR2_X1 U221 ( .A1(n84), .A2(n76), .ZN(\ab[2][10] ) );
  NOR2_X1 U222 ( .A1(n94), .A2(n76), .ZN(\ab[2][0] ) );
  NOR2_X1 U223 ( .A1(n85), .A2(n77), .ZN(\ab[1][9] ) );
  NOR2_X1 U224 ( .A1(n86), .A2(n77), .ZN(\ab[1][8] ) );
  NOR2_X1 U225 ( .A1(n87), .A2(n77), .ZN(\ab[1][7] ) );
  NOR2_X1 U226 ( .A1(n88), .A2(n77), .ZN(\ab[1][6] ) );
  NOR2_X1 U227 ( .A1(n89), .A2(n77), .ZN(\ab[1][5] ) );
  NOR2_X1 U228 ( .A1(n90), .A2(n77), .ZN(\ab[1][4] ) );
  NOR2_X1 U229 ( .A1(n91), .A2(n77), .ZN(\ab[1][3] ) );
  NOR2_X1 U230 ( .A1(n92), .A2(n77), .ZN(\ab[1][2] ) );
  NOR2_X1 U231 ( .A1(n93), .A2(n77), .ZN(\ab[1][1] ) );
  NOR2_X1 U232 ( .A1(n79), .A2(n77), .ZN(\ab[1][15] ) );
  NOR2_X1 U233 ( .A1(n80), .A2(n77), .ZN(\ab[1][14] ) );
  NOR2_X1 U234 ( .A1(n81), .A2(n77), .ZN(\ab[1][13] ) );
  NOR2_X1 U235 ( .A1(n82), .A2(n77), .ZN(\ab[1][12] ) );
  NOR2_X1 U236 ( .A1(n83), .A2(n77), .ZN(\ab[1][11] ) );
  NOR2_X1 U237 ( .A1(n84), .A2(n77), .ZN(\ab[1][10] ) );
  NOR2_X1 U238 ( .A1(n94), .A2(n77), .ZN(\ab[1][0] ) );
  NOR2_X1 U239 ( .A1(n85), .A2(n63), .ZN(\ab[15][9] ) );
  NOR2_X1 U240 ( .A1(n86), .A2(n63), .ZN(\ab[15][8] ) );
  NOR2_X1 U241 ( .A1(n87), .A2(n63), .ZN(\ab[15][7] ) );
  NOR2_X1 U242 ( .A1(n88), .A2(n63), .ZN(\ab[15][6] ) );
  NOR2_X1 U243 ( .A1(n89), .A2(n63), .ZN(\ab[15][5] ) );
  NOR2_X1 U244 ( .A1(n90), .A2(n63), .ZN(\ab[15][4] ) );
  NOR2_X1 U245 ( .A1(n91), .A2(n63), .ZN(\ab[15][3] ) );
  NOR2_X1 U246 ( .A1(n92), .A2(n63), .ZN(\ab[15][2] ) );
  NOR2_X1 U247 ( .A1(n93), .A2(n63), .ZN(\ab[15][1] ) );
  NOR2_X1 U248 ( .A1(n79), .A2(n63), .ZN(\ab[15][15] ) );
  NOR2_X1 U249 ( .A1(n80), .A2(n63), .ZN(\ab[15][14] ) );
  NOR2_X1 U250 ( .A1(n81), .A2(n63), .ZN(\ab[15][13] ) );
  NOR2_X1 U251 ( .A1(n82), .A2(n63), .ZN(\ab[15][12] ) );
  NOR2_X1 U252 ( .A1(n83), .A2(n63), .ZN(\ab[15][11] ) );
  NOR2_X1 U253 ( .A1(n84), .A2(n63), .ZN(\ab[15][10] ) );
  NOR2_X1 U254 ( .A1(n94), .A2(n63), .ZN(\ab[15][0] ) );
  NOR2_X1 U255 ( .A1(n85), .A2(n64), .ZN(\ab[14][9] ) );
  NOR2_X1 U256 ( .A1(n86), .A2(n64), .ZN(\ab[14][8] ) );
  NOR2_X1 U257 ( .A1(n87), .A2(n64), .ZN(\ab[14][7] ) );
  NOR2_X1 U258 ( .A1(n88), .A2(n64), .ZN(\ab[14][6] ) );
  NOR2_X1 U259 ( .A1(n89), .A2(n64), .ZN(\ab[14][5] ) );
  NOR2_X1 U260 ( .A1(n90), .A2(n64), .ZN(\ab[14][4] ) );
  NOR2_X1 U261 ( .A1(n91), .A2(n64), .ZN(\ab[14][3] ) );
  NOR2_X1 U262 ( .A1(n92), .A2(n64), .ZN(\ab[14][2] ) );
  NOR2_X1 U263 ( .A1(n93), .A2(n64), .ZN(\ab[14][1] ) );
  NOR2_X1 U264 ( .A1(n79), .A2(n64), .ZN(\ab[14][15] ) );
  NOR2_X1 U265 ( .A1(n80), .A2(n64), .ZN(\ab[14][14] ) );
  NOR2_X1 U266 ( .A1(n81), .A2(n64), .ZN(\ab[14][13] ) );
  NOR2_X1 U267 ( .A1(n82), .A2(n64), .ZN(\ab[14][12] ) );
  NOR2_X1 U268 ( .A1(n83), .A2(n64), .ZN(\ab[14][11] ) );
  NOR2_X1 U269 ( .A1(n84), .A2(n64), .ZN(\ab[14][10] ) );
  NOR2_X1 U270 ( .A1(n94), .A2(n64), .ZN(\ab[14][0] ) );
  NOR2_X1 U271 ( .A1(n85), .A2(n65), .ZN(\ab[13][9] ) );
  NOR2_X1 U272 ( .A1(n86), .A2(n65), .ZN(\ab[13][8] ) );
  NOR2_X1 U273 ( .A1(n87), .A2(n65), .ZN(\ab[13][7] ) );
  NOR2_X1 U274 ( .A1(n88), .A2(n65), .ZN(\ab[13][6] ) );
  NOR2_X1 U275 ( .A1(n89), .A2(n65), .ZN(\ab[13][5] ) );
  NOR2_X1 U276 ( .A1(n90), .A2(n65), .ZN(\ab[13][4] ) );
  NOR2_X1 U277 ( .A1(n91), .A2(n65), .ZN(\ab[13][3] ) );
  NOR2_X1 U278 ( .A1(n92), .A2(n65), .ZN(\ab[13][2] ) );
  NOR2_X1 U279 ( .A1(n93), .A2(n65), .ZN(\ab[13][1] ) );
  NOR2_X1 U280 ( .A1(n79), .A2(n65), .ZN(\ab[13][15] ) );
  NOR2_X1 U281 ( .A1(n80), .A2(n65), .ZN(\ab[13][14] ) );
  NOR2_X1 U282 ( .A1(n81), .A2(n65), .ZN(\ab[13][13] ) );
  NOR2_X1 U283 ( .A1(n82), .A2(n65), .ZN(\ab[13][12] ) );
  NOR2_X1 U284 ( .A1(n83), .A2(n65), .ZN(\ab[13][11] ) );
  NOR2_X1 U285 ( .A1(n84), .A2(n65), .ZN(\ab[13][10] ) );
  NOR2_X1 U286 ( .A1(n94), .A2(n65), .ZN(\ab[13][0] ) );
  NOR2_X1 U287 ( .A1(n85), .A2(n66), .ZN(\ab[12][9] ) );
  NOR2_X1 U288 ( .A1(n86), .A2(n66), .ZN(\ab[12][8] ) );
  NOR2_X1 U289 ( .A1(n87), .A2(n66), .ZN(\ab[12][7] ) );
  NOR2_X1 U290 ( .A1(n88), .A2(n66), .ZN(\ab[12][6] ) );
  NOR2_X1 U291 ( .A1(n89), .A2(n66), .ZN(\ab[12][5] ) );
  NOR2_X1 U292 ( .A1(n90), .A2(n66), .ZN(\ab[12][4] ) );
  NOR2_X1 U293 ( .A1(n91), .A2(n66), .ZN(\ab[12][3] ) );
  NOR2_X1 U294 ( .A1(n92), .A2(n66), .ZN(\ab[12][2] ) );
  NOR2_X1 U295 ( .A1(n93), .A2(n66), .ZN(\ab[12][1] ) );
  NOR2_X1 U296 ( .A1(n79), .A2(n66), .ZN(\ab[12][15] ) );
  NOR2_X1 U297 ( .A1(n80), .A2(n66), .ZN(\ab[12][14] ) );
  NOR2_X1 U298 ( .A1(n81), .A2(n66), .ZN(\ab[12][13] ) );
  NOR2_X1 U299 ( .A1(n82), .A2(n66), .ZN(\ab[12][12] ) );
  NOR2_X1 U300 ( .A1(n83), .A2(n66), .ZN(\ab[12][11] ) );
  NOR2_X1 U301 ( .A1(n84), .A2(n66), .ZN(\ab[12][10] ) );
  NOR2_X1 U302 ( .A1(n94), .A2(n66), .ZN(\ab[12][0] ) );
  NOR2_X1 U303 ( .A1(n85), .A2(n67), .ZN(\ab[11][9] ) );
  NOR2_X1 U304 ( .A1(n86), .A2(n67), .ZN(\ab[11][8] ) );
  NOR2_X1 U305 ( .A1(n87), .A2(n67), .ZN(\ab[11][7] ) );
  NOR2_X1 U306 ( .A1(n88), .A2(n67), .ZN(\ab[11][6] ) );
  NOR2_X1 U307 ( .A1(n89), .A2(n67), .ZN(\ab[11][5] ) );
  NOR2_X1 U308 ( .A1(n90), .A2(n67), .ZN(\ab[11][4] ) );
  NOR2_X1 U309 ( .A1(n91), .A2(n67), .ZN(\ab[11][3] ) );
  NOR2_X1 U310 ( .A1(n92), .A2(n67), .ZN(\ab[11][2] ) );
  NOR2_X1 U311 ( .A1(n93), .A2(n67), .ZN(\ab[11][1] ) );
  NOR2_X1 U312 ( .A1(n79), .A2(n67), .ZN(\ab[11][15] ) );
  NOR2_X1 U313 ( .A1(n80), .A2(n67), .ZN(\ab[11][14] ) );
  NOR2_X1 U314 ( .A1(n81), .A2(n67), .ZN(\ab[11][13] ) );
  NOR2_X1 U315 ( .A1(n82), .A2(n67), .ZN(\ab[11][12] ) );
  NOR2_X1 U316 ( .A1(n83), .A2(n67), .ZN(\ab[11][11] ) );
  NOR2_X1 U317 ( .A1(n84), .A2(n67), .ZN(\ab[11][10] ) );
  NOR2_X1 U318 ( .A1(n94), .A2(n67), .ZN(\ab[11][0] ) );
  NOR2_X1 U319 ( .A1(n85), .A2(n68), .ZN(\ab[10][9] ) );
  NOR2_X1 U320 ( .A1(n86), .A2(n68), .ZN(\ab[10][8] ) );
  NOR2_X1 U321 ( .A1(n87), .A2(n68), .ZN(\ab[10][7] ) );
  NOR2_X1 U322 ( .A1(n88), .A2(n68), .ZN(\ab[10][6] ) );
  NOR2_X1 U323 ( .A1(n89), .A2(n68), .ZN(\ab[10][5] ) );
  NOR2_X1 U324 ( .A1(n90), .A2(n68), .ZN(\ab[10][4] ) );
  NOR2_X1 U325 ( .A1(n91), .A2(n68), .ZN(\ab[10][3] ) );
  NOR2_X1 U326 ( .A1(n92), .A2(n68), .ZN(\ab[10][2] ) );
  NOR2_X1 U327 ( .A1(n93), .A2(n68), .ZN(\ab[10][1] ) );
  NOR2_X1 U328 ( .A1(n79), .A2(n68), .ZN(\ab[10][15] ) );
  NOR2_X1 U329 ( .A1(n80), .A2(n68), .ZN(\ab[10][14] ) );
  NOR2_X1 U330 ( .A1(n81), .A2(n68), .ZN(\ab[10][13] ) );
  NOR2_X1 U331 ( .A1(n82), .A2(n68), .ZN(\ab[10][12] ) );
  NOR2_X1 U332 ( .A1(n83), .A2(n68), .ZN(\ab[10][11] ) );
  NOR2_X1 U333 ( .A1(n84), .A2(n68), .ZN(\ab[10][10] ) );
  NOR2_X1 U334 ( .A1(n94), .A2(n68), .ZN(\ab[10][0] ) );
  NOR2_X1 U335 ( .A1(n85), .A2(n78), .ZN(\ab[0][9] ) );
  NOR2_X1 U336 ( .A1(n86), .A2(n78), .ZN(\ab[0][8] ) );
  NOR2_X1 U337 ( .A1(n87), .A2(n78), .ZN(\ab[0][7] ) );
  NOR2_X1 U338 ( .A1(n88), .A2(n78), .ZN(\ab[0][6] ) );
  NOR2_X1 U339 ( .A1(n89), .A2(n78), .ZN(\ab[0][5] ) );
  NOR2_X1 U340 ( .A1(n90), .A2(n78), .ZN(\ab[0][4] ) );
  NOR2_X1 U341 ( .A1(n91), .A2(n78), .ZN(\ab[0][3] ) );
  NOR2_X1 U342 ( .A1(n92), .A2(n78), .ZN(\ab[0][2] ) );
  NOR2_X1 U343 ( .A1(n93), .A2(n78), .ZN(\ab[0][1] ) );
  NOR2_X1 U344 ( .A1(n79), .A2(n78), .ZN(\ab[0][15] ) );
  NOR2_X1 U345 ( .A1(n80), .A2(n78), .ZN(\ab[0][14] ) );
  NOR2_X1 U346 ( .A1(n81), .A2(n78), .ZN(\ab[0][13] ) );
  NOR2_X1 U347 ( .A1(n82), .A2(n78), .ZN(\ab[0][12] ) );
  NOR2_X1 U348 ( .A1(n83), .A2(n78), .ZN(\ab[0][11] ) );
  NOR2_X1 U349 ( .A1(n84), .A2(n78), .ZN(\ab[0][10] ) );
  NOR2_X1 U350 ( .A1(n94), .A2(n78), .ZN(PRODUCT[0]) );
  multiplier_DW01_add_6 FS_1 ( .A({1'b0, n17, n25, n18, n26, n19, n27, n20, 
        n28, n21, n29, n22, n30, n23, n24, n61, \SUMB[15][0] , \A1[12] , 
        \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , 
        \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({n62, n46, n53, n47, 
        n54, n48, n55, n49, n56, n50, n57, n51, n58, n52, n59, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .CI(1'b0), .SUM(PRODUCT[31:2]) );
endmodule


module multiplier ( clk, reset, mul, a, b, done, working, result );
  input [0:31] a;
  input [0:31] b;
  output [0:63] result;
  input clk, reset, mul;
  output done, working;
  wire   N14, N15, N16, N43, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93,
         N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160,
         N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171,
         N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182,
         N183, N184, N185, N218, N219, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N314, N315, N316, N317, N318, N319, N320, N321, N322,
         N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333,
         N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344,
         N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366,
         N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377,
         N379, N380, N381, N382, N383, N384, N385, N386, N387, N388, N389,
         N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400,
         N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N412,
         N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, N423,
         N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434,
         N435, N436, N437, N438, N439, N440, N441, N442, N443, N445, N446,
         N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457,
         N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468,
         N469, N470, N471, N472, N473, N474, N475, N476, n33, n34, n35, n36,
         N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288,
         N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277,
         N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266,
         N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255,
         N254, N253, N252, N251, N250, N217, N216, N215, N214, N213, N212,
         N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201,
         N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190,
         N189, N188, N187, N186, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n37, n39, n40;
  wire   [0:2] CurrentState;
  wire   [0:31] L;
  wire   [0:31] Z;
  wire   [0:31] H;
  wire   [0:31] P1;
  wire   [0:31] P;
  wire   [0:31] P2;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46;

  AND2_X2 U9 ( .A1(N185), .A2(n39), .ZN(N476) );
  AND2_X2 U10 ( .A1(N184), .A2(n39), .ZN(N475) );
  AND2_X2 U11 ( .A1(N183), .A2(n39), .ZN(N474) );
  AND2_X2 U12 ( .A1(N182), .A2(n39), .ZN(N473) );
  AND2_X2 U13 ( .A1(N181), .A2(n39), .ZN(N472) );
  AND2_X2 U14 ( .A1(N180), .A2(n39), .ZN(N471) );
  AND2_X2 U15 ( .A1(N179), .A2(n39), .ZN(N470) );
  AND2_X2 U16 ( .A1(N178), .A2(n39), .ZN(N469) );
  AND2_X2 U17 ( .A1(N177), .A2(n39), .ZN(N468) );
  AND2_X2 U18 ( .A1(N176), .A2(n39), .ZN(N467) );
  AND2_X2 U19 ( .A1(N175), .A2(n11), .ZN(N466) );
  AND2_X2 U20 ( .A1(N174), .A2(n11), .ZN(N465) );
  AND2_X2 U21 ( .A1(N173), .A2(n11), .ZN(N464) );
  AND2_X2 U22 ( .A1(N172), .A2(n11), .ZN(N463) );
  AND2_X2 U23 ( .A1(N171), .A2(n11), .ZN(N462) );
  AND2_X2 U24 ( .A1(N170), .A2(n11), .ZN(N461) );
  AND2_X2 U25 ( .A1(N169), .A2(n11), .ZN(N460) );
  AND2_X2 U26 ( .A1(N168), .A2(n11), .ZN(N459) );
  AND2_X2 U27 ( .A1(N167), .A2(n11), .ZN(N458) );
  AND2_X2 U28 ( .A1(N166), .A2(n11), .ZN(N457) );
  AND2_X2 U29 ( .A1(N165), .A2(n11), .ZN(N456) );
  AND2_X2 U30 ( .A1(N164), .A2(n11), .ZN(N455) );
  AND2_X2 U31 ( .A1(N163), .A2(n11), .ZN(N454) );
  AND2_X2 U32 ( .A1(N162), .A2(n11), .ZN(N453) );
  AND2_X2 U33 ( .A1(N161), .A2(n11), .ZN(N452) );
  AND2_X2 U34 ( .A1(N160), .A2(n11), .ZN(N451) );
  AND2_X2 U35 ( .A1(N159), .A2(n11), .ZN(N450) );
  AND2_X2 U36 ( .A1(N158), .A2(n11), .ZN(N449) );
  AND2_X2 U37 ( .A1(N157), .A2(n11), .ZN(N448) );
  AND2_X2 U38 ( .A1(N156), .A2(n11), .ZN(N447) );
  AND2_X2 U39 ( .A1(N155), .A2(n11), .ZN(N446) );
  AND2_X2 U40 ( .A1(N154), .A2(n11), .ZN(N445) );
  AND2_X2 U42 ( .A1(N249), .A2(n12), .ZN(N443) );
  AND2_X2 U43 ( .A1(N248), .A2(n12), .ZN(N442) );
  AND2_X2 U44 ( .A1(N247), .A2(n12), .ZN(N441) );
  AND2_X2 U45 ( .A1(N246), .A2(n12), .ZN(N440) );
  AND2_X2 U46 ( .A1(N245), .A2(n12), .ZN(N439) );
  AND2_X2 U47 ( .A1(N244), .A2(n12), .ZN(N438) );
  AND2_X2 U48 ( .A1(N243), .A2(n12), .ZN(N437) );
  AND2_X2 U49 ( .A1(N242), .A2(n12), .ZN(N436) );
  AND2_X2 U50 ( .A1(N241), .A2(n12), .ZN(N435) );
  AND2_X2 U51 ( .A1(N240), .A2(n12), .ZN(N434) );
  AND2_X2 U52 ( .A1(N239), .A2(n12), .ZN(N433) );
  AND2_X2 U53 ( .A1(N238), .A2(n13), .ZN(N432) );
  AND2_X2 U54 ( .A1(N237), .A2(n13), .ZN(N431) );
  AND2_X2 U55 ( .A1(N236), .A2(n13), .ZN(N430) );
  AND2_X2 U56 ( .A1(N235), .A2(n13), .ZN(N429) );
  AND2_X2 U57 ( .A1(N234), .A2(n13), .ZN(N428) );
  AND2_X2 U58 ( .A1(N233), .A2(n13), .ZN(N427) );
  AND2_X2 U59 ( .A1(N232), .A2(n13), .ZN(N426) );
  AND2_X2 U60 ( .A1(N231), .A2(n13), .ZN(N425) );
  AND2_X2 U61 ( .A1(N230), .A2(n13), .ZN(N424) );
  AND2_X2 U62 ( .A1(N229), .A2(n13), .ZN(N423) );
  AND2_X2 U63 ( .A1(N228), .A2(n13), .ZN(N422) );
  AND2_X2 U64 ( .A1(N227), .A2(n14), .ZN(N421) );
  AND2_X2 U65 ( .A1(N226), .A2(n14), .ZN(N420) );
  AND2_X2 U66 ( .A1(N225), .A2(n14), .ZN(N419) );
  AND2_X2 U67 ( .A1(N224), .A2(n14), .ZN(N418) );
  AND2_X2 U68 ( .A1(N223), .A2(n14), .ZN(N417) );
  AND2_X2 U69 ( .A1(N222), .A2(n14), .ZN(N416) );
  AND2_X2 U70 ( .A1(N221), .A2(n14), .ZN(N415) );
  AND2_X2 U71 ( .A1(N220), .A2(n14), .ZN(N414) );
  AND2_X2 U72 ( .A1(N219), .A2(n14), .ZN(N413) );
  AND2_X2 U73 ( .A1(N218), .A2(n14), .ZN(N412) );
  AND2_X2 U75 ( .A1(N153), .A2(n17), .ZN(N410) );
  AND2_X2 U76 ( .A1(N152), .A2(n17), .ZN(N409) );
  AND2_X2 U77 ( .A1(N151), .A2(n17), .ZN(N408) );
  AND2_X2 U78 ( .A1(N150), .A2(n17), .ZN(N407) );
  AND2_X2 U79 ( .A1(N149), .A2(n17), .ZN(N406) );
  AND2_X2 U80 ( .A1(N148), .A2(n17), .ZN(N405) );
  AND2_X2 U81 ( .A1(N147), .A2(n17), .ZN(N404) );
  AND2_X2 U82 ( .A1(N146), .A2(n17), .ZN(N403) );
  AND2_X2 U83 ( .A1(N145), .A2(n17), .ZN(N402) );
  AND2_X2 U84 ( .A1(N144), .A2(n17), .ZN(N401) );
  AND2_X2 U85 ( .A1(N143), .A2(n16), .ZN(N400) );
  AND2_X2 U86 ( .A1(N142), .A2(n16), .ZN(N399) );
  AND2_X2 U87 ( .A1(N141), .A2(n16), .ZN(N398) );
  AND2_X2 U88 ( .A1(N140), .A2(n16), .ZN(N397) );
  AND2_X2 U89 ( .A1(N139), .A2(n16), .ZN(N396) );
  AND2_X2 U90 ( .A1(N138), .A2(n16), .ZN(N395) );
  AND2_X2 U91 ( .A1(N137), .A2(n16), .ZN(N394) );
  AND2_X2 U92 ( .A1(N136), .A2(n16), .ZN(N393) );
  AND2_X2 U93 ( .A1(N135), .A2(n16), .ZN(N392) );
  AND2_X2 U94 ( .A1(N134), .A2(n16), .ZN(N391) );
  AND2_X2 U95 ( .A1(N133), .A2(n16), .ZN(N390) );
  AND2_X2 U96 ( .A1(N132), .A2(n16), .ZN(N389) );
  AND2_X2 U97 ( .A1(N131), .A2(n16), .ZN(N388) );
  AND2_X2 U98 ( .A1(N130), .A2(n16), .ZN(N387) );
  AND2_X2 U99 ( .A1(N129), .A2(n16), .ZN(N386) );
  AND2_X2 U100 ( .A1(N128), .A2(n16), .ZN(N385) );
  AND2_X2 U101 ( .A1(N127), .A2(n16), .ZN(N384) );
  AND2_X2 U102 ( .A1(N126), .A2(n16), .ZN(N383) );
  AND2_X2 U103 ( .A1(N125), .A2(n16), .ZN(N382) );
  AND2_X2 U104 ( .A1(N124), .A2(n16), .ZN(N381) );
  AND2_X2 U105 ( .A1(N123), .A2(n16), .ZN(N380) );
  AND2_X2 U106 ( .A1(N122), .A2(n16), .ZN(N379) );
  DFF_X2 \CurrentState_reg[2]  ( .D(N14), .CK(clk), .Q(CurrentState[2]), .QN(
        n4) );
  DFF_X2 \CurrentState_reg[0]  ( .D(N16), .CK(clk), .Q(CurrentState[0]), .QN(
        n5) );
  DFF_X2 \CurrentState_reg[1]  ( .D(N15), .CK(clk), .Q(CurrentState[1]) );
  DLH_X2 \P2_reg[15]  ( .G(n17), .D(N121), .Q(P2[15]) );
  DLH_X2 \P2_reg[16]  ( .G(n17), .D(N120), .Q(P2[16]) );
  DLH_X2 \P2_reg[17]  ( .G(n15), .D(N119), .Q(P2[17]) );
  DLH_X2 \P2_reg[18]  ( .G(n15), .D(N118), .Q(P2[18]) );
  DLH_X2 \P2_reg[19]  ( .G(n15), .D(N117), .Q(P2[19]) );
  DLH_X2 \P2_reg[20]  ( .G(n15), .D(N116), .Q(P2[20]) );
  DLH_X2 \P2_reg[21]  ( .G(n15), .D(N115), .Q(P2[21]) );
  DLH_X2 \P2_reg[22]  ( .G(n15), .D(N114), .Q(P2[22]) );
  DLH_X2 \P2_reg[23]  ( .G(n15), .D(N113), .Q(P2[23]) );
  DLH_X2 \P2_reg[24]  ( .G(n15), .D(N112), .Q(P2[24]) );
  DLH_X2 \P2_reg[25]  ( .G(n15), .D(N111), .Q(P2[25]) );
  DLH_X2 \P2_reg[26]  ( .G(n15), .D(N110), .Q(P2[26]) );
  DLH_X2 \P2_reg[27]  ( .G(n15), .D(N109), .Q(P2[27]) );
  DLH_X2 \P2_reg[28]  ( .G(n15), .D(N108), .Q(P2[28]) );
  DLH_X2 \P2_reg[29]  ( .G(n15), .D(N107), .Q(P2[29]) );
  DLH_X2 \P2_reg[30]  ( .G(n15), .D(N106), .Q(P2[30]) );
  DLH_X2 \P2_reg[31]  ( .G(n15), .D(N105), .Q(P2[31]) );
  DLH_X2 done_reg ( .G(n8), .D(n18), .Q(done) );
  DLH_X2 \P_reg[0]  ( .G(n22), .D(N476), .Q(P[0]) );
  DLH_X2 \P_reg[1]  ( .G(n22), .D(N475), .Q(P[1]) );
  DLH_X2 \P_reg[2]  ( .G(n22), .D(N474), .Q(P[2]) );
  DLH_X2 \P_reg[3]  ( .G(n22), .D(N473), .Q(P[3]) );
  DLH_X2 \P_reg[4]  ( .G(n22), .D(N472), .Q(P[4]) );
  DLH_X2 \P_reg[5]  ( .G(n22), .D(N471), .Q(P[5]) );
  DLH_X2 \P_reg[6]  ( .G(n22), .D(N470), .Q(P[6]) );
  DLH_X2 \P_reg[7]  ( .G(n22), .D(N469), .Q(P[7]) );
  DLH_X2 \P_reg[8]  ( .G(n22), .D(N468), .Q(P[8]) );
  DLH_X2 \P_reg[9]  ( .G(n22), .D(N467), .Q(P[9]) );
  DLH_X2 \P_reg[10]  ( .G(n22), .D(N466), .Q(P[10]) );
  DLH_X2 \P_reg[11]  ( .G(n23), .D(N465), .Q(P[11]) );
  DLH_X2 \P_reg[12]  ( .G(n23), .D(N464), .Q(P[12]) );
  DLH_X2 \P_reg[13]  ( .G(n23), .D(N463), .Q(P[13]) );
  DLH_X2 \P_reg[14]  ( .G(n23), .D(N462), .Q(P[14]) );
  DLH_X2 \P_reg[15]  ( .G(n23), .D(N461), .Q(P[15]) );
  DLH_X2 \P_reg[16]  ( .G(n23), .D(N460), .Q(P[16]) );
  DLH_X2 \P_reg[17]  ( .G(n23), .D(N459), .Q(P[17]) );
  DLH_X2 \P_reg[18]  ( .G(n23), .D(N458), .Q(P[18]) );
  DLH_X2 \P_reg[19]  ( .G(n23), .D(N457), .Q(P[19]) );
  DLH_X2 \P_reg[20]  ( .G(n23), .D(N456), .Q(P[20]) );
  DLH_X2 \P_reg[21]  ( .G(n23), .D(N455), .Q(P[21]) );
  DLH_X2 \P_reg[22]  ( .G(n24), .D(N454), .Q(P[22]) );
  DLH_X2 \P_reg[23]  ( .G(n24), .D(N453), .Q(P[23]) );
  DLH_X2 \P_reg[24]  ( .G(n24), .D(N452), .Q(P[24]) );
  DLH_X2 \P_reg[25]  ( .G(n24), .D(N451), .Q(P[25]) );
  DLH_X2 \P_reg[26]  ( .G(n24), .D(N450), .Q(P[26]) );
  DLH_X2 \P_reg[27]  ( .G(n24), .D(N449), .Q(P[27]) );
  DLH_X2 \P_reg[28]  ( .G(n24), .D(N448), .Q(P[28]) );
  DLH_X2 \P_reg[29]  ( .G(n24), .D(N447), .Q(P[29]) );
  DLH_X2 \P_reg[30]  ( .G(n24), .D(N446), .Q(P[30]) );
  DLH_X2 \P_reg[31]  ( .G(n24), .D(N445), .Q(P[31]) );
  DLH_X2 \P1_reg[15]  ( .G(N43), .D(N104), .Q(P1[15]) );
  DLH_X2 \P1_reg[16]  ( .G(N43), .D(N103), .Q(P1[16]) );
  DLH_X2 \P1_reg[17]  ( .G(N43), .D(N102), .Q(P1[17]) );
  DLH_X2 \P1_reg[18]  ( .G(N43), .D(N101), .Q(P1[18]) );
  DLH_X2 \P1_reg[19]  ( .G(N43), .D(N100), .Q(P1[19]) );
  DLH_X2 \P1_reg[20]  ( .G(N43), .D(N99), .Q(P1[20]) );
  DLH_X2 \P1_reg[21]  ( .G(N43), .D(N98), .Q(P1[21]) );
  DLH_X2 \P1_reg[22]  ( .G(N43), .D(N97), .Q(P1[22]) );
  DLH_X2 \P1_reg[23]  ( .G(N43), .D(N96), .Q(P1[23]) );
  DLH_X2 \P1_reg[24]  ( .G(N43), .D(N95), .Q(P1[24]) );
  DLH_X2 \P1_reg[25]  ( .G(N43), .D(N94), .Q(P1[25]) );
  DLH_X2 \P1_reg[26]  ( .G(N43), .D(N93), .Q(P1[26]) );
  DLH_X2 \P1_reg[27]  ( .G(N43), .D(N92), .Q(P1[27]) );
  DLH_X2 \P1_reg[28]  ( .G(N43), .D(N91), .Q(P1[28]) );
  DLH_X2 \P1_reg[29]  ( .G(n32), .D(N90), .Q(P1[29]) );
  DLH_X2 \P1_reg[30]  ( .G(n32), .D(N89), .Q(P1[30]) );
  DLH_X2 \P1_reg[31]  ( .G(n32), .D(N88), .Q(P1[31]) );
  DLH_X2 \L_reg[0]  ( .G(n28), .D(N410), .Q(L[0]) );
  DLH_X2 \L_reg[1]  ( .G(n28), .D(N409), .Q(L[1]) );
  DLH_X2 \L_reg[2]  ( .G(n28), .D(N408), .Q(L[2]) );
  DLH_X2 \L_reg[3]  ( .G(n28), .D(N407), .Q(L[3]) );
  DLH_X2 \L_reg[4]  ( .G(n28), .D(N406), .Q(L[4]) );
  DLH_X2 \L_reg[5]  ( .G(n28), .D(N405), .Q(L[5]) );
  DLH_X2 \L_reg[6]  ( .G(n28), .D(N404), .Q(L[6]) );
  DLH_X2 \L_reg[7]  ( .G(n28), .D(N403), .Q(L[7]) );
  DLH_X2 \L_reg[8]  ( .G(n28), .D(N402), .Q(L[8]) );
  DLH_X2 \L_reg[9]  ( .G(n28), .D(N401), .Q(L[9]) );
  DLH_X2 \L_reg[10]  ( .G(n28), .D(N400), .Q(L[10]) );
  DLH_X2 \L_reg[11]  ( .G(n29), .D(N399), .Q(L[11]) );
  DLH_X2 \L_reg[12]  ( .G(n29), .D(N398), .Q(L[12]) );
  DLH_X2 \L_reg[13]  ( .G(n29), .D(N397), .Q(L[13]) );
  DLH_X2 \L_reg[14]  ( .G(n29), .D(N396), .Q(L[14]) );
  DLH_X2 \L_reg[15]  ( .G(n29), .D(N395), .Q(L[15]) );
  DLH_X2 \L_reg[16]  ( .G(n29), .D(N394), .Q(L[16]) );
  DLH_X2 \L_reg[17]  ( .G(n29), .D(N393), .Q(L[17]) );
  DLH_X2 \L_reg[18]  ( .G(n29), .D(N392), .Q(L[18]) );
  DLH_X2 \L_reg[19]  ( .G(n29), .D(N391), .Q(L[19]) );
  DLH_X2 \L_reg[20]  ( .G(n29), .D(N390), .Q(L[20]) );
  DLH_X2 \L_reg[21]  ( .G(n29), .D(N389), .Q(L[21]) );
  DLH_X2 \L_reg[22]  ( .G(n30), .D(N388), .Q(L[22]) );
  DLH_X2 \L_reg[23]  ( .G(n30), .D(N387), .Q(L[23]) );
  DLH_X2 \L_reg[24]  ( .G(n30), .D(N386), .Q(L[24]) );
  DLH_X2 \L_reg[25]  ( .G(n30), .D(N385), .Q(L[25]) );
  DLH_X2 \L_reg[26]  ( .G(n30), .D(N384), .Q(L[26]) );
  DLH_X2 \L_reg[27]  ( .G(n30), .D(N383), .Q(L[27]) );
  DLH_X2 \L_reg[28]  ( .G(n30), .D(N382), .Q(L[28]) );
  DLH_X2 \L_reg[29]  ( .G(n30), .D(N381), .Q(L[29]) );
  DLH_X2 \L_reg[30]  ( .G(n30), .D(N380), .Q(L[30]) );
  DLH_X2 \L_reg[31]  ( .G(n30), .D(N379), .Q(L[31]) );
  DLH_X2 \Z_reg[0]  ( .G(n25), .D(N443), .Q(Z[0]) );
  DLH_X2 \Z_reg[1]  ( .G(n25), .D(N442), .Q(Z[1]) );
  DLH_X2 \Z_reg[2]  ( .G(n25), .D(N441), .Q(Z[2]) );
  DLH_X2 \Z_reg[3]  ( .G(n25), .D(N440), .Q(Z[3]) );
  DLH_X2 \Z_reg[4]  ( .G(n25), .D(N439), .Q(Z[4]) );
  DLH_X2 \Z_reg[5]  ( .G(n25), .D(N438), .Q(Z[5]) );
  DLH_X2 \Z_reg[6]  ( .G(n25), .D(N437), .Q(Z[6]) );
  DLH_X2 \Z_reg[7]  ( .G(n25), .D(N436), .Q(Z[7]) );
  DLH_X2 \Z_reg[8]  ( .G(n25), .D(N435), .Q(Z[8]) );
  DLH_X2 \Z_reg[9]  ( .G(n25), .D(N434), .Q(Z[9]) );
  DLH_X2 \Z_reg[10]  ( .G(n25), .D(N433), .Q(Z[10]) );
  DLH_X2 \Z_reg[11]  ( .G(n26), .D(N432), .Q(Z[11]) );
  DLH_X2 \Z_reg[12]  ( .G(n26), .D(N431), .Q(Z[12]) );
  DLH_X2 \Z_reg[13]  ( .G(n26), .D(N430), .Q(Z[13]) );
  DLH_X2 \Z_reg[14]  ( .G(n26), .D(N429), .Q(Z[14]) );
  DLH_X2 \Z_reg[15]  ( .G(n26), .D(N428), .Q(Z[15]) );
  DLH_X2 \Z_reg[16]  ( .G(n26), .D(N427), .Q(Z[16]) );
  DLH_X2 \Z_reg[17]  ( .G(n26), .D(N426), .Q(Z[17]) );
  DLH_X2 \Z_reg[18]  ( .G(n26), .D(N425), .Q(Z[18]) );
  DLH_X2 \Z_reg[19]  ( .G(n26), .D(N424), .Q(Z[19]) );
  DLH_X2 \Z_reg[20]  ( .G(n26), .D(N423), .Q(Z[20]) );
  DLH_X2 \Z_reg[21]  ( .G(n26), .D(N422), .Q(Z[21]) );
  DLH_X2 \Z_reg[22]  ( .G(n27), .D(N421), .Q(Z[22]) );
  DLH_X2 \Z_reg[23]  ( .G(n27), .D(N420), .Q(Z[23]) );
  DLH_X2 \Z_reg[24]  ( .G(n27), .D(N419), .Q(Z[24]) );
  DLH_X2 \Z_reg[25]  ( .G(n27), .D(N418), .Q(Z[25]) );
  DLH_X2 \Z_reg[26]  ( .G(n27), .D(N417), .Q(Z[26]) );
  DLH_X2 \Z_reg[27]  ( .G(n27), .D(N416), .Q(Z[27]) );
  DLH_X2 \Z_reg[28]  ( .G(n27), .D(N415), .Q(Z[28]) );
  DLH_X2 \Z_reg[29]  ( .G(n27), .D(N414), .Q(Z[29]) );
  DLH_X2 \Z_reg[30]  ( .G(n27), .D(N413), .Q(Z[30]) );
  DLH_X2 \Z_reg[31]  ( .G(n27), .D(N412), .Q(Z[31]) );
  DLH_X2 \result_reg[0]  ( .G(n18), .D(N377), .Q(result[0]) );
  DLH_X2 \result_reg[1]  ( .G(n21), .D(N376), .Q(result[1]) );
  DLH_X2 \result_reg[2]  ( .G(n21), .D(N375), .Q(result[2]) );
  DLH_X2 \result_reg[3]  ( .G(n21), .D(N374), .Q(result[3]) );
  DLH_X2 \result_reg[4]  ( .G(n21), .D(N373), .Q(result[4]) );
  DLH_X2 \result_reg[5]  ( .G(n21), .D(N372), .Q(result[5]) );
  DLH_X2 \result_reg[6]  ( .G(n21), .D(N371), .Q(result[6]) );
  DLH_X2 \result_reg[7]  ( .G(n21), .D(N370), .Q(result[7]) );
  DLH_X2 \result_reg[8]  ( .G(n21), .D(N369), .Q(result[8]) );
  DLH_X2 \result_reg[9]  ( .G(n21), .D(N368), .Q(result[9]) );
  DLH_X2 \result_reg[10]  ( .G(n21), .D(N367), .Q(result[10]) );
  DLH_X2 \result_reg[11]  ( .G(n21), .D(N366), .Q(result[11]) );
  DLH_X2 \result_reg[12]  ( .G(n21), .D(N365), .Q(result[12]) );
  DLH_X2 \result_reg[13]  ( .G(n21), .D(N364), .Q(result[13]) );
  DLH_X2 \result_reg[14]  ( .G(n21), .D(N363), .Q(result[14]) );
  DLH_X2 \result_reg[15]  ( .G(n21), .D(N362), .Q(result[15]) );
  DLH_X2 \result_reg[16]  ( .G(n20), .D(N361), .Q(result[16]) );
  DLH_X2 \result_reg[17]  ( .G(n20), .D(N360), .Q(result[17]) );
  DLH_X2 \result_reg[18]  ( .G(n20), .D(N359), .Q(result[18]) );
  DLH_X2 \result_reg[19]  ( .G(n20), .D(N358), .Q(result[19]) );
  DLH_X2 \result_reg[20]  ( .G(n20), .D(N357), .Q(result[20]) );
  DLH_X2 \result_reg[21]  ( .G(n20), .D(N356), .Q(result[21]) );
  DLH_X2 \result_reg[22]  ( .G(n20), .D(N355), .Q(result[22]) );
  DLH_X2 \result_reg[23]  ( .G(n20), .D(N354), .Q(result[23]) );
  DLH_X2 \result_reg[24]  ( .G(n20), .D(N353), .Q(result[24]) );
  DLH_X2 \result_reg[25]  ( .G(n20), .D(N352), .Q(result[25]) );
  DLH_X2 \result_reg[26]  ( .G(n20), .D(N351), .Q(result[26]) );
  DLH_X2 \result_reg[27]  ( .G(n20), .D(N350), .Q(result[27]) );
  DLH_X2 \result_reg[28]  ( .G(n20), .D(N349), .Q(result[28]) );
  DLH_X2 \result_reg[29]  ( .G(n20), .D(N348), .Q(result[29]) );
  DLH_X2 \result_reg[30]  ( .G(n20), .D(N347), .Q(result[30]) );
  DLH_X2 \result_reg[31]  ( .G(n20), .D(N346), .Q(result[31]) );
  DLH_X2 \result_reg[32]  ( .G(n20), .D(N345), .Q(result[32]) );
  DLH_X2 \result_reg[33]  ( .G(n19), .D(N344), .Q(result[33]) );
  DLH_X2 \result_reg[34]  ( .G(n19), .D(N343), .Q(result[34]) );
  DLH_X2 \result_reg[35]  ( .G(n19), .D(N342), .Q(result[35]) );
  DLH_X2 \result_reg[36]  ( .G(n19), .D(N341), .Q(result[36]) );
  DLH_X2 \result_reg[37]  ( .G(n19), .D(N340), .Q(result[37]) );
  DLH_X2 \result_reg[38]  ( .G(n19), .D(N339), .Q(result[38]) );
  DLH_X2 \result_reg[39]  ( .G(n19), .D(N338), .Q(result[39]) );
  DLH_X2 \result_reg[40]  ( .G(n19), .D(N337), .Q(result[40]) );
  DLH_X2 \result_reg[41]  ( .G(n19), .D(N336), .Q(result[41]) );
  DLH_X2 \result_reg[42]  ( .G(n19), .D(N335), .Q(result[42]) );
  DLH_X2 \result_reg[43]  ( .G(n19), .D(N334), .Q(result[43]) );
  DLH_X2 \result_reg[44]  ( .G(n19), .D(N333), .Q(result[44]) );
  DLH_X2 \result_reg[45]  ( .G(n19), .D(N332), .Q(result[45]) );
  DLH_X2 \result_reg[46]  ( .G(n19), .D(N331), .Q(result[46]) );
  DLH_X2 \result_reg[47]  ( .G(n19), .D(N330), .Q(result[47]) );
  DLH_X2 \result_reg[48]  ( .G(n19), .D(N329), .Q(result[48]) );
  DLH_X2 \result_reg[49]  ( .G(n19), .D(N328), .Q(result[49]) );
  DLH_X2 \result_reg[50]  ( .G(n18), .D(N327), .Q(result[50]) );
  DLH_X2 \result_reg[51]  ( .G(n18), .D(N326), .Q(result[51]) );
  DLH_X2 \result_reg[52]  ( .G(n18), .D(N325), .Q(result[52]) );
  DLH_X2 \result_reg[53]  ( .G(n18), .D(N324), .Q(result[53]) );
  DLH_X2 \result_reg[54]  ( .G(n18), .D(N323), .Q(result[54]) );
  DLH_X2 \result_reg[55]  ( .G(n18), .D(N322), .Q(result[55]) );
  DLH_X2 \result_reg[56]  ( .G(n18), .D(N321), .Q(result[56]) );
  DLH_X2 \result_reg[57]  ( .G(n18), .D(N320), .Q(result[57]) );
  DLH_X2 \result_reg[58]  ( .G(n18), .D(N319), .Q(result[58]) );
  DLH_X2 \result_reg[59]  ( .G(n18), .D(N318), .Q(result[59]) );
  DLH_X2 \result_reg[60]  ( .G(n18), .D(N317), .Q(result[60]) );
  DLH_X2 \result_reg[61]  ( .G(n18), .D(N316), .Q(result[61]) );
  DLH_X2 \result_reg[62]  ( .G(n18), .D(N315), .Q(result[62]) );
  DLH_X2 \result_reg[63]  ( .G(n18), .D(N314), .Q(result[63]) );
  DLH_X2 \H_reg[0]  ( .G(n32), .D(N87), .Q(H[0]) );
  DLH_X2 \H_reg[1]  ( .G(n32), .D(N86), .Q(H[1]) );
  DLH_X2 \H_reg[2]  ( .G(n32), .D(N85), .Q(H[2]) );
  DLH_X2 \H_reg[3]  ( .G(n32), .D(N84), .Q(H[3]) );
  DLH_X2 \H_reg[4]  ( .G(n32), .D(N83), .Q(H[4]) );
  DLH_X2 \H_reg[5]  ( .G(n32), .D(N82), .Q(H[5]) );
  DLH_X2 \H_reg[6]  ( .G(n32), .D(N81), .Q(H[6]) );
  DLH_X2 \H_reg[7]  ( .G(n32), .D(N80), .Q(H[7]) );
  DLH_X2 \H_reg[8]  ( .G(n32), .D(N79), .Q(H[8]) );
  DLH_X2 \H_reg[9]  ( .G(n32), .D(N78), .Q(H[9]) );
  DLH_X2 \H_reg[10]  ( .G(n32), .D(N77), .Q(H[10]) );
  DLH_X2 \H_reg[11]  ( .G(n32), .D(N76), .Q(H[11]) );
  DLH_X2 \H_reg[12]  ( .G(n32), .D(N75), .Q(H[12]) );
  DLH_X2 \H_reg[13]  ( .G(n32), .D(N74), .Q(H[13]) );
  DLH_X2 \H_reg[14]  ( .G(n32), .D(N73), .Q(H[14]) );
  DLH_X2 \H_reg[15]  ( .G(n31), .D(N72), .Q(H[15]) );
  DLH_X2 \H_reg[16]  ( .G(n31), .D(N71), .Q(H[16]) );
  DLH_X2 \H_reg[17]  ( .G(n32), .D(N70), .Q(H[17]) );
  DLH_X2 \H_reg[18]  ( .G(n31), .D(N69), .Q(H[18]) );
  DLH_X2 \H_reg[19]  ( .G(n31), .D(N68), .Q(H[19]) );
  DLH_X2 \H_reg[20]  ( .G(n31), .D(N67), .Q(H[20]) );
  DLH_X2 \H_reg[21]  ( .G(n31), .D(N66), .Q(H[21]) );
  DLH_X2 \H_reg[22]  ( .G(n31), .D(N65), .Q(H[22]) );
  DLH_X2 \H_reg[23]  ( .G(n31), .D(N64), .Q(H[23]) );
  DLH_X2 \H_reg[24]  ( .G(n31), .D(N63), .Q(H[24]) );
  DLH_X2 \H_reg[25]  ( .G(n31), .D(N62), .Q(H[25]) );
  DLH_X2 \H_reg[26]  ( .G(n31), .D(N61), .Q(H[26]) );
  DLH_X2 \H_reg[27]  ( .G(n31), .D(N60), .Q(H[27]) );
  DLH_X2 \H_reg[28]  ( .G(n31), .D(N59), .Q(H[28]) );
  DLH_X2 \H_reg[29]  ( .G(n31), .D(N58), .Q(H[29]) );
  DLH_X2 \H_reg[30]  ( .G(n31), .D(N57), .Q(H[30]) );
  DLH_X2 \H_reg[31]  ( .G(n31), .D(N56), .Q(H[31]) );
  OR3_X4 U3 ( .A1(CurrentState[0]), .A2(CurrentState[1]), .A3(n4), .ZN(n3) );
  OR3_X4 U4 ( .A1(CurrentState[1]), .A2(CurrentState[2]), .A3(n5), .ZN(n6) );
  NOR2_X2 U5 ( .A1(N43), .A2(n17), .ZN(n7) );
  INV_X4 U6 ( .A(n7), .ZN(n29) );
  INV_X4 U41 ( .A(n7), .ZN(n28) );
  INV_X4 U74 ( .A(n7), .ZN(n30) );
  INV_X4 U107 ( .A(n35), .ZN(n11) );
  INV_X4 U108 ( .A(n6), .ZN(n19) );
  INV_X4 U109 ( .A(n6), .ZN(n20) );
  INV_X4 U110 ( .A(n3), .ZN(n16) );
  INV_X4 U111 ( .A(n6), .ZN(n21) );
  INV_X4 U112 ( .A(n9), .ZN(n26) );
  INV_X4 U113 ( .A(n9), .ZN(n25) );
  INV_X4 U114 ( .A(n10), .ZN(n23) );
  INV_X4 U115 ( .A(n10), .ZN(n22) );
  INV_X4 U116 ( .A(n9), .ZN(n27) );
  INV_X4 U117 ( .A(n10), .ZN(n24) );
  INV_X4 U118 ( .A(n33), .ZN(n13) );
  INV_X4 U119 ( .A(n33), .ZN(n12) );
  INV_X4 U120 ( .A(n33), .ZN(n14) );
  OR2_X2 U121 ( .A1(n18), .A2(n31), .ZN(n8) );
  INV_X4 U122 ( .A(n3), .ZN(n17) );
  NOR2_X2 U123 ( .A1(n33), .A2(n40), .ZN(N16) );
  NOR2_X2 U124 ( .A1(n34), .A2(n40), .ZN(N15) );
  NOR2_X2 U125 ( .A1(n15), .A2(n11), .ZN(n34) );
  INV_X4 U126 ( .A(n3), .ZN(n15) );
  AND2_X2 U127 ( .A1(n37), .A2(n33), .ZN(n9) );
  AND2_X2 U128 ( .A1(n37), .A2(n35), .ZN(n10) );
  INV_X4 U129 ( .A(n37), .ZN(n32) );
  INV_X4 U130 ( .A(n37), .ZN(n31) );
  INV_X4 U131 ( .A(N43), .ZN(n37) );
  INV_X4 U132 ( .A(n6), .ZN(n18) );
  NAND3_X2 U133 ( .A1(CurrentState[2]), .A2(n5), .A3(CurrentState[1]), .ZN(n33) );
  AOI21_X2 U134 ( .B1(n35), .B2(n36), .A(n40), .ZN(N14) );
  NAND3_X2 U135 ( .A1(n5), .A2(n4), .A3(mul), .ZN(n36) );
  NAND3_X2 U136 ( .A1(n5), .A2(n4), .A3(CurrentState[1]), .ZN(n35) );
  NOR3_X2 U137 ( .A1(CurrentState[1]), .A2(CurrentState[2]), .A3(
        CurrentState[0]), .ZN(N43) );
  INV_X4 U168 ( .A(n35), .ZN(n39) );
  INV_X4 U169 ( .A(reset), .ZN(n40) );
  multiplier_DW01_add_0 add_85 ( .A({1'b0, b[0:15]}), .B({1'b0, b[16:31]}), 
        .CI(1'b0), .SUM({N121, N120, N119, N118, N117, N116, N115, N114, N113, 
        N112, N111, N110, N109, N108, N107, N106, N105}) );
  multiplier_DW01_add_1 add_77 ( .A({1'b0, a[0:15]}), .B({1'b0, a[16:31]}), 
        .CI(1'b0), .SUM({N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, 
        N94, N93, N92, N91, N90, N89, N88}) );
  multiplier_DW01_add_3 add_1_root_add_0_root_add_98_2 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, L}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, Z, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, N298, N297, N296, 
        N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, 
        N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, 
        N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, 
        N259, N258, N257, N256, N255, N254, N253, N252, N251, N250}) );
  multiplier_DW01_add_2 add_0_root_add_0_root_add_98_2 ( .A({Z, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N298, N297, 
        N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, 
        N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, 
        N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, 
        N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250}), 
        .CI(1'b0), .SUM({N377, N376, N375, N374, N373, N372, N371, N370, N369, 
        N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, 
        N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, 
        N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, 
        N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, 
        N320, N319, N318, N317, N316, N315, N314}) );
  multiplier_DW01_sub_1 sub_1_root_sub_0_root_sub_94_2 ( .A(P), .B(L), .CI(
        1'b0), .DIFF({N217, N216, N215, N214, N213, N212, N211, N210, N209, 
        N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, 
        N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186}) );
  multiplier_DW01_sub_0 sub_0_root_sub_0_root_sub_94_2 ( .A({N217, N216, N215, 
        N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, 
        N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, 
        N190, N189, N188, N187, N186}), .B(H), .CI(1'b0), .DIFF({N249, N248, 
        N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, 
        N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, 
        N223, N222, N221, N220, N219, N218}) );
  multiplier_DW02_mult_0 mult_90 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, P1[15:31]}), .B(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, P2[15:31]}), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, N185, N184, N183, 
        N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, 
        N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, 
        N158, N157, N156, N155, N154}) );
  multiplier_DW02_mult_1 mult_76 ( .A(a[0:15]), .B(b[0:15]), .TC(1'b0), 
        .PRODUCT({N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, 
        N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, 
        N61, N60, N59, N58, N57, N56}) );
  multiplier_DW02_mult_2 mult_86 ( .A(a[16:31]), .B(b[16:31]), .TC(1'b0), 
        .PRODUCT({N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, 
        N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, 
        N131, N130, N129, N128, N127, N126, N125, N124, N123, N122}) );
endmodule


module mux_1_968 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_967 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_966 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_965 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_964 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_963 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_962 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_961 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_960 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_959 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_958 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_957 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_956 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_955 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_954 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_953 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_952 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_951 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_950 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_949 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_948 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_947 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_946 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_945 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_944 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_943 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_942 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_941 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_940 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_939 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_938 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_937 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n2;

  AND2_X4 U1 ( .A1(x), .A2(n2), .ZN(z) );
  INV_X4 U2 ( .A(sel), .ZN(n2) );
endmodule


module mux_1_936 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_935 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_934 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_933 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_932 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n5;

  AOI22_X2 U1 ( .A1(x), .A2(n2), .B1(y), .B2(n1), .ZN(n5) );
  INV_X4 U2 ( .A(n2), .ZN(n1) );
  INV_X4 U3 ( .A(sel), .ZN(n2) );
  INV_X4 U4 ( .A(n5), .ZN(z) );
endmodule


module mux_1_931 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_930 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_929 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_928 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_927 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_926 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_925 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_924 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_923 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_922 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_921 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_920 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n2, n5;

  AOI22_X2 U1 ( .A1(x), .A2(n2), .B1(y), .B2(n1), .ZN(n5) );
  INV_X4 U2 ( .A(n2), .ZN(n1) );
  INV_X4 U3 ( .A(sel), .ZN(n2) );
  INV_X4 U4 ( .A(n5), .ZN(z) );
endmodule


module mux_1_919 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_918 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_917 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_916 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_915 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_914 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_913 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_912 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_911 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_910 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_909 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_908 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_907 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_906 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_905 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux2to1_64bit ( X, Y, sel, Z );
  input [0:63] X;
  input [0:63] Y;
  output [0:63] Z;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  INV_X4 U1 ( .A(n8), .ZN(n6) );
  INV_X4 U2 ( .A(n8), .ZN(n5) );
  INV_X4 U3 ( .A(n1), .ZN(n4) );
  INV_X4 U4 ( .A(n1), .ZN(n3) );
  INV_X4 U5 ( .A(n1), .ZN(n2) );
  INV_X4 U6 ( .A(n8), .ZN(n7) );
  INV_X4 U7 ( .A(sel), .ZN(n8) );
  INV_X4 U8 ( .A(sel), .ZN(n1) );
  mux_1_968 \MUX2TO1_NBIT[0].MUX  ( .x(X[0]), .y(1'b0), .sel(n2), .z(Z[0]) );
  mux_1_967 \MUX2TO1_NBIT[1].MUX  ( .x(X[1]), .y(1'b0), .sel(n2), .z(Z[1]) );
  mux_1_966 \MUX2TO1_NBIT[2].MUX  ( .x(X[2]), .y(1'b0), .sel(n2), .z(Z[2]) );
  mux_1_965 \MUX2TO1_NBIT[3].MUX  ( .x(X[3]), .y(1'b0), .sel(n2), .z(Z[3]) );
  mux_1_964 \MUX2TO1_NBIT[4].MUX  ( .x(X[4]), .y(1'b0), .sel(n2), .z(Z[4]) );
  mux_1_963 \MUX2TO1_NBIT[5].MUX  ( .x(X[5]), .y(1'b0), .sel(n2), .z(Z[5]) );
  mux_1_962 \MUX2TO1_NBIT[6].MUX  ( .x(X[6]), .y(1'b0), .sel(n2), .z(Z[6]) );
  mux_1_961 \MUX2TO1_NBIT[7].MUX  ( .x(X[7]), .y(1'b0), .sel(n2), .z(Z[7]) );
  mux_1_960 \MUX2TO1_NBIT[8].MUX  ( .x(X[8]), .y(1'b0), .sel(n2), .z(Z[8]) );
  mux_1_959 \MUX2TO1_NBIT[9].MUX  ( .x(X[9]), .y(1'b0), .sel(n2), .z(Z[9]) );
  mux_1_958 \MUX2TO1_NBIT[10].MUX  ( .x(X[10]), .y(1'b0), .sel(n2), .z(Z[10])
         );
  mux_1_957 \MUX2TO1_NBIT[11].MUX  ( .x(X[11]), .y(1'b0), .sel(n2), .z(Z[11])
         );
  mux_1_956 \MUX2TO1_NBIT[12].MUX  ( .x(X[12]), .y(1'b0), .sel(n3), .z(Z[12])
         );
  mux_1_955 \MUX2TO1_NBIT[13].MUX  ( .x(X[13]), .y(1'b0), .sel(n3), .z(Z[13])
         );
  mux_1_954 \MUX2TO1_NBIT[14].MUX  ( .x(X[14]), .y(1'b0), .sel(n3), .z(Z[14])
         );
  mux_1_953 \MUX2TO1_NBIT[15].MUX  ( .x(X[15]), .y(1'b0), .sel(n3), .z(Z[15])
         );
  mux_1_952 \MUX2TO1_NBIT[16].MUX  ( .x(X[16]), .y(1'b0), .sel(n3), .z(Z[16])
         );
  mux_1_951 \MUX2TO1_NBIT[17].MUX  ( .x(X[17]), .y(1'b0), .sel(n3), .z(Z[17])
         );
  mux_1_950 \MUX2TO1_NBIT[18].MUX  ( .x(X[18]), .y(1'b0), .sel(n3), .z(Z[18])
         );
  mux_1_949 \MUX2TO1_NBIT[19].MUX  ( .x(X[19]), .y(1'b0), .sel(n3), .z(Z[19])
         );
  mux_1_948 \MUX2TO1_NBIT[20].MUX  ( .x(X[20]), .y(1'b0), .sel(n3), .z(Z[20])
         );
  mux_1_947 \MUX2TO1_NBIT[21].MUX  ( .x(X[21]), .y(1'b0), .sel(n3), .z(Z[21])
         );
  mux_1_946 \MUX2TO1_NBIT[22].MUX  ( .x(X[22]), .y(1'b0), .sel(n3), .z(Z[22])
         );
  mux_1_945 \MUX2TO1_NBIT[23].MUX  ( .x(X[23]), .y(1'b0), .sel(n3), .z(Z[23])
         );
  mux_1_944 \MUX2TO1_NBIT[24].MUX  ( .x(X[24]), .y(1'b0), .sel(n4), .z(Z[24])
         );
  mux_1_943 \MUX2TO1_NBIT[25].MUX  ( .x(X[25]), .y(1'b0), .sel(n4), .z(Z[25])
         );
  mux_1_942 \MUX2TO1_NBIT[26].MUX  ( .x(X[26]), .y(1'b0), .sel(n4), .z(Z[26])
         );
  mux_1_941 \MUX2TO1_NBIT[27].MUX  ( .x(X[27]), .y(1'b0), .sel(n4), .z(Z[27])
         );
  mux_1_940 \MUX2TO1_NBIT[28].MUX  ( .x(X[28]), .y(1'b0), .sel(n4), .z(Z[28])
         );
  mux_1_939 \MUX2TO1_NBIT[29].MUX  ( .x(X[29]), .y(1'b0), .sel(n4), .z(Z[29])
         );
  mux_1_938 \MUX2TO1_NBIT[30].MUX  ( .x(X[30]), .y(1'b0), .sel(n4), .z(Z[30])
         );
  mux_1_937 \MUX2TO1_NBIT[31].MUX  ( .x(X[31]), .y(1'b0), .sel(n4), .z(Z[31])
         );
  mux_1_936 \MUX2TO1_NBIT[32].MUX  ( .x(X[32]), .y(Y[32]), .sel(n4), .z(Z[32])
         );
  mux_1_935 \MUX2TO1_NBIT[33].MUX  ( .x(X[33]), .y(Y[33]), .sel(n4), .z(Z[33])
         );
  mux_1_934 \MUX2TO1_NBIT[34].MUX  ( .x(X[34]), .y(Y[34]), .sel(n4), .z(Z[34])
         );
  mux_1_933 \MUX2TO1_NBIT[35].MUX  ( .x(X[35]), .y(Y[35]), .sel(n4), .z(Z[35])
         );
  mux_1_932 \MUX2TO1_NBIT[36].MUX  ( .x(X[36]), .y(Y[36]), .sel(n5), .z(Z[36])
         );
  mux_1_931 \MUX2TO1_NBIT[37].MUX  ( .x(X[37]), .y(Y[37]), .sel(n5), .z(Z[37])
         );
  mux_1_930 \MUX2TO1_NBIT[38].MUX  ( .x(X[38]), .y(Y[38]), .sel(n5), .z(Z[38])
         );
  mux_1_929 \MUX2TO1_NBIT[39].MUX  ( .x(X[39]), .y(Y[39]), .sel(n5), .z(Z[39])
         );
  mux_1_928 \MUX2TO1_NBIT[40].MUX  ( .x(X[40]), .y(Y[40]), .sel(n5), .z(Z[40])
         );
  mux_1_927 \MUX2TO1_NBIT[41].MUX  ( .x(X[41]), .y(Y[41]), .sel(n5), .z(Z[41])
         );
  mux_1_926 \MUX2TO1_NBIT[42].MUX  ( .x(X[42]), .y(Y[42]), .sel(n5), .z(Z[42])
         );
  mux_1_925 \MUX2TO1_NBIT[43].MUX  ( .x(X[43]), .y(Y[43]), .sel(n5), .z(Z[43])
         );
  mux_1_924 \MUX2TO1_NBIT[44].MUX  ( .x(X[44]), .y(Y[44]), .sel(n5), .z(Z[44])
         );
  mux_1_923 \MUX2TO1_NBIT[45].MUX  ( .x(X[45]), .y(Y[45]), .sel(n5), .z(Z[45])
         );
  mux_1_922 \MUX2TO1_NBIT[46].MUX  ( .x(X[46]), .y(Y[46]), .sel(n5), .z(Z[46])
         );
  mux_1_921 \MUX2TO1_NBIT[47].MUX  ( .x(X[47]), .y(Y[47]), .sel(n5), .z(Z[47])
         );
  mux_1_920 \MUX2TO1_NBIT[48].MUX  ( .x(X[48]), .y(Y[48]), .sel(n6), .z(Z[48])
         );
  mux_1_919 \MUX2TO1_NBIT[49].MUX  ( .x(X[49]), .y(Y[49]), .sel(n6), .z(Z[49])
         );
  mux_1_918 \MUX2TO1_NBIT[50].MUX  ( .x(X[50]), .y(Y[50]), .sel(n6), .z(Z[50])
         );
  mux_1_917 \MUX2TO1_NBIT[51].MUX  ( .x(X[51]), .y(Y[51]), .sel(n6), .z(Z[51])
         );
  mux_1_916 \MUX2TO1_NBIT[52].MUX  ( .x(X[52]), .y(Y[52]), .sel(n6), .z(Z[52])
         );
  mux_1_915 \MUX2TO1_NBIT[53].MUX  ( .x(X[53]), .y(Y[53]), .sel(n6), .z(Z[53])
         );
  mux_1_914 \MUX2TO1_NBIT[54].MUX  ( .x(X[54]), .y(Y[54]), .sel(n6), .z(Z[54])
         );
  mux_1_913 \MUX2TO1_NBIT[55].MUX  ( .x(X[55]), .y(Y[55]), .sel(n6), .z(Z[55])
         );
  mux_1_912 \MUX2TO1_NBIT[56].MUX  ( .x(X[56]), .y(Y[56]), .sel(n6), .z(Z[56])
         );
  mux_1_911 \MUX2TO1_NBIT[57].MUX  ( .x(X[57]), .y(Y[57]), .sel(n6), .z(Z[57])
         );
  mux_1_910 \MUX2TO1_NBIT[58].MUX  ( .x(X[58]), .y(Y[58]), .sel(n6), .z(Z[58])
         );
  mux_1_909 \MUX2TO1_NBIT[59].MUX  ( .x(X[59]), .y(Y[59]), .sel(n6), .z(Z[59])
         );
  mux_1_908 \MUX2TO1_NBIT[60].MUX  ( .x(X[60]), .y(Y[60]), .sel(n7), .z(Z[60])
         );
  mux_1_907 \MUX2TO1_NBIT[61].MUX  ( .x(X[61]), .y(Y[61]), .sel(n7), .z(Z[61])
         );
  mux_1_906 \MUX2TO1_NBIT[62].MUX  ( .x(X[62]), .y(Y[62]), .sel(n7), .z(Z[62])
         );
  mux_1_905 \MUX2TO1_NBIT[63].MUX  ( .x(X[63]), .y(Y[63]), .sel(n7), .z(Z[63])
         );
endmodule


module zero_0 ( X, z );
  input [0:31] X;
  output z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  NAND4_X2 U2 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n2) );
  NOR4_X2 U3 ( .A1(X[23]), .A2(X[22]), .A3(X[21]), .A4(X[20]), .ZN(n6) );
  NOR4_X2 U4 ( .A1(X[1]), .A2(X[19]), .A3(X[18]), .A4(X[17]), .ZN(n5) );
  NOR4_X2 U5 ( .A1(X[16]), .A2(X[15]), .A3(X[14]), .A4(X[13]), .ZN(n4) );
  NOR4_X2 U6 ( .A1(X[12]), .A2(X[11]), .A3(X[10]), .A4(X[0]), .ZN(n3) );
  NAND4_X2 U7 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n1) );
  NOR4_X2 U8 ( .A1(X[9]), .A2(X[8]), .A3(X[7]), .A4(X[6]), .ZN(n10) );
  NOR4_X2 U9 ( .A1(X[5]), .A2(X[4]), .A3(X[3]), .A4(X[31]), .ZN(n9) );
  NOR4_X2 U10 ( .A1(X[30]), .A2(X[2]), .A3(X[29]), .A4(X[28]), .ZN(n8) );
  NOR4_X2 U11 ( .A1(X[27]), .A2(X[26]), .A3(X[25]), .A4(X[24]), .ZN(n7) );
  NOR2_X2 U1 ( .A1(n1), .A2(n2), .ZN(z) );
endmodule


module check_branch ( busA, aluZero, branchZero, branch, jump, leap );
  input [0:31] busA;
  input aluZero, branchZero, branch, jump;
  output leap;
  wire   zeroBit, n2, n3;

  XNOR2_X2 U2 ( .A(zeroBit), .B(branchZero), .ZN(n3) );
  AOI21_X2 U1 ( .B1(n3), .B2(branch), .A(jump), .ZN(n2) );
  INV_X4 U3 ( .A(n2), .ZN(leap) );
  zero_0 ZERO_A ( .X(busA), .z(zeroBit) );
endmodule


module mux_1_904 ( x, y, sel, z );
  input x, y, sel;
  output z;


  BUF_X32 U1 ( .A(y), .Z(z) );
endmodule


module extend_16to32 ( x, sign, Z );
  input [0:15] x;
  output [0:31] Z;
  input sign;
  wire   Z_0, n18;
  assign Z[0] = Z_0;

  mux_1_904 SELECT_EXTEND ( .x(1'b0), .y(x[0]), .sel(1'b1), .z(Z_0) );
  BUF_X32 U3 ( .A(x[15]), .Z(Z[31]) );
  BUF_X32 U4 ( .A(x[14]), .Z(Z[30]) );
  BUF_X32 U5 ( .A(x[13]), .Z(Z[29]) );
  BUF_X32 U6 ( .A(x[12]), .Z(Z[28]) );
  BUF_X32 U7 ( .A(x[11]), .Z(Z[27]) );
  BUF_X32 U8 ( .A(x[10]), .Z(Z[26]) );
  BUF_X32 U9 ( .A(x[9]), .Z(Z[25]) );
  BUF_X32 U10 ( .A(x[8]), .Z(Z[24]) );
  BUF_X32 U11 ( .A(x[7]), .Z(Z[23]) );
  BUF_X32 U12 ( .A(x[6]), .Z(Z[22]) );
  BUF_X32 U13 ( .A(x[5]), .Z(Z[21]) );
  BUF_X32 U14 ( .A(x[4]), .Z(Z[20]) );
  BUF_X32 U15 ( .A(x[3]), .Z(Z[19]) );
  BUF_X32 U16 ( .A(x[2]), .Z(Z[18]) );
  BUF_X32 U17 ( .A(x[1]), .Z(Z[17]) );
  BUF_X32 U18 ( .A(x[0]), .Z(Z[16]) );
  INV_X32 U19 ( .A(Z_0), .ZN(n18) );
  INV_X32 U20 ( .A(n18), .ZN(Z[1]) );
  INV_X32 U21 ( .A(n18), .ZN(Z[2]) );
  INV_X32 U22 ( .A(n18), .ZN(Z[3]) );
  INV_X32 U23 ( .A(n18), .ZN(Z[4]) );
  INV_X32 U24 ( .A(n18), .ZN(Z[5]) );
  INV_X32 U25 ( .A(n18), .ZN(Z[6]) );
  INV_X32 U26 ( .A(n18), .ZN(Z[7]) );
  INV_X32 U27 ( .A(n18), .ZN(Z[8]) );
  INV_X32 U28 ( .A(n18), .ZN(Z[9]) );
  INV_X32 U29 ( .A(n18), .ZN(Z[10]) );
  INV_X32 U30 ( .A(n18), .ZN(Z[11]) );
  INV_X32 U31 ( .A(n18), .ZN(Z[12]) );
  INV_X32 U32 ( .A(n18), .ZN(Z[13]) );
  INV_X32 U33 ( .A(n18), .ZN(Z[14]) );
  INV_X32 U34 ( .A(n18), .ZN(Z[15]) );
endmodule


module mux_1_903 ( x, y, sel, z );
  input x, y, sel;
  output z;


  BUF_X4 U1 ( .A(y), .Z(z) );
endmodule


module extend_26to32 ( x, sign, Z );
  input [0:25] x;
  output [0:31] Z;
  input sign;
  wire   Z_0;
  assign Z[0] = Z_0;

  mux_1_903 SELECT_EXTEND ( .x(1'b0), .y(x[0]), .sel(1'b1), .z(Z_0) );
  BUF_X32 U3 ( .A(x[25]), .Z(Z[31]) );
  BUF_X32 U4 ( .A(x[24]), .Z(Z[30]) );
  BUF_X32 U5 ( .A(x[23]), .Z(Z[29]) );
  BUF_X32 U6 ( .A(x[22]), .Z(Z[28]) );
  BUF_X32 U7 ( .A(x[21]), .Z(Z[27]) );
  BUF_X32 U8 ( .A(x[20]), .Z(Z[26]) );
  BUF_X32 U9 ( .A(x[19]), .Z(Z[25]) );
  BUF_X32 U10 ( .A(x[18]), .Z(Z[24]) );
  BUF_X32 U11 ( .A(x[17]), .Z(Z[23]) );
  BUF_X32 U12 ( .A(x[16]), .Z(Z[22]) );
  BUF_X32 U13 ( .A(x[15]), .Z(Z[21]) );
  BUF_X32 U14 ( .A(x[14]), .Z(Z[20]) );
  BUF_X32 U15 ( .A(x[13]), .Z(Z[19]) );
  BUF_X32 U16 ( .A(x[12]), .Z(Z[18]) );
  BUF_X32 U17 ( .A(x[11]), .Z(Z[17]) );
  BUF_X32 U18 ( .A(x[10]), .Z(Z[16]) );
  BUF_X32 U19 ( .A(x[9]), .Z(Z[15]) );
  BUF_X32 U20 ( .A(x[8]), .Z(Z[14]) );
  BUF_X32 U21 ( .A(x[7]), .Z(Z[13]) );
  BUF_X32 U22 ( .A(x[6]), .Z(Z[12]) );
  BUF_X32 U23 ( .A(x[5]), .Z(Z[11]) );
  BUF_X32 U24 ( .A(x[4]), .Z(Z[10]) );
  BUF_X32 U25 ( .A(x[3]), .Z(Z[9]) );
  BUF_X32 U26 ( .A(x[2]), .Z(Z[8]) );
  BUF_X32 U27 ( .A(x[1]), .Z(Z[7]) );
  BUF_X32 U28 ( .A(x[0]), .Z(Z[6]) );
  BUF_X32 U29 ( .A(Z_0), .Z(Z[1]) );
  BUF_X32 U30 ( .A(Z_0), .Z(Z[2]) );
  BUF_X32 U31 ( .A(Z_0), .Z(Z[3]) );
  BUF_X32 U32 ( .A(Z_0), .Z(Z[4]) );
  BUF_X32 U33 ( .A(Z_0), .Z(Z[5]) );
endmodule


module mux_1_902 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_901 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_900 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_899 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_898 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_897 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_896 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_895 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_894 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_893 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_892 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_891 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_890 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_889 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_888 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_887 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_886 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_885 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_884 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_883 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_882 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_881 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_880 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_879 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_878 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_877 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_876 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_875 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_874 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_873 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_872 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux_1_871 ( x, y, sel, z );
  input x, y, sel;
  output z;
  wire   n1, n4;

  AOI22_X2 U1 ( .A1(x), .A2(n1), .B1(y), .B2(sel), .ZN(n4) );
  INV_X4 U2 ( .A(sel), .ZN(n1) );
  INV_X4 U3 ( .A(n4), .ZN(z) );
endmodule


module mux2to1_32bit_28 ( X, Y, sel, Z );
  input [0:31] X;
  input [0:31] Y;
  output [0:31] Z;
  input sel;
  wire   n1, n2, n3;

  INV_X4 U1 ( .A(n3), .ZN(n2) );
  INV_X4 U2 ( .A(n3), .ZN(n1) );
  INV_X4 U3 ( .A(sel), .ZN(n3) );
  mux_1_902 \MUX2TO1_32BIT[0].MUX  ( .x(X[0]), .y(Y[0]), .sel(n1), .z(Z[0]) );
  mux_1_901 \MUX2TO1_32BIT[1].MUX  ( .x(X[1]), .y(Y[1]), .sel(n1), .z(Z[1]) );
  mux_1_900 \MUX2TO1_32BIT[2].MUX  ( .x(X[2]), .y(Y[2]), .sel(n1), .z(Z[2]) );
  mux_1_899 \MUX2TO1_32BIT[3].MUX  ( .x(X[3]), .y(Y[3]), .sel(n1), .z(Z[3]) );
  mux_1_898 \MUX2TO1_32BIT[4].MUX  ( .x(X[4]), .y(Y[4]), .sel(n1), .z(Z[4]) );
  mux_1_897 \MUX2TO1_32BIT[5].MUX  ( .x(X[5]), .y(Y[5]), .sel(n1), .z(Z[5]) );
  mux_1_896 \MUX2TO1_32BIT[6].MUX  ( .x(X[6]), .y(Y[6]), .sel(n1), .z(Z[6]) );
  mux_1_895 \MUX2TO1_32BIT[7].MUX  ( .x(X[7]), .y(Y[7]), .sel(n1), .z(Z[7]) );
  mux_1_894 \MUX2TO1_32BIT[8].MUX  ( .x(X[8]), .y(Y[8]), .sel(n1), .z(Z[8]) );
  mux_1_893 \MUX2TO1_32BIT[9].MUX  ( .x(X[9]), .y(Y[9]), .sel(n1), .z(Z[9]) );
  mux_1_892 \MUX2TO1_32BIT[10].MUX  ( .x(X[10]), .y(Y[10]), .sel(n1), .z(Z[10]) );
  mux_1_891 \MUX2TO1_32BIT[11].MUX  ( .x(X[11]), .y(Y[11]), .sel(n1), .z(Z[11]) );
  mux_1_890 \MUX2TO1_32BIT[12].MUX  ( .x(X[12]), .y(Y[12]), .sel(n2), .z(Z[12]) );
  mux_1_889 \MUX2TO1_32BIT[13].MUX  ( .x(X[13]), .y(Y[13]), .sel(n2), .z(Z[13]) );
  mux_1_888 \MUX2TO1_32BIT[14].MUX  ( .x(X[14]), .y(Y[14]), .sel(n2), .z(Z[14]) );
  mux_1_887 \MUX2TO1_32BIT[15].MUX  ( .x(X[15]), .y(Y[15]), .sel(n2), .z(Z[15]) );
  mux_1_886 \MUX2TO1_32BIT[16].MUX  ( .x(X[16]), .y(Y[16]), .sel(n2), .z(Z[16]) );
  mux_1_885 \MUX2TO1_32BIT[17].MUX  ( .x(X[17]), .y(Y[17]), .sel(n2), .z(Z[17]) );
  mux_1_884 \MUX2TO1_32BIT[18].MUX  ( .x(X[18]), .y(Y[18]), .sel(n2), .z(Z[18]) );
  mux_1_883 \MUX2TO1_32BIT[19].MUX  ( .x(X[19]), .y(Y[19]), .sel(n2), .z(Z[19]) );
  mux_1_882 \MUX2TO1_32BIT[20].MUX  ( .x(X[20]), .y(Y[20]), .sel(n2), .z(Z[20]) );
  mux_1_881 \MUX2TO1_32BIT[21].MUX  ( .x(X[21]), .y(Y[21]), .sel(n2), .z(Z[21]) );
  mux_1_880 \MUX2TO1_32BIT[22].MUX  ( .x(X[22]), .y(Y[22]), .sel(n2), .z(Z[22]) );
  mux_1_879 \MUX2TO1_32BIT[23].MUX  ( .x(X[23]), .y(Y[23]), .sel(n2), .z(Z[23]) );
  mux_1_878 \MUX2TO1_32BIT[24].MUX  ( .x(X[24]), .y(Y[24]), .sel(sel), .z(
        Z[24]) );
  mux_1_877 \MUX2TO1_32BIT[25].MUX  ( .x(X[25]), .y(Y[25]), .sel(sel), .z(
        Z[25]) );
  mux_1_876 \MUX2TO1_32BIT[26].MUX  ( .x(X[26]), .y(Y[26]), .sel(sel), .z(
        Z[26]) );
  mux_1_875 \MUX2TO1_32BIT[27].MUX  ( .x(X[27]), .y(Y[27]), .sel(sel), .z(
        Z[27]) );
  mux_1_874 \MUX2TO1_32BIT[28].MUX  ( .x(X[28]), .y(Y[28]), .sel(sel), .z(
        Z[28]) );
  mux_1_873 \MUX2TO1_32BIT[29].MUX  ( .x(X[29]), .y(Y[29]), .sel(sel), .z(
        Z[29]) );
  mux_1_872 \MUX2TO1_32BIT[30].MUX  ( .x(X[30]), .y(Y[30]), .sel(sel), .z(
        Z[30]) );
  mux_1_871 \MUX2TO1_32BIT[31].MUX  ( .x(X[31]), .y(Y[31]), .sel(sel), .z(
        Z[31]) );
endmodule


module execute ( nextPC_in, opA_in, opB_in, offset26_in, offset16_in, 
        destReg_in, PCtoReg_in, RegToPC_in, jump_in, branch_in, branchZero_in, 
        RType_in, RegWrite_in, MemToReg_in, MemWrite_in, loadSign_in, mul_in, 
        DSize_in, ALUCtrl_in, memVal_in, f1_in, f2_in, fDestReg_in, FPRType_in, 
        FPRegWrite_in, movfp2i_in, movi2fp_in, clk, reset, nextPC_out, 
        aluResult_out, leapAddr_out, destReg_out, leap_out, PCtoReg_out, 
        RegToPC_out, RegWrite_out, MemToReg_out, MemWrite_out, loadSign_out, 
        DSize_out, memVal_out, stall_out, fDestReg_out, fbusW, FPRegWrite_out, 
        mul_out );
  input [0:31] nextPC_in;
  input [0:31] opA_in;
  input [0:31] opB_in;
  input [0:25] offset26_in;
  input [0:15] offset16_in;
  input [0:4] destReg_in;
  input [0:1] DSize_in;
  input [0:3] ALUCtrl_in;
  input [0:31] memVal_in;
  input [0:31] f1_in;
  input [0:31] f2_in;
  input [0:4] fDestReg_in;
  output [0:31] nextPC_out;
  output [0:31] aluResult_out;
  output [0:31] leapAddr_out;
  output [0:4] destReg_out;
  output [0:1] DSize_out;
  output [0:31] memVal_out;
  output [0:4] fDestReg_out;
  output [0:63] fbusW;
  input PCtoReg_in, RegToPC_in, jump_in, branch_in, branchZero_in, RType_in,
         RegWrite_in, MemToReg_in, MemWrite_in, loadSign_in, mul_in,
         FPRType_in, FPRegWrite_in, movfp2i_in, movi2fp_in, clk, reset;
  output leap_out, PCtoReg_out, RegToPC_out, RegWrite_out, MemToReg_out,
         MemWrite_out, loadSign_out, stall_out, FPRegWrite_out, mul_out;
  wire   mul_done, n2;
  wire   [0:31] not_mul_result;
  wire   [0:63] mul_result_long;
  wire   [0:31] imm16_32;
  wire   [0:31] imm26_32;

  NOR2_X2 U5 ( .A1(mul_done), .A2(n2), .ZN(stall_out) );
  INV_X4 U6 ( .A(mul_in), .ZN(n2) );
  alu alu_ex ( .A(opA_in), .B(opB_in), .ctrl(ALUCtrl_in), .ALUout(
        not_mul_result) );
  mux2to1_32bit_0 CHOOSE_FP_OR_NOTMUL ( .X(not_mul_result), .Y(f1_in), .sel(
        movfp2i_in), .Z(aluResult_out) );
  multiplier mul_ex ( .clk(clk), .reset(reset), .mul(mul_in), .a(f1_in), .b(
        f2_in), .done(mul_done), .result(mul_result_long) );
  mux2to1_64bit CHOOSE_MULT_OR_INT ( .X(mul_result_long), .Y({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, opA_in}), .sel(movi2fp_in), .Z(fbusW) );
  check_branch decide_if_leap ( .busA(opA_in), .aluZero(1'b0), .branchZero(
        branchZero_in), .branch(branch_in), .jump(jump_in), .leap(leap_out) );
  extend_16to32 EXTEND_IMM16 ( .x(offset16_in), .sign(1'b1), .Z(imm16_32) );
  extend_26to32 EXTEND_IMM26 ( .x(offset26_in), .sign(1'b1), .Z(imm26_32) );
  mux2to1_32bit_28 CHOOSE_IMMEDIATE ( .X(imm26_32), .Y(imm16_32), .sel(
        branch_in), .Z(leapAddr_out) );
  BUF_X32 U8 ( .A(mul_in), .Z(mul_out) );
  BUF_X32 U9 ( .A(FPRegWrite_in), .Z(FPRegWrite_out) );
  BUF_X32 U10 ( .A(fDestReg_in[4]), .Z(fDestReg_out[4]) );
  BUF_X32 U11 ( .A(fDestReg_in[3]), .Z(fDestReg_out[3]) );
  BUF_X32 U12 ( .A(fDestReg_in[2]), .Z(fDestReg_out[2]) );
  BUF_X32 U13 ( .A(fDestReg_in[1]), .Z(fDestReg_out[1]) );
  BUF_X32 U14 ( .A(fDestReg_in[0]), .Z(fDestReg_out[0]) );
  BUF_X32 U15 ( .A(memVal_in[31]), .Z(memVal_out[31]) );
  BUF_X32 U16 ( .A(memVal_in[30]), .Z(memVal_out[30]) );
  BUF_X32 U17 ( .A(memVal_in[29]), .Z(memVal_out[29]) );
  BUF_X32 U18 ( .A(memVal_in[28]), .Z(memVal_out[28]) );
  BUF_X32 U19 ( .A(memVal_in[27]), .Z(memVal_out[27]) );
  BUF_X32 U20 ( .A(memVal_in[26]), .Z(memVal_out[26]) );
  BUF_X32 U21 ( .A(memVal_in[25]), .Z(memVal_out[25]) );
  BUF_X32 U22 ( .A(memVal_in[24]), .Z(memVal_out[24]) );
  BUF_X32 U23 ( .A(memVal_in[23]), .Z(memVal_out[23]) );
  BUF_X32 U24 ( .A(memVal_in[22]), .Z(memVal_out[22]) );
  BUF_X32 U25 ( .A(memVal_in[21]), .Z(memVal_out[21]) );
  BUF_X32 U26 ( .A(memVal_in[20]), .Z(memVal_out[20]) );
  BUF_X32 U27 ( .A(memVal_in[19]), .Z(memVal_out[19]) );
  BUF_X32 U28 ( .A(memVal_in[18]), .Z(memVal_out[18]) );
  BUF_X32 U29 ( .A(memVal_in[17]), .Z(memVal_out[17]) );
  BUF_X32 U30 ( .A(memVal_in[16]), .Z(memVal_out[16]) );
  BUF_X32 U31 ( .A(memVal_in[15]), .Z(memVal_out[15]) );
  BUF_X32 U32 ( .A(memVal_in[14]), .Z(memVal_out[14]) );
  BUF_X32 U33 ( .A(memVal_in[13]), .Z(memVal_out[13]) );
  BUF_X32 U34 ( .A(memVal_in[12]), .Z(memVal_out[12]) );
  BUF_X32 U35 ( .A(memVal_in[11]), .Z(memVal_out[11]) );
  BUF_X32 U36 ( .A(memVal_in[10]), .Z(memVal_out[10]) );
  BUF_X32 U37 ( .A(memVal_in[9]), .Z(memVal_out[9]) );
  BUF_X32 U38 ( .A(memVal_in[8]), .Z(memVal_out[8]) );
  BUF_X32 U39 ( .A(memVal_in[7]), .Z(memVal_out[7]) );
  BUF_X32 U40 ( .A(memVal_in[6]), .Z(memVal_out[6]) );
  BUF_X32 U41 ( .A(memVal_in[5]), .Z(memVal_out[5]) );
  BUF_X32 U42 ( .A(memVal_in[4]), .Z(memVal_out[4]) );
  BUF_X32 U43 ( .A(memVal_in[3]), .Z(memVal_out[3]) );
  BUF_X32 U44 ( .A(memVal_in[2]), .Z(memVal_out[2]) );
  BUF_X32 U45 ( .A(memVal_in[1]), .Z(memVal_out[1]) );
  BUF_X32 U46 ( .A(memVal_in[0]), .Z(memVal_out[0]) );
  BUF_X32 U47 ( .A(DSize_in[1]), .Z(DSize_out[1]) );
  BUF_X32 U48 ( .A(DSize_in[0]), .Z(DSize_out[0]) );
  BUF_X32 U49 ( .A(loadSign_in), .Z(loadSign_out) );
  BUF_X32 U50 ( .A(MemWrite_in), .Z(MemWrite_out) );
  BUF_X32 U51 ( .A(MemToReg_in), .Z(MemToReg_out) );
  BUF_X32 U52 ( .A(RegWrite_in), .Z(RegWrite_out) );
  BUF_X32 U53 ( .A(RegToPC_in), .Z(RegToPC_out) );
  BUF_X32 U54 ( .A(PCtoReg_in), .Z(PCtoReg_out) );
  BUF_X32 U55 ( .A(destReg_in[4]), .Z(destReg_out[4]) );
  BUF_X32 U56 ( .A(destReg_in[3]), .Z(destReg_out[3]) );
  BUF_X32 U57 ( .A(destReg_in[2]), .Z(destReg_out[2]) );
  BUF_X32 U58 ( .A(destReg_in[1]), .Z(destReg_out[1]) );
  BUF_X32 U59 ( .A(destReg_in[0]), .Z(destReg_out[0]) );
  BUF_X32 U60 ( .A(nextPC_in[31]), .Z(nextPC_out[31]) );
  BUF_X32 U61 ( .A(nextPC_in[30]), .Z(nextPC_out[30]) );
  BUF_X32 U62 ( .A(nextPC_in[29]), .Z(nextPC_out[29]) );
  BUF_X32 U63 ( .A(nextPC_in[28]), .Z(nextPC_out[28]) );
  BUF_X32 U64 ( .A(nextPC_in[27]), .Z(nextPC_out[27]) );
  BUF_X32 U65 ( .A(nextPC_in[26]), .Z(nextPC_out[26]) );
  BUF_X32 U66 ( .A(nextPC_in[25]), .Z(nextPC_out[25]) );
  BUF_X32 U67 ( .A(nextPC_in[24]), .Z(nextPC_out[24]) );
  BUF_X32 U68 ( .A(nextPC_in[23]), .Z(nextPC_out[23]) );
  BUF_X32 U69 ( .A(nextPC_in[22]), .Z(nextPC_out[22]) );
  BUF_X32 U70 ( .A(nextPC_in[21]), .Z(nextPC_out[21]) );
  BUF_X32 U71 ( .A(nextPC_in[20]), .Z(nextPC_out[20]) );
  BUF_X32 U72 ( .A(nextPC_in[19]), .Z(nextPC_out[19]) );
  BUF_X32 U73 ( .A(nextPC_in[18]), .Z(nextPC_out[18]) );
  BUF_X32 U74 ( .A(nextPC_in[17]), .Z(nextPC_out[17]) );
  BUF_X32 U75 ( .A(nextPC_in[16]), .Z(nextPC_out[16]) );
  BUF_X32 U76 ( .A(nextPC_in[15]), .Z(nextPC_out[15]) );
  BUF_X32 U77 ( .A(nextPC_in[14]), .Z(nextPC_out[14]) );
  BUF_X32 U78 ( .A(nextPC_in[13]), .Z(nextPC_out[13]) );
  BUF_X32 U79 ( .A(nextPC_in[12]), .Z(nextPC_out[12]) );
  BUF_X32 U80 ( .A(nextPC_in[11]), .Z(nextPC_out[11]) );
  BUF_X32 U81 ( .A(nextPC_in[10]), .Z(nextPC_out[10]) );
  BUF_X32 U82 ( .A(nextPC_in[9]), .Z(nextPC_out[9]) );
  BUF_X32 U83 ( .A(nextPC_in[8]), .Z(nextPC_out[8]) );
  BUF_X32 U84 ( .A(nextPC_in[7]), .Z(nextPC_out[7]) );
  BUF_X32 U85 ( .A(nextPC_in[6]), .Z(nextPC_out[6]) );
  BUF_X32 U86 ( .A(nextPC_in[5]), .Z(nextPC_out[5]) );
  BUF_X32 U87 ( .A(nextPC_in[4]), .Z(nextPC_out[4]) );
  BUF_X32 U88 ( .A(nextPC_in[3]), .Z(nextPC_out[3]) );
  BUF_X32 U89 ( .A(nextPC_in[2]), .Z(nextPC_out[2]) );
  BUF_X32 U90 ( .A(nextPC_in[1]), .Z(nextPC_out[1]) );
  BUF_X32 U91 ( .A(nextPC_in[0]), .Z(nextPC_out[0]) );
endmodule

