
module pipeline_processor ( clk, reset, DMEM_BUS_OUT, DMEM_BUS_IN, 
        IMEM_BUS_OUT, IMEM_BUS_IN );
  output [0:66] DMEM_BUS_OUT;
  input [0:31] DMEM_BUS_IN;
  output [0:31] IMEM_BUS_OUT;
  input [0:31] IMEM_BUS_IN;
  input clk, reset;
  wire   DSize_ex_out_0_, EXEC_MEM_IN_250, EXEC_MEM_OUT_109, EXEC_MEM_OUT_110,
         EXEC_MEM_OUT_111, EXEC_MEM_OUT_112, EXEC_MEM_OUT_113,
         EXEC_MEM_OUT_114, EXEC_MEM_OUT_115, EXEC_MEM_OUT_116,
         EXEC_MEM_OUT_117, EXEC_MEM_OUT_118, EXEC_MEM_OUT_119,
         EXEC_MEM_OUT_120, EXEC_MEM_OUT_121, EXEC_MEM_OUT_122,
         EXEC_MEM_OUT_123, EXEC_MEM_OUT_124, EXEC_MEM_OUT_125,
         EXEC_MEM_OUT_126, EXEC_MEM_OUT_127, EXEC_MEM_OUT_128,
         EXEC_MEM_OUT_129, EXEC_MEM_OUT_130, EXEC_MEM_OUT_131,
         EXEC_MEM_OUT_132, EXEC_MEM_OUT_133, EXEC_MEM_OUT_134,
         EXEC_MEM_OUT_135, EXEC_MEM_OUT_136, EXEC_MEM_OUT_137,
         EXEC_MEM_OUT_138, EXEC_MEM_OUT_139, EXEC_MEM_OUT_140,
         EXEC_MEM_OUT_141, RegWrite_wb_out, EXEC_STAGE_mul_done,
         EXEC_STAGE_mul_ex_N479, EXEC_STAGE_mul_ex_N476,
         EXEC_STAGE_mul_ex_N475, EXEC_STAGE_mul_ex_N474,
         EXEC_STAGE_mul_ex_N473, EXEC_STAGE_mul_ex_N472,
         EXEC_STAGE_mul_ex_N471, EXEC_STAGE_mul_ex_N470,
         EXEC_STAGE_mul_ex_N469, EXEC_STAGE_mul_ex_N468,
         EXEC_STAGE_mul_ex_N467, EXEC_STAGE_mul_ex_N466,
         EXEC_STAGE_mul_ex_N465, EXEC_STAGE_mul_ex_N464,
         EXEC_STAGE_mul_ex_N463, EXEC_STAGE_mul_ex_N462,
         EXEC_STAGE_mul_ex_N461, EXEC_STAGE_mul_ex_N460,
         EXEC_STAGE_mul_ex_N459, EXEC_STAGE_mul_ex_N458,
         EXEC_STAGE_mul_ex_N457, EXEC_STAGE_mul_ex_N456,
         EXEC_STAGE_mul_ex_N455, EXEC_STAGE_mul_ex_N454,
         EXEC_STAGE_mul_ex_N453, EXEC_STAGE_mul_ex_N452,
         EXEC_STAGE_mul_ex_N451, EXEC_STAGE_mul_ex_N450,
         EXEC_STAGE_mul_ex_N449, EXEC_STAGE_mul_ex_N448,
         EXEC_STAGE_mul_ex_N447, EXEC_STAGE_mul_ex_N446,
         EXEC_STAGE_mul_ex_N445, EXEC_STAGE_mul_ex_N444,
         EXEC_STAGE_mul_ex_N443, EXEC_STAGE_mul_ex_N442,
         EXEC_STAGE_mul_ex_N441, EXEC_STAGE_mul_ex_N440,
         EXEC_STAGE_mul_ex_N439, EXEC_STAGE_mul_ex_N438,
         EXEC_STAGE_mul_ex_N437, EXEC_STAGE_mul_ex_N436,
         EXEC_STAGE_mul_ex_N435, EXEC_STAGE_mul_ex_N434,
         EXEC_STAGE_mul_ex_N433, EXEC_STAGE_mul_ex_N432,
         EXEC_STAGE_mul_ex_N431, EXEC_STAGE_mul_ex_N430,
         EXEC_STAGE_mul_ex_N429, EXEC_STAGE_mul_ex_N428,
         EXEC_STAGE_mul_ex_N427, EXEC_STAGE_mul_ex_N426,
         EXEC_STAGE_mul_ex_N425, EXEC_STAGE_mul_ex_N424,
         EXEC_STAGE_mul_ex_N423, EXEC_STAGE_mul_ex_N422,
         EXEC_STAGE_mul_ex_N421, EXEC_STAGE_mul_ex_N420,
         EXEC_STAGE_mul_ex_N419, EXEC_STAGE_mul_ex_N418,
         EXEC_STAGE_mul_ex_N417, EXEC_STAGE_mul_ex_N416,
         EXEC_STAGE_mul_ex_N415, EXEC_STAGE_mul_ex_N414,
         EXEC_STAGE_mul_ex_N413, EXEC_STAGE_mul_ex_N412,
         EXEC_STAGE_mul_ex_N411, EXEC_STAGE_mul_ex_N410,
         EXEC_STAGE_mul_ex_N409, EXEC_STAGE_mul_ex_N408,
         EXEC_STAGE_mul_ex_N407, EXEC_STAGE_mul_ex_N406,
         EXEC_STAGE_mul_ex_N405, EXEC_STAGE_mul_ex_N404,
         EXEC_STAGE_mul_ex_N403, EXEC_STAGE_mul_ex_N402,
         EXEC_STAGE_mul_ex_N401, EXEC_STAGE_mul_ex_N400,
         EXEC_STAGE_mul_ex_N399, EXEC_STAGE_mul_ex_N398,
         EXEC_STAGE_mul_ex_N397, EXEC_STAGE_mul_ex_N396,
         EXEC_STAGE_mul_ex_N395, EXEC_STAGE_mul_ex_N394,
         EXEC_STAGE_mul_ex_N393, EXEC_STAGE_mul_ex_N392,
         EXEC_STAGE_mul_ex_N391, EXEC_STAGE_mul_ex_N390,
         EXEC_STAGE_mul_ex_N389, EXEC_STAGE_mul_ex_N388,
         EXEC_STAGE_mul_ex_N387, EXEC_STAGE_mul_ex_N386,
         EXEC_STAGE_mul_ex_N385, EXEC_STAGE_mul_ex_N384,
         EXEC_STAGE_mul_ex_N383, EXEC_STAGE_mul_ex_N382,
         EXEC_STAGE_mul_ex_N381, EXEC_STAGE_mul_ex_N380,
         EXEC_STAGE_mul_ex_N379, EXEC_STAGE_mul_ex_N378,
         EXEC_STAGE_mul_ex_N377, EXEC_STAGE_mul_ex_N376,
         EXEC_STAGE_mul_ex_N375, EXEC_STAGE_mul_ex_N374,
         EXEC_STAGE_mul_ex_N373, EXEC_STAGE_mul_ex_N372,
         EXEC_STAGE_mul_ex_N371, EXEC_STAGE_mul_ex_N370,
         EXEC_STAGE_mul_ex_N369, EXEC_STAGE_mul_ex_N368,
         EXEC_STAGE_mul_ex_N367, EXEC_STAGE_mul_ex_N366,
         EXEC_STAGE_mul_ex_N365, EXEC_STAGE_mul_ex_N364,
         EXEC_STAGE_mul_ex_N363, EXEC_STAGE_mul_ex_N362,
         EXEC_STAGE_mul_ex_N361, EXEC_STAGE_mul_ex_N360,
         EXEC_STAGE_mul_ex_N359, EXEC_STAGE_mul_ex_N358,
         EXEC_STAGE_mul_ex_N357, EXEC_STAGE_mul_ex_N356,
         EXEC_STAGE_mul_ex_N355, EXEC_STAGE_mul_ex_N354,
         EXEC_STAGE_mul_ex_N353, EXEC_STAGE_mul_ex_N352,
         EXEC_STAGE_mul_ex_N351, EXEC_STAGE_mul_ex_N350,
         EXEC_STAGE_mul_ex_N349, EXEC_STAGE_mul_ex_N348,
         EXEC_STAGE_mul_ex_N347, EXEC_STAGE_mul_ex_N346,
         EXEC_STAGE_mul_ex_N345, EXEC_STAGE_mul_ex_N344,
         EXEC_STAGE_mul_ex_N343, EXEC_STAGE_mul_ex_N342,
         EXEC_STAGE_mul_ex_N341, EXEC_STAGE_mul_ex_N340,
         EXEC_STAGE_mul_ex_N339, EXEC_STAGE_mul_ex_N338,
         EXEC_STAGE_mul_ex_N337, EXEC_STAGE_mul_ex_N336,
         EXEC_STAGE_mul_ex_N335, EXEC_STAGE_mul_ex_N334,
         EXEC_STAGE_mul_ex_N333, EXEC_STAGE_mul_ex_N332,
         EXEC_STAGE_mul_ex_N331, EXEC_STAGE_mul_ex_N330,
         EXEC_STAGE_mul_ex_N329, EXEC_STAGE_mul_ex_N328,
         EXEC_STAGE_mul_ex_N327, EXEC_STAGE_mul_ex_N326,
         EXEC_STAGE_mul_ex_N325, EXEC_STAGE_mul_ex_N324,
         EXEC_STAGE_mul_ex_N323, EXEC_STAGE_mul_ex_N322,
         EXEC_STAGE_mul_ex_N321, EXEC_STAGE_mul_ex_N320,
         EXEC_STAGE_mul_ex_N319, EXEC_STAGE_mul_ex_N318,
         EXEC_STAGE_mul_ex_N317, EXEC_STAGE_mul_ex_N316,
         EXEC_STAGE_mul_ex_N315, EXEC_STAGE_mul_ex_N314,
         EXEC_STAGE_mul_ex_N249, EXEC_STAGE_mul_ex_N248,
         EXEC_STAGE_mul_ex_N247, EXEC_STAGE_mul_ex_N246,
         EXEC_STAGE_mul_ex_N245, EXEC_STAGE_mul_ex_N244,
         EXEC_STAGE_mul_ex_N243, EXEC_STAGE_mul_ex_N242,
         EXEC_STAGE_mul_ex_N241, EXEC_STAGE_mul_ex_N240,
         EXEC_STAGE_mul_ex_N239, EXEC_STAGE_mul_ex_N238,
         EXEC_STAGE_mul_ex_N237, EXEC_STAGE_mul_ex_N236,
         EXEC_STAGE_mul_ex_N235, EXEC_STAGE_mul_ex_N234,
         EXEC_STAGE_mul_ex_N233, EXEC_STAGE_mul_ex_N232,
         EXEC_STAGE_mul_ex_N231, EXEC_STAGE_mul_ex_N230,
         EXEC_STAGE_mul_ex_N229, EXEC_STAGE_mul_ex_N228,
         EXEC_STAGE_mul_ex_N227, EXEC_STAGE_mul_ex_N226,
         EXEC_STAGE_mul_ex_N225, EXEC_STAGE_mul_ex_N224,
         EXEC_STAGE_mul_ex_N223, EXEC_STAGE_mul_ex_N222,
         EXEC_STAGE_mul_ex_N221, EXEC_STAGE_mul_ex_N220,
         EXEC_STAGE_mul_ex_N219, EXEC_STAGE_mul_ex_N218,
         EXEC_STAGE_mul_ex_N185, EXEC_STAGE_mul_ex_N184,
         EXEC_STAGE_mul_ex_N183, EXEC_STAGE_mul_ex_N182,
         EXEC_STAGE_mul_ex_N181, EXEC_STAGE_mul_ex_N180,
         EXEC_STAGE_mul_ex_N179, EXEC_STAGE_mul_ex_N178,
         EXEC_STAGE_mul_ex_N177, EXEC_STAGE_mul_ex_N176,
         EXEC_STAGE_mul_ex_N175, EXEC_STAGE_mul_ex_N174,
         EXEC_STAGE_mul_ex_N173, EXEC_STAGE_mul_ex_N172,
         EXEC_STAGE_mul_ex_N171, EXEC_STAGE_mul_ex_N170,
         EXEC_STAGE_mul_ex_N169, EXEC_STAGE_mul_ex_N168,
         EXEC_STAGE_mul_ex_N167, EXEC_STAGE_mul_ex_N166,
         EXEC_STAGE_mul_ex_N165, EXEC_STAGE_mul_ex_N164,
         EXEC_STAGE_mul_ex_N163, EXEC_STAGE_mul_ex_N162,
         EXEC_STAGE_mul_ex_N161, EXEC_STAGE_mul_ex_N160,
         EXEC_STAGE_mul_ex_N159, EXEC_STAGE_mul_ex_N158,
         EXEC_STAGE_mul_ex_N157, EXEC_STAGE_mul_ex_N156,
         EXEC_STAGE_mul_ex_N155, EXEC_STAGE_mul_ex_N154,
         EXEC_STAGE_mul_ex_N119, EXEC_STAGE_mul_ex_N118,
         EXEC_STAGE_mul_ex_N117, EXEC_STAGE_mul_ex_N116,
         EXEC_STAGE_mul_ex_N115, EXEC_STAGE_mul_ex_N114,
         EXEC_STAGE_mul_ex_N113, EXEC_STAGE_mul_ex_N112,
         EXEC_STAGE_mul_ex_N111, EXEC_STAGE_mul_ex_N110,
         EXEC_STAGE_mul_ex_N109, EXEC_STAGE_mul_ex_N108,
         EXEC_STAGE_mul_ex_N107, EXEC_STAGE_mul_ex_N106,
         EXEC_STAGE_mul_ex_N105, EXEC_STAGE_mul_ex_N104,
         EXEC_STAGE_mul_ex_N103, EXEC_STAGE_mul_ex_N102,
         EXEC_STAGE_mul_ex_N101, EXEC_STAGE_mul_ex_N100, EXEC_STAGE_mul_ex_N99,
         EXEC_STAGE_mul_ex_N98, EXEC_STAGE_mul_ex_N97, EXEC_STAGE_mul_ex_N96,
         EXEC_STAGE_mul_ex_N95, EXEC_STAGE_mul_ex_N94, EXEC_STAGE_mul_ex_N93,
         EXEC_STAGE_mul_ex_N92, EXEC_STAGE_mul_ex_N91, EXEC_STAGE_mul_ex_N90,
         EXEC_STAGE_mul_ex_N89, EXEC_STAGE_mul_ex_N88, EXEC_STAGE_mul_ex_N87,
         EXEC_STAGE_mul_ex_N86, EXEC_STAGE_mul_ex_N85, EXEC_STAGE_mul_ex_N84,
         EXEC_STAGE_mul_ex_N83, EXEC_STAGE_mul_ex_N82, EXEC_STAGE_mul_ex_N81,
         EXEC_STAGE_mul_ex_N80, EXEC_STAGE_mul_ex_N79, EXEC_STAGE_mul_ex_N78,
         EXEC_STAGE_mul_ex_N77, EXEC_STAGE_mul_ex_N76, EXEC_STAGE_mul_ex_N75,
         EXEC_STAGE_mul_ex_N74, EXEC_STAGE_mul_ex_N73, EXEC_STAGE_mul_ex_N72,
         EXEC_STAGE_mul_ex_N71, EXEC_STAGE_mul_ex_N70, EXEC_STAGE_mul_ex_N69,
         EXEC_STAGE_mul_ex_N68, EXEC_STAGE_mul_ex_N67, EXEC_STAGE_mul_ex_N66,
         EXEC_STAGE_mul_ex_N65, EXEC_STAGE_mul_ex_N64, EXEC_STAGE_mul_ex_N63,
         EXEC_STAGE_mul_ex_N62, EXEC_STAGE_mul_ex_N61, EXEC_STAGE_mul_ex_N60,
         EXEC_STAGE_mul_ex_N59, EXEC_STAGE_mul_ex_N58, EXEC_STAGE_mul_ex_N57,
         EXEC_STAGE_mul_ex_N56, EXEC_STAGE_mul_ex_Z_31_,
         EXEC_STAGE_mul_ex_Z_30_, EXEC_STAGE_mul_ex_Z_29_,
         EXEC_STAGE_mul_ex_Z_28_, EXEC_STAGE_mul_ex_Z_27_,
         EXEC_STAGE_mul_ex_Z_26_, EXEC_STAGE_mul_ex_Z_25_,
         EXEC_STAGE_mul_ex_Z_24_, EXEC_STAGE_mul_ex_Z_23_,
         EXEC_STAGE_mul_ex_Z_22_, EXEC_STAGE_mul_ex_Z_21_,
         EXEC_STAGE_mul_ex_Z_20_, EXEC_STAGE_mul_ex_Z_19_,
         EXEC_STAGE_mul_ex_Z_18_, EXEC_STAGE_mul_ex_Z_17_,
         EXEC_STAGE_mul_ex_Z_16_, EXEC_STAGE_mul_ex_Z_15_,
         EXEC_STAGE_mul_ex_Z_14_, EXEC_STAGE_mul_ex_Z_13_,
         EXEC_STAGE_mul_ex_Z_12_, EXEC_STAGE_mul_ex_Z_11_,
         EXEC_STAGE_mul_ex_Z_10_, EXEC_STAGE_mul_ex_Z_9_,
         EXEC_STAGE_mul_ex_Z_8_, EXEC_STAGE_mul_ex_Z_7_,
         EXEC_STAGE_mul_ex_Z_6_, EXEC_STAGE_mul_ex_Z_5_,
         EXEC_STAGE_mul_ex_Z_4_, EXEC_STAGE_mul_ex_Z_3_,
         EXEC_STAGE_mul_ex_Z_2_, EXEC_STAGE_mul_ex_Z_1_,
         EXEC_STAGE_mul_ex_Z_0_, EXEC_STAGE_mul_ex_L_31_,
         EXEC_STAGE_mul_ex_L_30_, EXEC_STAGE_mul_ex_L_29_,
         EXEC_STAGE_mul_ex_L_28_, EXEC_STAGE_mul_ex_L_27_,
         EXEC_STAGE_mul_ex_L_26_, EXEC_STAGE_mul_ex_L_25_,
         EXEC_STAGE_mul_ex_L_24_, EXEC_STAGE_mul_ex_L_23_,
         EXEC_STAGE_mul_ex_L_22_, EXEC_STAGE_mul_ex_L_21_,
         EXEC_STAGE_mul_ex_L_20_, EXEC_STAGE_mul_ex_L_19_,
         EXEC_STAGE_mul_ex_L_18_, EXEC_STAGE_mul_ex_L_17_,
         EXEC_STAGE_mul_ex_L_16_, EXEC_STAGE_mul_ex_L_15_,
         EXEC_STAGE_mul_ex_L_14_, EXEC_STAGE_mul_ex_L_13_,
         EXEC_STAGE_mul_ex_L_12_, EXEC_STAGE_mul_ex_L_11_,
         EXEC_STAGE_mul_ex_L_10_, EXEC_STAGE_mul_ex_L_9_,
         EXEC_STAGE_mul_ex_L_8_, EXEC_STAGE_mul_ex_L_7_,
         EXEC_STAGE_mul_ex_L_6_, EXEC_STAGE_mul_ex_L_5_,
         EXEC_STAGE_mul_ex_L_4_, EXEC_STAGE_mul_ex_L_3_,
         EXEC_STAGE_mul_ex_L_2_, EXEC_STAGE_mul_ex_L_1_,
         EXEC_STAGE_mul_ex_L_0_, EXEC_STAGE_mul_ex_N16, EXEC_STAGE_mul_ex_N15,
         EXEC_STAGE_mul_ex_N14, EXEC_STAGE_mul_ex_CurrentState_2_,
         EXEC_STAGE_mul_ex_CurrentState_1_, EXEC_STAGE_mul_ex_CurrentState_0_,
         MEM_WB_REG_MEM_WB_REG_N179, MEM_WB_REG_MEM_WB_REG_N178,
         MEM_WB_REG_MEM_WB_REG_N177, MEM_WB_REG_MEM_WB_REG_N176,
         MEM_WB_REG_MEM_WB_REG_N175, MEM_WB_REG_MEM_WB_REG_N174,
         MEM_WB_REG_MEM_WB_REG_N173, MEM_WB_REG_MEM_WB_REG_N172,
         MEM_WB_REG_MEM_WB_REG_N171, MEM_WB_REG_MEM_WB_REG_N170,
         MEM_WB_REG_MEM_WB_REG_N169, MEM_WB_REG_MEM_WB_REG_N168,
         MEM_WB_REG_MEM_WB_REG_N167, MEM_WB_REG_MEM_WB_REG_N166,
         MEM_WB_REG_MEM_WB_REG_N165, MEM_WB_REG_MEM_WB_REG_N163,
         MEM_WB_REG_MEM_WB_REG_N160, MEM_WB_REG_MEM_WB_REG_N158,
         MEM_WB_REG_MEM_WB_REG_N156, MEM_WB_REG_MEM_WB_REG_N152,
         MEM_WB_REG_MEM_WB_REG_N148, MEM_WB_REG_MEM_WB_REG_N147,
         MEM_WB_REG_MEM_WB_REG_N146, MEM_WB_REG_MEM_WB_REG_N145,
         MEM_WB_REG_MEM_WB_REG_N144, MEM_WB_REG_MEM_WB_REG_N78,
         MEM_WB_REG_MEM_WB_REG_N77, MEM_WB_REG_MEM_WB_REG_N76,
         MEM_WB_REG_MEM_WB_REG_N75, MEM_WB_REG_MEM_WB_REG_N66,
         MEM_WB_REG_MEM_WB_REG_N65, MEM_WB_REG_MEM_WB_REG_N64,
         MEM_WB_REG_MEM_WB_REG_N63, MEM_WB_REG_MEM_WB_REG_N62,
         MEM_WB_REG_MEM_WB_REG_N61, MEM_WB_REG_MEM_WB_REG_N60,
         MEM_WB_REG_MEM_WB_REG_N59, MEM_WB_REG_MEM_WB_REG_N58,
         MEM_WB_REG_MEM_WB_REG_N57, MEM_WB_REG_MEM_WB_REG_N56,
         MEM_WB_REG_MEM_WB_REG_N55, MEM_WB_REG_MEM_WB_REG_N54,
         MEM_WB_REG_MEM_WB_REG_N53, MEM_WB_REG_MEM_WB_REG_N52,
         MEM_WB_REG_MEM_WB_REG_N51, MEM_WB_REG_MEM_WB_REG_N50,
         MEM_WB_REG_MEM_WB_REG_N49, MEM_WB_REG_MEM_WB_REG_N48,
         MEM_WB_REG_MEM_WB_REG_N47, MEM_WB_REG_MEM_WB_REG_N46,
         MEM_WB_REG_MEM_WB_REG_N45, MEM_WB_REG_MEM_WB_REG_N44,
         MEM_WB_REG_MEM_WB_REG_N43, MEM_WB_REG_MEM_WB_REG_N42,
         MEM_WB_REG_MEM_WB_REG_N41, MEM_WB_REG_MEM_WB_REG_N40,
         MEM_WB_REG_MEM_WB_REG_N39, MEM_WB_REG_MEM_WB_REG_N38,
         MEM_WB_REG_MEM_WB_REG_N37, MEM_WB_REG_MEM_WB_REG_N36,
         MEM_WB_REG_MEM_WB_REG_N35, REG_FILE_reg_out_29__31_,
         REG_FILE_reg_out_29__30_, REG_FILE_reg_out_29__29_,
         REG_FILE_reg_out_29__28_, REG_FILE_reg_out_29__27_,
         REG_FILE_reg_out_29__26_, REG_FILE_reg_out_29__25_,
         REG_FILE_reg_out_29__24_, REG_FILE_reg_out_29__23_,
         REG_FILE_reg_out_29__22_, REG_FILE_reg_out_29__21_,
         REG_FILE_reg_out_29__20_, REG_FILE_reg_out_29__19_,
         REG_FILE_reg_out_29__18_, REG_FILE_reg_out_29__17_,
         REG_FILE_reg_out_29__16_, REG_FILE_reg_out_27__31_,
         REG_FILE_reg_out_27__30_, REG_FILE_reg_out_27__29_,
         REG_FILE_reg_out_27__28_, REG_FILE_reg_out_27__27_,
         REG_FILE_reg_out_27__26_, REG_FILE_reg_out_27__25_,
         REG_FILE_reg_out_27__24_, REG_FILE_reg_out_27__23_,
         REG_FILE_reg_out_27__22_, REG_FILE_reg_out_27__21_,
         REG_FILE_reg_out_27__20_, REG_FILE_reg_out_27__19_,
         REG_FILE_reg_out_27__18_, REG_FILE_reg_out_27__17_,
         REG_FILE_reg_out_27__16_, REG_FILE_reg_out_26__31_,
         REG_FILE_reg_out_26__30_, REG_FILE_reg_out_26__29_,
         REG_FILE_reg_out_26__28_, REG_FILE_reg_out_26__27_,
         REG_FILE_reg_out_26__26_, REG_FILE_reg_out_26__25_,
         REG_FILE_reg_out_26__24_, REG_FILE_reg_out_26__23_,
         REG_FILE_reg_out_26__22_, REG_FILE_reg_out_26__21_,
         REG_FILE_reg_out_26__20_, REG_FILE_reg_out_26__19_,
         REG_FILE_reg_out_26__18_, REG_FILE_reg_out_26__17_,
         REG_FILE_reg_out_26__16_, REG_FILE_reg_out_26__15_,
         REG_FILE_reg_out_26__14_, REG_FILE_reg_out_26__13_,
         REG_FILE_reg_out_26__12_, REG_FILE_reg_out_26__11_,
         REG_FILE_reg_out_26__10_, REG_FILE_reg_out_26__9_,
         REG_FILE_reg_out_26__8_, REG_FILE_reg_out_26__7_,
         REG_FILE_reg_out_26__6_, REG_FILE_reg_out_26__5_,
         REG_FILE_reg_out_26__4_, REG_FILE_reg_out_26__3_,
         REG_FILE_reg_out_26__2_, REG_FILE_reg_out_26__1_,
         REG_FILE_reg_out_26__0_, REG_FILE_reg_out_25__31_,
         REG_FILE_reg_out_25__30_, REG_FILE_reg_out_25__29_,
         REG_FILE_reg_out_25__28_, REG_FILE_reg_out_25__27_,
         REG_FILE_reg_out_25__26_, REG_FILE_reg_out_25__25_,
         REG_FILE_reg_out_25__24_, REG_FILE_reg_out_25__23_,
         REG_FILE_reg_out_25__22_, REG_FILE_reg_out_25__21_,
         REG_FILE_reg_out_25__20_, REG_FILE_reg_out_25__19_,
         REG_FILE_reg_out_25__18_, REG_FILE_reg_out_25__17_,
         REG_FILE_reg_out_25__16_, REG_FILE_reg_out_25__15_,
         REG_FILE_reg_out_25__14_, REG_FILE_reg_out_25__13_,
         REG_FILE_reg_out_25__12_, REG_FILE_reg_out_25__11_,
         REG_FILE_reg_out_25__10_, REG_FILE_reg_out_25__9_,
         REG_FILE_reg_out_25__8_, REG_FILE_reg_out_25__7_,
         REG_FILE_reg_out_25__6_, REG_FILE_reg_out_25__5_,
         REG_FILE_reg_out_25__4_, REG_FILE_reg_out_25__3_,
         REG_FILE_reg_out_25__2_, REG_FILE_reg_out_25__1_,
         REG_FILE_reg_out_25__0_, REG_FILE_reg_out_24__31_,
         REG_FILE_reg_out_22__30_, REG_FILE_reg_out_22__29_,
         REG_FILE_reg_out_22__28_, REG_FILE_reg_out_22__27_,
         REG_FILE_reg_out_22__26_, REG_FILE_reg_out_22__25_,
         REG_FILE_reg_out_22__24_, REG_FILE_reg_out_22__23_,
         REG_FILE_reg_out_22__22_, REG_FILE_reg_out_22__21_,
         REG_FILE_reg_out_22__20_, REG_FILE_reg_out_22__19_,
         REG_FILE_reg_out_22__18_, REG_FILE_reg_out_22__17_,
         REG_FILE_reg_out_22__16_, REG_FILE_reg_out_20__31_,
         REG_FILE_reg_out_20__30_, REG_FILE_reg_out_20__29_,
         REG_FILE_reg_out_20__28_, REG_FILE_reg_out_20__27_,
         REG_FILE_reg_out_20__26_, REG_FILE_reg_out_20__25_,
         REG_FILE_reg_out_20__24_, REG_FILE_reg_out_20__23_,
         REG_FILE_reg_out_20__22_, REG_FILE_reg_out_20__21_,
         REG_FILE_reg_out_20__20_, REG_FILE_reg_out_20__19_,
         REG_FILE_reg_out_20__18_, REG_FILE_reg_out_20__17_,
         REG_FILE_reg_out_20__16_, REG_FILE_reg_out_19__30_,
         REG_FILE_reg_out_19__29_, REG_FILE_reg_out_19__28_,
         REG_FILE_reg_out_19__27_, REG_FILE_reg_out_19__26_,
         REG_FILE_reg_out_19__25_, REG_FILE_reg_out_19__24_,
         REG_FILE_reg_out_19__23_, REG_FILE_reg_out_19__22_,
         REG_FILE_reg_out_19__21_, REG_FILE_reg_out_19__20_,
         REG_FILE_reg_out_19__19_, REG_FILE_reg_out_19__18_,
         REG_FILE_reg_out_19__17_, REG_FILE_reg_out_19__16_,
         REG_FILE_reg_out_19__15_, REG_FILE_reg_out_19__14_,
         REG_FILE_reg_out_19__13_, REG_FILE_reg_out_19__12_,
         REG_FILE_reg_out_19__11_, REG_FILE_reg_out_19__10_,
         REG_FILE_reg_out_19__9_, REG_FILE_reg_out_19__8_,
         REG_FILE_reg_out_19__7_, REG_FILE_reg_out_19__6_,
         REG_FILE_reg_out_19__5_, REG_FILE_reg_out_19__4_,
         REG_FILE_reg_out_19__3_, REG_FILE_reg_out_19__2_,
         REG_FILE_reg_out_19__1_, REG_FILE_reg_out_19__0_,
         REG_FILE_reg_out_18__31_, REG_FILE_reg_out_17__31_,
         REG_FILE_reg_out_17__30_, REG_FILE_reg_out_17__29_,
         REG_FILE_reg_out_17__28_, REG_FILE_reg_out_17__27_,
         REG_FILE_reg_out_17__26_, REG_FILE_reg_out_17__25_,
         REG_FILE_reg_out_17__24_, REG_FILE_reg_out_17__23_,
         REG_FILE_reg_out_17__22_, REG_FILE_reg_out_17__21_,
         REG_FILE_reg_out_17__20_, REG_FILE_reg_out_17__19_,
         REG_FILE_reg_out_17__18_, REG_FILE_reg_out_17__17_,
         REG_FILE_reg_out_17__16_, REG_FILE_reg_out_17__15_,
         REG_FILE_reg_out_17__14_, REG_FILE_reg_out_17__13_,
         REG_FILE_reg_out_17__12_, REG_FILE_reg_out_17__11_,
         REG_FILE_reg_out_17__10_, REG_FILE_reg_out_17__9_,
         REG_FILE_reg_out_17__8_, REG_FILE_reg_out_17__7_,
         REG_FILE_reg_out_17__6_, REG_FILE_reg_out_17__5_,
         REG_FILE_reg_out_17__4_, REG_FILE_reg_out_17__3_,
         REG_FILE_reg_out_17__2_, REG_FILE_reg_out_17__1_,
         REG_FILE_reg_out_17__0_, REG_FILE_reg_out_15__31_,
         REG_FILE_reg_out_15__15_, REG_FILE_reg_out_15__14_,
         REG_FILE_reg_out_15__13_, REG_FILE_reg_out_15__12_,
         REG_FILE_reg_out_15__11_, REG_FILE_reg_out_15__10_,
         REG_FILE_reg_out_15__9_, REG_FILE_reg_out_15__8_,
         REG_FILE_reg_out_15__7_, REG_FILE_reg_out_15__6_,
         REG_FILE_reg_out_15__5_, REG_FILE_reg_out_15__4_,
         REG_FILE_reg_out_15__3_, REG_FILE_reg_out_15__2_,
         REG_FILE_reg_out_15__1_, REG_FILE_reg_out_15__0_,
         REG_FILE_reg_out_14__31_, REG_FILE_reg_out_14__30_,
         REG_FILE_reg_out_14__29_, REG_FILE_reg_out_14__28_,
         REG_FILE_reg_out_14__27_, REG_FILE_reg_out_14__26_,
         REG_FILE_reg_out_14__25_, REG_FILE_reg_out_14__24_,
         REG_FILE_reg_out_14__23_, REG_FILE_reg_out_14__22_,
         REG_FILE_reg_out_14__21_, REG_FILE_reg_out_14__20_,
         REG_FILE_reg_out_14__19_, REG_FILE_reg_out_14__18_,
         REG_FILE_reg_out_14__17_, REG_FILE_reg_out_14__16_,
         REG_FILE_reg_out_13__31_, REG_FILE_reg_out_13__30_,
         REG_FILE_reg_out_13__29_, REG_FILE_reg_out_13__28_,
         REG_FILE_reg_out_13__27_, REG_FILE_reg_out_13__26_,
         REG_FILE_reg_out_13__25_, REG_FILE_reg_out_13__24_,
         REG_FILE_reg_out_13__23_, REG_FILE_reg_out_13__22_,
         REG_FILE_reg_out_13__21_, REG_FILE_reg_out_13__20_,
         REG_FILE_reg_out_13__19_, REG_FILE_reg_out_13__18_,
         REG_FILE_reg_out_13__17_, REG_FILE_reg_out_13__16_,
         REG_FILE_reg_out_13__15_, REG_FILE_reg_out_13__14_,
         REG_FILE_reg_out_13__13_, REG_FILE_reg_out_13__12_,
         REG_FILE_reg_out_13__11_, REG_FILE_reg_out_13__10_,
         REG_FILE_reg_out_13__9_, REG_FILE_reg_out_13__8_,
         REG_FILE_reg_out_13__7_, REG_FILE_reg_out_13__6_,
         REG_FILE_reg_out_13__5_, REG_FILE_reg_out_13__4_,
         REG_FILE_reg_out_13__3_, REG_FILE_reg_out_13__2_,
         REG_FILE_reg_out_13__1_, REG_FILE_reg_out_13__0_,
         REG_FILE_reg_out_12__31_, REG_FILE_reg_out_12__30_,
         REG_FILE_reg_out_12__29_, REG_FILE_reg_out_12__28_,
         REG_FILE_reg_out_12__27_, REG_FILE_reg_out_12__26_,
         REG_FILE_reg_out_12__25_, REG_FILE_reg_out_12__24_,
         REG_FILE_reg_out_12__23_, REG_FILE_reg_out_12__22_,
         REG_FILE_reg_out_12__21_, REG_FILE_reg_out_12__20_,
         REG_FILE_reg_out_12__19_, REG_FILE_reg_out_12__18_,
         REG_FILE_reg_out_12__17_, REG_FILE_reg_out_12__16_,
         REG_FILE_reg_out_12__15_, REG_FILE_reg_out_12__14_,
         REG_FILE_reg_out_12__13_, REG_FILE_reg_out_12__12_,
         REG_FILE_reg_out_12__11_, REG_FILE_reg_out_12__10_,
         REG_FILE_reg_out_12__9_, REG_FILE_reg_out_12__8_,
         REG_FILE_reg_out_12__7_, REG_FILE_reg_out_12__6_,
         REG_FILE_reg_out_12__5_, REG_FILE_reg_out_12__4_,
         REG_FILE_reg_out_12__3_, REG_FILE_reg_out_12__2_,
         REG_FILE_reg_out_12__1_, REG_FILE_reg_out_12__0_,
         REG_FILE_reg_out_11__30_, REG_FILE_reg_out_11__29_,
         REG_FILE_reg_out_11__28_, REG_FILE_reg_out_11__27_,
         REG_FILE_reg_out_11__26_, REG_FILE_reg_out_11__25_,
         REG_FILE_reg_out_11__24_, REG_FILE_reg_out_11__23_,
         REG_FILE_reg_out_11__22_, REG_FILE_reg_out_11__21_,
         REG_FILE_reg_out_11__20_, REG_FILE_reg_out_11__19_,
         REG_FILE_reg_out_11__18_, REG_FILE_reg_out_11__17_,
         REG_FILE_reg_out_11__16_, REG_FILE_reg_out_9__15_,
         REG_FILE_reg_out_9__13_, REG_FILE_reg_out_9__11_,
         REG_FILE_reg_out_9__10_, REG_FILE_reg_out_9__9_,
         REG_FILE_reg_out_9__6_, REG_FILE_reg_out_9__4_,
         REG_FILE_reg_out_9__3_, REG_FILE_reg_out_7__30_,
         REG_FILE_reg_out_7__29_, REG_FILE_reg_out_7__28_,
         REG_FILE_reg_out_7__27_, REG_FILE_reg_out_7__26_,
         REG_FILE_reg_out_7__25_, REG_FILE_reg_out_7__24_,
         REG_FILE_reg_out_7__23_, REG_FILE_reg_out_7__22_,
         REG_FILE_reg_out_7__21_, REG_FILE_reg_out_7__20_,
         REG_FILE_reg_out_7__19_, REG_FILE_reg_out_7__18_,
         REG_FILE_reg_out_7__17_, REG_FILE_reg_out_7__16_,
         REG_FILE_reg_out_6__31_, REG_FILE_reg_out_6__30_,
         REG_FILE_reg_out_6__29_, REG_FILE_reg_out_6__28_,
         REG_FILE_reg_out_6__27_, REG_FILE_reg_out_6__26_,
         REG_FILE_reg_out_6__25_, REG_FILE_reg_out_6__24_,
         REG_FILE_reg_out_6__23_, REG_FILE_reg_out_6__22_,
         REG_FILE_reg_out_6__21_, REG_FILE_reg_out_6__20_,
         REG_FILE_reg_out_6__19_, REG_FILE_reg_out_6__18_,
         REG_FILE_reg_out_6__17_, REG_FILE_reg_out_6__16_,
         REG_FILE_reg_out_5__30_, REG_FILE_reg_out_5__29_,
         REG_FILE_reg_out_5__28_, REG_FILE_reg_out_5__27_,
         REG_FILE_reg_out_5__26_, REG_FILE_reg_out_5__25_,
         REG_FILE_reg_out_5__24_, REG_FILE_reg_out_5__23_,
         REG_FILE_reg_out_5__22_, REG_FILE_reg_out_5__21_,
         REG_FILE_reg_out_5__20_, REG_FILE_reg_out_5__19_,
         REG_FILE_reg_out_5__18_, REG_FILE_reg_out_5__17_,
         REG_FILE_reg_out_5__16_, REG_FILE_reg_out_4__31_,
         REG_FILE_reg_out_4__30_, REG_FILE_reg_out_4__29_,
         REG_FILE_reg_out_4__28_, REG_FILE_reg_out_4__27_,
         REG_FILE_reg_out_4__26_, REG_FILE_reg_out_4__25_,
         REG_FILE_reg_out_4__24_, REG_FILE_reg_out_4__23_,
         REG_FILE_reg_out_4__22_, REG_FILE_reg_out_4__21_,
         REG_FILE_reg_out_4__20_, REG_FILE_reg_out_4__19_,
         REG_FILE_reg_out_4__18_, REG_FILE_reg_out_4__17_,
         REG_FILE_reg_out_4__16_, REG_FILE_reg_out_4__15_,
         REG_FILE_reg_out_4__14_, REG_FILE_reg_out_4__13_,
         REG_FILE_reg_out_4__12_, REG_FILE_reg_out_4__11_,
         REG_FILE_reg_out_4__10_, REG_FILE_reg_out_4__9_,
         REG_FILE_reg_out_4__8_, REG_FILE_reg_out_4__7_,
         REG_FILE_reg_out_4__6_, REG_FILE_reg_out_4__5_,
         REG_FILE_reg_out_4__4_, REG_FILE_reg_out_4__3_,
         REG_FILE_reg_out_4__2_, REG_FILE_reg_out_4__1_,
         REG_FILE_reg_out_4__0_, REG_FILE_reg_out_3__15_,
         REG_FILE_reg_out_3__14_, REG_FILE_reg_out_3__13_,
         REG_FILE_reg_out_3__12_, REG_FILE_reg_out_3__11_,
         REG_FILE_reg_out_3__10_, REG_FILE_reg_out_3__9_,
         REG_FILE_reg_out_3__8_, REG_FILE_reg_out_3__7_,
         REG_FILE_reg_out_3__6_, REG_FILE_reg_out_3__5_,
         REG_FILE_reg_out_3__4_, REG_FILE_reg_out_3__3_,
         REG_FILE_reg_out_3__2_, REG_FILE_reg_out_3__1_,
         REG_FILE_reg_out_3__0_, REG_FILE_reg_out_1__30_,
         REG_FILE_reg_out_1__29_, REG_FILE_reg_out_1__28_,
         REG_FILE_reg_out_1__27_, REG_FILE_reg_out_1__26_,
         REG_FILE_reg_out_1__25_, REG_FILE_reg_out_1__24_,
         REG_FILE_reg_out_1__23_, REG_FILE_reg_out_1__22_,
         REG_FILE_reg_out_1__21_, REG_FILE_reg_out_1__20_,
         REG_FILE_reg_out_1__19_, REG_FILE_reg_out_1__18_,
         REG_FILE_reg_out_1__17_, REG_FILE_reg_out_1__16_,
         REG_FILE_reg_out_0__31_, REG_FILE_reg_out_0__15_,
         REG_FILE_reg_out_0__14_, REG_FILE_reg_out_0__13_,
         REG_FILE_reg_out_0__12_, REG_FILE_reg_out_0__11_,
         REG_FILE_reg_out_0__10_, REG_FILE_reg_out_0__9_,
         REG_FILE_reg_out_0__8_, REG_FILE_reg_out_0__7_,
         REG_FILE_reg_out_0__6_, REG_FILE_reg_out_0__5_,
         REG_FILE_reg_out_0__4_, REG_FILE_reg_out_0__3_,
         REG_FILE_reg_out_0__2_, REG_FILE_reg_out_0__1_,
         REG_FILE_reg_out_0__0_, FP_REG_FILE_reg_out_30__31_,
         FP_REG_FILE_reg_out_30__30_, FP_REG_FILE_reg_out_30__29_,
         FP_REG_FILE_reg_out_30__28_, FP_REG_FILE_reg_out_30__27_,
         FP_REG_FILE_reg_out_30__26_, FP_REG_FILE_reg_out_30__25_,
         FP_REG_FILE_reg_out_30__24_, FP_REG_FILE_reg_out_30__23_,
         FP_REG_FILE_reg_out_30__22_, FP_REG_FILE_reg_out_30__21_,
         FP_REG_FILE_reg_out_30__20_, FP_REG_FILE_reg_out_30__19_,
         FP_REG_FILE_reg_out_30__18_, FP_REG_FILE_reg_out_30__17_,
         FP_REG_FILE_reg_out_30__16_, FP_REG_FILE_reg_out_30__15_,
         FP_REG_FILE_reg_out_30__14_, FP_REG_FILE_reg_out_30__13_,
         FP_REG_FILE_reg_out_30__12_, FP_REG_FILE_reg_out_30__11_,
         FP_REG_FILE_reg_out_30__10_, FP_REG_FILE_reg_out_30__9_,
         FP_REG_FILE_reg_out_30__8_, FP_REG_FILE_reg_out_30__7_,
         FP_REG_FILE_reg_out_30__6_, FP_REG_FILE_reg_out_30__5_,
         FP_REG_FILE_reg_out_30__4_, FP_REG_FILE_reg_out_30__3_,
         FP_REG_FILE_reg_out_30__2_, FP_REG_FILE_reg_out_30__1_,
         FP_REG_FILE_reg_out_30__0_, FP_REG_FILE_reg_out_29__31_,
         FP_REG_FILE_reg_out_29__30_, FP_REG_FILE_reg_out_29__29_,
         FP_REG_FILE_reg_out_29__28_, FP_REG_FILE_reg_out_29__27_,
         FP_REG_FILE_reg_out_29__26_, FP_REG_FILE_reg_out_29__25_,
         FP_REG_FILE_reg_out_29__24_, FP_REG_FILE_reg_out_29__23_,
         FP_REG_FILE_reg_out_29__22_, FP_REG_FILE_reg_out_29__21_,
         FP_REG_FILE_reg_out_29__20_, FP_REG_FILE_reg_out_29__19_,
         FP_REG_FILE_reg_out_29__18_, FP_REG_FILE_reg_out_29__17_,
         FP_REG_FILE_reg_out_29__16_, FP_REG_FILE_reg_out_29__15_,
         FP_REG_FILE_reg_out_29__14_, FP_REG_FILE_reg_out_29__13_,
         FP_REG_FILE_reg_out_29__12_, FP_REG_FILE_reg_out_29__11_,
         FP_REG_FILE_reg_out_29__10_, FP_REG_FILE_reg_out_29__9_,
         FP_REG_FILE_reg_out_29__8_, FP_REG_FILE_reg_out_29__7_,
         FP_REG_FILE_reg_out_29__6_, FP_REG_FILE_reg_out_29__5_,
         FP_REG_FILE_reg_out_29__4_, FP_REG_FILE_reg_out_29__3_,
         FP_REG_FILE_reg_out_29__2_, FP_REG_FILE_reg_out_29__1_,
         FP_REG_FILE_reg_out_29__0_, FP_REG_FILE_reg_out_28__31_,
         FP_REG_FILE_reg_out_28__30_, FP_REG_FILE_reg_out_28__29_,
         FP_REG_FILE_reg_out_28__28_, FP_REG_FILE_reg_out_28__27_,
         FP_REG_FILE_reg_out_28__26_, FP_REG_FILE_reg_out_28__25_,
         FP_REG_FILE_reg_out_28__24_, FP_REG_FILE_reg_out_28__23_,
         FP_REG_FILE_reg_out_28__22_, FP_REG_FILE_reg_out_28__21_,
         FP_REG_FILE_reg_out_28__20_, FP_REG_FILE_reg_out_28__19_,
         FP_REG_FILE_reg_out_28__18_, FP_REG_FILE_reg_out_28__17_,
         FP_REG_FILE_reg_out_28__16_, FP_REG_FILE_reg_out_28__15_,
         FP_REG_FILE_reg_out_28__14_, FP_REG_FILE_reg_out_28__13_,
         FP_REG_FILE_reg_out_28__12_, FP_REG_FILE_reg_out_28__11_,
         FP_REG_FILE_reg_out_28__10_, FP_REG_FILE_reg_out_28__9_,
         FP_REG_FILE_reg_out_28__8_, FP_REG_FILE_reg_out_28__7_,
         FP_REG_FILE_reg_out_28__6_, FP_REG_FILE_reg_out_28__5_,
         FP_REG_FILE_reg_out_28__4_, FP_REG_FILE_reg_out_28__3_,
         FP_REG_FILE_reg_out_28__2_, FP_REG_FILE_reg_out_28__1_,
         FP_REG_FILE_reg_out_28__0_, FP_REG_FILE_reg_out_27__31_,
         FP_REG_FILE_reg_out_27__30_, FP_REG_FILE_reg_out_27__29_,
         FP_REG_FILE_reg_out_27__28_, FP_REG_FILE_reg_out_27__27_,
         FP_REG_FILE_reg_out_27__26_, FP_REG_FILE_reg_out_27__25_,
         FP_REG_FILE_reg_out_27__24_, FP_REG_FILE_reg_out_27__23_,
         FP_REG_FILE_reg_out_27__22_, FP_REG_FILE_reg_out_27__21_,
         FP_REG_FILE_reg_out_27__20_, FP_REG_FILE_reg_out_27__19_,
         FP_REG_FILE_reg_out_27__18_, FP_REG_FILE_reg_out_27__17_,
         FP_REG_FILE_reg_out_27__16_, FP_REG_FILE_reg_out_27__15_,
         FP_REG_FILE_reg_out_27__14_, FP_REG_FILE_reg_out_27__13_,
         FP_REG_FILE_reg_out_27__12_, FP_REG_FILE_reg_out_27__11_,
         FP_REG_FILE_reg_out_27__10_, FP_REG_FILE_reg_out_27__9_,
         FP_REG_FILE_reg_out_27__8_, FP_REG_FILE_reg_out_27__7_,
         FP_REG_FILE_reg_out_27__6_, FP_REG_FILE_reg_out_27__5_,
         FP_REG_FILE_reg_out_27__4_, FP_REG_FILE_reg_out_27__3_,
         FP_REG_FILE_reg_out_27__2_, FP_REG_FILE_reg_out_27__1_,
         FP_REG_FILE_reg_out_27__0_, FP_REG_FILE_reg_out_25__31_,
         FP_REG_FILE_reg_out_25__30_, FP_REG_FILE_reg_out_25__29_,
         FP_REG_FILE_reg_out_25__28_, FP_REG_FILE_reg_out_25__27_,
         FP_REG_FILE_reg_out_25__26_, FP_REG_FILE_reg_out_25__25_,
         FP_REG_FILE_reg_out_25__24_, FP_REG_FILE_reg_out_25__23_,
         FP_REG_FILE_reg_out_25__22_, FP_REG_FILE_reg_out_25__21_,
         FP_REG_FILE_reg_out_25__20_, FP_REG_FILE_reg_out_25__19_,
         FP_REG_FILE_reg_out_25__18_, FP_REG_FILE_reg_out_25__17_,
         FP_REG_FILE_reg_out_25__16_, FP_REG_FILE_reg_out_25__15_,
         FP_REG_FILE_reg_out_25__14_, FP_REG_FILE_reg_out_25__13_,
         FP_REG_FILE_reg_out_25__12_, FP_REG_FILE_reg_out_25__11_,
         FP_REG_FILE_reg_out_25__10_, FP_REG_FILE_reg_out_25__9_,
         FP_REG_FILE_reg_out_25__8_, FP_REG_FILE_reg_out_25__7_,
         FP_REG_FILE_reg_out_25__6_, FP_REG_FILE_reg_out_25__5_,
         FP_REG_FILE_reg_out_25__4_, FP_REG_FILE_reg_out_25__3_,
         FP_REG_FILE_reg_out_25__2_, FP_REG_FILE_reg_out_25__1_,
         FP_REG_FILE_reg_out_25__0_, FP_REG_FILE_reg_out_24__31_,
         FP_REG_FILE_reg_out_24__30_, FP_REG_FILE_reg_out_24__29_,
         FP_REG_FILE_reg_out_24__28_, FP_REG_FILE_reg_out_24__27_,
         FP_REG_FILE_reg_out_24__26_, FP_REG_FILE_reg_out_24__25_,
         FP_REG_FILE_reg_out_24__24_, FP_REG_FILE_reg_out_24__23_,
         FP_REG_FILE_reg_out_24__22_, FP_REG_FILE_reg_out_24__21_,
         FP_REG_FILE_reg_out_24__20_, FP_REG_FILE_reg_out_24__19_,
         FP_REG_FILE_reg_out_24__18_, FP_REG_FILE_reg_out_24__17_,
         FP_REG_FILE_reg_out_24__16_, FP_REG_FILE_reg_out_24__15_,
         FP_REG_FILE_reg_out_24__14_, FP_REG_FILE_reg_out_24__13_,
         FP_REG_FILE_reg_out_24__12_, FP_REG_FILE_reg_out_24__11_,
         FP_REG_FILE_reg_out_24__10_, FP_REG_FILE_reg_out_24__9_,
         FP_REG_FILE_reg_out_24__8_, FP_REG_FILE_reg_out_24__7_,
         FP_REG_FILE_reg_out_24__6_, FP_REG_FILE_reg_out_24__5_,
         FP_REG_FILE_reg_out_24__4_, FP_REG_FILE_reg_out_24__3_,
         FP_REG_FILE_reg_out_24__2_, FP_REG_FILE_reg_out_24__1_,
         FP_REG_FILE_reg_out_24__0_, FP_REG_FILE_reg_out_23__31_,
         FP_REG_FILE_reg_out_23__30_, FP_REG_FILE_reg_out_23__29_,
         FP_REG_FILE_reg_out_23__28_, FP_REG_FILE_reg_out_23__27_,
         FP_REG_FILE_reg_out_23__26_, FP_REG_FILE_reg_out_23__25_,
         FP_REG_FILE_reg_out_23__24_, FP_REG_FILE_reg_out_23__23_,
         FP_REG_FILE_reg_out_23__22_, FP_REG_FILE_reg_out_23__21_,
         FP_REG_FILE_reg_out_23__20_, FP_REG_FILE_reg_out_23__19_,
         FP_REG_FILE_reg_out_23__18_, FP_REG_FILE_reg_out_23__17_,
         FP_REG_FILE_reg_out_23__16_, FP_REG_FILE_reg_out_23__15_,
         FP_REG_FILE_reg_out_23__14_, FP_REG_FILE_reg_out_23__13_,
         FP_REG_FILE_reg_out_23__12_, FP_REG_FILE_reg_out_23__11_,
         FP_REG_FILE_reg_out_23__10_, FP_REG_FILE_reg_out_23__9_,
         FP_REG_FILE_reg_out_23__8_, FP_REG_FILE_reg_out_23__7_,
         FP_REG_FILE_reg_out_23__6_, FP_REG_FILE_reg_out_23__5_,
         FP_REG_FILE_reg_out_23__4_, FP_REG_FILE_reg_out_23__3_,
         FP_REG_FILE_reg_out_23__2_, FP_REG_FILE_reg_out_23__1_,
         FP_REG_FILE_reg_out_23__0_, FP_REG_FILE_reg_out_20__31_,
         FP_REG_FILE_reg_out_20__30_, FP_REG_FILE_reg_out_20__29_,
         FP_REG_FILE_reg_out_20__28_, FP_REG_FILE_reg_out_20__27_,
         FP_REG_FILE_reg_out_20__26_, FP_REG_FILE_reg_out_20__25_,
         FP_REG_FILE_reg_out_20__24_, FP_REG_FILE_reg_out_20__23_,
         FP_REG_FILE_reg_out_20__22_, FP_REG_FILE_reg_out_20__21_,
         FP_REG_FILE_reg_out_20__20_, FP_REG_FILE_reg_out_20__19_,
         FP_REG_FILE_reg_out_20__18_, FP_REG_FILE_reg_out_20__17_,
         FP_REG_FILE_reg_out_20__16_, FP_REG_FILE_reg_out_20__15_,
         FP_REG_FILE_reg_out_20__14_, FP_REG_FILE_reg_out_20__13_,
         FP_REG_FILE_reg_out_20__12_, FP_REG_FILE_reg_out_20__11_,
         FP_REG_FILE_reg_out_20__10_, FP_REG_FILE_reg_out_20__9_,
         FP_REG_FILE_reg_out_20__8_, FP_REG_FILE_reg_out_20__7_,
         FP_REG_FILE_reg_out_20__6_, FP_REG_FILE_reg_out_20__5_,
         FP_REG_FILE_reg_out_20__4_, FP_REG_FILE_reg_out_20__3_,
         FP_REG_FILE_reg_out_20__2_, FP_REG_FILE_reg_out_20__1_,
         FP_REG_FILE_reg_out_20__0_, FP_REG_FILE_reg_out_19__31_,
         FP_REG_FILE_reg_out_19__30_, FP_REG_FILE_reg_out_19__29_,
         FP_REG_FILE_reg_out_19__28_, FP_REG_FILE_reg_out_19__27_,
         FP_REG_FILE_reg_out_19__26_, FP_REG_FILE_reg_out_19__25_,
         FP_REG_FILE_reg_out_19__24_, FP_REG_FILE_reg_out_19__23_,
         FP_REG_FILE_reg_out_19__22_, FP_REG_FILE_reg_out_19__21_,
         FP_REG_FILE_reg_out_19__20_, FP_REG_FILE_reg_out_19__19_,
         FP_REG_FILE_reg_out_19__18_, FP_REG_FILE_reg_out_19__17_,
         FP_REG_FILE_reg_out_19__16_, FP_REG_FILE_reg_out_19__15_,
         FP_REG_FILE_reg_out_19__14_, FP_REG_FILE_reg_out_19__13_,
         FP_REG_FILE_reg_out_19__12_, FP_REG_FILE_reg_out_19__11_,
         FP_REG_FILE_reg_out_19__10_, FP_REG_FILE_reg_out_19__9_,
         FP_REG_FILE_reg_out_19__8_, FP_REG_FILE_reg_out_19__7_,
         FP_REG_FILE_reg_out_19__6_, FP_REG_FILE_reg_out_19__5_,
         FP_REG_FILE_reg_out_19__4_, FP_REG_FILE_reg_out_19__3_,
         FP_REG_FILE_reg_out_19__2_, FP_REG_FILE_reg_out_19__1_,
         FP_REG_FILE_reg_out_19__0_, FP_REG_FILE_reg_out_18__31_,
         FP_REG_FILE_reg_out_18__30_, FP_REG_FILE_reg_out_18__29_,
         FP_REG_FILE_reg_out_18__28_, FP_REG_FILE_reg_out_18__27_,
         FP_REG_FILE_reg_out_18__26_, FP_REG_FILE_reg_out_18__25_,
         FP_REG_FILE_reg_out_18__24_, FP_REG_FILE_reg_out_18__23_,
         FP_REG_FILE_reg_out_18__22_, FP_REG_FILE_reg_out_18__21_,
         FP_REG_FILE_reg_out_18__20_, FP_REG_FILE_reg_out_18__19_,
         FP_REG_FILE_reg_out_18__18_, FP_REG_FILE_reg_out_18__17_,
         FP_REG_FILE_reg_out_18__16_, FP_REG_FILE_reg_out_18__15_,
         FP_REG_FILE_reg_out_18__14_, FP_REG_FILE_reg_out_18__13_,
         FP_REG_FILE_reg_out_18__12_, FP_REG_FILE_reg_out_18__11_,
         FP_REG_FILE_reg_out_18__10_, FP_REG_FILE_reg_out_18__9_,
         FP_REG_FILE_reg_out_18__8_, FP_REG_FILE_reg_out_18__7_,
         FP_REG_FILE_reg_out_18__6_, FP_REG_FILE_reg_out_18__5_,
         FP_REG_FILE_reg_out_18__4_, FP_REG_FILE_reg_out_18__3_,
         FP_REG_FILE_reg_out_18__2_, FP_REG_FILE_reg_out_18__1_,
         FP_REG_FILE_reg_out_18__0_, FP_REG_FILE_reg_out_17__31_,
         FP_REG_FILE_reg_out_17__30_, FP_REG_FILE_reg_out_17__29_,
         FP_REG_FILE_reg_out_17__28_, FP_REG_FILE_reg_out_17__27_,
         FP_REG_FILE_reg_out_17__26_, FP_REG_FILE_reg_out_17__25_,
         FP_REG_FILE_reg_out_17__24_, FP_REG_FILE_reg_out_17__23_,
         FP_REG_FILE_reg_out_17__22_, FP_REG_FILE_reg_out_17__21_,
         FP_REG_FILE_reg_out_17__20_, FP_REG_FILE_reg_out_17__19_,
         FP_REG_FILE_reg_out_17__18_, FP_REG_FILE_reg_out_17__17_,
         FP_REG_FILE_reg_out_17__16_, FP_REG_FILE_reg_out_17__15_,
         FP_REG_FILE_reg_out_17__14_, FP_REG_FILE_reg_out_17__13_,
         FP_REG_FILE_reg_out_17__12_, FP_REG_FILE_reg_out_17__11_,
         FP_REG_FILE_reg_out_17__10_, FP_REG_FILE_reg_out_17__9_,
         FP_REG_FILE_reg_out_17__8_, FP_REG_FILE_reg_out_17__7_,
         FP_REG_FILE_reg_out_17__6_, FP_REG_FILE_reg_out_17__5_,
         FP_REG_FILE_reg_out_17__4_, FP_REG_FILE_reg_out_17__3_,
         FP_REG_FILE_reg_out_17__2_, FP_REG_FILE_reg_out_17__1_,
         FP_REG_FILE_reg_out_17__0_, FP_REG_FILE_reg_out_16__10_,
         FP_REG_FILE_reg_out_16__9_, FP_REG_FILE_reg_out_16__8_,
         FP_REG_FILE_reg_out_16__7_, FP_REG_FILE_reg_out_16__6_,
         FP_REG_FILE_reg_out_16__5_, FP_REG_FILE_reg_out_16__4_,
         FP_REG_FILE_reg_out_16__3_, FP_REG_FILE_reg_out_16__2_,
         FP_REG_FILE_reg_out_16__1_, FP_REG_FILE_reg_out_16__0_,
         FP_REG_FILE_reg_out_15__31_, FP_REG_FILE_reg_out_15__30_,
         FP_REG_FILE_reg_out_15__29_, FP_REG_FILE_reg_out_15__28_,
         FP_REG_FILE_reg_out_15__27_, FP_REG_FILE_reg_out_15__26_,
         FP_REG_FILE_reg_out_15__25_, FP_REG_FILE_reg_out_15__24_,
         FP_REG_FILE_reg_out_15__23_, FP_REG_FILE_reg_out_15__22_,
         FP_REG_FILE_reg_out_15__21_, FP_REG_FILE_reg_out_15__20_,
         FP_REG_FILE_reg_out_15__19_, FP_REG_FILE_reg_out_15__18_,
         FP_REG_FILE_reg_out_15__17_, FP_REG_FILE_reg_out_15__16_,
         FP_REG_FILE_reg_out_15__15_, FP_REG_FILE_reg_out_15__14_,
         FP_REG_FILE_reg_out_15__13_, FP_REG_FILE_reg_out_15__12_,
         FP_REG_FILE_reg_out_15__11_, FP_REG_FILE_reg_out_15__10_,
         FP_REG_FILE_reg_out_15__9_, FP_REG_FILE_reg_out_15__8_,
         FP_REG_FILE_reg_out_15__7_, FP_REG_FILE_reg_out_15__6_,
         FP_REG_FILE_reg_out_15__5_, FP_REG_FILE_reg_out_15__4_,
         FP_REG_FILE_reg_out_15__3_, FP_REG_FILE_reg_out_15__2_,
         FP_REG_FILE_reg_out_15__1_, FP_REG_FILE_reg_out_15__0_,
         FP_REG_FILE_reg_out_14__31_, FP_REG_FILE_reg_out_14__30_,
         FP_REG_FILE_reg_out_14__29_, FP_REG_FILE_reg_out_14__28_,
         FP_REG_FILE_reg_out_14__27_, FP_REG_FILE_reg_out_14__26_,
         FP_REG_FILE_reg_out_14__25_, FP_REG_FILE_reg_out_14__24_,
         FP_REG_FILE_reg_out_14__23_, FP_REG_FILE_reg_out_14__22_,
         FP_REG_FILE_reg_out_14__21_, FP_REG_FILE_reg_out_14__20_,
         FP_REG_FILE_reg_out_14__19_, FP_REG_FILE_reg_out_14__18_,
         FP_REG_FILE_reg_out_14__17_, FP_REG_FILE_reg_out_14__16_,
         FP_REG_FILE_reg_out_14__15_, FP_REG_FILE_reg_out_14__14_,
         FP_REG_FILE_reg_out_14__13_, FP_REG_FILE_reg_out_14__12_,
         FP_REG_FILE_reg_out_14__11_, FP_REG_FILE_reg_out_14__10_,
         FP_REG_FILE_reg_out_14__9_, FP_REG_FILE_reg_out_14__8_,
         FP_REG_FILE_reg_out_14__7_, FP_REG_FILE_reg_out_14__6_,
         FP_REG_FILE_reg_out_14__5_, FP_REG_FILE_reg_out_14__4_,
         FP_REG_FILE_reg_out_14__3_, FP_REG_FILE_reg_out_14__2_,
         FP_REG_FILE_reg_out_14__1_, FP_REG_FILE_reg_out_14__0_,
         FP_REG_FILE_reg_out_13__31_, FP_REG_FILE_reg_out_13__30_,
         FP_REG_FILE_reg_out_13__29_, FP_REG_FILE_reg_out_13__28_,
         FP_REG_FILE_reg_out_13__27_, FP_REG_FILE_reg_out_13__26_,
         FP_REG_FILE_reg_out_13__25_, FP_REG_FILE_reg_out_13__24_,
         FP_REG_FILE_reg_out_13__23_, FP_REG_FILE_reg_out_13__22_,
         FP_REG_FILE_reg_out_13__21_, FP_REG_FILE_reg_out_13__20_,
         FP_REG_FILE_reg_out_13__19_, FP_REG_FILE_reg_out_13__18_,
         FP_REG_FILE_reg_out_13__17_, FP_REG_FILE_reg_out_13__16_,
         FP_REG_FILE_reg_out_13__15_, FP_REG_FILE_reg_out_13__14_,
         FP_REG_FILE_reg_out_13__13_, FP_REG_FILE_reg_out_13__12_,
         FP_REG_FILE_reg_out_13__11_, FP_REG_FILE_reg_out_13__10_,
         FP_REG_FILE_reg_out_13__9_, FP_REG_FILE_reg_out_13__8_,
         FP_REG_FILE_reg_out_13__7_, FP_REG_FILE_reg_out_13__6_,
         FP_REG_FILE_reg_out_13__5_, FP_REG_FILE_reg_out_13__4_,
         FP_REG_FILE_reg_out_13__3_, FP_REG_FILE_reg_out_13__2_,
         FP_REG_FILE_reg_out_13__1_, FP_REG_FILE_reg_out_13__0_,
         FP_REG_FILE_reg_out_12__31_, FP_REG_FILE_reg_out_12__30_,
         FP_REG_FILE_reg_out_12__29_, FP_REG_FILE_reg_out_12__28_,
         FP_REG_FILE_reg_out_12__27_, FP_REG_FILE_reg_out_12__26_,
         FP_REG_FILE_reg_out_12__25_, FP_REG_FILE_reg_out_12__24_,
         FP_REG_FILE_reg_out_12__23_, FP_REG_FILE_reg_out_12__22_,
         FP_REG_FILE_reg_out_12__21_, FP_REG_FILE_reg_out_12__20_,
         FP_REG_FILE_reg_out_12__19_, FP_REG_FILE_reg_out_12__18_,
         FP_REG_FILE_reg_out_12__17_, FP_REG_FILE_reg_out_12__16_,
         FP_REG_FILE_reg_out_12__15_, FP_REG_FILE_reg_out_12__14_,
         FP_REG_FILE_reg_out_12__13_, FP_REG_FILE_reg_out_12__12_,
         FP_REG_FILE_reg_out_12__11_, FP_REG_FILE_reg_out_12__10_,
         FP_REG_FILE_reg_out_12__9_, FP_REG_FILE_reg_out_12__8_,
         FP_REG_FILE_reg_out_12__7_, FP_REG_FILE_reg_out_12__6_,
         FP_REG_FILE_reg_out_12__5_, FP_REG_FILE_reg_out_12__4_,
         FP_REG_FILE_reg_out_12__3_, FP_REG_FILE_reg_out_12__2_,
         FP_REG_FILE_reg_out_12__1_, FP_REG_FILE_reg_out_12__0_,
         FP_REG_FILE_reg_out_11__31_, FP_REG_FILE_reg_out_11__30_,
         FP_REG_FILE_reg_out_11__29_, FP_REG_FILE_reg_out_11__28_,
         FP_REG_FILE_reg_out_11__27_, FP_REG_FILE_reg_out_11__26_,
         FP_REG_FILE_reg_out_11__25_, FP_REG_FILE_reg_out_11__24_,
         FP_REG_FILE_reg_out_11__23_, FP_REG_FILE_reg_out_11__22_,
         FP_REG_FILE_reg_out_11__21_, FP_REG_FILE_reg_out_11__20_,
         FP_REG_FILE_reg_out_11__19_, FP_REG_FILE_reg_out_11__18_,
         FP_REG_FILE_reg_out_11__17_, FP_REG_FILE_reg_out_11__16_,
         FP_REG_FILE_reg_out_11__15_, FP_REG_FILE_reg_out_11__14_,
         FP_REG_FILE_reg_out_11__13_, FP_REG_FILE_reg_out_11__12_,
         FP_REG_FILE_reg_out_11__11_, FP_REG_FILE_reg_out_11__10_,
         FP_REG_FILE_reg_out_11__9_, FP_REG_FILE_reg_out_11__8_,
         FP_REG_FILE_reg_out_11__7_, FP_REG_FILE_reg_out_11__6_,
         FP_REG_FILE_reg_out_11__5_, FP_REG_FILE_reg_out_11__4_,
         FP_REG_FILE_reg_out_11__3_, FP_REG_FILE_reg_out_11__2_,
         FP_REG_FILE_reg_out_11__1_, FP_REG_FILE_reg_out_11__0_,
         FP_REG_FILE_reg_out_10__31_, FP_REG_FILE_reg_out_10__30_,
         FP_REG_FILE_reg_out_10__29_, FP_REG_FILE_reg_out_10__28_,
         FP_REG_FILE_reg_out_10__27_, FP_REG_FILE_reg_out_10__26_,
         FP_REG_FILE_reg_out_10__25_, FP_REG_FILE_reg_out_10__24_,
         FP_REG_FILE_reg_out_10__23_, FP_REG_FILE_reg_out_10__22_,
         FP_REG_FILE_reg_out_10__21_, FP_REG_FILE_reg_out_10__20_,
         FP_REG_FILE_reg_out_10__19_, FP_REG_FILE_reg_out_10__18_,
         FP_REG_FILE_reg_out_10__17_, FP_REG_FILE_reg_out_10__16_,
         FP_REG_FILE_reg_out_10__15_, FP_REG_FILE_reg_out_10__14_,
         FP_REG_FILE_reg_out_10__13_, FP_REG_FILE_reg_out_10__12_,
         FP_REG_FILE_reg_out_10__11_, FP_REG_FILE_reg_out_10__10_,
         FP_REG_FILE_reg_out_10__9_, FP_REG_FILE_reg_out_10__8_,
         FP_REG_FILE_reg_out_10__7_, FP_REG_FILE_reg_out_10__6_,
         FP_REG_FILE_reg_out_10__5_, FP_REG_FILE_reg_out_10__4_,
         FP_REG_FILE_reg_out_10__3_, FP_REG_FILE_reg_out_10__2_,
         FP_REG_FILE_reg_out_10__1_, FP_REG_FILE_reg_out_10__0_,
         FP_REG_FILE_reg_out_9__31_, FP_REG_FILE_reg_out_9__30_,
         FP_REG_FILE_reg_out_9__29_, FP_REG_FILE_reg_out_9__28_,
         FP_REG_FILE_reg_out_9__27_, FP_REG_FILE_reg_out_9__26_,
         FP_REG_FILE_reg_out_9__25_, FP_REG_FILE_reg_out_9__24_,
         FP_REG_FILE_reg_out_9__23_, FP_REG_FILE_reg_out_9__22_,
         FP_REG_FILE_reg_out_9__21_, FP_REG_FILE_reg_out_9__20_,
         FP_REG_FILE_reg_out_9__19_, FP_REG_FILE_reg_out_9__18_,
         FP_REG_FILE_reg_out_9__17_, FP_REG_FILE_reg_out_9__16_,
         FP_REG_FILE_reg_out_9__15_, FP_REG_FILE_reg_out_9__14_,
         FP_REG_FILE_reg_out_9__13_, FP_REG_FILE_reg_out_9__12_,
         FP_REG_FILE_reg_out_9__11_, FP_REG_FILE_reg_out_9__10_,
         FP_REG_FILE_reg_out_9__9_, FP_REG_FILE_reg_out_9__8_,
         FP_REG_FILE_reg_out_9__7_, FP_REG_FILE_reg_out_9__6_,
         FP_REG_FILE_reg_out_9__5_, FP_REG_FILE_reg_out_9__4_,
         FP_REG_FILE_reg_out_9__3_, FP_REG_FILE_reg_out_9__2_,
         FP_REG_FILE_reg_out_9__1_, FP_REG_FILE_reg_out_9__0_,
         FP_REG_FILE_reg_out_5__31_, FP_REG_FILE_reg_out_5__30_,
         FP_REG_FILE_reg_out_5__29_, FP_REG_FILE_reg_out_5__28_,
         FP_REG_FILE_reg_out_5__27_, FP_REG_FILE_reg_out_5__26_,
         FP_REG_FILE_reg_out_5__25_, FP_REG_FILE_reg_out_5__24_,
         FP_REG_FILE_reg_out_5__23_, FP_REG_FILE_reg_out_5__22_,
         FP_REG_FILE_reg_out_5__21_, FP_REG_FILE_reg_out_5__20_,
         FP_REG_FILE_reg_out_5__19_, FP_REG_FILE_reg_out_5__18_,
         FP_REG_FILE_reg_out_5__17_, FP_REG_FILE_reg_out_5__16_,
         FP_REG_FILE_reg_out_5__15_, FP_REG_FILE_reg_out_5__14_,
         FP_REG_FILE_reg_out_5__13_, FP_REG_FILE_reg_out_5__12_,
         FP_REG_FILE_reg_out_5__11_, FP_REG_FILE_reg_out_5__10_,
         FP_REG_FILE_reg_out_5__9_, FP_REG_FILE_reg_out_5__8_,
         FP_REG_FILE_reg_out_5__7_, FP_REG_FILE_reg_out_5__6_,
         FP_REG_FILE_reg_out_5__5_, FP_REG_FILE_reg_out_5__4_,
         FP_REG_FILE_reg_out_5__3_, FP_REG_FILE_reg_out_5__2_,
         FP_REG_FILE_reg_out_5__1_, FP_REG_FILE_reg_out_5__0_,
         FP_REG_FILE_reg_out_4__31_, FP_REG_FILE_reg_out_4__30_,
         FP_REG_FILE_reg_out_4__29_, FP_REG_FILE_reg_out_4__28_,
         FP_REG_FILE_reg_out_4__27_, FP_REG_FILE_reg_out_4__26_,
         FP_REG_FILE_reg_out_4__25_, FP_REG_FILE_reg_out_4__24_,
         FP_REG_FILE_reg_out_4__23_, FP_REG_FILE_reg_out_4__22_,
         FP_REG_FILE_reg_out_4__21_, FP_REG_FILE_reg_out_4__20_,
         FP_REG_FILE_reg_out_4__19_, FP_REG_FILE_reg_out_4__18_,
         FP_REG_FILE_reg_out_4__17_, FP_REG_FILE_reg_out_4__16_,
         FP_REG_FILE_reg_out_4__15_, FP_REG_FILE_reg_out_4__14_,
         FP_REG_FILE_reg_out_4__13_, FP_REG_FILE_reg_out_4__12_,
         FP_REG_FILE_reg_out_4__11_, FP_REG_FILE_reg_out_4__10_,
         FP_REG_FILE_reg_out_4__9_, FP_REG_FILE_reg_out_4__8_,
         FP_REG_FILE_reg_out_4__7_, FP_REG_FILE_reg_out_4__6_,
         FP_REG_FILE_reg_out_4__5_, FP_REG_FILE_reg_out_4__4_,
         FP_REG_FILE_reg_out_4__3_, FP_REG_FILE_reg_out_4__2_,
         FP_REG_FILE_reg_out_4__1_, FP_REG_FILE_reg_out_4__0_,
         FP_REG_FILE_reg_out_3__31_, FP_REG_FILE_reg_out_3__30_,
         FP_REG_FILE_reg_out_3__29_, FP_REG_FILE_reg_out_3__28_,
         FP_REG_FILE_reg_out_3__27_, FP_REG_FILE_reg_out_3__26_,
         FP_REG_FILE_reg_out_3__25_, FP_REG_FILE_reg_out_3__24_,
         FP_REG_FILE_reg_out_3__23_, FP_REG_FILE_reg_out_3__22_,
         FP_REG_FILE_reg_out_3__21_, FP_REG_FILE_reg_out_3__20_,
         FP_REG_FILE_reg_out_3__19_, FP_REG_FILE_reg_out_3__18_,
         FP_REG_FILE_reg_out_3__17_, FP_REG_FILE_reg_out_3__16_,
         FP_REG_FILE_reg_out_3__15_, FP_REG_FILE_reg_out_3__14_,
         FP_REG_FILE_reg_out_3__13_, FP_REG_FILE_reg_out_3__12_,
         FP_REG_FILE_reg_out_3__11_, FP_REG_FILE_reg_out_3__10_,
         FP_REG_FILE_reg_out_3__9_, FP_REG_FILE_reg_out_3__8_,
         FP_REG_FILE_reg_out_3__7_, FP_REG_FILE_reg_out_3__6_,
         FP_REG_FILE_reg_out_3__5_, FP_REG_FILE_reg_out_3__4_,
         FP_REG_FILE_reg_out_3__3_, FP_REG_FILE_reg_out_3__2_,
         FP_REG_FILE_reg_out_3__1_, FP_REG_FILE_reg_out_3__0_,
         FP_REG_FILE_reg_out_2__31_, FP_REG_FILE_reg_out_2__30_,
         FP_REG_FILE_reg_out_2__29_, FP_REG_FILE_reg_out_2__28_,
         FP_REG_FILE_reg_out_2__27_, FP_REG_FILE_reg_out_2__26_,
         FP_REG_FILE_reg_out_2__25_, FP_REG_FILE_reg_out_2__24_,
         FP_REG_FILE_reg_out_2__23_, FP_REG_FILE_reg_out_2__22_,
         FP_REG_FILE_reg_out_2__21_, FP_REG_FILE_reg_out_2__20_,
         FP_REG_FILE_reg_out_2__19_, FP_REG_FILE_reg_out_2__18_,
         FP_REG_FILE_reg_out_2__17_, FP_REG_FILE_reg_out_2__16_,
         FP_REG_FILE_reg_out_2__15_, FP_REG_FILE_reg_out_2__14_,
         FP_REG_FILE_reg_out_2__13_, FP_REG_FILE_reg_out_2__12_,
         FP_REG_FILE_reg_out_2__11_, FP_REG_FILE_reg_out_2__10_,
         FP_REG_FILE_reg_out_2__9_, FP_REG_FILE_reg_out_2__8_,
         FP_REG_FILE_reg_out_2__7_, FP_REG_FILE_reg_out_2__6_,
         FP_REG_FILE_reg_out_2__5_, FP_REG_FILE_reg_out_2__4_,
         FP_REG_FILE_reg_out_2__3_, FP_REG_FILE_reg_out_2__2_,
         FP_REG_FILE_reg_out_2__1_, FP_REG_FILE_reg_out_2__0_,
         FP_REG_FILE_reg_out_1__31_, FP_REG_FILE_reg_out_1__30_,
         FP_REG_FILE_reg_out_1__29_, FP_REG_FILE_reg_out_1__28_,
         FP_REG_FILE_reg_out_1__27_, FP_REG_FILE_reg_out_1__26_,
         FP_REG_FILE_reg_out_1__25_, FP_REG_FILE_reg_out_1__24_,
         FP_REG_FILE_reg_out_1__23_, FP_REG_FILE_reg_out_1__22_,
         FP_REG_FILE_reg_out_1__21_, FP_REG_FILE_reg_out_1__20_,
         FP_REG_FILE_reg_out_1__19_, FP_REG_FILE_reg_out_1__18_,
         FP_REG_FILE_reg_out_1__17_, FP_REG_FILE_reg_out_1__16_,
         FP_REG_FILE_reg_out_1__15_, FP_REG_FILE_reg_out_1__14_,
         FP_REG_FILE_reg_out_1__13_, FP_REG_FILE_reg_out_1__12_,
         FP_REG_FILE_reg_out_1__11_, FP_REG_FILE_reg_out_1__10_,
         FP_REG_FILE_reg_out_1__9_, FP_REG_FILE_reg_out_1__8_,
         FP_REG_FILE_reg_out_1__7_, FP_REG_FILE_reg_out_1__6_,
         FP_REG_FILE_reg_out_1__5_, FP_REG_FILE_reg_out_1__4_,
         FP_REG_FILE_reg_out_1__3_, FP_REG_FILE_reg_out_1__2_,
         FP_REG_FILE_reg_out_1__1_, FP_REG_FILE_reg_out_1__0_,
         FP_REG_FILE_reg_out_0__31_, FP_REG_FILE_reg_out_0__30_,
         FP_REG_FILE_reg_out_0__29_, FP_REG_FILE_reg_out_0__28_,
         FP_REG_FILE_reg_out_0__27_, FP_REG_FILE_reg_out_0__26_,
         FP_REG_FILE_reg_out_0__25_, FP_REG_FILE_reg_out_0__24_,
         FP_REG_FILE_reg_out_0__23_, FP_REG_FILE_reg_out_0__22_,
         FP_REG_FILE_reg_out_0__21_, FP_REG_FILE_reg_out_0__20_,
         FP_REG_FILE_reg_out_0__19_, FP_REG_FILE_reg_out_0__18_,
         FP_REG_FILE_reg_out_0__17_, FP_REG_FILE_reg_out_0__16_,
         FP_REG_FILE_reg_out_0__15_, FP_REG_FILE_reg_out_0__14_,
         FP_REG_FILE_reg_out_0__13_, FP_REG_FILE_reg_out_0__12_,
         FP_REG_FILE_reg_out_0__11_, FP_REG_FILE_reg_out_0__10_,
         FP_REG_FILE_reg_out_0__9_, FP_REG_FILE_reg_out_0__8_,
         FP_REG_FILE_reg_out_0__7_, FP_REG_FILE_reg_out_0__6_,
         FP_REG_FILE_reg_out_0__5_, FP_REG_FILE_reg_out_0__4_,
         FP_REG_FILE_reg_out_0__3_, FP_REG_FILE_reg_out_0__2_,
         FP_REG_FILE_reg_out_0__1_, FP_REG_FILE_reg_out_0__0_,
         IF_STAGE_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         n27, n94, n95, n129, n164, n200, n201, n235, n272, n342, n376, n581,
         n616, n651, n685, n719, n787, n924, n959, n1028, n1135, n1236, n1238,
         n1240, n1242, n1244, n1248, n1250, n1252, n1254, n1256, n1258, n1260,
         n1262, n1264, n1266, n1270, n1271, n1290, n1291, n1292, n1293, n1294,
         n1295, n1298, n1301, n1306, n1307, n1308, n1313, n1316, n1317, n1320,
         n1338, n1345, n1348, n1351, n1358, n1433, n1434, n1435, n1436, n1437,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1487, n1719, n1746,
         n1790, n1830, n1831, n1832, n1833, n1834, n1837, n1842, n1858, n1859,
         n1860, n1861, n1866, n1871, n1875, n1880, n1881, n1882, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1895, n1896, n1897, n1898, n1901,
         n1902, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1915, n1916,
         n1917, n1918, n1921, n1922, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1935, n1936, n1937, n1938, n1941, n1942, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1956, n1957, n1958, n1959, n1962, n1963,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1976, n1977, n1978,
         n1979, n1982, n1983, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1996, n1997, n1998, n1999, n2002, n2003, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2016, n2017, n2018, n2019, n2022, n2023, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2036, n2037, n2038, n2039,
         n2042, n2043, n2046, n2048, n2049, n2050, n2051, n2056, n2057, n2058,
         n2059, n2062, n2063, n2066, n2068, n2069, n2070, n2071, n2076, n2077,
         n2078, n2079, n2082, n2083, n2086, n2088, n2089, n2090, n2091, n2096,
         n2097, n2098, n2099, n2102, n2103, n2106, n2108, n2109, n2110, n2111,
         n2116, n2117, n2118, n2119, n2122, n2123, n2126, n2128, n2129, n2130,
         n2131, n2136, n2137, n2138, n2139, n2142, n2143, n2147, n2149, n2150,
         n2151, n2152, n2157, n2158, n2159, n2160, n2163, n2164, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2177, n2178, n2179, n2180, n2182,
         n2184, n2185, n2188, n2189, n2193, n2194, n2195, n2196, n2198, n2201,
         n2202, n2204, n2206, n2211, n2212, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2231, n2232, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2251, n2252, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2271, n2272, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2291, n2292, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2311, n2312, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2331, n2332, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2351, n2352, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2372,
         n2373, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2392, n2393, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2412, n2413, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2432, n2433, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2452, n2453, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2472, n2473,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2492, n2493, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2506, n2508, n2509, n2511, n2513, n2514, n2515, n2517, n2522, n2524,
         n2527, n2528, n2530, n2531, n2532, n2533, n2536, n2538, n2539, n2555,
         n2557, n2559, n2562, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2577, n2584, n2598, n2602, n2603, n2608, n2619, n2626,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2641, n2644,
         n2650, n2651, n2652, n2655, n2659, n2662, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2675, n2678, n2684, n2685, n2686, n2689,
         n2693, n2696, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2709, n2712, n2718, n2719, n2720, n2723, n2727, n2730, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2743, n2746, n2752, n2753,
         n2754, n2757, n2761, n2764, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2777, n2780, n2786, n2787, n2788, n2791, n2795, n2798,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2811, n2814,
         n2820, n2821, n2822, n2825, n2829, n2832, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2845, n2848, n2854, n2855, n2856, n2859,
         n2863, n2866, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2880, n2883, n2889, n2890, n2891, n2894, n2898, n2901, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2914, n2917, n2923, n2924,
         n2925, n2928, n2932, n2935, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2948, n2951, n2957, n2958, n2959, n2962, n2966, n2969,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2982, n2985,
         n2991, n2992, n2993, n2996, n3000, n3003, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3016, n3019, n3025, n3026, n3027, n3030,
         n3034, n3037, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3050, n3053, n3059, n3060, n3061, n3064, n3068, n3071, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3084, n3087, n3093, n3094,
         n3095, n3098, n3102, n3105, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3118, n3121, n3127, n3128, n3129, n3132, n3136, n3139,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3152, n3155,
         n3161, n3162, n3163, n3166, n3170, n3173, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3186, n3189, n3195, n3196, n3197, n3200,
         n3204, n3207, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3221, n3224, n3230, n3231, n3232, n3235, n3239, n3242, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3255, n3258, n3264,
         n3265, n3266, n3269, n3273, n3276, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3289, n3292, n3298, n3299, n3300, n3303, n3307,
         n3310, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3323,
         n3326, n3332, n3333, n3334, n3337, n3341, n3344, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3357, n3360, n3366, n3367, n3368,
         n3371, n3375, n3378, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3391, n3394, n3400, n3401, n3402, n3405, n3409, n3412, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3425, n3428, n3434,
         n3435, n3436, n3439, n3443, n3446, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3459, n3462, n3468, n3469, n3470, n3473, n3477,
         n3480, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3493,
         n3496, n3502, n3503, n3504, n3507, n3511, n3514, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3527, n3530, n3536, n3537, n3538,
         n3541, n3545, n3548, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3562, n3565, n3571, n3572, n3573, n3576, n3580, n3583, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3596, n3599, n3605,
         n3606, n3607, n3610, n3614, n3617, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3630, n3633, n3639, n3640, n3641, n3644, n3648,
         n3651, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3664,
         n3674, n3684, n3685, n3686, n3689, n3695, n3699, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3714, n3720, n3738, n3739, n3743,
         n3750, n3755, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3775, n3782, n3783, n3785, n3788, n3789, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3804, n3811, n3812, n3814,
         n3817, n3818, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3833, n3840, n3841, n3843, n3846, n3847, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3862, n3869, n3870, n3872,
         n3875, n3876, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3891, n3898, n3899, n3901, n3904, n3905, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3921, n3928, n3929, n3931,
         n3934, n3935, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3950, n3957, n3958, n3960, n3963, n3964, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3979, n3986, n3987, n3989,
         n3992, n3993, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4008, n4015, n4016, n4018, n4021, n4022, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4037, n4044, n4045, n4047,
         n4050, n4051, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4066, n4073, n4074, n4076, n4079, n4080, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4095, n4102, n4103, n4105,
         n4108, n4109, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4124, n4131, n4132, n4134, n4137, n4138, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4153, n4160, n4161, n4163,
         n4166, n4167, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4182, n4189, n4190, n4192, n4195, n4196, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4212, n4219, n4220, n4222,
         n4225, n4226, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4241, n4248, n4249, n4251, n4254, n4255, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4270, n4277, n4278, n4280,
         n4283, n4284, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4299, n4306, n4307, n4309, n4312, n4313, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4328, n4335, n4336, n4338,
         n4341, n4342, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4357, n4364, n4365, n4367, n4370, n4371, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4386, n4393, n4394, n4396,
         n4399, n4400, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4415, n4422, n4423, n4425, n4428, n4429, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4444, n4451, n4452, n4454,
         n4457, n4458, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4473, n4480, n4481, n4483, n4486, n4487, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4503, n4510, n4511, n4513,
         n4516, n4517, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4532, n4539, n4540, n4542, n4545, n4546, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4561, n4568, n4569, n4571,
         n4574, n4575, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4590, n4597, n4598, n4600, n4603, n4604, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4619, n4626, n4627, n4629,
         n4632, n4633, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4650, n4659, n4660, n4662, n4665, n4666, n4674, n4685, n5463,
         n5464, n5466, n5467, n5478, n5482, n5484, n5499, n5506, n5513, n5516,
         n5518, n5520, n5529, n5535, n5546, n5549, n5555, n5558, n5586, n5588,
         n5590, n5595, n5597, n5603, n5606, n5608, n5612, n5614, n5630, n5662,
         n5663, n5664, n5667, n5668, n5669, n5670, n5673, n5675, n5676, n5679,
         n5680, n5684, n5717, n5718, n5721, n5723, n5724, n5727, n5729, n5732,
         n5764, n5767, n5769, n5770, n5773, n5774, n5776, n5777, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5815, n5816, n5818, n5851, n5853, n5886, n5888,
         n5890, n5891, n5893, n5895, n5897, n5899, n5901, n5903, n5905, n5907,
         n5909, n5910, n6625, n6741, n6744, n6746, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6756, n6757, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6889, n6890, n6891, n6892, n6893, n7279, n7280, n7283,
         n7284, n7286, n7288, n7289, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7519, n7520, n7521, n7522, n7523,
         n7526, n7527, n7528, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7582, n7583, n7584, n7586, n7587, n7588, n7589, n7590,
         n7592, n7593, n7594, n7595, n7596, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7622, n7623, n7624, n7626,
         n7627, n7628, n7629, n7630, n7632, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7904, n7905, n7906, n7909, n7910,
         n7911, n7912, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7980, n7981, n7982, n7983, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7999,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8020, n10104,
         n10105, n10106, EXEC_STAGE_mul_ex_N153, EXEC_STAGE_mul_ex_N152,
         EXEC_STAGE_mul_ex_N151, EXEC_STAGE_mul_ex_N150,
         EXEC_STAGE_mul_ex_N149, EXEC_STAGE_mul_ex_N148,
         EXEC_STAGE_mul_ex_N147, EXEC_STAGE_mul_ex_N146,
         EXEC_STAGE_mul_ex_N145, EXEC_STAGE_mul_ex_N144,
         EXEC_STAGE_mul_ex_N143, EXEC_STAGE_mul_ex_N142,
         EXEC_STAGE_mul_ex_N141, EXEC_STAGE_mul_ex_N140,
         EXEC_STAGE_mul_ex_N139, EXEC_STAGE_mul_ex_N138,
         EXEC_STAGE_mul_ex_N137, EXEC_STAGE_mul_ex_N136,
         EXEC_STAGE_mul_ex_N135, EXEC_STAGE_mul_ex_N134,
         EXEC_STAGE_mul_ex_N133, EXEC_STAGE_mul_ex_N132,
         EXEC_STAGE_mul_ex_N131, EXEC_STAGE_mul_ex_N130,
         EXEC_STAGE_mul_ex_N129, EXEC_STAGE_mul_ex_N128,
         EXEC_STAGE_mul_ex_N127, EXEC_STAGE_mul_ex_N126,
         EXEC_STAGE_mul_ex_N125, EXEC_STAGE_mul_ex_N124,
         EXEC_STAGE_mul_ex_N123, EXEC_STAGE_mul_ex_N122,
         EXEC_STAGE_mul_ex_N121, EXEC_STAGE_mul_ex_N120,
         EXEC_STAGE_mul_ex_N217, EXEC_STAGE_mul_ex_N216,
         EXEC_STAGE_mul_ex_N215, EXEC_STAGE_mul_ex_N214,
         EXEC_STAGE_mul_ex_N213, EXEC_STAGE_mul_ex_N212,
         EXEC_STAGE_mul_ex_N211, EXEC_STAGE_mul_ex_N210,
         EXEC_STAGE_mul_ex_N209, EXEC_STAGE_mul_ex_N208,
         EXEC_STAGE_mul_ex_N207, EXEC_STAGE_mul_ex_N206,
         EXEC_STAGE_mul_ex_N205, EXEC_STAGE_mul_ex_N204,
         EXEC_STAGE_mul_ex_N203, EXEC_STAGE_mul_ex_N202,
         EXEC_STAGE_mul_ex_N201, EXEC_STAGE_mul_ex_N200,
         EXEC_STAGE_mul_ex_N199, EXEC_STAGE_mul_ex_N198,
         EXEC_STAGE_mul_ex_N197, EXEC_STAGE_mul_ex_N196,
         EXEC_STAGE_mul_ex_N195, EXEC_STAGE_mul_ex_N194,
         EXEC_STAGE_mul_ex_N193, EXEC_STAGE_mul_ex_N192,
         EXEC_STAGE_mul_ex_N191, EXEC_STAGE_mul_ex_N190,
         EXEC_STAGE_mul_ex_N189, EXEC_STAGE_mul_ex_N188,
         EXEC_STAGE_mul_ex_N187, EXEC_STAGE_mul_ex_N186,
         EXEC_STAGE_mul_ex_N298, EXEC_STAGE_mul_ex_N297,
         EXEC_STAGE_mul_ex_N296, EXEC_STAGE_mul_ex_N295,
         EXEC_STAGE_mul_ex_N294, EXEC_STAGE_mul_ex_N293,
         EXEC_STAGE_mul_ex_N292, EXEC_STAGE_mul_ex_N291,
         EXEC_STAGE_mul_ex_N290, EXEC_STAGE_mul_ex_N289,
         EXEC_STAGE_mul_ex_N288, EXEC_STAGE_mul_ex_N287,
         EXEC_STAGE_mul_ex_N286, EXEC_STAGE_mul_ex_N285,
         EXEC_STAGE_mul_ex_N284, EXEC_STAGE_mul_ex_N283,
         EXEC_STAGE_mul_ex_N282, EXEC_STAGE_mul_ex_N281,
         EXEC_STAGE_mul_ex_N280, EXEC_STAGE_mul_ex_N279,
         EXEC_STAGE_mul_ex_N278, EXEC_STAGE_mul_ex_N277,
         EXEC_STAGE_mul_ex_N276, EXEC_STAGE_mul_ex_N275,
         EXEC_STAGE_mul_ex_N274, EXEC_STAGE_mul_ex_N273,
         EXEC_STAGE_mul_ex_N272, EXEC_STAGE_mul_ex_N271,
         EXEC_STAGE_mul_ex_N270, EXEC_STAGE_mul_ex_N269,
         EXEC_STAGE_mul_ex_N268, EXEC_STAGE_mul_ex_N267,
         EXEC_STAGE_mul_ex_N266, EXEC_STAGE_mul_ex_N265,
         EXEC_STAGE_mul_ex_N264, EXEC_STAGE_mul_ex_N263,
         EXEC_STAGE_mul_ex_N262, EXEC_STAGE_mul_ex_N261,
         EXEC_STAGE_mul_ex_N260, EXEC_STAGE_mul_ex_N259,
         EXEC_STAGE_mul_ex_N258, EXEC_STAGE_mul_ex_N257,
         EXEC_STAGE_mul_ex_N256, EXEC_STAGE_mul_ex_N255,
         EXEC_STAGE_mul_ex_N254, EXEC_STAGE_mul_ex_N253,
         EXEC_STAGE_mul_ex_N252, EXEC_STAGE_mul_ex_N251,
         EXEC_STAGE_mul_ex_N250, net137185, net137303, net137317, net137343,
         net137549, net137550, net137569, net139967, net222300, net222304,
         net222353, net222497, net222531, net222628, net222629, net222642,
         net222698, net222980, net222982, net223077, net223078, net223079,
         net223104, net223109, net223324, net223365, net223368, net223439,
         net223440, net223586, net223589, net223591, net223662, net223664,
         net223665, net223666, net223740, net223741, net223742, net223743,
         net223794, net223796, net223797, net223985, net224151, net224170,
         net224171, net224173, net224174, net224180, net224182, net224402,
         net224492, net224493, net224658, net224699, net224704, net224707,
         net224710, net224711, net224713, net224816, net224837, net224838,
         net224839, net224840, net224844, net224845, net224846, net224848,
         net224850, net224853, net224952, net224953, net225075, net225076,
         net225077, net225160, net225162, net225163, net225172, net225183,
         net225184, net225185, net225186, net225187, net225188, net225191,
         net225192, net225194, net225195, net225196, net225198, net225212,
         net225214, net225448, net225449, net225526, net225527, net225529,
         net225681, net225777, net225780, net225821, net225823, net225889,
         net225890, net225892, net225894, net225906, net225908, net226995,
         net227002, net227008, net227014, net227015, net227019, net227020,
         net227024, net227026, net227035, net227040, net227041, net227042,
         net227043, net227045, net227046, net227047, net227052, net227058,
         net227062, net227067, net227070, net227071, net227073, net227077,
         net227081, net227084, net227094, net227095, net227106, net227108,
         net227110, net227115, net227116, net227117, net227121, net227122,
         net227135, net227137, net227142, net227143, net227148, net227149,
         net227150, net227159, net227160, net227163, net227164, net227165,
         net227166, net227167, net227169, net227170, net227174, net227175,
         net227176, net227177, net227180, net227182, net227183, net227186,
         net227187, net227188, net227189, net227190, net227192, net227197,
         net227198, net227202, net227213, net227214, net227216, net227217,
         net227219, net227224, net227225, net227226, net227232, net227233,
         net227236, net227239, net227240, net227241, net227242, net227243,
         net227245, net227246, net227247, net227248, net227256, net227265,
         net227269, net227276, net227277, net227282, net230393, net230387,
         net230383, net230381, net230379, net230377, net230373, net231353,
         net231349, net231345, net231341, net231339, net231337, net231335,
         net231333, net231331, net231325, net231323, net231321, net231319,
         net231317, net231315, net231313, net231311, net231309, net231307,
         net231305, net231303, net231301, net231297, net231295, net231293,
         net231291, net231289, net231283, net231279, net231277, net231275,
         net231273, net231271, net231263, net231261, net231259, net231257,
         net231255, net231253, net231251, net231249, net231247, net231245,
         net231243, net231241, net231239, net231237, net231235, net231233,
         net231231, net231229, net231227, net231225, net231223, net231221,
         net231217, net231211, net231357, net231615, net231915, net232817,
         net232816, net232877, net232881, net233102, net233124, net233133,
         net233142, net233156, net233181, net233216, net233233, net233242,
         net239032, net239031, net239030, net239035, net239082, net239083,
         net239150, net239221, net239220, net239254, net239329, net239344,
         net239371, net239370, net239374, net239379, net239390, net239415,
         net239414, net239424, net239454, net239459, net239473, net239475,
         net239496, net239507, net239508, net239528, net239527, net239555,
         net239554, net239553, net239557, net239572, net239598, net239597,
         net239621, net239628, net239627, net239631, net239630, net239667,
         net239669, net239674, net239673, net239678, net239718, net239737,
         net239744, net239756, net239767, net239774, net239776, net239782,
         net239805, net239806, net239816, net239815, net239823, net239825,
         net239828, net239846, net227201, net227158, net227153, net227119,
         net224491, net224404, net227065, net227064, net227053, net227048,
         net225210, net225209, net239356, net227231, net227230, net227229,
         net227157, net227156, net227075, net239404, net233131, net227145,
         net227144, net227136, net224403, net227044, net239761, net239722,
         net227207, net225201, net239533, net227191, net239017, net227072,
         net227068, net227063, net225893, net225824, net227128, net227098,
         net225453, net225452, net239380, net233078, net227033, net227013,
         net227012, net227010, net227009, net224847, net224843, net224842,
         net224841, net231361, net231359, net231355, net231329, net230403,
         net230399, net225206, net225203, net225202, net139963, net227271,
         net227270, net227254, net223444, net227086, net227079, net225684,
         net225528, net233106, net225207, net225204, net224709, net224708,
         net239477, net227275, net227274, net227262, net227261, net227259,
         net227199, net223442, net223366, net227208, net227205, net227204,
         net224181, net227107, net227102, net227101, net227093, net225450,
         net227139, net227105, net227104, net227103, net224955, net224954,
         net224661, net224660, net233241, net227290, net227090, net227089,
         net227088, net227087, net227069, net225778, net239616, net233180,
         net233141, net227255, net227221, net227220, net227200, net223663,
         net223447, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12037, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12982, n12983, n12984, n12985, n12987, n12988, n12989, n12990,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13108, n13109, n13110, n13111, n13112, n13113, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         EXEC_STAGE_mul_ex_add_88_n2, EXEC_STAGE_mul_ex_add_88_2_n2,
         EXEC_STAGE_mul_ex_mult_88_n100, EXEC_STAGE_mul_ex_mult_88_n99,
         EXEC_STAGE_mul_ex_mult_88_n98, EXEC_STAGE_mul_ex_mult_88_n97,
         EXEC_STAGE_mul_ex_mult_88_n96, EXEC_STAGE_mul_ex_mult_88_n95,
         EXEC_STAGE_mul_ex_mult_88_n94, EXEC_STAGE_mul_ex_mult_88_n93,
         EXEC_STAGE_mul_ex_mult_88_n92, EXEC_STAGE_mul_ex_mult_88_n91,
         EXEC_STAGE_mul_ex_mult_88_n90, EXEC_STAGE_mul_ex_mult_88_n89,
         EXEC_STAGE_mul_ex_mult_88_n88, EXEC_STAGE_mul_ex_mult_88_n87,
         EXEC_STAGE_mul_ex_mult_88_n86, EXEC_STAGE_mul_ex_mult_88_n85,
         EXEC_STAGE_mul_ex_mult_88_n84, EXEC_STAGE_mul_ex_mult_88_n83,
         EXEC_STAGE_mul_ex_mult_88_n82, EXEC_STAGE_mul_ex_mult_88_n81,
         EXEC_STAGE_mul_ex_mult_88_n80, EXEC_STAGE_mul_ex_mult_88_n79,
         EXEC_STAGE_mul_ex_mult_88_n78, EXEC_STAGE_mul_ex_mult_88_n77,
         EXEC_STAGE_mul_ex_mult_88_n76, EXEC_STAGE_mul_ex_mult_88_n75,
         EXEC_STAGE_mul_ex_mult_88_n74, EXEC_STAGE_mul_ex_mult_88_n73,
         EXEC_STAGE_mul_ex_mult_88_n72, EXEC_STAGE_mul_ex_mult_88_n71,
         EXEC_STAGE_mul_ex_mult_88_n70, EXEC_STAGE_mul_ex_mult_88_n69,
         EXEC_STAGE_mul_ex_mult_88_n68, EXEC_STAGE_mul_ex_mult_88_n67,
         EXEC_STAGE_mul_ex_mult_88_n66, EXEC_STAGE_mul_ex_mult_88_n65,
         EXEC_STAGE_mul_ex_mult_88_n63, EXEC_STAGE_mul_ex_mult_88_n62,
         EXEC_STAGE_mul_ex_mult_88_n61, EXEC_STAGE_mul_ex_mult_88_n60,
         EXEC_STAGE_mul_ex_mult_88_n59, EXEC_STAGE_mul_ex_mult_88_n58,
         EXEC_STAGE_mul_ex_mult_88_n57, EXEC_STAGE_mul_ex_mult_88_n56,
         EXEC_STAGE_mul_ex_mult_88_n55, EXEC_STAGE_mul_ex_mult_88_n54,
         EXEC_STAGE_mul_ex_mult_88_n53, EXEC_STAGE_mul_ex_mult_88_n52,
         EXEC_STAGE_mul_ex_mult_88_n51, EXEC_STAGE_mul_ex_mult_88_n50,
         EXEC_STAGE_mul_ex_mult_88_n49, EXEC_STAGE_mul_ex_mult_88_n48,
         EXEC_STAGE_mul_ex_mult_88_n47, EXEC_STAGE_mul_ex_mult_88_n46,
         EXEC_STAGE_mul_ex_mult_88_n45, EXEC_STAGE_mul_ex_mult_88_n44,
         EXEC_STAGE_mul_ex_mult_88_n43, EXEC_STAGE_mul_ex_mult_88_n42,
         EXEC_STAGE_mul_ex_mult_88_n41, EXEC_STAGE_mul_ex_mult_88_n40,
         EXEC_STAGE_mul_ex_mult_88_n39, EXEC_STAGE_mul_ex_mult_88_n38,
         EXEC_STAGE_mul_ex_mult_88_n37, EXEC_STAGE_mul_ex_mult_88_n36,
         EXEC_STAGE_mul_ex_mult_88_n35, EXEC_STAGE_mul_ex_mult_88_n34,
         EXEC_STAGE_mul_ex_mult_88_n33, EXEC_STAGE_mul_ex_mult_88_n32,
         EXEC_STAGE_mul_ex_mult_88_n31, EXEC_STAGE_mul_ex_mult_88_n30,
         EXEC_STAGE_mul_ex_mult_88_n29, EXEC_STAGE_mul_ex_mult_88_n28,
         EXEC_STAGE_mul_ex_mult_88_n27, EXEC_STAGE_mul_ex_mult_88_n26,
         EXEC_STAGE_mul_ex_mult_88_n25, EXEC_STAGE_mul_ex_mult_88_n24,
         EXEC_STAGE_mul_ex_mult_88_n23, EXEC_STAGE_mul_ex_mult_88_n22,
         EXEC_STAGE_mul_ex_mult_88_n21, EXEC_STAGE_mul_ex_mult_88_n20,
         EXEC_STAGE_mul_ex_mult_88_n19, EXEC_STAGE_mul_ex_mult_88_n18,
         EXEC_STAGE_mul_ex_mult_88_n17, EXEC_STAGE_mul_ex_mult_88_n16,
         EXEC_STAGE_mul_ex_mult_88_n15, EXEC_STAGE_mul_ex_mult_88_n14,
         EXEC_STAGE_mul_ex_mult_88_n13, EXEC_STAGE_mul_ex_mult_88_n12,
         EXEC_STAGE_mul_ex_mult_88_n11, EXEC_STAGE_mul_ex_mult_88_n10,
         EXEC_STAGE_mul_ex_mult_88_n9, EXEC_STAGE_mul_ex_mult_88_n8,
         EXEC_STAGE_mul_ex_mult_88_n7, EXEC_STAGE_mul_ex_mult_88_n6,
         EXEC_STAGE_mul_ex_mult_88_n5, EXEC_STAGE_mul_ex_mult_88_n4,
         EXEC_STAGE_mul_ex_mult_88_n3, EXEC_STAGE_mul_ex_mult_88_A1_0_,
         EXEC_STAGE_mul_ex_mult_88_A1_1_, EXEC_STAGE_mul_ex_mult_88_A1_2_,
         EXEC_STAGE_mul_ex_mult_88_A1_3_, EXEC_STAGE_mul_ex_mult_88_A1_4_,
         EXEC_STAGE_mul_ex_mult_88_A1_5_, EXEC_STAGE_mul_ex_mult_88_A1_6_,
         EXEC_STAGE_mul_ex_mult_88_A1_7_, EXEC_STAGE_mul_ex_mult_88_A1_8_,
         EXEC_STAGE_mul_ex_mult_88_A1_9_, EXEC_STAGE_mul_ex_mult_88_A1_10_,
         EXEC_STAGE_mul_ex_mult_88_A1_11_, EXEC_STAGE_mul_ex_mult_88_A1_12_,
         EXEC_STAGE_mul_ex_mult_88_A1_13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_2__1_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_2__2_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_2__3_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_2__4_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_2__5_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_2__6_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_2__7_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_2__8_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_2__9_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_2__10_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_2__11_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_2__12_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_2__13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_2__14_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_2__15_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_3__1_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_3__2_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_3__3_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_3__4_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_3__5_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_3__6_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_3__7_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_3__8_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_3__9_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_3__10_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_3__11_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_3__12_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_3__13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_3__14_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_3__15_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_4__1_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_4__2_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_4__3_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_4__4_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_4__5_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_4__6_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_4__7_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_4__8_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_4__9_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_4__10_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_4__11_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_4__12_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_4__13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_4__14_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_4__15_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_5__1_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_5__2_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_5__3_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_5__4_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_5__5_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_5__6_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_5__7_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_5__8_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_5__9_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_5__10_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_5__11_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_5__12_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_5__13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_5__14_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_5__15_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_6__1_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_6__2_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_6__3_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_6__4_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_6__5_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_6__6_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_6__7_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_6__8_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_6__9_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_6__10_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_6__11_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_6__12_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_6__13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_6__14_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_6__15_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_7__1_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_7__2_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_7__3_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_7__4_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_7__5_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_7__6_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_7__7_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_7__8_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_7__9_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_7__10_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_7__11_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_7__12_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_7__13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_7__14_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_7__15_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_8__1_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_8__2_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_8__3_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_8__4_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_8__5_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_8__6_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_8__7_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_8__8_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_8__9_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_8__10_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_8__11_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_8__12_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_8__13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_8__14_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_8__15_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_9__1_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_9__2_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_9__3_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_9__4_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_9__5_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_9__6_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_9__7_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_9__8_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_9__9_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_9__10_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_9__11_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_9__12_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_9__13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_9__14_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_9__15_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_10__1_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_10__2_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_10__3_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_10__4_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_10__5_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_10__6_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_10__7_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_10__8_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_10__9_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_10__10_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_10__11_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_10__12_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_10__13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_10__14_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_10__15_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_11__1_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_11__2_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_11__3_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_11__4_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_11__5_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_11__6_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_11__7_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_11__8_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_11__9_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_11__10_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_11__11_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_11__12_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_11__13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_11__14_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_11__15_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_12__1_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_12__2_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_12__3_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_12__4_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_12__5_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_12__6_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_12__7_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_12__8_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_12__9_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_12__10_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_12__11_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_12__12_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_12__13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_12__14_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_12__15_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_13__1_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_13__2_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_13__3_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_13__4_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_13__5_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_13__6_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_13__7_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_13__8_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_13__9_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_13__10_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_13__11_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_13__12_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_13__13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_13__14_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_13__15_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_14__1_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_14__2_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_14__3_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_14__4_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_14__5_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_14__6_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_14__7_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_14__8_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_14__9_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_14__10_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_14__11_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_14__12_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_14__13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_14__14_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_14__15_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_15__1_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_15__2_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_15__3_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_15__4_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_15__5_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_15__6_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_15__7_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_15__8_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_15__9_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_15__10_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_15__11_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_15__12_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_15__13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_15__14_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_15__15_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__0_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__1_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__2_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__3_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__4_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__5_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__6_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__7_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__8_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__9_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__10_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__11_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__12_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__13_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__14_,
         EXEC_STAGE_mul_ex_mult_88_SUMB_16__15_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__0_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__1_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__2_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__3_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__4_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__5_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__6_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__7_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__8_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__9_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__10_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__11_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__12_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__13_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__14_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_2__15_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__0_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__1_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__2_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__3_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__4_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__5_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__6_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__7_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__8_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__9_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__10_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__11_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__12_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__13_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__14_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_3__15_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__0_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__1_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__2_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__3_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__4_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__5_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__6_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__7_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__8_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__9_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__10_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__11_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__12_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__13_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__14_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_4__15_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__0_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__1_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__2_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__3_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__4_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__5_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__6_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__7_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__8_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__9_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__10_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__11_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__12_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__13_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__14_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_5__15_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__0_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__1_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__2_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__3_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__4_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__5_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__6_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__7_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__8_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__9_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__10_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__11_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__12_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__13_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__14_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_6__15_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__0_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__1_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__2_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__3_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__4_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__5_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__6_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__7_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__8_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__9_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__10_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__11_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__12_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__13_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__14_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_7__15_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__0_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__1_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__2_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__3_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__4_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__5_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__6_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__7_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__8_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__9_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__10_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__11_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__12_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__13_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__14_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_8__15_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__0_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__1_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__2_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__3_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__4_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__5_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__6_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__7_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__8_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__9_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__10_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__11_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__12_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__13_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__14_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_9__15_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__0_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__1_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__2_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__3_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__4_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__5_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__6_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__7_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__8_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__9_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__10_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__11_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__12_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__13_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__14_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_10__15_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__0_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__1_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__2_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__3_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__4_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__5_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__6_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__7_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__8_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__9_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__10_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__11_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__12_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__13_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__14_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_11__15_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__0_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__1_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__2_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__3_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__4_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__5_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__6_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__7_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__8_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__9_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__10_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__11_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__12_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__13_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__14_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_12__15_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__0_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__1_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__2_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__3_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__4_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__5_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__6_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__7_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__8_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__9_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__10_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__11_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__12_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__13_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__14_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_13__15_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__0_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__1_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__2_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__3_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__4_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__5_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__6_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__7_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__8_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__9_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__10_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__11_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__12_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__13_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__14_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_14__15_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__0_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__1_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__2_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__3_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__4_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__5_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__6_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__7_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__8_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__9_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__10_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__11_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__12_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__13_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__14_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_15__15_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__0_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__1_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__2_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__3_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__4_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__5_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__6_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__7_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__8_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__9_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__10_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__11_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__12_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__13_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__14_,
         EXEC_STAGE_mul_ex_mult_88_CARRYB_16__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_0__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_1__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_2__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_3__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_4__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_5__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_6__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_7__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_8__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_9__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_10__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_11__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_12__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_13__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_14__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_15__16_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__0_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__1_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__2_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__3_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__4_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__5_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__6_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__7_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__8_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__9_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__10_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__11_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__12_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__13_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__14_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__15_,
         EXEC_STAGE_mul_ex_mult_88_ab_16__16_,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n65,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n64,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n63,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n62,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n61,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n60,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n59,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n58,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n57,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n56,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n55,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n54,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n53,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n52,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n51,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n50,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n49,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n48,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n47,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n46,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n45,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n44,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n43,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n42,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n41,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n40,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n39,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n38,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n37,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n36,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n35,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n34,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n33,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n32,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n31,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n30,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n29,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n28,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n27,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n26,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n25,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n24,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n23,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n22,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n21,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n20,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n19,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n18,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n17,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n16,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n15,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n14,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n13,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n12,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n11,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n10, EXEC_STAGE_mul_ex_mult_88_FS_1_n9,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n8, EXEC_STAGE_mul_ex_mult_88_FS_1_n7,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n6, EXEC_STAGE_mul_ex_mult_88_FS_1_n5,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n4, EXEC_STAGE_mul_ex_mult_88_FS_1_n3,
         EXEC_STAGE_mul_ex_mult_88_FS_1_n1,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n33,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n32,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n31,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n30,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n29,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n28,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n27,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n26,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n25,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n24,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n23,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n22,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n21,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n20,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n19,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n18,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n17,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n16,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n15,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n14,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n13,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n12,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n11,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n10,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n9,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n8,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n7,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n6,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n5,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n4,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n3,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n2,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n1,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n33,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n32,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n31,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n30,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n29,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n28,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n27,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n26,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n25,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n24,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n23,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n22,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n21,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n20,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n19,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n18,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n17,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n16,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n15,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n14,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n13,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n12,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n11,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n10,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n9,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n8,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n7,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n6,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n5,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n4,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n3,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n2,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n1,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n33,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n17,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n16,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n15,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n14,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n13,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n12,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n11,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n10,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n8,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n7,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n6,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n5,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n4,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n3,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n2,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_18_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_19_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_20_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_21_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_22_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_23_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_24_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_25_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_26_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_27_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_28_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_29_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_30_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_31_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_32_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n25,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n24,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n23,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n22,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n21,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n20,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n19,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n18,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n17,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n6,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n5,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n4,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n3,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n2,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n1,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_34_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_35_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_36_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_37_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_38_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_39_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_40_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_41_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_42_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_43_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_44_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_45_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_46_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_47_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_48_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_49_,
         EXEC_STAGE_mul_ex_mult_84_n94, EXEC_STAGE_mul_ex_mult_84_n93,
         EXEC_STAGE_mul_ex_mult_84_n92, EXEC_STAGE_mul_ex_mult_84_n91,
         EXEC_STAGE_mul_ex_mult_84_n90, EXEC_STAGE_mul_ex_mult_84_n89,
         EXEC_STAGE_mul_ex_mult_84_n88, EXEC_STAGE_mul_ex_mult_84_n87,
         EXEC_STAGE_mul_ex_mult_84_n86, EXEC_STAGE_mul_ex_mult_84_n85,
         EXEC_STAGE_mul_ex_mult_84_n84, EXEC_STAGE_mul_ex_mult_84_n83,
         EXEC_STAGE_mul_ex_mult_84_n82, EXEC_STAGE_mul_ex_mult_84_n81,
         EXEC_STAGE_mul_ex_mult_84_n80, EXEC_STAGE_mul_ex_mult_84_n79,
         EXEC_STAGE_mul_ex_mult_84_n78, EXEC_STAGE_mul_ex_mult_84_n77,
         EXEC_STAGE_mul_ex_mult_84_n76, EXEC_STAGE_mul_ex_mult_84_n75,
         EXEC_STAGE_mul_ex_mult_84_n74, EXEC_STAGE_mul_ex_mult_84_n73,
         EXEC_STAGE_mul_ex_mult_84_n72, EXEC_STAGE_mul_ex_mult_84_n71,
         EXEC_STAGE_mul_ex_mult_84_n70, EXEC_STAGE_mul_ex_mult_84_n69,
         EXEC_STAGE_mul_ex_mult_84_n68, EXEC_STAGE_mul_ex_mult_84_n67,
         EXEC_STAGE_mul_ex_mult_84_n66, EXEC_STAGE_mul_ex_mult_84_n65,
         EXEC_STAGE_mul_ex_mult_84_n64, EXEC_STAGE_mul_ex_mult_84_n63,
         EXEC_STAGE_mul_ex_mult_84_n62, EXEC_STAGE_mul_ex_mult_84_n61,
         EXEC_STAGE_mul_ex_mult_84_n59, EXEC_STAGE_mul_ex_mult_84_n58,
         EXEC_STAGE_mul_ex_mult_84_n57, EXEC_STAGE_mul_ex_mult_84_n56,
         EXEC_STAGE_mul_ex_mult_84_n55, EXEC_STAGE_mul_ex_mult_84_n54,
         EXEC_STAGE_mul_ex_mult_84_n53, EXEC_STAGE_mul_ex_mult_84_n52,
         EXEC_STAGE_mul_ex_mult_84_n51, EXEC_STAGE_mul_ex_mult_84_n50,
         EXEC_STAGE_mul_ex_mult_84_n49, EXEC_STAGE_mul_ex_mult_84_n48,
         EXEC_STAGE_mul_ex_mult_84_n47, EXEC_STAGE_mul_ex_mult_84_n46,
         EXEC_STAGE_mul_ex_mult_84_n45, EXEC_STAGE_mul_ex_mult_84_n44,
         EXEC_STAGE_mul_ex_mult_84_n43, EXEC_STAGE_mul_ex_mult_84_n42,
         EXEC_STAGE_mul_ex_mult_84_n41, EXEC_STAGE_mul_ex_mult_84_n40,
         EXEC_STAGE_mul_ex_mult_84_n39, EXEC_STAGE_mul_ex_mult_84_n38,
         EXEC_STAGE_mul_ex_mult_84_n37, EXEC_STAGE_mul_ex_mult_84_n36,
         EXEC_STAGE_mul_ex_mult_84_n35, EXEC_STAGE_mul_ex_mult_84_n34,
         EXEC_STAGE_mul_ex_mult_84_n33, EXEC_STAGE_mul_ex_mult_84_n32,
         EXEC_STAGE_mul_ex_mult_84_n31, EXEC_STAGE_mul_ex_mult_84_n30,
         EXEC_STAGE_mul_ex_mult_84_n29, EXEC_STAGE_mul_ex_mult_84_n28,
         EXEC_STAGE_mul_ex_mult_84_n27, EXEC_STAGE_mul_ex_mult_84_n26,
         EXEC_STAGE_mul_ex_mult_84_n25, EXEC_STAGE_mul_ex_mult_84_n24,
         EXEC_STAGE_mul_ex_mult_84_n23, EXEC_STAGE_mul_ex_mult_84_n22,
         EXEC_STAGE_mul_ex_mult_84_n21, EXEC_STAGE_mul_ex_mult_84_n20,
         EXEC_STAGE_mul_ex_mult_84_n19, EXEC_STAGE_mul_ex_mult_84_n18,
         EXEC_STAGE_mul_ex_mult_84_n17, EXEC_STAGE_mul_ex_mult_84_n16,
         EXEC_STAGE_mul_ex_mult_84_n15, EXEC_STAGE_mul_ex_mult_84_n14,
         EXEC_STAGE_mul_ex_mult_84_n13, EXEC_STAGE_mul_ex_mult_84_n12,
         EXEC_STAGE_mul_ex_mult_84_n11, EXEC_STAGE_mul_ex_mult_84_n10,
         EXEC_STAGE_mul_ex_mult_84_n9, EXEC_STAGE_mul_ex_mult_84_n8,
         EXEC_STAGE_mul_ex_mult_84_n7, EXEC_STAGE_mul_ex_mult_84_n6,
         EXEC_STAGE_mul_ex_mult_84_n5, EXEC_STAGE_mul_ex_mult_84_n4,
         EXEC_STAGE_mul_ex_mult_84_n3, EXEC_STAGE_mul_ex_mult_84_A1_0_,
         EXEC_STAGE_mul_ex_mult_84_A1_1_, EXEC_STAGE_mul_ex_mult_84_A1_2_,
         EXEC_STAGE_mul_ex_mult_84_A1_3_, EXEC_STAGE_mul_ex_mult_84_A1_4_,
         EXEC_STAGE_mul_ex_mult_84_A1_5_, EXEC_STAGE_mul_ex_mult_84_A1_6_,
         EXEC_STAGE_mul_ex_mult_84_A1_7_, EXEC_STAGE_mul_ex_mult_84_A1_8_,
         EXEC_STAGE_mul_ex_mult_84_A1_9_, EXEC_STAGE_mul_ex_mult_84_A1_10_,
         EXEC_STAGE_mul_ex_mult_84_A1_11_, EXEC_STAGE_mul_ex_mult_84_A1_12_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_2__1_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_2__2_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_2__3_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_2__4_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_2__5_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_2__6_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_2__7_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_2__8_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_2__9_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_2__10_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_2__11_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_2__12_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_2__13_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_2__14_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_3__1_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_3__2_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_3__3_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_3__4_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_3__5_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_3__6_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_3__7_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_3__8_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_3__9_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_3__10_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_3__11_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_3__12_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_3__13_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_3__14_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_4__1_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_4__2_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_4__3_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_4__4_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_4__5_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_4__6_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_4__7_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_4__8_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_4__9_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_4__10_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_4__11_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_4__12_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_4__13_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_4__14_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_5__1_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_5__2_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_5__3_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_5__4_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_5__5_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_5__6_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_5__7_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_5__8_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_5__9_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_5__10_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_5__11_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_5__12_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_5__13_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_5__14_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_6__1_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_6__2_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_6__3_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_6__4_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_6__5_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_6__6_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_6__7_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_6__8_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_6__9_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_6__10_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_6__11_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_6__12_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_6__13_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_6__14_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_7__1_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_7__2_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_7__3_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_7__4_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_7__5_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_7__6_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_7__7_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_7__8_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_7__9_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_7__10_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_7__11_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_7__12_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_7__13_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_7__14_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_8__1_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_8__2_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_8__3_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_8__4_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_8__5_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_8__6_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_8__7_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_8__8_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_8__9_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_8__10_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_8__11_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_8__12_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_8__13_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_8__14_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_9__1_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_9__2_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_9__3_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_9__4_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_9__5_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_9__6_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_9__7_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_9__8_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_9__9_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_9__10_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_9__11_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_9__12_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_9__13_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_9__14_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_10__1_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_10__2_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_10__3_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_10__4_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_10__5_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_10__6_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_10__7_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_10__8_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_10__9_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_10__10_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_10__11_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_10__12_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_10__13_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_10__14_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_11__1_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_11__2_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_11__3_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_11__4_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_11__5_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_11__6_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_11__7_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_11__8_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_11__9_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_11__10_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_11__11_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_11__12_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_11__13_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_11__14_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_12__1_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_12__2_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_12__3_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_12__4_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_12__5_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_12__6_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_12__7_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_12__8_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_12__9_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_12__10_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_12__11_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_12__12_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_12__13_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_12__14_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_13__1_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_13__2_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_13__3_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_13__4_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_13__5_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_13__6_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_13__7_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_13__8_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_13__9_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_13__10_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_13__11_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_13__12_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_13__13_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_13__14_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_14__1_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_14__2_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_14__3_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_14__4_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_14__5_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_14__6_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_14__7_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_14__8_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_14__9_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_14__10_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_14__11_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_14__12_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_14__13_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_14__14_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_15__0_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_15__1_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_15__2_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_15__3_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_15__4_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_15__5_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_15__6_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_15__7_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_15__8_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_15__9_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_15__10_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_15__11_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_15__12_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_15__13_,
         EXEC_STAGE_mul_ex_mult_84_SUMB_15__14_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_2__0_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_2__1_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_2__2_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_2__3_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_2__4_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_2__5_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_2__6_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_2__7_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_2__8_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_2__9_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_2__10_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_2__11_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_2__12_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_2__13_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_2__14_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_3__0_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_3__1_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_3__2_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_3__3_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_3__4_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_3__5_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_3__6_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_3__7_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_3__8_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_3__9_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_3__10_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_3__11_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_3__12_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_3__13_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_3__14_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_4__0_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_4__1_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_4__2_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_4__3_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_4__4_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_4__5_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_4__6_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_4__7_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_4__8_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_4__9_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_4__10_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_4__11_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_4__12_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_4__13_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_4__14_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_5__0_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_5__1_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_5__2_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_5__3_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_5__4_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_5__5_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_5__6_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_5__7_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_5__8_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_5__9_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_5__10_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_5__11_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_5__12_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_5__13_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_5__14_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_6__0_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_6__1_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_6__2_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_6__3_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_6__4_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_6__5_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_6__6_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_6__7_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_6__8_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_6__9_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_6__10_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_6__11_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_6__12_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_6__13_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_6__14_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_7__0_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_7__1_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_7__2_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_7__3_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_7__4_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_7__5_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_7__6_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_7__7_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_7__8_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_7__9_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_7__10_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_7__11_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_7__12_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_7__13_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_7__14_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_8__0_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_8__1_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_8__2_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_8__3_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_8__4_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_8__5_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_8__6_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_8__7_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_8__8_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_8__9_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_8__10_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_8__11_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_8__12_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_8__13_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_8__14_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_9__0_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_9__1_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_9__2_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_9__3_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_9__4_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_9__5_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_9__6_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_9__7_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_9__8_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_9__9_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_9__10_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_9__11_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_9__12_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_9__13_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_9__14_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_10__0_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_10__1_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_10__2_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_10__3_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_10__4_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_10__5_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_10__6_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_10__7_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_10__8_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_10__9_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_10__10_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_10__11_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_10__12_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_10__13_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_10__14_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_11__0_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_11__1_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_11__2_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_11__3_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_11__4_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_11__5_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_11__6_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_11__7_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_11__8_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_11__9_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_11__10_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_11__11_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_11__12_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_11__13_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_11__14_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_12__0_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_12__1_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_12__2_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_12__3_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_12__4_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_12__5_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_12__6_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_12__7_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_12__8_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_12__9_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_12__10_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_12__11_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_12__12_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_12__13_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_12__14_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_13__0_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_13__1_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_13__2_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_13__3_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_13__4_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_13__5_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_13__6_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_13__7_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_13__8_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_13__9_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_13__10_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_13__11_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_13__12_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_13__13_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_13__14_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_14__0_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_14__1_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_14__2_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_14__3_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_14__4_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_14__5_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_14__6_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_14__7_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_14__8_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_14__9_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_14__10_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_14__11_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_14__12_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_14__13_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_14__14_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_15__0_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_15__1_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_15__2_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_15__3_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_15__4_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_15__5_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_15__6_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_15__7_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_15__8_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_15__9_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_15__10_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_15__11_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_15__12_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_15__13_,
         EXEC_STAGE_mul_ex_mult_84_CARRYB_15__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_0__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_0__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_0__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_0__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_0__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_0__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_0__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_0__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_0__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_0__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_0__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_0__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_0__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_0__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_0__15_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__0_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_1__15_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__0_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_2__15_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__0_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_3__15_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__0_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_4__15_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__0_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_5__15_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__0_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_6__15_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__0_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_7__15_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__0_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_8__15_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__0_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_9__15_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__0_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_10__15_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__0_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_11__15_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__0_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_12__15_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__0_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_13__15_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__0_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_14__15_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__0_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__1_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__2_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__3_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__4_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__5_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__6_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__7_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__8_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__9_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__10_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__11_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__12_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__13_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__14_,
         EXEC_STAGE_mul_ex_mult_84_ab_15__15_,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n70,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n69,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n68,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n67,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n66,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n65,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n64,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n63,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n62,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n61,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n60,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n59,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n58,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n57,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n56,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n55,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n54,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n53,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n52,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n51,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n50,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n49,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n48,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n47,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n46,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n45,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n44,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n43,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n42,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n41,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n40,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n39,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n38,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n37,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n36,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n35,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n34,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n33,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n32,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n31,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n30,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n29,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n28,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n27,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n26,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n25,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n24,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n23,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n22,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n21,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n20,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n19,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n18,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n17,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n16,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n15,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n14,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n13,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n12,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n11,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n10, EXEC_STAGE_mul_ex_mult_84_FS_1_n9,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n8, EXEC_STAGE_mul_ex_mult_84_FS_1_n7,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n6, EXEC_STAGE_mul_ex_mult_84_FS_1_n5,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n4, EXEC_STAGE_mul_ex_mult_84_FS_1_n3,
         EXEC_STAGE_mul_ex_mult_84_FS_1_n1, EXEC_STAGE_mul_ex_mult_76_n94,
         EXEC_STAGE_mul_ex_mult_76_n93, EXEC_STAGE_mul_ex_mult_76_n92,
         EXEC_STAGE_mul_ex_mult_76_n91, EXEC_STAGE_mul_ex_mult_76_n90,
         EXEC_STAGE_mul_ex_mult_76_n89, EXEC_STAGE_mul_ex_mult_76_n88,
         EXEC_STAGE_mul_ex_mult_76_n87, EXEC_STAGE_mul_ex_mult_76_n86,
         EXEC_STAGE_mul_ex_mult_76_n85, EXEC_STAGE_mul_ex_mult_76_n84,
         EXEC_STAGE_mul_ex_mult_76_n83, EXEC_STAGE_mul_ex_mult_76_n82,
         EXEC_STAGE_mul_ex_mult_76_n81, EXEC_STAGE_mul_ex_mult_76_n80,
         EXEC_STAGE_mul_ex_mult_76_n79, EXEC_STAGE_mul_ex_mult_76_n78,
         EXEC_STAGE_mul_ex_mult_76_n77, EXEC_STAGE_mul_ex_mult_76_n76,
         EXEC_STAGE_mul_ex_mult_76_n75, EXEC_STAGE_mul_ex_mult_76_n74,
         EXEC_STAGE_mul_ex_mult_76_n73, EXEC_STAGE_mul_ex_mult_76_n72,
         EXEC_STAGE_mul_ex_mult_76_n71, EXEC_STAGE_mul_ex_mult_76_n70,
         EXEC_STAGE_mul_ex_mult_76_n69, EXEC_STAGE_mul_ex_mult_76_n68,
         EXEC_STAGE_mul_ex_mult_76_n67, EXEC_STAGE_mul_ex_mult_76_n66,
         EXEC_STAGE_mul_ex_mult_76_n65, EXEC_STAGE_mul_ex_mult_76_n64,
         EXEC_STAGE_mul_ex_mult_76_n63, EXEC_STAGE_mul_ex_mult_76_n62,
         EXEC_STAGE_mul_ex_mult_76_n61, EXEC_STAGE_mul_ex_mult_76_n60,
         EXEC_STAGE_mul_ex_mult_76_n59, EXEC_STAGE_mul_ex_mult_76_n58,
         EXEC_STAGE_mul_ex_mult_76_n57, EXEC_STAGE_mul_ex_mult_76_n56,
         EXEC_STAGE_mul_ex_mult_76_n55, EXEC_STAGE_mul_ex_mult_76_n54,
         EXEC_STAGE_mul_ex_mult_76_n53, EXEC_STAGE_mul_ex_mult_76_n52,
         EXEC_STAGE_mul_ex_mult_76_n51, EXEC_STAGE_mul_ex_mult_76_n50,
         EXEC_STAGE_mul_ex_mult_76_n49, EXEC_STAGE_mul_ex_mult_76_n48,
         EXEC_STAGE_mul_ex_mult_76_n47, EXEC_STAGE_mul_ex_mult_76_n45,
         EXEC_STAGE_mul_ex_mult_76_n44, EXEC_STAGE_mul_ex_mult_76_n43,
         EXEC_STAGE_mul_ex_mult_76_n42, EXEC_STAGE_mul_ex_mult_76_n41,
         EXEC_STAGE_mul_ex_mult_76_n40, EXEC_STAGE_mul_ex_mult_76_n39,
         EXEC_STAGE_mul_ex_mult_76_n38, EXEC_STAGE_mul_ex_mult_76_n37,
         EXEC_STAGE_mul_ex_mult_76_n36, EXEC_STAGE_mul_ex_mult_76_n35,
         EXEC_STAGE_mul_ex_mult_76_n34, EXEC_STAGE_mul_ex_mult_76_n33,
         EXEC_STAGE_mul_ex_mult_76_n32, EXEC_STAGE_mul_ex_mult_76_n31,
         EXEC_STAGE_mul_ex_mult_76_n30, EXEC_STAGE_mul_ex_mult_76_n29,
         EXEC_STAGE_mul_ex_mult_76_n28, EXEC_STAGE_mul_ex_mult_76_n27,
         EXEC_STAGE_mul_ex_mult_76_n26, EXEC_STAGE_mul_ex_mult_76_n25,
         EXEC_STAGE_mul_ex_mult_76_n24, EXEC_STAGE_mul_ex_mult_76_n23,
         EXEC_STAGE_mul_ex_mult_76_n22, EXEC_STAGE_mul_ex_mult_76_n21,
         EXEC_STAGE_mul_ex_mult_76_n20, EXEC_STAGE_mul_ex_mult_76_n19,
         EXEC_STAGE_mul_ex_mult_76_n18, EXEC_STAGE_mul_ex_mult_76_n17,
         EXEC_STAGE_mul_ex_mult_76_n16, EXEC_STAGE_mul_ex_mult_76_n15,
         EXEC_STAGE_mul_ex_mult_76_n14, EXEC_STAGE_mul_ex_mult_76_n13,
         EXEC_STAGE_mul_ex_mult_76_n12, EXEC_STAGE_mul_ex_mult_76_n11,
         EXEC_STAGE_mul_ex_mult_76_n10, EXEC_STAGE_mul_ex_mult_76_n9,
         EXEC_STAGE_mul_ex_mult_76_n8, EXEC_STAGE_mul_ex_mult_76_n7,
         EXEC_STAGE_mul_ex_mult_76_n6, EXEC_STAGE_mul_ex_mult_76_n5,
         EXEC_STAGE_mul_ex_mult_76_n4, EXEC_STAGE_mul_ex_mult_76_n3,
         EXEC_STAGE_mul_ex_mult_76_A1_0_, EXEC_STAGE_mul_ex_mult_76_A1_1_,
         EXEC_STAGE_mul_ex_mult_76_A1_2_, EXEC_STAGE_mul_ex_mult_76_A1_3_,
         EXEC_STAGE_mul_ex_mult_76_A1_4_, EXEC_STAGE_mul_ex_mult_76_A1_5_,
         EXEC_STAGE_mul_ex_mult_76_A1_6_, EXEC_STAGE_mul_ex_mult_76_A1_7_,
         EXEC_STAGE_mul_ex_mult_76_A1_8_, EXEC_STAGE_mul_ex_mult_76_A1_9_,
         EXEC_STAGE_mul_ex_mult_76_A1_10_, EXEC_STAGE_mul_ex_mult_76_A1_11_,
         EXEC_STAGE_mul_ex_mult_76_A1_12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__0_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__15_,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n70,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n69,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n68,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n67,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n66,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n65,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n64,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n63,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n62,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n61,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n60,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n59,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n58,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n57,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n56,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n55,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n54,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n53,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n52,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n51,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n50,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n49,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n48,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n47,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n46,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n45,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n44,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n43,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n42,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n41,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n40,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n39,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n38,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n37,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n36,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n35,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n34,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n33,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n32,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n31,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n30,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n29,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n28,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n27,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n26,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n25,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n24,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n23,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n22,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n21,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n20,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n19,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n18,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n17,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n16,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n15,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n14,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n13,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n12,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n11,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n10, EXEC_STAGE_mul_ex_mult_76_FS_1_n9,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n8, EXEC_STAGE_mul_ex_mult_76_FS_1_n7,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n6, EXEC_STAGE_mul_ex_mult_76_FS_1_n5,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n4, EXEC_STAGE_mul_ex_mult_76_FS_1_n3,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n1;
  wire   [24:37] IF_ID_OUT;
  wire   [0:9] offset_26_id;
  wire   [32:276] ID_EXEC_OUT;
  wire   [0:31] nextPC_ex_out;
  wire   [102:105] EXEC_MEM_IN;
  wire   [0:178] MEM_WB_OUT;
  wire   [0:4] destReg_wb_out;
  wire   [16:31] ID_STAGE_imm16_aluA;
  wire   [6:31] EXEC_STAGE_imm26_32;
  wire   [16:31] EXEC_STAGE_imm16_32;
  wire   [0:63] EXEC_STAGE_mul_result_long;
  wire   [0:31] EXEC_STAGE_mul_ex_P;
  wire   [0:31] EXEC_STAGE_mul_ex_H;
  wire   [16:31] WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf;
  wire   [15:2] EXEC_STAGE_mul_ex_add_88_carry;
  wire   [15:2] EXEC_STAGE_mul_ex_add_88_2_carry;
  wire   [31:1] sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry;
  wire   [31:1] sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry;

  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_235_ ( .D(n8020), .CK(clk), .RN(n13914), 
        .Q(ID_EXEC_OUT[235]), .QN(n10815) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_100_ ( .D(n19151), .CK(clk), .RN(
        n13882), .Q(DMEM_BUS_OUT[31]), .QN(n11990) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_141_ ( .D(n8018), .CK(clk), .RN(
        n13891), .Q(EXEC_MEM_OUT_141), .QN(n10157) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_98_ ( .D(n8014), .CK(clk), .RN(n13932), 
        .Q(MEM_WB_OUT[98]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_97_ ( .D(n8013), .CK(clk), .RN(n13881), 
        .Q(MEM_WB_OUT[97]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_96_ ( .D(n8012), .CK(clk), .RN(n13932), 
        .Q(MEM_WB_OUT[96]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_79_ ( .D(n8011), .CK(clk), .RN(n13881), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[26]), .QN(n12220) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_148_ ( .D(n7996), .CK(clk), .RN(n13897), 
        .Q(ID_EXEC_OUT[148]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_57_ ( .D(n7992), .CK(clk), .RN(n13887), 
        .QN(n12300) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_96_ ( .D(n7969), .CK(clk), .RN(n13922), 
        .Q(EXEC_STAGE_imm26_32[6]), .QN(n12217) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_97_ ( .D(n7966), .CK(clk), .RN(n13891), 
        .Q(EXEC_STAGE_imm26_32[7]), .QN(n12218) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_98_ ( .D(n7963), .CK(clk), .RN(n13922), 
        .Q(EXEC_STAGE_imm26_32[8]), .QN(n12057) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_99_ ( .D(n7960), .CK(clk), .RN(n13885), 
        .Q(EXEC_STAGE_imm26_32[9]), .QN(n12056) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_100_ ( .D(n7957), .CK(clk), .RN(n13881), 
        .Q(EXEC_STAGE_imm26_32[10]), .QN(n12055) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_103_ ( .D(n7952), .CK(clk), .RN(n13905), 
        .Q(EXEC_STAGE_imm26_32[13]), .QN(n12214) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_104_ ( .D(n7949), .CK(clk), .RN(n13916), 
        .Q(EXEC_STAGE_imm26_32[14]), .QN(n12054) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_105_ ( .D(n7946), .CK(clk), .RN(n13909), 
        .QN(n12065) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_268_ ( .D(n7944), .CK(clk), .RN(n13892), 
        .QN(n10935) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_180_ ( .D(n7943), .CK(clk), .RN(
        n13907), .QN(n12198) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_108_ ( .D(n7942), .CK(clk), .RN(n13887), .Q(MEM_WB_OUT[108]), .QN(n10845) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_122_ ( .D(n7941), .CK(clk), .RN(n13889), 
        .Q(EXEC_STAGE_imm16_32[16]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_106_ ( .D(n7940), .CK(clk), .RN(n13919), 
        .Q(EXEC_STAGE_imm26_32[16]), .QN(n12058) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_107_ ( .D(n7938), .CK(clk), .RN(n13890), 
        .Q(EXEC_STAGE_imm26_32[17]), .QN(n11569) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_123_ ( .D(n7937), .CK(clk), .RN(n13913), 
        .Q(EXEC_STAGE_imm16_32[17]), .QN(n12566) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_269_ ( .D(n7936), .CK(clk), .RN(n13920), 
        .QN(n10936) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_181_ ( .D(n7935), .CK(clk), .RN(
        n13902), .QN(n12199) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_109_ ( .D(n7934), .CK(clk), .RN(n13925), .Q(MEM_WB_OUT[109]), .QN(n10802) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_108_ ( .D(n7932), .CK(clk), .RN(n13897), 
        .QN(n12072) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_124_ ( .D(n7931), .CK(clk), .RN(n13909), 
        .QN(n12551) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_270_ ( .D(n7930), .CK(clk), .RN(n13919), 
        .QN(n10937) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_182_ ( .D(n7929), .CK(clk), .RN(
        n13907), .QN(n12200) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_110_ ( .D(n7928), .CK(clk), .RN(n13925), .Q(MEM_WB_OUT[110]), .QN(n10353) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_271_ ( .D(n7924), .CK(clk), .RN(n13892), 
        .QN(n10938) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_183_ ( .D(n7923), .CK(clk), .RN(
        n13902), .QN(n12201) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_111_ ( .D(n7922), .CK(clk), .RN(n13884), .Q(MEM_WB_OUT[111]), .QN(n10817) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_272_ ( .D(n7918), .CK(clk), .RN(n13919), 
        .QN(n10939) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_184_ ( .D(n7917), .CK(clk), .RN(
        n13907), .QN(n12202) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_112_ ( .D(n7916), .CK(clk), .RN(n13925), .Q(MEM_WB_OUT[112]), .QN(n10947) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_152_ ( .D(n7905), .CK(clk), .RN(n13914), 
        .QN(n10933) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_106_ ( .D(n7904), .CK(clk), .RN(
        n13923), .Q(MEM_WB_REG_MEM_WB_REG_N75), .QN(n12522) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_145_ ( .D(n7900), .CK(clk), .RN(n13914), 
        .Q(ID_EXEC_OUT[145]), .QN(n12136) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_144_ ( .D(n7898), .CK(clk), .RN(n13897), 
        .Q(EXEC_MEM_IN[102]), .QN(n10948) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_150_ ( .D(n7896), .CK(clk), .RN(n13914), 
        .QN(n12064) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_138_ ( .D(n7893), .CK(clk), .RN(n13913), 
        .QN(n12182) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_139_ ( .D(n7890), .CK(clk), .RN(n13897), 
        .QN(n12306) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_140_ ( .D(n7887), .CK(clk), .RN(n13897), 
        .QN(n12183) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_141_ ( .D(n7884), .CK(clk), .RN(n13914), 
        .QN(n12307) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_143_ ( .D(n7881), .CK(clk), .RN(n13914), 
        .QN(n12197) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_101_ ( .D(n7880), .CK(clk), .RN(
        n13897), .Q(MEM_WB_REG_MEM_WB_REG_N78), .QN(n11543) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_147_ ( .D(n7878), .CK(clk), .RN(n13914), 
        .QN(n12212) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_151_ ( .D(n7877), .CK(clk), .RN(n13897), 
        .Q(EXEC_MEM_IN[105]), .QN(n13142) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_142_ ( .D(n7876), .CK(clk), .RN(n13897), 
        .QN(n12184) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_275_ ( .D(n7873), .CK(clk), .RN(n13919), 
        .Q(ID_EXEC_OUT[275]), .QN(n12017) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_149_ ( .D(n7872), .CK(clk), .RN(n13914), 
        .QN(n12051) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_276_ ( .D(n7869), .CK(clk), .RN(n13892), 
        .Q(ID_EXEC_OUT[276]), .QN(n10906) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_84_ ( .D(n7864), .CK(clk), .RN(n13881), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[31]), .QN(n12050) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_85_ ( .D(n7863), .CK(clk), .RN(n13932), 
        .Q(MEM_WB_OUT[85]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_86_ ( .D(n7862), .CK(clk), .RN(n13881), 
        .Q(MEM_WB_OUT[86]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_87_ ( .D(n7861), .CK(clk), .RN(n13932), 
        .Q(MEM_WB_OUT[87]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_88_ ( .D(n7860), .CK(clk), .RN(n13881), 
        .Q(MEM_WB_OUT[88]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_89_ ( .D(n7859), .CK(clk), .RN(n13932), 
        .Q(MEM_WB_OUT[89]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_90_ ( .D(n7858), .CK(clk), .RN(n13932), 
        .Q(MEM_WB_OUT[90]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_91_ ( .D(n7857), .CK(clk), .RN(n13881), 
        .Q(MEM_WB_OUT[91]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_93_ ( .D(n7855), .CK(clk), .RN(n13881), 
        .Q(MEM_WB_OUT[93]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_94_ ( .D(n7854), .CK(clk), .RN(n13932), 
        .Q(MEM_WB_OUT[94]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_274_ ( .D(n7852), .CK(clk), .RN(n13892), 
        .QN(n11102) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_249_ ( .D(n7851), .CK(clk), .RN(
        n13910), .QN(n12203) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_177_ ( .D(n7850), .CK(clk), .RN(n13884), .QN(n10365) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_154_ ( .D(n7849), .CK(clk), .RN(n13914), 
        .Q(DSize_ex_out_0_), .QN(n11542) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_107_ ( .D(n7848), .CK(clk), .RN(
        n13895), .Q(DMEM_BUS_OUT[65]), .QN(n10781) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_155_ ( .D(n7846), .CK(clk), .RN(n13896), 
        .QN(n12052) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_108_ ( .D(n7845), .CK(clk), .RN(
        n13912), .Q(DMEM_BUS_OUT[66]), .QN(n11471) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_156_ ( .D(n7843), .CK(clk), .RN(n13914), 
        .Q(ID_EXEC_OUT[156]), .QN(n10236) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_157_ ( .D(n7842), .CK(clk), .RN(n13896), 
        .Q(ID_EXEC_OUT[157]), .QN(n11915) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_101_ ( .D(n7838), .CK(clk), .RN(n13906), 
        .Q(EXEC_STAGE_imm26_32[11]), .QN(n12215) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_102_ ( .D(n7836), .CK(clk), .RN(n13923), 
        .Q(EXEC_STAGE_imm26_32[12]), .QN(n12216) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_105_ ( .D(n7835), .CK(clk), .RN(
        n13919), .Q(DMEM_BUS_OUT[64]), .QN(n12601) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_140_ ( .D(n7834), .CK(clk), .RN(
        n13906), .Q(EXEC_MEM_OUT_140), .QN(n11505) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_31_ ( .D(n7833), .CK(clk), .RN(n13889), 
        .QN(n11111) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_31_ ( .D(n7831), .CK(clk), .RN(
        n13911), .QN(n11109) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_31_ ( .D(n7830), .CK(clk), .RN(n13884), 
        .Q(MEM_WB_OUT[31]), .QN(n12538) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_191_ ( .D(n7829), .CK(clk), .RN(n13895), 
        .Q(ID_EXEC_OUT[191]), .QN(n11537) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_95_ ( .D(n7828), .CK(clk), .RN(n13898), 
        .Q(ID_EXEC_OUT[95]), .QN(n12275) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_63_ ( .D(n7827), .CK(clk), .RN(n13920), 
        .Q(ID_EXEC_OUT[63]), .QN(n12550) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_173_ ( .D(n7826), .CK(clk), .RN(
        n13907), .Q(DMEM_BUS_OUT[63]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_185_ ( .D(n19193), .CK(clk), .RN(
        n13902), .Q(MEM_WB_REG_MEM_WB_REG_N66) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_113_ ( .D(n19277), .CK(clk), .RN(
        n13911), .Q(MEM_WB_OUT[113]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_186_ ( .D(n19194), .CK(clk), .RN(
        n13908), .Q(MEM_WB_REG_MEM_WB_REG_N65) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_114_ ( .D(n19276), .CK(clk), .RN(
        n13925), .Q(MEM_WB_OUT[114]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_187_ ( .D(n19195), .CK(clk), .RN(
        n13902), .Q(MEM_WB_REG_MEM_WB_REG_N64) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_115_ ( .D(n19275), .CK(clk), .RN(
        n13893), .Q(MEM_WB_OUT[115]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_188_ ( .D(n19196), .CK(clk), .RN(
        n13908), .Q(MEM_WB_REG_MEM_WB_REG_N63) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_116_ ( .D(n19274), .CK(clk), .RN(
        n13926), .Q(MEM_WB_OUT[116]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_189_ ( .D(n19197), .CK(clk), .RN(
        n13902), .Q(MEM_WB_REG_MEM_WB_REG_N62) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_117_ ( .D(n19273), .CK(clk), .RN(
        n13896), .Q(MEM_WB_OUT[117]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_190_ ( .D(n19198), .CK(clk), .RN(
        n13902), .Q(MEM_WB_REG_MEM_WB_REG_N61) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_118_ ( .D(n19272), .CK(clk), .RN(
        n13926), .Q(MEM_WB_OUT[118]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_191_ ( .D(n19199), .CK(clk), .RN(
        n13908), .Q(MEM_WB_REG_MEM_WB_REG_N60) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_119_ ( .D(n19271), .CK(clk), .RN(
        n13898), .Q(MEM_WB_OUT[119]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_192_ ( .D(n19200), .CK(clk), .RN(
        n13902), .Q(MEM_WB_REG_MEM_WB_REG_N59) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_120_ ( .D(n19270), .CK(clk), .RN(
        n13914), .Q(MEM_WB_OUT[120]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_193_ ( .D(n19201), .CK(clk), .RN(
        n13908), .Q(MEM_WB_REG_MEM_WB_REG_N58) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_121_ ( .D(n19269), .CK(clk), .RN(
        n13926), .Q(MEM_WB_OUT[121]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_194_ ( .D(n19202), .CK(clk), .RN(
        n13902), .Q(MEM_WB_REG_MEM_WB_REG_N57) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_122_ ( .D(n19268), .CK(clk), .RN(
        n13915), .Q(MEM_WB_OUT[122]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_195_ ( .D(n19203), .CK(clk), .RN(
        n13908), .Q(MEM_WB_REG_MEM_WB_REG_N56) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_123_ ( .D(n19267), .CK(clk), .RN(
        n13926), .Q(MEM_WB_OUT[123]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_196_ ( .D(n19204), .CK(clk), .RN(
        n13902), .Q(MEM_WB_REG_MEM_WB_REG_N55) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_124_ ( .D(n19266), .CK(clk), .RN(
        n13917), .Q(MEM_WB_OUT[124]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_197_ ( .D(n19205), .CK(clk), .RN(
        n13908), .Q(MEM_WB_REG_MEM_WB_REG_N54) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_125_ ( .D(n19265), .CK(clk), .RN(
        n13926), .Q(MEM_WB_OUT[125]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_198_ ( .D(n19206), .CK(clk), .RN(
        n13902), .Q(MEM_WB_REG_MEM_WB_REG_N53) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_126_ ( .D(n19264), .CK(clk), .RN(
        n13918), .Q(MEM_WB_OUT[126]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_199_ ( .D(n19207), .CK(clk), .RN(
        n13908), .Q(MEM_WB_REG_MEM_WB_REG_N52) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_127_ ( .D(n19263), .CK(clk), .RN(
        n13926), .Q(MEM_WB_OUT[127]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_200_ ( .D(n19208), .CK(clk), .RN(
        n13901), .Q(MEM_WB_REG_MEM_WB_REG_N51) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_128_ ( .D(n19262), .CK(clk), .RN(
        n13883), .Q(MEM_WB_OUT[128]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_201_ ( .D(n19209), .CK(clk), .RN(
        n13908), .Q(MEM_WB_REG_MEM_WB_REG_N50) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_129_ ( .D(n19261), .CK(clk), .RN(
        n13926), .Q(MEM_WB_OUT[129]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_202_ ( .D(n19210), .CK(clk), .RN(
        n13901), .Q(MEM_WB_REG_MEM_WB_REG_N49) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_130_ ( .D(n19260), .CK(clk), .RN(
        n13926), .Q(MEM_WB_OUT[130]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_203_ ( .D(n19211), .CK(clk), .RN(
        n13908), .Q(MEM_WB_REG_MEM_WB_REG_N48) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_131_ ( .D(n19259), .CK(clk), .RN(
        n13886), .Q(MEM_WB_OUT[131]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_204_ ( .D(n19212), .CK(clk), .RN(
        n13901), .Q(MEM_WB_REG_MEM_WB_REG_N47) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_132_ ( .D(n19258), .CK(clk), .RN(
        n13926), .Q(MEM_WB_OUT[132]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_205_ ( .D(n19213), .CK(clk), .RN(
        n13908), .Q(MEM_WB_REG_MEM_WB_REG_N46) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_133_ ( .D(n19257), .CK(clk), .RN(
        n13886), .Q(MEM_WB_OUT[133]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_206_ ( .D(n19214), .CK(clk), .RN(
        n13901), .Q(MEM_WB_REG_MEM_WB_REG_N45) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_134_ ( .D(n19256), .CK(clk), .RN(
        n13926), .Q(MEM_WB_OUT[134]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_207_ ( .D(n19215), .CK(clk), .RN(
        n13909), .Q(MEM_WB_REG_MEM_WB_REG_N44) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_135_ ( .D(n19255), .CK(clk), .RN(
        n13886), .Q(MEM_WB_OUT[135]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_208_ ( .D(n19216), .CK(clk), .RN(
        n13901), .Q(MEM_WB_REG_MEM_WB_REG_N43) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_136_ ( .D(n19254), .CK(clk), .RN(
        n13926), .Q(MEM_WB_OUT[136]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_209_ ( .D(n19217), .CK(clk), .RN(
        n13909), .Q(MEM_WB_REG_MEM_WB_REG_N42) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_137_ ( .D(n19253), .CK(clk), .RN(
        n13886), .Q(MEM_WB_OUT[137]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_210_ ( .D(n19218), .CK(clk), .RN(
        n13909), .Q(MEM_WB_REG_MEM_WB_REG_N41) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_138_ ( .D(n19252), .CK(clk), .RN(
        n13927), .Q(MEM_WB_OUT[138]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_211_ ( .D(n19219), .CK(clk), .RN(
        n13901), .Q(MEM_WB_REG_MEM_WB_REG_N40) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_139_ ( .D(n19251), .CK(clk), .RN(
        n13886), .Q(MEM_WB_OUT[139]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_212_ ( .D(n19220), .CK(clk), .RN(
        n13909), .Q(MEM_WB_REG_MEM_WB_REG_N39) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_140_ ( .D(n19250), .CK(clk), .RN(
        n13886), .Q(MEM_WB_OUT[140]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_213_ ( .D(n19221), .CK(clk), .RN(
        n13901), .Q(MEM_WB_REG_MEM_WB_REG_N38) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_141_ ( .D(n19249), .CK(clk), .RN(
        n13927), .Q(MEM_WB_OUT[141]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_214_ ( .D(n19222), .CK(clk), .RN(
        n13909), .Q(MEM_WB_REG_MEM_WB_REG_N37) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_142_ ( .D(n19248), .CK(clk), .RN(
        n13886), .Q(MEM_WB_OUT[142]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_215_ ( .D(n19223), .CK(clk), .RN(
        n13901), .Q(MEM_WB_REG_MEM_WB_REG_N36) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_143_ ( .D(n19247), .CK(clk), .RN(
        n13927), .Q(MEM_WB_OUT[143]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_216_ ( .D(n19224), .CK(clk), .RN(
        n13909), .Q(MEM_WB_REG_MEM_WB_REG_N35) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_144_ ( .D(n19246), .CK(clk), .RN(
        n13886), .Q(MEM_WB_OUT[144]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_248_ ( .D(n7761), .CK(clk), .RN(
        n13899), .QN(n12176) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_250_ ( .D(n7759), .CK(clk), .RN(
        n13911), .QN(n12204) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_178_ ( .D(n7758), .CK(clk), .RN(n13928), .Q(MEM_WB_OUT[178]), .QN(n12978) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_204_ ( .D(n7757), .CK(clk), .RN(n13894), 
        .Q(ID_EXEC_OUT[204]), .QN(n11960) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_69_ ( .D(n7756), .CK(clk), .RN(
        n13898), .Q(DMEM_BUS_OUT[0]), .QN(n10825) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_37_ ( .D(n7755), .CK(clk), .RN(n13883), 
        .Q(MEM_WB_OUT[37]), .QN(n12040) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_217_ ( .D(n7754), .CK(clk), .RN(
        n13901), .QN(n12178) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_87_ ( .D(n7752), .CK(clk), .RN(
        n13898), .Q(DMEM_BUS_OUT[18]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_55_ ( .D(n19230), .CK(clk), .RN(n13883), .Q(MEM_WB_OUT[55]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_235_ ( .D(n7750), .CK(clk), .RN(
        n13900), .QN(n12164) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_222_ ( .D(n7748), .CK(clk), .RN(n13926), 
        .Q(ID_EXEC_OUT[222]), .QN(n10814) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_254_ ( .D(n7747), .CK(clk), .RN(n13903), 
        .Q(ID_EXEC_OUT[254]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_99_ ( .D(n7746), .CK(clk), .RN(
        n13910), .Q(DMEM_BUS_OUT[30]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_67_ ( .D(n7745), .CK(clk), .RN(n13931), 
        .Q(MEM_WB_OUT[67]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_139_ ( .D(n7744), .CK(clk), .RN(
        n13906), .Q(EXEC_MEM_OUT_139), .QN(n11504) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_30_ ( .D(n7743), .CK(clk), .RN(n13923), 
        .QN(n11110) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_30_ ( .D(n7741), .CK(clk), .RN(
        n13899), .QN(n11108) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_30_ ( .D(n7740), .CK(clk), .RN(n13929), 
        .Q(MEM_WB_OUT[30]), .QN(n12537) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_190_ ( .D(n7739), .CK(clk), .RN(n13916), 
        .Q(ID_EXEC_OUT[190]), .QN(n11536) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_172_ ( .D(n7738), .CK(clk), .RN(
        n13903), .Q(DMEM_BUS_OUT[62]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_94_ ( .D(n7737), .CK(clk), .RN(n13922), 
        .Q(ID_EXEC_OUT[94]), .QN(n11562) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_62_ ( .D(n7736), .CK(clk), .RN(n13890), 
        .Q(ID_EXEC_OUT[62]), .QN(n12549) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_247_ ( .D(n7735), .CK(clk), .RN(
        n13910), .QN(n12175) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_234_ ( .D(n7733), .CK(clk), .RN(n13918), 
        .Q(ID_EXEC_OUT[234]), .QN(n11937) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_266_ ( .D(n7732), .CK(clk), .RN(n13892), 
        .Q(ID_EXEC_OUT[266]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_66_ ( .D(n7730), .CK(clk), .RN(n13882), 
        .Q(MEM_WB_OUT[66]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_138_ ( .D(n7729), .CK(clk), .RN(
        n13900), .Q(EXEC_MEM_OUT_138) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_29_ ( .D(n7728), .CK(clk), .RN(n13923), 
        .QN(n12310) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_29_ ( .D(n7726), .CK(clk), .RN(
        n13899), .QN(n11115) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_29_ ( .D(n7725), .CK(clk), .RN(n13929), 
        .Q(MEM_WB_OUT[29]), .QN(n12499) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_189_ ( .D(n7724), .CK(clk), .RN(n13916), 
        .Q(ID_EXEC_OUT[189]), .QN(n11535) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_171_ ( .D(n7723), .CK(clk), .RN(
        n13907), .Q(DMEM_BUS_OUT[61]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_93_ ( .D(n7722), .CK(clk), .RN(n13896), 
        .Q(ID_EXEC_OUT[93]), .QN(n11571) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_61_ ( .D(n7721), .CK(clk), .RN(n13920), 
        .Q(ID_EXEC_OUT[61]), .QN(n12301) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_246_ ( .D(n7720), .CK(clk), .RN(
        n13899), .QN(n12174) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_233_ ( .D(n7718), .CK(clk), .RN(n13918), 
        .Q(ID_EXEC_OUT[233]), .QN(n10823) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_265_ ( .D(n7717), .CK(clk), .RN(n13902), 
        .Q(ID_EXEC_OUT[265]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_62_ ( .D(n7715), .CK(clk), .RN(n13882), 
        .Q(MEM_WB_OUT[62]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_242_ ( .D(n7714), .CK(clk), .RN(
        n13900), .QN(n12299) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_229_ ( .D(n7712), .CK(clk), .RN(n13918), 
        .Q(ID_EXEC_OUT[229]), .QN(n11933) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_261_ ( .D(n7711), .CK(clk), .RN(n13930), 
        .Q(ID_EXEC_OUT[261]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_64_ ( .D(n7709), .CK(clk), .RN(n13882), 
        .Q(MEM_WB_OUT[64]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_244_ ( .D(n7708), .CK(clk), .RN(
        n13899), .QN(n12172) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_231_ ( .D(n7706), .CK(clk), .RN(n13908), 
        .Q(ID_EXEC_OUT[231]), .QN(n10819) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_263_ ( .D(n7705), .CK(clk), .RN(n13926), 
        .Q(ID_EXEC_OUT[263]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_243_ ( .D(n7702), .CK(clk), .RN(
        n13910), .QN(n12171) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_230_ ( .D(n7700), .CK(clk), .RN(n13918), 
        .Q(ID_EXEC_OUT[230]), .QN(n11936) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_262_ ( .D(n7699), .CK(clk), .RN(n13893), 
        .Q(ID_EXEC_OUT[262]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_61_ ( .D(n7697), .CK(clk), .RN(n13930), 
        .Q(MEM_WB_OUT[61]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_65_ ( .D(n7695), .CK(clk), .RN(n13931), 
        .Q(MEM_WB_OUT[65]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_137_ ( .D(n7694), .CK(clk), .RN(
        n13906), .Q(EXEC_MEM_OUT_137) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_28_ ( .D(n7693), .CK(clk), .RN(n13889), 
        .QN(n12192) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_28_ ( .D(n7691), .CK(clk), .RN(
        n13911), .Q(MEM_WB_REG_MEM_WB_REG_N152), .QN(n12523) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_28_ ( .D(n19241), .CK(clk), .RN(n13884), .Q(MEM_WB_OUT[28]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_188_ ( .D(n7689), .CK(clk), .RN(n13895), 
        .Q(ID_EXEC_OUT[188]), .QN(n11534) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_170_ ( .D(n7688), .CK(clk), .RN(
        n13903), .Q(DMEM_BUS_OUT[60]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_92_ ( .D(n7687), .CK(clk), .RN(n13922), 
        .Q(ID_EXEC_OUT[92]), .QN(n11280) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_60_ ( .D(n7686), .CK(clk), .RN(n13890), 
        .Q(ID_EXEC_OUT[60]), .QN(n12231) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_136_ ( .D(n7685), .CK(clk), .RN(
        n13901), .Q(EXEC_MEM_OUT_136) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_27_ ( .D(n7684), .CK(clk), .RN(n13923), 
        .QN(n19321) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_27_ ( .D(n7682), .CK(clk), .RN(
        n13899), .QN(n11107) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_27_ ( .D(n7681), .CK(clk), .RN(n13929), 
        .Q(MEM_WB_OUT[27]), .QN(n12224) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_187_ ( .D(n7680), .CK(clk), .RN(n13916), 
        .Q(ID_EXEC_OUT[187]), .QN(n11533) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_169_ ( .D(n7679), .CK(clk), .RN(
        n13903), .Q(DMEM_BUS_OUT[59]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_91_ ( .D(n7678), .CK(clk), .RN(n13893), 
        .Q(ID_EXEC_OUT[91]), .QN(n11563) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_59_ ( .D(n7677), .CK(clk), .RN(n13890), 
        .Q(ID_EXEC_OUT[59]), .QN(n12230) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_26_ ( .D(n7676), .CK(clk), .RN(n13889), 
        .QN(n12191) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_26_ ( .D(n7674), .CK(clk), .RN(
        n13911), .QN(n11114) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_26_ ( .D(n7673), .CK(clk), .RN(n13884), 
        .Q(MEM_WB_OUT[26]), .QN(n12536) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_186_ ( .D(n7672), .CK(clk), .RN(n13895), 
        .Q(ID_EXEC_OUT[186]), .QN(n11532) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_168_ ( .D(n7671), .CK(clk), .RN(
        n13907), .Q(DMEM_BUS_OUT[58]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_90_ ( .D(n7670), .CK(clk), .RN(n13922), 
        .Q(ID_EXEC_OUT[90]), .QN(n11561) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_58_ ( .D(n7669), .CK(clk), .RN(n13920), 
        .Q(ID_EXEC_OUT[58]), .QN(n12525) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_135_ ( .D(n7668), .CK(clk), .RN(
        n13905), .Q(EXEC_MEM_OUT_135), .QN(n12316) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_25_ ( .D(n7667), .CK(clk), .RN(n13923), 
        .QN(n19322) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_25_ ( .D(n7665), .CK(clk), .RN(
        n13899), .QN(n12308) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_25_ ( .D(n7664), .CK(clk), .RN(n13929), 
        .Q(MEM_WB_OUT[25]), .QN(n11136) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_185_ ( .D(n7663), .CK(clk), .RN(n13916), 
        .Q(ID_EXEC_OUT[185]), .QN(n11531) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_167_ ( .D(n7662), .CK(clk), .RN(
        n13903), .Q(DMEM_BUS_OUT[57]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_89_ ( .D(n7661), .CK(clk), .RN(n13922), 
        .Q(ID_EXEC_OUT[89]), .QN(n11570) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_57_ ( .D(n7660), .CK(clk), .RN(n13891), 
        .Q(ID_EXEC_OUT[57]), .QN(n12524) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_134_ ( .D(n7659), .CK(clk), .RN(
        n13902), .Q(EXEC_MEM_OUT_134), .QN(n11477) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_24_ ( .D(n7658), .CK(clk), .RN(n13889), 
        .Q(IF_ID_OUT[24]), .QN(n12500) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_24_ ( .D(n19289), .CK(clk), .RN(
        n13899), .Q(MEM_WB_REG_MEM_WB_REG_N156) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_24_ ( .D(n19242), .CK(clk), .RN(n13884), .Q(MEM_WB_OUT[24]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_184_ ( .D(n7654), .CK(clk), .RN(n13895), 
        .Q(ID_EXEC_OUT[184]), .QN(n11530) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_166_ ( .D(n7653), .CK(clk), .RN(
        n13907), .Q(DMEM_BUS_OUT[56]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_88_ ( .D(n7652), .CK(clk), .RN(n13886), 
        .Q(ID_EXEC_OUT[88]), .QN(n11560) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_56_ ( .D(n7651), .CK(clk), .RN(n13920), 
        .Q(ID_EXEC_OUT[56]), .QN(n12548) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_133_ ( .D(n7650), .CK(clk), .RN(
        n13905), .Q(EXEC_MEM_OUT_133), .QN(n11476) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_245_ ( .D(n7649), .CK(clk), .RN(
        n13910), .QN(n12173) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_232_ ( .D(n7647), .CK(clk), .RN(n13918), 
        .Q(ID_EXEC_OUT[232]), .QN(n11981) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_264_ ( .D(n7646), .CK(clk), .RN(n13892), 
        .Q(ID_EXEC_OUT[264]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_132_ ( .D(n7643), .CK(clk), .RN(
        n13890), .Q(EXEC_MEM_OUT_132) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_23_ ( .D(n7642), .CK(clk), .RN(n13923), 
        .QN(n19323) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_23_ ( .D(n7640), .CK(clk), .RN(
        n13910), .QN(n11106) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_23_ ( .D(n7639), .CK(clk), .RN(n13929), 
        .Q(MEM_WB_OUT[23]), .QN(n12535) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_183_ ( .D(n7638), .CK(clk), .RN(n13916), 
        .Q(ID_EXEC_OUT[183]), .QN(n11529) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_165_ ( .D(n7637), .CK(clk), .RN(
        n13903), .Q(DMEM_BUS_OUT[55]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_87_ ( .D(n7636), .CK(clk), .RN(n13922), 
        .Q(ID_EXEC_OUT[87]), .QN(n12543) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_55_ ( .D(n7635), .CK(clk), .RN(n13891), 
        .Q(ID_EXEC_OUT[55]), .QN(n12211) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_56_ ( .D(n19229), .CK(clk), .RN(n13930), .Q(MEM_WB_OUT[56]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_52_ ( .D(n19232), .CK(clk), .RN(n13930), .Q(MEM_WB_OUT[52]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_232_ ( .D(n7630), .CK(clk), .RN(
        n13910), .QN(n12161) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_219_ ( .D(n7628), .CK(clk), .RN(n13894), 
        .Q(ID_EXEC_OUT[219]), .QN(n10822) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_251_ ( .D(n7627), .CK(clk), .RN(n13893), 
        .Q(ID_EXEC_OUT[251]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_59_ ( .D(n19226), .CK(clk), .RN(n13882), .Q(MEM_WB_OUT[59]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_131_ ( .D(n7624), .CK(clk), .RN(
        n13905), .Q(EXEC_MEM_OUT_131), .QN(n11475) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_22_ ( .D(n7623), .CK(clk), .RN(n13889), 
        .QN(n19324) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_22_ ( .D(n19290), .CK(clk), .RN(
        n13900), .Q(MEM_WB_REG_MEM_WB_REG_N158) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_22_ ( .D(n19243), .CK(clk), .RN(n13884), .Q(MEM_WB_OUT[22]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_182_ ( .D(n7619), .CK(clk), .RN(n13895), 
        .Q(ID_EXEC_OUT[182]), .QN(n11528) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_164_ ( .D(n7618), .CK(clk), .RN(
        n13907), .Q(DMEM_BUS_OUT[54]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_86_ ( .D(n7617), .CK(clk), .RN(n13903), 
        .Q(ID_EXEC_OUT[86]), .QN(n11478) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_54_ ( .D(n7616), .CK(clk), .RN(n13920), 
        .Q(ID_EXEC_OUT[54]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_83_ ( .D(n7615), .CK(clk), .RN(
        n13898), .Q(DMEM_BUS_OUT[14]), .QN(n11968) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_51_ ( .D(n7614), .CK(clk), .RN(n13883), 
        .Q(MEM_WB_OUT[51]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_231_ ( .D(n7613), .CK(clk), .RN(
        n13900), .QN(n12160) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_218_ ( .D(n7611), .CK(clk), .RN(n13917), 
        .Q(ID_EXEC_OUT[218]), .QN(n11940) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_250_ ( .D(n7610), .CK(clk), .RN(n13907), 
        .Q(ID_EXEC_OUT[250]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_90_ ( .D(n7609), .CK(clk), .RN(
        n13924), .Q(DMEM_BUS_OUT[21]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_58_ ( .D(n19227), .CK(clk), .RN(n13930), .Q(MEM_WB_OUT[58]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_130_ ( .D(n7607), .CK(clk), .RN(
        n13905), .Q(EXEC_MEM_OUT_130) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_21_ ( .D(n7606), .CK(clk), .RN(n13923), 
        .QN(n19325) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_21_ ( .D(n7604), .CK(clk), .RN(
        n13909), .QN(n11105) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_21_ ( .D(n7603), .CK(clk), .RN(n13929), 
        .Q(MEM_WB_OUT[21]), .QN(n12547) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_181_ ( .D(n7602), .CK(clk), .RN(n13915), 
        .Q(ID_EXEC_OUT[181]), .QN(n11527) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_163_ ( .D(n7601), .CK(clk), .RN(
        n13903), .Q(DMEM_BUS_OUT[53]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_85_ ( .D(n7600), .CK(clk), .RN(n13921), 
        .Q(ID_EXEC_OUT[85]), .QN(n12521) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_53_ ( .D(n7599), .CK(clk), .RN(n13891), 
        .Q(ID_EXEC_OUT[53]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_82_ ( .D(n7598), .CK(clk), .RN(
        n13912), .Q(DMEM_BUS_OUT[13]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_50_ ( .D(n19233), .CK(clk), .RN(n13930), .Q(MEM_WB_OUT[50]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_230_ ( .D(n7596), .CK(clk), .RN(
        n13910), .QN(n12159) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_217_ ( .D(n7594), .CK(clk), .RN(n13894), 
        .Q(ID_EXEC_OUT[217]), .QN(n11945) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_249_ ( .D(n7593), .CK(clk), .RN(n13922), 
        .Q(ID_EXEC_OUT[249]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_72_ ( .D(n7592), .CK(clk), .RN(
        n13898), .Q(DMEM_BUS_OUT[3]), .QN(n11964) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_40_ ( .D(n19239), .CK(clk), .RN(n13883), .Q(MEM_WB_OUT[40]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_220_ ( .D(n7590), .CK(clk), .RN(
        n13901), .QN(n12149) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_207_ ( .D(n7588), .CK(clk), .RN(n13917), 
        .Q(ID_EXEC_OUT[207]), .QN(n11930) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_239_ ( .D(n7587), .CK(clk), .RN(n13928), 
        .Q(ID_EXEC_OUT[239]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_57_ ( .D(n19228), .CK(clk), .RN(n13882), .Q(MEM_WB_OUT[57]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_129_ ( .D(n7584), .CK(clk), .RN(
        n13904), .Q(EXEC_MEM_OUT_129) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_20_ ( .D(n7583), .CK(clk), .RN(n13889), 
        .QN(n19326) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_20_ ( .D(n19291), .CK(clk), .RN(
        n13901), .Q(MEM_WB_REG_MEM_WB_REG_N160) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_20_ ( .D(n19244), .CK(clk), .RN(n13884), .Q(MEM_WB_OUT[20]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_180_ ( .D(n7579), .CK(clk), .RN(n13895), 
        .Q(ID_EXEC_OUT[180]), .QN(n11526) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_162_ ( .D(n7578), .CK(clk), .RN(
        n13907), .Q(DMEM_BUS_OUT[52]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_84_ ( .D(n7577), .CK(clk), .RN(n13894), 
        .Q(ID_EXEC_OUT[84]), .QN(n12520) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_52_ ( .D(n7576), .CK(clk), .RN(n13920), 
        .Q(ID_EXEC_OUT[52]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_128_ ( .D(n7575), .CK(clk), .RN(
        n13905), .Q(EXEC_MEM_OUT_128) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_19_ ( .D(n7574), .CK(clk), .RN(n13889), 
        .QN(n12190) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_19_ ( .D(n7572), .CK(clk), .RN(
        n13902), .QN(n11113) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_19_ ( .D(n7571), .CK(clk), .RN(n13884), 
        .Q(MEM_WB_OUT[19]), .QN(n12546) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_179_ ( .D(n7570), .CK(clk), .RN(n13895), 
        .Q(ID_EXEC_OUT[179]), .QN(n11525) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_161_ ( .D(n7569), .CK(clk), .RN(
        n13903), .Q(DMEM_BUS_OUT[51]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_83_ ( .D(n7568), .CK(clk), .RN(n13921), 
        .Q(ID_EXEC_OUT[83]), .QN(n12519) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_51_ ( .D(n7567), .CK(clk), .RN(n13891), 
        .Q(ID_EXEC_OUT[51]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_18_ ( .D(n7566), .CK(clk), .RN(n13923), 
        .QN(n12187) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_18_ ( .D(n7564), .CK(clk), .RN(
        n13908), .QN(n11104) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_18_ ( .D(n7563), .CK(clk), .RN(n13928), 
        .Q(MEM_WB_OUT[18]), .QN(n12545) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_178_ ( .D(n7562), .CK(clk), .RN(n13915), 
        .Q(ID_EXEC_OUT[178]), .QN(n11524) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_160_ ( .D(n7561), .CK(clk), .RN(
        n13907), .Q(DMEM_BUS_OUT[50]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_82_ ( .D(n7560), .CK(clk), .RN(n13911), 
        .Q(ID_EXEC_OUT[82]), .QN(n12518) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_50_ ( .D(n7559), .CK(clk), .RN(n13920), 
        .Q(ID_EXEC_OUT[50]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_127_ ( .D(n7558), .CK(clk), .RN(
        n13904), .Q(EXEC_MEM_OUT_127) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_73_ ( .D(n7557), .CK(clk), .RN(
        n13911), .Q(DMEM_BUS_OUT[4]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_41_ ( .D(n19238), .CK(clk), .RN(n13930), .Q(MEM_WB_OUT[41]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_113_ ( .D(n7555), .CK(clk), .RN(
        n13912), .Q(EXEC_MEM_OUT_113), .QN(n12126) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_4_ ( .D(n7554), .CK(clk), .RN(n13888), 
        .QN(n19327) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_4_ ( .D(n7553), .CK(clk), .RN(n13891), 
        .Q(nextPC_ex_out[4]), .QN(n11914) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_4_ ( .D(n7552), .CK(clk), .RN(
        n13911), .Q(MEM_WB_REG_MEM_WB_REG_N176), .QN(n11550) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_4_ ( .D(n7551), .CK(clk), .RN(n13883), 
        .Q(MEM_WB_OUT[4]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_36_ ( .D(n7550), .CK(clk), .RN(n13919), 
        .Q(ID_EXEC_OUT[36]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_68_ ( .D(n7549), .CK(clk), .RN(n13890), 
        .Q(ID_EXEC_OUT[68]), .QN(n12516) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_164_ ( .D(n7548), .CK(clk), .RN(n13896), 
        .Q(ID_EXEC_OUT[164]), .QN(n11523) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_112_ ( .D(n7547), .CK(clk), .RN(
        n13904), .Q(EXEC_MEM_OUT_112), .QN(n12125) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_2_ ( .D(n7546), .CK(clk), .RN(n13889), 
        .QN(n12304) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_2_ ( .D(n7545), .CK(clk), .RN(n13892), 
        .Q(nextPC_ex_out[2]), .QN(n10358) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_2_ ( .D(n7544), .CK(clk), .RN(
        n13911), .Q(MEM_WB_REG_MEM_WB_REG_N178), .QN(n11548) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_2_ ( .D(n7543), .CK(clk), .RN(n13884), 
        .Q(MEM_WB_OUT[2]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_111_ ( .D(n7542), .CK(clk), .RN(
        n13916), .Q(EXEC_MEM_OUT_111), .QN(n12124) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_1_ ( .D(n7541), .CK(clk), .RN(n13923), 
        .QN(n12303) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_1_ ( .D(n7540), .CK(clk), .RN(n13894), 
        .Q(nextPC_ex_out[1]), .QN(n10362) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_1_ ( .D(n7539), .CK(clk), .RN(
        n13908), .Q(MEM_WB_REG_MEM_WB_REG_N179), .QN(n11547) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_1_ ( .D(n7538), .CK(clk), .RN(n13929), 
        .Q(MEM_WB_OUT[1]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_33_ ( .D(n7537), .CK(clk), .RN(n13892), 
        .Q(ID_EXEC_OUT[33]), .QN(n12206) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_65_ ( .D(n7536), .CK(clk), .RN(n13921), 
        .Q(ID_EXEC_OUT[65]), .QN(n12515) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_161_ ( .D(n7535), .CK(clk), .RN(n13915), 
        .Q(ID_EXEC_OUT[161]), .QN(n11522) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_218_ ( .D(n7534), .CK(clk), .RN(
        n13909), .QN(n12147) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_205_ ( .D(n7532), .CK(clk), .RN(n13917), 
        .Q(ID_EXEC_OUT[205]), .QN(n11939) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_237_ ( .D(n7531), .CK(clk), .RN(n13927), 
        .Q(ID_EXEC_OUT[237]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_86_ ( .D(n7530), .CK(clk), .RN(
        n13912), .Q(DMEM_BUS_OUT[17]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_54_ ( .D(n19231), .CK(clk), .RN(n13930), .Q(MEM_WB_OUT[54]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_126_ ( .D(n7528), .CK(clk), .RN(
        n13905), .Q(EXEC_MEM_OUT_126) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_17_ ( .D(n7527), .CK(clk), .RN(n13889), 
        .QN(n12186) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_17_ ( .D(n7526), .CK(clk), .RN(n13915), 
        .Q(nextPC_ex_out[17]), .QN(n11995) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_17_ ( .D(net139967), .CK(clk), 
        .RN(n13902), .Q(MEM_WB_REG_MEM_WB_REG_N163) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_17_ ( .D(n19245), .CK(clk), .RN(n13884), .Q(MEM_WB_OUT[17]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_49_ ( .D(n7523), .CK(clk), .RN(n13920), 
        .Q(ID_EXEC_OUT[49]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_81_ ( .D(n7522), .CK(clk), .RN(n13921), 
        .Q(ID_EXEC_OUT[81]), .QN(n12517) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_177_ ( .D(n7521), .CK(clk), .RN(n13895), 
        .Q(ID_EXEC_OUT[177]), .QN(n11521) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_159_ ( .D(n7520), .CK(clk), .RN(
        n13907), .Q(DMEM_BUS_OUT[49]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_78_ ( .D(n7519), .CK(clk), .RN(
        n13898), .Q(DMEM_BUS_OUT[9]), .QN(n11977) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_46_ ( .D(n19236), .CK(clk), .RN(n13883), .Q(MEM_WB_OUT[46]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_118_ ( .D(n7517), .CK(clk), .RN(
        n13904), .Q(EXEC_MEM_OUT_118), .QN(n10946) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_9_ ( .D(n7516), .CK(clk), .RN(n13925), 
        .QN(net137185) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_9_ ( .D(n7515), .CK(clk), .RN(n13922), 
        .Q(nextPC_ex_out[9]), .QN(n11920) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_9_ ( .D(n7514), .CK(clk), .RN(
        n13895), .Q(MEM_WB_REG_MEM_WB_REG_N171), .QN(n11540) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_9_ ( .D(n7513), .CK(clk), .RN(n13932), 
        .Q(MEM_WB_OUT[9]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_41_ ( .D(n7512), .CK(clk), .RN(n13919), 
        .Q(ID_EXEC_OUT[41]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_73_ ( .D(n7511), .CK(clk), .RN(n13890), 
        .Q(ID_EXEC_OUT[73]), .QN(n12514) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_169_ ( .D(n7510), .CK(clk), .RN(n13915), 
        .Q(ID_EXEC_OUT[169]), .QN(n11520) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_117_ ( .D(n7509), .CK(clk), .RN(
        n13905), .Q(EXEC_MEM_OUT_117) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_8_ ( .D(n7508), .CK(clk), .RN(n13887), 
        .QN(n12196) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_8_ ( .D(n7507), .CK(clk), .RN(n13884), 
        .Q(nextPC_ex_out[8]), .QN(n10357) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_8_ ( .D(n7506), .CK(clk), .RN(
        n13912), .Q(MEM_WB_REG_MEM_WB_REG_N172), .QN(n11554) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_8_ ( .D(n7505), .CK(clk), .RN(n13881), 
        .Q(MEM_WB_OUT[8]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_116_ ( .D(n7504), .CK(clk), .RN(
        n13904), .Q(EXEC_MEM_OUT_116) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_6_ ( .D(n7503), .CK(clk), .RN(n13887), 
        .QN(n12194) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_6_ ( .D(n7502), .CK(clk), .RN(n13890), 
        .Q(nextPC_ex_out[6]), .QN(n10356) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_6_ ( .D(n7501), .CK(clk), .RN(
        n13911), .Q(MEM_WB_REG_MEM_WB_REG_N174), .QN(n11552) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_6_ ( .D(n7500), .CK(clk), .RN(n13882), 
        .Q(MEM_WB_OUT[6]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_115_ ( .D(n7499), .CK(clk), .RN(
        n13905), .Q(EXEC_MEM_OUT_115), .QN(n12123) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_5_ ( .D(n7498), .CK(clk), .RN(n13924), 
        .QN(n12193) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_5_ ( .D(n7497), .CK(clk), .RN(n13920), 
        .Q(nextPC_ex_out[5]), .QN(n10355) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_5_ ( .D(n7496), .CK(clk), .RN(
        n13899), .Q(MEM_WB_REG_MEM_WB_REG_N175), .QN(n11551) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_5_ ( .D(n7495), .CK(clk), .RN(n13930), 
        .Q(MEM_WB_OUT[5]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_114_ ( .D(n7494), .CK(clk), .RN(
        n13904), .Q(EXEC_MEM_OUT_114) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_3_ ( .D(n7493), .CK(clk), .RN(n13924), 
        .QN(n12305) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_3_ ( .D(n7491), .CK(clk), .RN(
        n13899), .Q(MEM_WB_REG_MEM_WB_REG_N177), .QN(n11549) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_3_ ( .D(n7490), .CK(clk), .RN(n13929), 
        .Q(MEM_WB_OUT[3]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_35_ ( .D(n7489), .CK(clk), .RN(n13892), 
        .Q(ID_EXEC_OUT[35]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_67_ ( .D(n7488), .CK(clk), .RN(n13921), 
        .Q(ID_EXEC_OUT[67]), .QN(n12513) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_163_ ( .D(n7487), .CK(clk), .RN(n13915), 
        .Q(ID_EXEC_OUT[163]), .QN(n11519) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_71_ ( .D(n19149), .CK(clk), .RN(
        n13911), .Q(DMEM_BUS_OUT[2]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_39_ ( .D(n19240), .CK(clk), .RN(n13883), .Q(MEM_WB_OUT[39]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_34_ ( .D(n7484), .CK(clk), .RN(n13919), 
        .Q(ID_EXEC_OUT[34]), .QN(n12541) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_66_ ( .D(n7483), .CK(clk), .RN(n13890), 
        .Q(ID_EXEC_OUT[66]), .QN(n12512) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_162_ ( .D(n7482), .CK(clk), .RN(n13896), 
        .Q(ID_EXEC_OUT[162]), .QN(n11518) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_219_ ( .D(n7481), .CK(clk), .RN(
        n13901), .QN(n12148) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_206_ ( .D(n7479), .CK(clk), .RN(n13894), 
        .Q(ID_EXEC_OUT[206]), .QN(n11943) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_238_ ( .D(n7478), .CK(clk), .RN(n13918), 
        .Q(ID_EXEC_OUT[238]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_53_ ( .D(n7476), .CK(clk), .RN(n13883), 
        .Q(MEM_WB_OUT[53]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_125_ ( .D(n7475), .CK(clk), .RN(
        n13904), .Q(EXEC_MEM_OUT_125) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_16_ ( .D(n7474), .CK(clk), .RN(n13922), 
        .QN(n12185) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_16_ ( .D(n7473), .CK(clk), .RN(n13896), 
        .Q(nextPC_ex_out[16]), .QN(n11928) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_16_ ( .D(n7472), .CK(clk), .RN(
        n13907), .QN(n11103) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_16_ ( .D(n7471), .CK(clk), .RN(n13885), 
        .Q(MEM_WB_OUT[16]), .QN(n12223) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_48_ ( .D(n7470), .CK(clk), .RN(n13891), 
        .Q(ID_EXEC_OUT[48]), .QN(n12131) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_80_ ( .D(n7469), .CK(clk), .RN(n13883), 
        .Q(ID_EXEC_OUT[80]), .QN(n12320) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_176_ ( .D(n7468), .CK(clk), .RN(n13915), 
        .Q(ID_EXEC_OUT[176]), .QN(n11517) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_158_ ( .D(n7467), .CK(clk), .RN(
        n13903), .Q(DMEM_BUS_OUT[48]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_124_ ( .D(n7466), .CK(clk), .RN(
        n13905), .Q(EXEC_MEM_OUT_124), .QN(n11474) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_15_ ( .D(n7465), .CK(clk), .RN(n13889), 
        .QN(n12189) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_15_ ( .D(n7464), .CK(clk), .RN(n13914), 
        .Q(nextPC_ex_out[15]), .QN(n11955) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_15_ ( .D(n7463), .CK(clk), .RN(
        n13903), .Q(MEM_WB_REG_MEM_WB_REG_N165), .QN(n11546) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_47_ ( .D(n7461), .CK(clk), .RN(n13920), 
        .Q(ID_EXEC_OUT[47]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_79_ ( .D(n7460), .CK(clk), .RN(n13890), 
        .Q(ID_EXEC_OUT[79]), .QN(n12511) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_175_ ( .D(n7459), .CK(clk), .RN(n13896), 
        .Q(ID_EXEC_OUT[175]), .QN(n11516) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_157_ ( .D(n7458), .CK(clk), .RN(
        n13906), .Q(DMEM_BUS_OUT[47]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_14_ ( .D(n7457), .CK(clk), .RN(n13922), 
        .QN(n19328) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_14_ ( .D(n7456), .CK(clk), .RN(n13897), 
        .Q(nextPC_ex_out[14]), .QN(n11993) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_14_ ( .D(n7455), .CK(clk), .RN(
        n13906), .Q(MEM_WB_REG_MEM_WB_REG_N166), .QN(n11541) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_14_ ( .D(n7454), .CK(clk), .RN(n13886), 
        .Q(MEM_WB_OUT[14]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_46_ ( .D(n7453), .CK(clk), .RN(n13891), 
        .Q(ID_EXEC_OUT[46]), .QN(n12210) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_78_ ( .D(n7452), .CK(clk), .RN(n13921), 
        .Q(ID_EXEC_OUT[78]), .QN(n12510) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_174_ ( .D(n7451), .CK(clk), .RN(n13915), 
        .Q(ID_EXEC_OUT[174]), .QN(n11515) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_156_ ( .D(n7450), .CK(clk), .RN(
        n13903), .Q(DMEM_BUS_OUT[46]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_123_ ( .D(n7449), .CK(clk), .RN(
        n13904), .Q(EXEC_MEM_OUT_123) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_13_ ( .D(n7448), .CK(clk), .RN(n13889), 
        .QN(n19329) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_13_ ( .D(n7447), .CK(clk), .RN(n13914), 
        .Q(nextPC_ex_out[13]), .QN(n11934) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_13_ ( .D(n7446), .CK(clk), .RN(
        n13889), .Q(MEM_WB_REG_MEM_WB_REG_N167), .QN(n11539) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_13_ ( .D(n7445), .CK(clk), .RN(n13927), 
        .Q(MEM_WB_OUT[13]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_45_ ( .D(n7444), .CK(clk), .RN(n13920), 
        .Q(ID_EXEC_OUT[45]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_77_ ( .D(n7443), .CK(clk), .RN(n13890), 
        .Q(ID_EXEC_OUT[77]), .QN(n12509) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_173_ ( .D(n7442), .CK(clk), .RN(n13896), 
        .Q(ID_EXEC_OUT[173]), .QN(n11514) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_155_ ( .D(n7441), .CK(clk), .RN(
        n13906), .Q(DMEM_BUS_OUT[45]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_122_ ( .D(n7440), .CK(clk), .RN(
        n13905), .Q(EXEC_MEM_OUT_122) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_233_ ( .D(n7439), .CK(clk), .RN(
        n13900), .QN(n12162) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_220_ ( .D(n7437), .CK(clk), .RN(n13917), 
        .Q(ID_EXEC_OUT[220]), .QN(n10813) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_252_ ( .D(n7436), .CK(clk), .RN(n13901), 
        .Q(ID_EXEC_OUT[252]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_81_ ( .D(n7435), .CK(clk), .RN(
        n13898), .Q(DMEM_BUS_OUT[12]), .QN(n11987) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_49_ ( .D(n7434), .CK(clk), .RN(n13930), 
        .Q(MEM_WB_OUT[49]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_121_ ( .D(n7433), .CK(clk), .RN(
        n13904), .Q(EXEC_MEM_OUT_121) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_12_ ( .D(n7432), .CK(clk), .RN(n13922), 
        .QN(n12188) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_12_ ( .D(n7431), .CK(clk), .RN(n13907), 
        .Q(nextPC_ex_out[12]), .QN(n11921) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_12_ ( .D(n7430), .CK(clk), .RN(
        n13905), .Q(MEM_WB_REG_MEM_WB_REG_N168), .QN(n11545) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_12_ ( .D(n7429), .CK(clk), .RN(n13894), 
        .Q(MEM_WB_OUT[12]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_44_ ( .D(n7428), .CK(clk), .RN(n13891), 
        .Q(ID_EXEC_OUT[44]), .QN(n12209) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_76_ ( .D(n7427), .CK(clk), .RN(n13921), 
        .Q(ID_EXEC_OUT[76]), .QN(n12508) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_172_ ( .D(n7426), .CK(clk), .RN(n13915), 
        .Q(ID_EXEC_OUT[172]), .QN(n11513) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_154_ ( .D(n7425), .CK(clk), .RN(
        n13903), .Q(DMEM_BUS_OUT[44]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_120_ ( .D(n7424), .CK(clk), .RN(
        n13905), .Q(EXEC_MEM_OUT_120), .QN(n11473) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_11_ ( .D(n7423), .CK(clk), .RN(n13889), 
        .QN(n19330) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_11_ ( .D(n7422), .CK(clk), .RN(n13913), 
        .Q(nextPC_ex_out[11]), .QN(n12018) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_11_ ( .D(n7421), .CK(clk), .RN(
        n13904), .Q(MEM_WB_REG_MEM_WB_REG_N169), .QN(n11538) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_11_ ( .D(n7420), .CK(clk), .RN(n13926), 
        .Q(MEM_WB_OUT[11]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_10_ ( .D(n7419), .CK(clk), .RN(n13922), 
        .QN(n19331) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_10_ ( .D(n7418), .CK(clk), .RN(n13882), 
        .Q(nextPC_ex_out[10]), .QN(n11919) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_10_ ( .D(n7417), .CK(clk), .RN(
        n13881), .Q(MEM_WB_REG_MEM_WB_REG_N170), .QN(n11544) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_10_ ( .D(n7416), .CK(clk), .RN(n13929), 
        .Q(MEM_WB_OUT[10]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_119_ ( .D(n7415), .CK(clk), .RN(
        n13905), .Q(EXEC_MEM_OUT_119) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_7_ ( .D(n7414), .CK(clk), .RN(n13925), 
        .QN(n12195) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_7_ ( .D(n7413), .CK(clk), .RN(n13921), 
        .Q(nextPC_ex_out[7]), .QN(n10366) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_7_ ( .D(n7412), .CK(clk), .RN(
        n13898), .Q(MEM_WB_REG_MEM_WB_REG_N173), .QN(n11553) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_7_ ( .D(n7411), .CK(clk), .RN(n13931), 
        .Q(MEM_WB_OUT[7]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_39_ ( .D(n7410), .CK(clk), .RN(n13891), 
        .Q(ID_EXEC_OUT[39]), .QN(n12179) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_71_ ( .D(n7409), .CK(clk), .RN(n13890), 
        .Q(ID_EXEC_OUT[71]), .QN(n12507) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_167_ ( .D(n7408), .CK(clk), .RN(n13915), 
        .Q(ID_EXEC_OUT[167]), .QN(n11512) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_224_ ( .D(n7407), .CK(clk), .RN(
        n13900), .QN(n12153) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_211_ ( .D(n7405), .CK(clk), .RN(n13894), 
        .Q(ID_EXEC_OUT[211]), .QN(n11957) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_243_ ( .D(n7404), .CK(clk), .RN(n13918), 
        .Q(ID_EXEC_OUT[243]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_48_ ( .D(n19234), .CK(clk), .RN(n13883), .Q(MEM_WB_OUT[48]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_43_ ( .D(n7401), .CK(clk), .RN(n13920), 
        .Q(ID_EXEC_OUT[43]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_75_ ( .D(n7400), .CK(clk), .RN(n13890), 
        .Q(ID_EXEC_OUT[75]), .QN(n12506) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_171_ ( .D(n7399), .CK(clk), .RN(n13896), 
        .Q(ID_EXEC_OUT[171]), .QN(n11511) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_153_ ( .D(n7398), .CK(clk), .RN(
        n13906), .Q(DMEM_BUS_OUT[43]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_228_ ( .D(n7397), .CK(clk), .RN(
        n13900), .QN(n12157) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_215_ ( .D(n7395), .CK(clk), .RN(n13894), 
        .Q(ID_EXEC_OUT[215]), .QN(n11942) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_247_ ( .D(n7394), .CK(clk), .RN(n13918), 
        .Q(ID_EXEC_OUT[247]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_79_ ( .D(n7393), .CK(clk), .RN(
        n13912), .Q(DMEM_BUS_OUT[10]), .QN(n11966) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_47_ ( .D(n19235), .CK(clk), .RN(n13930), .Q(MEM_WB_OUT[47]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_42_ ( .D(n7391), .CK(clk), .RN(n13891), 
        .Q(ID_EXEC_OUT[42]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_74_ ( .D(n7390), .CK(clk), .RN(n13921), 
        .Q(ID_EXEC_OUT[74]), .QN(n12505) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_170_ ( .D(n7389), .CK(clk), .RN(n13915), 
        .Q(ID_EXEC_OUT[170]), .QN(n11510) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_152_ ( .D(n7388), .CK(clk), .RN(
        n13903), .Q(DMEM_BUS_OUT[42]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_227_ ( .D(n7387), .CK(clk), .RN(
        n13909), .QN(n12156) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_214_ ( .D(n7385), .CK(clk), .RN(n13917), 
        .Q(ID_EXEC_OUT[214]), .QN(n11958) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_246_ ( .D(n7384), .CK(clk), .RN(n13893), 
        .Q(ID_EXEC_OUT[246]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_77_ ( .D(n7383), .CK(clk), .RN(
        n13912), .Q(DMEM_BUS_OUT[8]), .QN(n11986) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_45_ ( .D(n7382), .CK(clk), .RN(n13930), 
        .Q(MEM_WB_OUT[45]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_40_ ( .D(n7381), .CK(clk), .RN(n13891), 
        .Q(ID_EXEC_OUT[40]), .QN(n12208) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_72_ ( .D(n7380), .CK(clk), .RN(n13921), 
        .Q(ID_EXEC_OUT[72]), .QN(n12504) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_168_ ( .D(n7379), .CK(clk), .RN(n13896), 
        .Q(ID_EXEC_OUT[168]), .QN(n11509) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_225_ ( .D(n7378), .CK(clk), .RN(
        n13909), .QN(n12154) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_212_ ( .D(n7376), .CK(clk), .RN(n13917), 
        .Q(ID_EXEC_OUT[212]), .QN(n10820) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_244_ ( .D(n7375), .CK(clk), .RN(n13893), 
        .Q(ID_EXEC_OUT[244]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_75_ ( .D(n7374), .CK(clk), .RN(
        n13912), .Q(DMEM_BUS_OUT[6]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_43_ ( .D(n19237), .CK(clk), .RN(n13930), .Q(MEM_WB_OUT[43]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_38_ ( .D(n7372), .CK(clk), .RN(n13919), 
        .Q(ID_EXEC_OUT[38]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_70_ ( .D(n7371), .CK(clk), .RN(n13921), 
        .Q(ID_EXEC_OUT[70]), .QN(n12503) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_166_ ( .D(n7370), .CK(clk), .RN(n13896), 
        .Q(ID_EXEC_OUT[166]), .QN(n11508) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_76_ ( .D(n7369), .CK(clk), .RN(
        n13898), .Q(DMEM_BUS_OUT[7]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_44_ ( .D(n7368), .CK(clk), .RN(n13883), 
        .Q(MEM_WB_OUT[44]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_74_ ( .D(n7367), .CK(clk), .RN(
        n13898), .Q(DMEM_BUS_OUT[5]), .QN(n11967) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_42_ ( .D(n7366), .CK(clk), .RN(n13883), 
        .Q(MEM_WB_OUT[42]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_37_ ( .D(n7365), .CK(clk), .RN(n13891), 
        .Q(ID_EXEC_OUT[37]), .QN(n12207) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_69_ ( .D(n7364), .CK(clk), .RN(n13921), 
        .Q(ID_EXEC_OUT[69]), .QN(n12502) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_165_ ( .D(n7363), .CK(clk), .RN(n13915), 
        .Q(ID_EXEC_OUT[165]), .QN(n11507) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_222_ ( .D(n7362), .CK(clk), .RN(
        n13900), .QN(n12151) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_209_ ( .D(n7360), .CK(clk), .RN(n13917), 
        .Q(ID_EXEC_OUT[209]), .QN(n11931) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_241_ ( .D(n7359), .CK(clk), .RN(n13918), 
        .Q(ID_EXEC_OUT[241]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_147_ ( .D(n7358), .CK(clk), .RN(
        n13908), .Q(DMEM_BUS_OUT[37]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_149_ ( .D(n7357), .CK(clk), .RN(
        n13906), .Q(DMEM_BUS_OUT[39]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_223_ ( .D(n7356), .CK(clk), .RN(
        n13909), .QN(n12152) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_210_ ( .D(n7354), .CK(clk), .RN(n13917), 
        .Q(ID_EXEC_OUT[210]), .QN(n11941) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_242_ ( .D(n7353), .CK(clk), .RN(n13893), 
        .Q(ID_EXEC_OUT[242]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_148_ ( .D(n7352), .CK(clk), .RN(
        n13906), .Q(DMEM_BUS_OUT[38]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_150_ ( .D(n7351), .CK(clk), .RN(
        n13907), .Q(DMEM_BUS_OUT[40]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_229_ ( .D(n7350), .CK(clk), .RN(
        n13910), .QN(n12158) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_216_ ( .D(n7348), .CK(clk), .RN(n13917), 
        .Q(ID_EXEC_OUT[216]), .QN(n10821) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_248_ ( .D(n7347), .CK(clk), .RN(n13893), 
        .Q(ID_EXEC_OUT[248]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_144_ ( .D(n7346), .CK(clk), .RN(
        n13906), .Q(DMEM_BUS_OUT[34]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_226_ ( .D(n7345), .CK(clk), .RN(
        n13900), .QN(n12155) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_213_ ( .D(n7343), .CK(clk), .RN(n13894), 
        .Q(ID_EXEC_OUT[213]), .QN(n11961) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_245_ ( .D(n7342), .CK(clk), .RN(n13918), 
        .Q(ID_EXEC_OUT[245]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_151_ ( .D(n7341), .CK(clk), .RN(
        n13906), .Q(DMEM_BUS_OUT[41]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_234_ ( .D(n7340), .CK(clk), .RN(
        n13910), .QN(n12163) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_221_ ( .D(n7338), .CK(clk), .RN(n13917), 
        .Q(ID_EXEC_OUT[221]), .QN(n11935) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_253_ ( .D(n7337), .CK(clk), .RN(n13893), 
        .Q(ID_EXEC_OUT[253]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_70_ ( .D(n19150), .CK(clk), .RN(
        n13898), .Q(DMEM_BUS_OUT[1]), .QN(n10826) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_38_ ( .D(n7335), .CK(clk), .RN(n13929), 
        .Q(MEM_WB_OUT[38]), .QN(n12180) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_143_ ( .D(n7334), .CK(clk), .RN(
        n13910), .Q(DMEM_BUS_OUT[33]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_110_ ( .D(n7333), .CK(clk), .RN(
        n13904), .Q(EXEC_MEM_OUT_110), .QN(n12122) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_0_ ( .D(n7331), .CK(clk), .RN(n13888), 
        .Q(nextPC_ex_out[0]), .QN(n10243) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_0_ ( .D(n7330), .CK(clk), .RN(
        n13929), .QN(n11112) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_0_ ( .D(n7329), .CK(clk), .RN(n13887), 
        .Q(MEM_WB_OUT[0]), .QN(n12534) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_32_ ( .D(n7328), .CK(clk), .RN(n13919), 
        .Q(ID_EXEC_OUT[32]), .QN(n12229) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_64_ ( .D(n7327), .CK(clk), .RN(n13890), 
        .Q(ID_EXEC_OUT[64]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_160_ ( .D(n7326), .CK(clk), .RN(n13896), 
        .Q(ID_EXEC_OUT[160]), .QN(n11506) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_109_ ( .D(n7325), .CK(clk), .RN(
        n13904), .Q(EXEC_MEM_OUT_109) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_221_ ( .D(n7324), .CK(clk), .RN(
        n13909), .QN(n12150) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_208_ ( .D(n7322), .CK(clk), .RN(n13894), 
        .Q(ID_EXEC_OUT[208]), .QN(n11944) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_240_ ( .D(n7321), .CK(clk), .RN(n13930), 
        .Q(ID_EXEC_OUT[240]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_146_ ( .D(n7320), .CK(clk), .RN(
        n13906), .Q(DMEM_BUS_OUT[36]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_237_ ( .D(n7319), .CK(clk), .RN(
        n13900), .QN(n12166) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_224_ ( .D(n7317), .CK(clk), .RN(n13922), 
        .Q(ID_EXEC_OUT[224]), .QN(n10812) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_256_ ( .D(n7316), .CK(clk), .RN(n13904), 
        .Q(ID_EXEC_OUT[256]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_145_ ( .D(n7315), .CK(clk), .RN(
        n13909), .Q(DMEM_BUS_OUT[35]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_238_ ( .D(n7314), .CK(clk), .RN(
        n13910), .QN(n12167) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_225_ ( .D(n7312), .CK(clk), .RN(n13917), 
        .Q(ID_EXEC_OUT[225]), .QN(n11956) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_257_ ( .D(n7311), .CK(clk), .RN(n13893), 
        .Q(ID_EXEC_OUT[257]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_239_ ( .D(n7310), .CK(clk), .RN(
        n13900), .QN(n12168) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_226_ ( .D(n7308), .CK(clk), .RN(n13921), 
        .Q(ID_EXEC_OUT[226]), .QN(n10818) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_258_ ( .D(n7307), .CK(clk), .RN(n13921), 
        .Q(ID_EXEC_OUT[258]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_236_ ( .D(n7306), .CK(clk), .RN(
        n13910), .QN(n12165) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_223_ ( .D(n7304), .CK(clk), .RN(n13917), 
        .Q(ID_EXEC_OUT[223]), .QN(n11959) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_255_ ( .D(n7303), .CK(clk), .RN(n13893), 
        .Q(ID_EXEC_OUT[255]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_240_ ( .D(n7302), .CK(clk), .RN(
        n13900), .QN(n12169) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_227_ ( .D(n7300), .CK(clk), .RN(n13918), 
        .Q(ID_EXEC_OUT[227]), .QN(n11932) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_259_ ( .D(n7299), .CK(clk), .RN(n13893), 
        .Q(ID_EXEC_OUT[259]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_241_ ( .D(n7298), .CK(clk), .RN(
        n13910), .QN(n12170) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_228_ ( .D(n7296), .CK(clk), .RN(n13920), 
        .Q(ID_EXEC_OUT[228]), .QN(n10811) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_260_ ( .D(n7295), .CK(clk), .RN(n13893), 
        .Q(ID_EXEC_OUT[260]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_142_ ( .D(n7294), .CK(clk), .RN(
        n13906), .Q(DMEM_BUS_OUT[32]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_236_ ( .D(n7293), .CK(clk), .RN(n13918), 
        .Q(ID_EXEC_OUT[236]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_267_ ( .D(n7292), .CK(clk), .RN(n13900), 
        .Q(ID_EXEC_OUT[267]) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10291) );
  DFF_X2 EXEC_STAGE_mul_ex_CurrentState_reg_2_ ( .D(EXEC_STAGE_mul_ex_N14), 
        .CK(clk), .Q(EXEC_STAGE_mul_ex_CurrentState_2_) );
  DFF_X2 EXEC_STAGE_mul_ex_CurrentState_reg_1_ ( .D(EXEC_STAGE_mul_ex_N15), 
        .CK(clk), .Q(EXEC_STAGE_mul_ex_CurrentState_1_), .QN(n10543) );
  DFF_X2 EXEC_STAGE_mul_ex_CurrentState_reg_0_ ( .D(EXEC_STAGE_mul_ex_N16), 
        .CK(clk), .Q(EXEC_STAGE_mul_ex_CurrentState_0_), .QN(n10159) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_0_ ( .G(n13544), .D(
        EXEC_STAGE_mul_ex_N377), .Q(EXEC_STAGE_mul_result_long[0]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_1_ ( .G(n13544), .D(
        EXEC_STAGE_mul_ex_N376), .Q(EXEC_STAGE_mul_result_long[1]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_2_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N375), .Q(EXEC_STAGE_mul_result_long[2]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_3_ ( .G(n10106), .D(
        EXEC_STAGE_mul_ex_N374), .Q(EXEC_STAGE_mul_result_long[3]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_4_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N373), .Q(EXEC_STAGE_mul_result_long[4]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_5_ ( .G(n10106), .D(
        EXEC_STAGE_mul_ex_N372), .Q(EXEC_STAGE_mul_result_long[5]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_6_ ( .G(n10106), .D(
        EXEC_STAGE_mul_ex_N371), .Q(EXEC_STAGE_mul_result_long[6]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_7_ ( .G(n10106), .D(
        EXEC_STAGE_mul_ex_N370), .Q(EXEC_STAGE_mul_result_long[7]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_8_ ( .G(n13544), .D(
        EXEC_STAGE_mul_ex_N369), .Q(EXEC_STAGE_mul_result_long[8]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_9_ ( .G(n10106), .D(
        EXEC_STAGE_mul_ex_N368), .Q(EXEC_STAGE_mul_result_long[9]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_10_ ( .G(n10106), .D(
        EXEC_STAGE_mul_ex_N367), .Q(EXEC_STAGE_mul_result_long[10]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_11_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N366), .Q(EXEC_STAGE_mul_result_long[11]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_12_ ( .G(n13544), .D(
        EXEC_STAGE_mul_ex_N365), .Q(EXEC_STAGE_mul_result_long[12]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_13_ ( .G(n10106), .D(
        EXEC_STAGE_mul_ex_N364), .Q(EXEC_STAGE_mul_result_long[13]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_14_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N363), .Q(EXEC_STAGE_mul_result_long[14]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_15_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N362), .Q(EXEC_STAGE_mul_result_long[15]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_16_ ( .G(n10106), .D(
        EXEC_STAGE_mul_ex_N361), .Q(EXEC_STAGE_mul_result_long[16]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_17_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N360), .Q(EXEC_STAGE_mul_result_long[17]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_18_ ( .G(n10106), .D(
        EXEC_STAGE_mul_ex_N359), .Q(EXEC_STAGE_mul_result_long[18]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_19_ ( .G(n13544), .D(
        EXEC_STAGE_mul_ex_N358), .Q(EXEC_STAGE_mul_result_long[19]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_20_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N357), .Q(EXEC_STAGE_mul_result_long[20]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_21_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N356), .Q(EXEC_STAGE_mul_result_long[21]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_22_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N355), .Q(EXEC_STAGE_mul_result_long[22]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_23_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N354), .Q(EXEC_STAGE_mul_result_long[23]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_24_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N353), .Q(EXEC_STAGE_mul_result_long[24]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_25_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N352), .Q(EXEC_STAGE_mul_result_long[25]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_26_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N351), .Q(EXEC_STAGE_mul_result_long[26]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_27_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N350), .Q(EXEC_STAGE_mul_result_long[27]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_28_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N349), .Q(EXEC_STAGE_mul_result_long[28]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_29_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N348), .Q(EXEC_STAGE_mul_result_long[29]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_30_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N347), .Q(EXEC_STAGE_mul_result_long[30]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_31_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N346), .Q(EXEC_STAGE_mul_result_long[31]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_32_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N345), .Q(EXEC_STAGE_mul_result_long[32]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_33_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N344), .Q(EXEC_STAGE_mul_result_long[33]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_34_ ( .G(n10106), .D(
        EXEC_STAGE_mul_ex_N343), .Q(EXEC_STAGE_mul_result_long[34]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_35_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N342), .Q(EXEC_STAGE_mul_result_long[35]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_36_ ( .G(n10106), .D(
        EXEC_STAGE_mul_ex_N341), .Q(EXEC_STAGE_mul_result_long[36]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_37_ ( .G(n10106), .D(
        EXEC_STAGE_mul_ex_N340), .Q(EXEC_STAGE_mul_result_long[37]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_38_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N339), .Q(EXEC_STAGE_mul_result_long[38]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_39_ ( .G(n10106), .D(
        EXEC_STAGE_mul_ex_N338), .Q(EXEC_STAGE_mul_result_long[39]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_40_ ( .G(n13544), .D(
        EXEC_STAGE_mul_ex_N337), .Q(EXEC_STAGE_mul_result_long[40]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_41_ ( .G(n10106), .D(
        EXEC_STAGE_mul_ex_N336), .Q(EXEC_STAGE_mul_result_long[41]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_42_ ( .G(n13546), .D(
        EXEC_STAGE_mul_ex_N335), .Q(EXEC_STAGE_mul_result_long[42]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_43_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N334), .Q(EXEC_STAGE_mul_result_long[43]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_44_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N333), .Q(EXEC_STAGE_mul_result_long[44]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_45_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N332), .Q(EXEC_STAGE_mul_result_long[45]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_46_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N331), .Q(EXEC_STAGE_mul_result_long[46]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_47_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N330), .Q(EXEC_STAGE_mul_result_long[47]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_48_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N329), .Q(EXEC_STAGE_mul_result_long[48]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_49_ ( .G(n10106), .D(
        EXEC_STAGE_mul_ex_N328), .Q(EXEC_STAGE_mul_result_long[49]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_50_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N327), .Q(EXEC_STAGE_mul_result_long[50]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_51_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N326), .Q(EXEC_STAGE_mul_result_long[51]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_52_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N325), .Q(EXEC_STAGE_mul_result_long[52]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_53_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N324), .Q(EXEC_STAGE_mul_result_long[53]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_54_ ( .G(n13545), .D(
        EXEC_STAGE_mul_ex_N323), .Q(EXEC_STAGE_mul_result_long[54]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_55_ ( .G(n13544), .D(
        EXEC_STAGE_mul_ex_N322), .Q(EXEC_STAGE_mul_result_long[55]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_56_ ( .G(n13544), .D(
        EXEC_STAGE_mul_ex_N321), .Q(EXEC_STAGE_mul_result_long[56]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_57_ ( .G(n13544), .D(
        EXEC_STAGE_mul_ex_N320), .Q(EXEC_STAGE_mul_result_long[57]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_58_ ( .G(n13544), .D(
        EXEC_STAGE_mul_ex_N319), .Q(EXEC_STAGE_mul_result_long[58]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_59_ ( .G(n13544), .D(
        EXEC_STAGE_mul_ex_N318), .Q(EXEC_STAGE_mul_result_long[59]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_60_ ( .G(n13544), .D(
        EXEC_STAGE_mul_ex_N317), .Q(EXEC_STAGE_mul_result_long[60]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_61_ ( .G(n13544), .D(
        EXEC_STAGE_mul_ex_N316), .Q(EXEC_STAGE_mul_result_long[61]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_62_ ( .G(n13544), .D(
        EXEC_STAGE_mul_ex_N315), .Q(EXEC_STAGE_mul_result_long[62]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_63_ ( .G(n13544), .D(
        EXEC_STAGE_mul_ex_N314), .Q(EXEC_STAGE_mul_result_long[63]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_31_ ( .G(n13542), .D(EXEC_STAGE_mul_ex_N56), 
        .Q(EXEC_STAGE_mul_ex_H[31]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_30_ ( .G(n13542), .D(EXEC_STAGE_mul_ex_N57), 
        .Q(EXEC_STAGE_mul_ex_H[30]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_29_ ( .G(n13542), .D(EXEC_STAGE_mul_ex_N58), 
        .Q(EXEC_STAGE_mul_ex_H[29]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_28_ ( .G(n13542), .D(EXEC_STAGE_mul_ex_N59), 
        .Q(EXEC_STAGE_mul_ex_H[28]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_27_ ( .G(n13542), .D(EXEC_STAGE_mul_ex_N60), 
        .Q(EXEC_STAGE_mul_ex_H[27]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_26_ ( .G(n13542), .D(EXEC_STAGE_mul_ex_N61), 
        .Q(EXEC_STAGE_mul_ex_H[26]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_25_ ( .G(n13542), .D(EXEC_STAGE_mul_ex_N62), 
        .Q(EXEC_STAGE_mul_ex_H[25]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_24_ ( .G(n13542), .D(EXEC_STAGE_mul_ex_N63), 
        .Q(EXEC_STAGE_mul_ex_H[24]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_23_ ( .G(n13542), .D(EXEC_STAGE_mul_ex_N64), 
        .Q(EXEC_STAGE_mul_ex_H[23]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_22_ ( .G(n13542), .D(EXEC_STAGE_mul_ex_N65), 
        .Q(EXEC_STAGE_mul_ex_H[22]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_21_ ( .G(n13542), .D(EXEC_STAGE_mul_ex_N66), 
        .Q(EXEC_STAGE_mul_ex_H[21]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_20_ ( .G(n13543), .D(EXEC_STAGE_mul_ex_N67), 
        .Q(EXEC_STAGE_mul_ex_H[20]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_19_ ( .G(n13543), .D(EXEC_STAGE_mul_ex_N68), 
        .Q(EXEC_STAGE_mul_ex_H[19]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_18_ ( .G(n13543), .D(EXEC_STAGE_mul_ex_N69), 
        .Q(EXEC_STAGE_mul_ex_H[18]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_17_ ( .G(n13543), .D(EXEC_STAGE_mul_ex_N70), 
        .Q(EXEC_STAGE_mul_ex_H[17]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_16_ ( .G(n13543), .D(EXEC_STAGE_mul_ex_N71), 
        .Q(EXEC_STAGE_mul_ex_H[16]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_15_ ( .G(n13543), .D(EXEC_STAGE_mul_ex_N72), 
        .Q(EXEC_STAGE_mul_ex_H[15]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_14_ ( .G(n13543), .D(EXEC_STAGE_mul_ex_N73), 
        .Q(EXEC_STAGE_mul_ex_H[14]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_13_ ( .G(n13543), .D(EXEC_STAGE_mul_ex_N74), 
        .Q(EXEC_STAGE_mul_ex_H[13]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_12_ ( .G(n13543), .D(EXEC_STAGE_mul_ex_N75), 
        .Q(EXEC_STAGE_mul_ex_H[12]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_11_ ( .G(n13543), .D(EXEC_STAGE_mul_ex_N76), 
        .Q(EXEC_STAGE_mul_ex_H[11]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_10_ ( .G(n13543), .D(EXEC_STAGE_mul_ex_N77), 
        .Q(EXEC_STAGE_mul_ex_H[10]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_9_ ( .G(n19192), .D(EXEC_STAGE_mul_ex_N78), 
        .Q(EXEC_STAGE_mul_ex_H[9]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_8_ ( .G(n13543), .D(EXEC_STAGE_mul_ex_N79), 
        .Q(EXEC_STAGE_mul_ex_H[8]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_7_ ( .G(n13542), .D(EXEC_STAGE_mul_ex_N80), 
        .Q(EXEC_STAGE_mul_ex_H[7]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_6_ ( .G(n19192), .D(EXEC_STAGE_mul_ex_N81), 
        .Q(EXEC_STAGE_mul_ex_H[6]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_5_ ( .G(n13543), .D(EXEC_STAGE_mul_ex_N82), 
        .Q(EXEC_STAGE_mul_ex_H[5]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_4_ ( .G(n13542), .D(EXEC_STAGE_mul_ex_N83), 
        .Q(EXEC_STAGE_mul_ex_H[4]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_3_ ( .G(n19192), .D(EXEC_STAGE_mul_ex_N84), 
        .Q(EXEC_STAGE_mul_ex_H[3]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_2_ ( .G(n19192), .D(EXEC_STAGE_mul_ex_N85), 
        .Q(EXEC_STAGE_mul_ex_H[2]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_1_ ( .G(n19192), .D(EXEC_STAGE_mul_ex_N86), 
        .Q(EXEC_STAGE_mul_ex_H[1]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_0_ ( .G(n19192), .D(EXEC_STAGE_mul_ex_N87), 
        .Q(EXEC_STAGE_mul_ex_H[0]) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_31_ ( .G(n13868), .D(EXEC_STAGE_mul_ex_N412), 
        .Q(EXEC_STAGE_mul_ex_Z_31_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_30_ ( .G(n13868), .D(EXEC_STAGE_mul_ex_N413), 
        .Q(EXEC_STAGE_mul_ex_Z_30_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_29_ ( .G(n13868), .D(EXEC_STAGE_mul_ex_N414), 
        .Q(EXEC_STAGE_mul_ex_Z_29_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_28_ ( .G(n13868), .D(EXEC_STAGE_mul_ex_N415), 
        .Q(EXEC_STAGE_mul_ex_Z_28_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_27_ ( .G(n13868), .D(EXEC_STAGE_mul_ex_N416), 
        .Q(EXEC_STAGE_mul_ex_Z_27_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_26_ ( .G(n13868), .D(EXEC_STAGE_mul_ex_N417), 
        .Q(EXEC_STAGE_mul_ex_Z_26_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_25_ ( .G(n13868), .D(EXEC_STAGE_mul_ex_N418), 
        .Q(EXEC_STAGE_mul_ex_Z_25_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_24_ ( .G(n13868), .D(EXEC_STAGE_mul_ex_N419), 
        .Q(EXEC_STAGE_mul_ex_Z_24_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_23_ ( .G(n13868), .D(EXEC_STAGE_mul_ex_N420), 
        .Q(EXEC_STAGE_mul_ex_Z_23_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_22_ ( .G(n13868), .D(EXEC_STAGE_mul_ex_N421), 
        .Q(EXEC_STAGE_mul_ex_Z_22_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_21_ ( .G(n13868), .D(EXEC_STAGE_mul_ex_N422), 
        .Q(EXEC_STAGE_mul_ex_Z_21_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_20_ ( .G(n13869), .D(EXEC_STAGE_mul_ex_N423), 
        .Q(EXEC_STAGE_mul_ex_Z_20_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_19_ ( .G(n13869), .D(EXEC_STAGE_mul_ex_N424), 
        .Q(EXEC_STAGE_mul_ex_Z_19_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_18_ ( .G(n13869), .D(EXEC_STAGE_mul_ex_N425), 
        .Q(EXEC_STAGE_mul_ex_Z_18_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_17_ ( .G(n13869), .D(EXEC_STAGE_mul_ex_N426), 
        .Q(EXEC_STAGE_mul_ex_Z_17_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_16_ ( .G(n13869), .D(EXEC_STAGE_mul_ex_N427), 
        .Q(EXEC_STAGE_mul_ex_Z_16_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_15_ ( .G(n13869), .D(EXEC_STAGE_mul_ex_N428), 
        .Q(EXEC_STAGE_mul_ex_Z_15_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_14_ ( .G(n13869), .D(EXEC_STAGE_mul_ex_N429), 
        .Q(EXEC_STAGE_mul_ex_Z_14_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_13_ ( .G(n13869), .D(EXEC_STAGE_mul_ex_N430), 
        .Q(EXEC_STAGE_mul_ex_Z_13_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_12_ ( .G(n13869), .D(EXEC_STAGE_mul_ex_N431), 
        .Q(EXEC_STAGE_mul_ex_Z_12_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_11_ ( .G(n13869), .D(EXEC_STAGE_mul_ex_N432), 
        .Q(EXEC_STAGE_mul_ex_Z_11_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_10_ ( .G(n13869), .D(EXEC_STAGE_mul_ex_N433), 
        .Q(EXEC_STAGE_mul_ex_Z_10_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_9_ ( .G(n13868), .D(EXEC_STAGE_mul_ex_N434), 
        .Q(EXEC_STAGE_mul_ex_Z_9_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_8_ ( .G(EXEC_STAGE_mul_ex_N411), .D(
        EXEC_STAGE_mul_ex_N435), .Q(EXEC_STAGE_mul_ex_Z_8_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_7_ ( .G(n13869), .D(EXEC_STAGE_mul_ex_N436), 
        .Q(EXEC_STAGE_mul_ex_Z_7_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_6_ ( .G(n13869), .D(EXEC_STAGE_mul_ex_N437), 
        .Q(EXEC_STAGE_mul_ex_Z_6_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_5_ ( .G(n13868), .D(EXEC_STAGE_mul_ex_N438), 
        .Q(EXEC_STAGE_mul_ex_Z_5_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_4_ ( .G(EXEC_STAGE_mul_ex_N411), .D(
        EXEC_STAGE_mul_ex_N439), .Q(EXEC_STAGE_mul_ex_Z_4_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_3_ ( .G(EXEC_STAGE_mul_ex_N411), .D(
        EXEC_STAGE_mul_ex_N440), .Q(EXEC_STAGE_mul_ex_Z_3_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_2_ ( .G(EXEC_STAGE_mul_ex_N411), .D(
        EXEC_STAGE_mul_ex_N441), .Q(EXEC_STAGE_mul_ex_Z_2_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_1_ ( .G(EXEC_STAGE_mul_ex_N411), .D(
        EXEC_STAGE_mul_ex_N442), .Q(EXEC_STAGE_mul_ex_Z_1_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_0_ ( .G(EXEC_STAGE_mul_ex_N411), .D(
        EXEC_STAGE_mul_ex_N443), .Q(EXEC_STAGE_mul_ex_Z_0_) );
  DLH_X2 EXEC_STAGE_mul_ex_done_reg ( .G(EXEC_STAGE_mul_ex_N479), .D(n13544), 
        .Q(EXEC_STAGE_mul_done) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_0_ ( .G(EXEC_STAGE_mul_ex_N378), .D(
        EXEC_STAGE_mul_ex_N410), .Q(EXEC_STAGE_mul_ex_L_0_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_1_ ( .G(EXEC_STAGE_mul_ex_N378), .D(
        EXEC_STAGE_mul_ex_N409), .Q(EXEC_STAGE_mul_ex_L_1_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_2_ ( .G(EXEC_STAGE_mul_ex_N378), .D(
        EXEC_STAGE_mul_ex_N408), .Q(EXEC_STAGE_mul_ex_L_2_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_3_ ( .G(n13866), .D(EXEC_STAGE_mul_ex_N407), 
        .Q(EXEC_STAGE_mul_ex_L_3_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_4_ ( .G(EXEC_STAGE_mul_ex_N378), .D(
        EXEC_STAGE_mul_ex_N406), .Q(EXEC_STAGE_mul_ex_L_4_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_5_ ( .G(n13865), .D(EXEC_STAGE_mul_ex_N405), 
        .Q(EXEC_STAGE_mul_ex_L_5_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_6_ ( .G(n13866), .D(EXEC_STAGE_mul_ex_N404), 
        .Q(EXEC_STAGE_mul_ex_L_6_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_7_ ( .G(EXEC_STAGE_mul_ex_N378), .D(
        EXEC_STAGE_mul_ex_N403), .Q(EXEC_STAGE_mul_ex_L_7_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_8_ ( .G(n13865), .D(EXEC_STAGE_mul_ex_N402), 
        .Q(EXEC_STAGE_mul_ex_L_8_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_9_ ( .G(n13866), .D(EXEC_STAGE_mul_ex_N401), 
        .Q(EXEC_STAGE_mul_ex_L_9_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_10_ ( .G(EXEC_STAGE_mul_ex_N378), .D(
        EXEC_STAGE_mul_ex_N400), .Q(EXEC_STAGE_mul_ex_L_10_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_11_ ( .G(n13865), .D(EXEC_STAGE_mul_ex_N399), 
        .Q(EXEC_STAGE_mul_ex_L_11_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_12_ ( .G(n13865), .D(EXEC_STAGE_mul_ex_N398), 
        .Q(EXEC_STAGE_mul_ex_L_12_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_13_ ( .G(n13865), .D(EXEC_STAGE_mul_ex_N397), 
        .Q(EXEC_STAGE_mul_ex_L_13_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_14_ ( .G(n13865), .D(EXEC_STAGE_mul_ex_N396), 
        .Q(EXEC_STAGE_mul_ex_L_14_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_15_ ( .G(n13865), .D(EXEC_STAGE_mul_ex_N395), 
        .Q(EXEC_STAGE_mul_ex_L_15_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_16_ ( .G(n13865), .D(EXEC_STAGE_mul_ex_N394), 
        .Q(EXEC_STAGE_mul_ex_L_16_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_17_ ( .G(n13865), .D(EXEC_STAGE_mul_ex_N393), 
        .Q(EXEC_STAGE_mul_ex_L_17_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_18_ ( .G(n13865), .D(EXEC_STAGE_mul_ex_N392), 
        .Q(EXEC_STAGE_mul_ex_L_18_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_19_ ( .G(n13865), .D(EXEC_STAGE_mul_ex_N391), 
        .Q(EXEC_STAGE_mul_ex_L_19_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_20_ ( .G(n13865), .D(EXEC_STAGE_mul_ex_N390), 
        .Q(EXEC_STAGE_mul_ex_L_20_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_21_ ( .G(n13865), .D(EXEC_STAGE_mul_ex_N389), 
        .Q(EXEC_STAGE_mul_ex_L_21_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_22_ ( .G(n13866), .D(EXEC_STAGE_mul_ex_N388), 
        .Q(EXEC_STAGE_mul_ex_L_22_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_23_ ( .G(n13866), .D(EXEC_STAGE_mul_ex_N387), 
        .Q(EXEC_STAGE_mul_ex_L_23_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_24_ ( .G(n13866), .D(EXEC_STAGE_mul_ex_N386), 
        .Q(EXEC_STAGE_mul_ex_L_24_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_25_ ( .G(n13866), .D(EXEC_STAGE_mul_ex_N385), 
        .Q(EXEC_STAGE_mul_ex_L_25_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_26_ ( .G(n13866), .D(EXEC_STAGE_mul_ex_N384), 
        .Q(EXEC_STAGE_mul_ex_L_26_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_27_ ( .G(n13866), .D(EXEC_STAGE_mul_ex_N383), 
        .Q(EXEC_STAGE_mul_ex_L_27_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_28_ ( .G(n13866), .D(EXEC_STAGE_mul_ex_N382), 
        .Q(EXEC_STAGE_mul_ex_L_28_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_29_ ( .G(n13866), .D(EXEC_STAGE_mul_ex_N381), 
        .Q(EXEC_STAGE_mul_ex_L_29_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_30_ ( .G(n13866), .D(EXEC_STAGE_mul_ex_N380), 
        .Q(EXEC_STAGE_mul_ex_L_30_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_31_ ( .G(n13866), .D(EXEC_STAGE_mul_ex_N379), 
        .Q(EXEC_STAGE_mul_ex_L_31_) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_0_ ( .G(n13871), .D(EXEC_STAGE_mul_ex_N476), 
        .Q(EXEC_STAGE_mul_ex_P[0]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_1_ ( .G(n13871), .D(EXEC_STAGE_mul_ex_N475), 
        .Q(EXEC_STAGE_mul_ex_P[1]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_2_ ( .G(n13871), .D(EXEC_STAGE_mul_ex_N474), 
        .Q(EXEC_STAGE_mul_ex_P[2]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_3_ ( .G(n13871), .D(EXEC_STAGE_mul_ex_N473), 
        .Q(EXEC_STAGE_mul_ex_P[3]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_4_ ( .G(n13871), .D(EXEC_STAGE_mul_ex_N472), 
        .Q(EXEC_STAGE_mul_ex_P[4]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_5_ ( .G(n13871), .D(EXEC_STAGE_mul_ex_N471), 
        .Q(EXEC_STAGE_mul_ex_P[5]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_6_ ( .G(n13871), .D(EXEC_STAGE_mul_ex_N470), 
        .Q(EXEC_STAGE_mul_ex_P[6]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_7_ ( .G(n13871), .D(EXEC_STAGE_mul_ex_N469), 
        .Q(EXEC_STAGE_mul_ex_P[7]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_8_ ( .G(n13871), .D(EXEC_STAGE_mul_ex_N468), 
        .Q(EXEC_STAGE_mul_ex_P[8]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_9_ ( .G(n13871), .D(EXEC_STAGE_mul_ex_N467), 
        .Q(EXEC_STAGE_mul_ex_P[9]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_10_ ( .G(n13871), .D(EXEC_STAGE_mul_ex_N466), 
        .Q(EXEC_STAGE_mul_ex_P[10]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_11_ ( .G(n13872), .D(EXEC_STAGE_mul_ex_N465), 
        .Q(EXEC_STAGE_mul_ex_P[11]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_12_ ( .G(n13872), .D(EXEC_STAGE_mul_ex_N464), 
        .Q(EXEC_STAGE_mul_ex_P[12]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_13_ ( .G(n13872), .D(EXEC_STAGE_mul_ex_N463), 
        .Q(EXEC_STAGE_mul_ex_P[13]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_14_ ( .G(n13872), .D(EXEC_STAGE_mul_ex_N462), 
        .Q(EXEC_STAGE_mul_ex_P[14]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_15_ ( .G(n13872), .D(EXEC_STAGE_mul_ex_N461), 
        .Q(EXEC_STAGE_mul_ex_P[15]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_16_ ( .G(n13872), .D(EXEC_STAGE_mul_ex_N460), 
        .Q(EXEC_STAGE_mul_ex_P[16]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_17_ ( .G(n13872), .D(EXEC_STAGE_mul_ex_N459), 
        .Q(EXEC_STAGE_mul_ex_P[17]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_18_ ( .G(n13872), .D(EXEC_STAGE_mul_ex_N458), 
        .Q(EXEC_STAGE_mul_ex_P[18]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_19_ ( .G(n13872), .D(EXEC_STAGE_mul_ex_N457), 
        .Q(EXEC_STAGE_mul_ex_P[19]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_20_ ( .G(n13872), .D(EXEC_STAGE_mul_ex_N456), 
        .Q(EXEC_STAGE_mul_ex_P[20]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_21_ ( .G(n13872), .D(EXEC_STAGE_mul_ex_N455), 
        .Q(EXEC_STAGE_mul_ex_P[21]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_22_ ( .G(EXEC_STAGE_mul_ex_N444), .D(
        EXEC_STAGE_mul_ex_N454), .Q(EXEC_STAGE_mul_ex_P[22]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_23_ ( .G(n13871), .D(EXEC_STAGE_mul_ex_N453), 
        .Q(EXEC_STAGE_mul_ex_P[23]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_24_ ( .G(n13872), .D(EXEC_STAGE_mul_ex_N452), 
        .Q(EXEC_STAGE_mul_ex_P[24]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_25_ ( .G(EXEC_STAGE_mul_ex_N444), .D(
        EXEC_STAGE_mul_ex_N451), .Q(EXEC_STAGE_mul_ex_P[25]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_26_ ( .G(EXEC_STAGE_mul_ex_N444), .D(
        EXEC_STAGE_mul_ex_N450), .Q(EXEC_STAGE_mul_ex_P[26]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_27_ ( .G(EXEC_STAGE_mul_ex_N444), .D(
        EXEC_STAGE_mul_ex_N449), .Q(EXEC_STAGE_mul_ex_P[27]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_28_ ( .G(n13871), .D(EXEC_STAGE_mul_ex_N448), 
        .Q(EXEC_STAGE_mul_ex_P[28]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_29_ ( .G(n13872), .D(EXEC_STAGE_mul_ex_N447), 
        .Q(EXEC_STAGE_mul_ex_P[29]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_30_ ( .G(EXEC_STAGE_mul_ex_N444), .D(
        EXEC_STAGE_mul_ex_N446), .Q(EXEC_STAGE_mul_ex_P[30]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_31_ ( .G(EXEC_STAGE_mul_ex_N444), .D(
        EXEC_STAGE_mul_ex_N445), .Q(EXEC_STAGE_mul_ex_P[31]) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12824) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12079) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11846) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__31_), .QN(n12298) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10461) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__31_), .QN(n12177) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12025) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12920) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12785) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10530) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__31_), .QN(n11430) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10847) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__31_), .QN(n12081) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__31_), .QN(n12666) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__31_), .QN(n12643) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__31_), .QN(n10750) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12498) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10367) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10251) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__31_), .QN(n12062) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12411) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10257) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__31_), .QN(n11469) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__31_), .QN(n10718) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12919) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__31_), .QN(n10689) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__31_), .QN(n12063) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__31_), .QN(n12088) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__31_), .QN(n10766) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12412) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12766) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__31_), .QN(n12135) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__31_), .QN(n11739) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__31_), .QN(n11346) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__31_), .QN(n11749) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__31_), .QN(n11307) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10491) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__31_), .QN(n10608) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__31_), .QN(n11213) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__31_), .QN(n11172) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10430) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__31_), .QN(n11396) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__31_), .QN(n11273) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__31_), .QN(n11288) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__31_), .QN(n11774) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__31_), .QN(n11460) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__31_), .QN(n11036) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11495) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__31_), .QN(n11585) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__31_), .QN(n11243) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10229) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10460) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__31_), .QN(n11026) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__31_), .QN(n11337) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__31_), .QN(n11673) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11486) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__31_), .QN(n11609) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__31_), .QN(n10638) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__31_), .QN(n11015) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__31_), .QN(n10589) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11496) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__31_), .QN(n11135) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__31_), .QN(n11641) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__0_), .QN(n11617) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__0_), .QN(n12644) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10400) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__0_), .QN(n10719) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__0_), .QN(n11373) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10263) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__0_), .QN(n12667) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__0_), .QN(n11244) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__0_), .QN(n11347) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__0_), .QN(n10650) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10462) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__0_), .QN(n10639) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__0_), .QN(n12691) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__0_), .QN(n11184) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__0_), .QN(n11431) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__0_), .QN(n11143) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__0_), .QN(n11821) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12321) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12345) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__0_), .QN(n11597) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__0_), .QN(n12232) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__0_), .QN(n11214) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__0_), .QN(n10609) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10200) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__0_), .QN(n11784) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10431) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__0_), .QN(n10560) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__0_), .QN(n11795) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__0_), .QN(n11681) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__0_), .QN(n11308) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__0_), .QN(n11173) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__0_), .QN(n11649) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__18_), .QN(n12653) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10417) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__18_), .QN(n10737) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__18_), .QN(n11382) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10280) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__18_), .QN(n12676) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__18_), .QN(n11262) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__18_), .QN(n11296) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__18_), .QN(n10659) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10480) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__18_), .QN(n10597) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__18_), .QN(n12700) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__18_), .QN(n11202) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__18_), .QN(n11449) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__18_), .QN(n11161) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__18_), .QN(n11034) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12339) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12370) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__18_), .QN(n11606) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__18_), .QN(n12249) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__18_), .QN(n11232) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__18_), .QN(n10627) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10218) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__18_), .QN(n11013) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10449) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__18_), .QN(n10578) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__18_), .QN(n11024) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12371) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__18_), .QN(n11326) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__18_), .QN(n11124) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__18_), .QN(n11658) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__18_), .QN(n11626) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12823) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11880) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__30_), .QN(n11736) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__30_), .QN(n11820) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_5__30_), .QN(n10749) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__30_), .QN(n10791) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12049) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12918) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12784) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10529) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__30_), .QN(n11429) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10926) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__30_), .QN(n12270) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__30_), .QN(n12599) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__30_), .QN(n12584) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12497) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12765) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__30_), .QN(n10540) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10300) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__30_), .QN(n12146) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__30_), .QN(n11735) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__30_), .QN(n10348) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12496) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__30_), .QN(n10717) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12917) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11895) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__30_), .QN(n10800) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__30_), .QN(n11771) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__30_), .QN(n10765) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__30_), .QN(n11734) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12495) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11503) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__30_), .QN(n11738) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10429) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__30_), .QN(n11345) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__30_), .QN(n11395) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10290) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__30_), .QN(n11748) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__30_), .QN(n11272) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__30_), .QN(n11306) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__30_), .QN(n11287) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10490) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__30_), .QN(n10607) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__30_), .QN(n11773) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__30_), .QN(n11212) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__30_), .QN(n11459) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__30_), .QN(n11171) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__30_), .QN(n11035) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11485) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11493) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__30_), .QN(n11608) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__30_), .QN(n11584) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__30_), .QN(n11242) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__30_), .QN(n10637) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10228) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__30_), .QN(n11014) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10459) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__30_), .QN(n10588) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__30_), .QN(n11025) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11494) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__30_), .QN(n11336) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__30_), .QN(n11134) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__30_), .QN(n11672) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__30_), .QN(n11640) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12822) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11879) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__29_), .QN(n11733) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__29_), .QN(n11819) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_5__29_), .QN(n10748) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__29_), .QN(n10790) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12048) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12916) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12783) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10528) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__29_), .QN(n11428) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10925) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__29_), .QN(n12269) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__29_), .QN(n12598) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__29_), .QN(n12583) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12494) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12764) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__29_), .QN(n10539) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10299) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__29_), .QN(n12145) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__29_), .QN(n11732) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__29_), .QN(n10347) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12493) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__29_), .QN(n10716) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12915) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11894) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__29_), .QN(n10799) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__29_), .QN(n11770) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__29_), .QN(n10764) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__29_), .QN(n11731) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12492) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11502) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__29_), .QN(n12665) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10428) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__29_), .QN(n11344) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__29_), .QN(n11393) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10289) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__29_), .QN(n12688) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__29_), .QN(n11271) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__29_), .QN(n11305) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__29_), .QN(n11286) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10489) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__29_), .QN(n10606) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__29_), .QN(n12712) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__29_), .QN(n11211) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__29_), .QN(n11458) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__29_), .QN(n11170) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__29_), .QN(n12121) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11484) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11492) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__29_), .QN(n12626) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__29_), .QN(n12614) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__29_), .QN(n11241) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__29_), .QN(n10636) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10227) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__29_), .QN(n12099) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10458) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__29_), .QN(n10587) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__29_), .QN(n12110) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12078) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__29_), .QN(n11335) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__29_), .QN(n11133) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__29_), .QN(n11670) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__29_), .QN(n11638) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__25_), .QN(n12661) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10424) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__25_), .QN(n11340) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__25_), .QN(n11389) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10285) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__25_), .QN(n12684) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__25_), .QN(n11267) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__25_), .QN(n11301) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__25_), .QN(n11282) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10485) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__25_), .QN(n10602) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__25_), .QN(n12708) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__25_), .QN(n11207) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__25_), .QN(n11454) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__25_), .QN(n11166) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__25_), .QN(n12117) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11480) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11488) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__25_), .QN(n12622) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__25_), .QN(n12610) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__25_), .QN(n11237) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__25_), .QN(n10632) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10223) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__25_), .QN(n12095) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10454) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__25_), .QN(n10583) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__25_), .QN(n12106) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12074) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__25_), .QN(n11331) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__25_), .QN(n11129) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__25_), .QN(n11666) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__25_), .QN(n11634) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__27_), .QN(n12663) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10426) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__27_), .QN(n11342) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__27_), .QN(n11391) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10287) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__27_), .QN(n12686) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__27_), .QN(n11269) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__27_), .QN(n11303) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__27_), .QN(n11284) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10487) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__27_), .QN(n10604) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__27_), .QN(n12710) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__27_), .QN(n11209) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__27_), .QN(n11456) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__27_), .QN(n11168) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__27_), .QN(n12119) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11482) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11490) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__27_), .QN(n12624) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__27_), .QN(n12612) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__27_), .QN(n11239) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__27_), .QN(n10634) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10225) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__27_), .QN(n12097) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10456) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__27_), .QN(n10585) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__27_), .QN(n12108) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12076) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__27_), .QN(n11333) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__27_), .QN(n11131) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__27_), .QN(n11668) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__27_), .QN(n11636) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__26_), .QN(n12662) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10425) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__26_), .QN(n11341) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__26_), .QN(n11390) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10286) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__26_), .QN(n12685) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__26_), .QN(n11268) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__26_), .QN(n11302) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__26_), .QN(n11283) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10486) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__26_), .QN(n10603) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__26_), .QN(n12709) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__26_), .QN(n11208) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__26_), .QN(n11455) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__26_), .QN(n11167) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__26_), .QN(n12118) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11481) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11489) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__26_), .QN(n12623) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__26_), .QN(n12611) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__26_), .QN(n11238) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__26_), .QN(n10633) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10224) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__26_), .QN(n12096) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10455) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__26_), .QN(n10584) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__26_), .QN(n12107) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12075) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__26_), .QN(n11332) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__26_), .QN(n11130) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__26_), .QN(n11667) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__26_), .QN(n11635) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[28]), .QN(n12553) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12821) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11878) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__28_), .QN(n11730) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__28_), .QN(n11818) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_5__28_), .QN(n10747) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__28_), .QN(n10789) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12047) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12914) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12782) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10527) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__28_), .QN(n11427) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10924) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__28_), .QN(n12268) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__28_), .QN(n12597) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__28_), .QN(n12582) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12491) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12763) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__28_), .QN(n10538) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10298) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__28_), .QN(n12144) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__28_), .QN(n11729) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__28_), .QN(n10346) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12490) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__28_), .QN(n12278) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12913) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11893) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__28_), .QN(n10798) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__28_), .QN(n11769) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__28_), .QN(n10763) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__28_), .QN(n11728) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12489) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11501) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12820) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11877) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__27_), .QN(n11727) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__27_), .QN(n11817) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_5__27_), .QN(n10746) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__27_), .QN(n10788) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12046) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12912) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12781) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10526) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__27_), .QN(n11426) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10923) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__27_), .QN(n12267) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__27_), .QN(n12596) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__27_), .QN(n12581) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12488) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12762) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__27_), .QN(n10537) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10297) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__27_), .QN(n12143) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__27_), .QN(n11726) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__27_), .QN(n10345) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12487) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__27_), .QN(n10715) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12911) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11892) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__27_), .QN(n10797) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__27_), .QN(n11768) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__27_), .QN(n10762) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__27_), .QN(n11725) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12486) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11500) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12819) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11876) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__26_), .QN(n11724) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__26_), .QN(n11816) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_5__26_), .QN(n10745) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__26_), .QN(n10787) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12045) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12910) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12780) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10525) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__26_), .QN(n11425) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10922) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__26_), .QN(n12266) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__26_), .QN(n12595) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__26_), .QN(n12580) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12485) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12761) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__26_), .QN(n10536) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10296) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__26_), .QN(n12142) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__26_), .QN(n11723) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__26_), .QN(n10344) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12484) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__26_), .QN(n12277) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12909) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11891) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__26_), .QN(n10796) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__26_), .QN(n11767) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__26_), .QN(n10761) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__26_), .QN(n11722) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12483) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11499) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12818) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11875) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__25_), .QN(n11721) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__25_), .QN(n11815) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_5__25_), .QN(n10744) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__25_), .QN(n10786) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12044) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12908) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12779) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10524) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__25_), .QN(n11424) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10921) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__25_), .QN(n12265) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__25_), .QN(n12594) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__25_), .QN(n12579) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12482) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12760) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__25_), .QN(n10535) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10295) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__25_), .QN(n12141) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__25_), .QN(n11720) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__25_), .QN(n10343) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12481) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__25_), .QN(n10714) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12907) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11890) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__25_), .QN(n10795) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__25_), .QN(n11766) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__25_), .QN(n10760) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__25_), .QN(n11719) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12480) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11498) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12817) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11874) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__24_), .QN(n11718) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__24_), .QN(n11814) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_5__24_), .QN(n10743) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__24_), .QN(n10785) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12043) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12906) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12778) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10523) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__24_), .QN(n11423) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10920) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__24_), .QN(n12264) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__24_), .QN(n12593) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__24_), .QN(n12578) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12479) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12759) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__24_), .QN(n10534) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10294) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__24_), .QN(n12140) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__24_), .QN(n11717) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__24_), .QN(n10342) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12478) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__24_), .QN(n10713) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12905) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11889) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__24_), .QN(n10794) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__24_), .QN(n11765) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__24_), .QN(n10759) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__24_), .QN(n11716) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12477) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11497) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__28_), .QN(n12664) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10427) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__28_), .QN(n11343) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__28_), .QN(n11392) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10288) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__28_), .QN(n12687) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__28_), .QN(n11270) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__28_), .QN(n11304) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__28_), .QN(n11285) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10488) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__28_), .QN(n10605) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__28_), .QN(n12711) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__28_), .QN(n11210) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__28_), .QN(n11457) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__28_), .QN(n11169) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__28_), .QN(n12120) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11483) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11491) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__28_), .QN(n12625) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__28_), .QN(n12613) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__28_), .QN(n11240) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__28_), .QN(n10635) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10226) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__28_), .QN(n12098) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10457) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__28_), .QN(n10586) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__28_), .QN(n12109) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12077) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__28_), .QN(n11334) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__28_), .QN(n11132) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__28_), .QN(n11669) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__28_), .QN(n11637) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12816) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11873) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__23_), .QN(n11715) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__23_), .QN(n11813) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_5__23_), .QN(n10742) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__23_), .QN(n10784) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12042) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12904) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12777) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10522) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__23_), .QN(n11422) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10919) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__23_), .QN(n12263) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__23_), .QN(n12592) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__23_), .QN(n12577) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12476) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12758) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__23_), .QN(n10533) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10293) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__23_), .QN(n12139) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__23_), .QN(n11714) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__23_), .QN(n10341) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12475) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__23_), .QN(n10712) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12903) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11888) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__23_), .QN(n10793) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__23_), .QN(n11764) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__23_), .QN(n10758) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__23_), .QN(n11713) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12474) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12410) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__15_), .QN(n12650) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10414) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__15_), .QN(n10734) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__15_), .QN(n11379) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10277) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__15_), .QN(n12673) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__15_), .QN(n11259) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__15_), .QN(n11293) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__15_), .QN(n10656) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10477) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__15_), .QN(n10594) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__15_), .QN(n12697) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__15_), .QN(n11199) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__15_), .QN(n11446) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__15_), .QN(n11158) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__15_), .QN(n11031) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12336) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12364) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__15_), .QN(n11603) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__15_), .QN(n12246) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__15_), .QN(n11229) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__15_), .QN(n10624) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10215) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__15_), .QN(n11010) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10446) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__15_), .QN(n10575) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__15_), .QN(n11021) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12365) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__15_), .QN(n11323) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__15_), .QN(n11121) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__15_), .QN(n11655) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__15_), .QN(n11623) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12814) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12213) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__22_), .QN(n11712) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__22_), .QN(n11812) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_5__22_), .QN(n10741) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__22_), .QN(n10783) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10321) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12902) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12250) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10521) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__22_), .QN(n11421) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10918) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__22_), .QN(n12262) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__22_), .QN(n12591) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__22_), .QN(n12576) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12473) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11872) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__22_), .QN(n10324) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10292) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__22_), .QN(n12138) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__22_), .QN(n11711) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__22_), .QN(n10340) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12472) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__22_), .QN(n10711) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12901) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12815) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__22_), .QN(n10792) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__22_), .QN(n11763) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__22_), .QN(n10757) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__22_), .QN(n11710) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12471) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12409) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__14_), .QN(n12649) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10413) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__14_), .QN(n10733) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__14_), .QN(n11378) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10276) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__14_), .QN(n12672) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__14_), .QN(n11258) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__14_), .QN(n11292) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__14_), .QN(n10655) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10476) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__14_), .QN(n10593) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__14_), .QN(n12696) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__14_), .QN(n11198) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__14_), .QN(n11445) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__14_), .QN(n11157) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__14_), .QN(n11030) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12335) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12362) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__14_), .QN(n11602) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__14_), .QN(n12245) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__14_), .QN(n11228) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__14_), .QN(n10623) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10214) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__14_), .QN(n11009) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10445) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__14_), .QN(n10574) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__14_), .QN(n11020) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12363) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__14_), .QN(n11322) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__14_), .QN(n11120) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__14_), .QN(n11654) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__14_), .QN(n11622) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12812) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11870) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__21_), .QN(n11709) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__21_), .QN(n11811) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_5__21_), .QN(n11420) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__21_), .QN(n11577) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10320) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12900) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11869) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10932) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__21_), .QN(n12295) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10502) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__21_), .QN(n11279) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__21_), .QN(n12590) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__21_), .QN(n12575) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12470) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11871) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__21_), .QN(n10234) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10503) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__21_), .QN(n11101) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__21_), .QN(n11708) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__21_), .QN(n10772) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12469) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__21_), .QN(n10710) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12899) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12813) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__21_), .QN(n11582) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__21_), .QN(n11762) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__21_), .QN(n10756) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__21_), .QN(n11707) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12468) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12408) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__13_), .QN(n12648) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10412) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__13_), .QN(n10732) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__13_), .QN(n11377) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10275) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__13_), .QN(n12671) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__13_), .QN(n11257) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__13_), .QN(n11291) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__13_), .QN(n10654) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10475) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__13_), .QN(n10592) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__13_), .QN(n12695) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__13_), .QN(n11197) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__13_), .QN(n11444) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__13_), .QN(n11156) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__13_), .QN(n11029) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12334) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12360) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__13_), .QN(n11601) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__13_), .QN(n12244) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__13_), .QN(n11227) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__13_), .QN(n10622) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10213) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__13_), .QN(n11008) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10444) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__13_), .QN(n10573) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__13_), .QN(n11019) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12361) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__13_), .QN(n11321) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__13_), .QN(n11119) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__13_), .QN(n11653) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__13_), .QN(n11621) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__3_), .QN(n11740) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10402) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__3_), .QN(n10722) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__3_), .QN(n11397) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10265) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__3_), .QN(n11750) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__3_), .QN(n11247) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__3_), .QN(n11350) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__3_), .QN(n10666) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10465) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__3_), .QN(n10642) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__3_), .QN(n11775) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__3_), .QN(n11187) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__3_), .QN(n11434) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__3_), .QN(n11146) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__3_), .QN(n11825) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12324) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12348) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__3_), .QN(n11610) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__3_), .QN(n12234) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__3_), .QN(n11217) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__3_), .QN(n10612) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10203) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__3_), .QN(n11788) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10434) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__3_), .QN(n10563) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__3_), .QN(n11799) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__3_), .QN(n11685) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__3_), .QN(n11311) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__3_), .QN(n11176) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__3_), .QN(n11674) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__3_), .QN(n11642) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12810) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11867) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__20_), .QN(n11706) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__20_), .QN(n11810) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_5__20_), .QN(n11419) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__20_), .QN(n11576) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10319) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12898) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11866) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10931) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__20_), .QN(n12294) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10500) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__20_), .QN(n11278) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__20_), .QN(n12589) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__20_), .QN(n12574) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12467) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11868) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__20_), .QN(n10233) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10501) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__20_), .QN(n11100) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__20_), .QN(n11705) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__20_), .QN(n10771) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12466) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__20_), .QN(n10709) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12897) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12811) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__20_), .QN(n11581) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__20_), .QN(n11761) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__20_), .QN(n10755) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__20_), .QN(n11704) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12465) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12407) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12808) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11864) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__19_), .QN(n11703) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__19_), .QN(n11809) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_5__19_), .QN(n11418) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__19_), .QN(n11575) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10318) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12896) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12757) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10930) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__19_), .QN(n12293) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10498) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__19_), .QN(n11277) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__19_), .QN(n12588) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__19_), .QN(n12573) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12464) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11865) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__19_), .QN(n10232) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10499) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__19_), .QN(n11099) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__19_), .QN(n11702) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__19_), .QN(n10770) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12463) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__19_), .QN(n10708) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12895) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12809) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__19_), .QN(n11580) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__19_), .QN(n11760) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__19_), .QN(n10754) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__19_), .QN(n11701) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12462) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12406) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12806) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11862) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__18_), .QN(n11700) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__18_), .QN(n11808) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_5__18_), .QN(n11417) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__18_), .QN(n11574) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10317) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12894) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12756) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10929) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__18_), .QN(n12292) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10496) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__18_), .QN(n11276) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__18_), .QN(n12587) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__18_), .QN(n12572) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12461) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11863) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__18_), .QN(n10231) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10497) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__18_), .QN(n11098) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__18_), .QN(n11699) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__18_), .QN(n10769) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12460) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__18_), .QN(n10707) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12893) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12807) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__18_), .QN(n11579) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__18_), .QN(n11759) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__18_), .QN(n10753) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__18_), .QN(n11698) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12459) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12405) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[4]) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__4_), .QN(n12805) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11861) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12744) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12456) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10305) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__4_), .QN(n10704) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__4_), .QN(n11005) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12892) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12755) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10509) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12457) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10878) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10879) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__4_), .QN(n10677) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__4_), .QN(n10339) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12736) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12455) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10256) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10389) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12951) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10384) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__4_), .QN(n12087) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12891) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__4_), .QN(n12642) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12890) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__4_), .QN(n11407) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12458) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__4_), .QN(n10981) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__4_), .QN(n11361) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10249) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12889) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__4_), .QN(n12391) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[3]) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[2]) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12804) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11860) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11839) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12385) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10302) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__1_), .QN(n10703) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__1_), .QN(n11004) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12888) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12768) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10506) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12386) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10872) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10873) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__1_), .QN(n10674) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__1_), .QN(n10338) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12735) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12454) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10868) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10386) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12938) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10381) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__1_), .QN(n12086) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12887) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__1_), .QN(n12641) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12886) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__1_), .QN(n11404) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11882) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__1_), .QN(n10980) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__1_), .QN(n11358) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10246) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12885) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__1_), .QN(n12384) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__1_), .QN(n12655) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10913) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__1_), .QN(n10720) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__1_), .QN(n12284) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10399) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__1_), .QN(n12678) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__1_), .QN(n11245) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__1_), .QN(n11348) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__1_), .QN(n12271) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10463) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__1_), .QN(n10640) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__1_), .QN(n12702) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__1_), .QN(n11185) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__1_), .QN(n11432) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__1_), .QN(n11144) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__1_), .QN(n11823) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12322) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12346) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__1_), .QN(n12616) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__1_), .QN(n12604) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__1_), .QN(n11215) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__1_), .QN(n10610) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10201) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__1_), .QN(n11786) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10432) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__1_), .QN(n10561) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__1_), .QN(n11797) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__1_), .QN(n11683) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__1_), .QN(n11309) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__1_), .QN(n11174) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__1_), .QN(n11660) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__1_), .QN(n11628) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12802) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11858) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__17_), .QN(n11697) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__17_), .QN(n11807) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_5__17_), .QN(n11416) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__17_), .QN(n11783) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10316) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12884) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12754) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10928) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__17_), .QN(n12291) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10494) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__17_), .QN(n11275) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__17_), .QN(n12586) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__17_), .QN(n12571) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12453) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11859) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__17_), .QN(n10230) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10495) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__17_), .QN(n11274) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__17_), .QN(n11696) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__17_), .QN(n10768) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12452) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__17_), .QN(n10706) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12883) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12803) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__17_), .QN(n11782) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__17_), .QN(n11758) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__17_), .QN(n10752) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__17_), .QN(n11695) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12451) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12404) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__9_), .QN(n12801) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11857) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12743) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12448) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10310) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__9_), .QN(n10702) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__9_), .QN(n11003) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12882) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12753) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10514) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12449) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10892) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10893) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__9_), .QN(n10682) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__9_), .QN(n10337) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12734) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12447) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10255) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10390) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12950) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10851) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__9_), .QN(n12085) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12881) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__9_), .QN(n12640) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12880) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__9_), .QN(n11408) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12450) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__9_), .QN(n10979) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__9_), .QN(n11366) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10375) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12879) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__9_), .QN(n12398) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[5]) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__3_), .QN(n12800) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11856) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12742) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12444) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10304) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__3_), .QN(n10701) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__3_), .QN(n11002) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12878) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12752) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10508) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12445) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10876) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10877) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__3_), .QN(n10676) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__3_), .QN(n10336) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12733) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12443) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10254) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10388) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12949) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10383) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__3_), .QN(n12084) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12877) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__3_), .QN(n12639) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12876) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__3_), .QN(n11406) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12446) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__3_), .QN(n10978) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__3_), .QN(n11360) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10248) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12875) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__3_), .QN(n12390) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12799) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11855) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11840) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12388) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10303) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__2_), .QN(n10700) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__2_), .QN(n11001) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12874) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12769) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10507) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12389) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10874) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10875) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__2_), .QN(n10675) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__2_), .QN(n10335) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12732) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12442) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10867) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10387) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12939) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10382) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__2_), .QN(n12083) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12873) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__2_), .QN(n12638) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12872) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__2_), .QN(n11405) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11883) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__2_), .QN(n10977) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__2_), .QN(n11359) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10247) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12871) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__2_), .QN(n12387) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__2_), .QN(n11737) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10401) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__2_), .QN(n10721) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__2_), .QN(n11394) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10264) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__2_), .QN(n11747) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__2_), .QN(n11246) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__2_), .QN(n11349) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__2_), .QN(n10665) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10464) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__2_), .QN(n10641) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__2_), .QN(n11772) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__2_), .QN(n11186) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__2_), .QN(n11433) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__2_), .QN(n11145) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__2_), .QN(n11824) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12323) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12347) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__2_), .QN(n11607) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__2_), .QN(n12233) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__2_), .QN(n11216) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__2_), .QN(n10611) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10202) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__2_), .QN(n11787) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10433) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__2_), .QN(n10562) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__2_), .QN(n11798) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__2_), .QN(n11684) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__2_), .QN(n11310) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__2_), .QN(n11175) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__2_), .QN(n11671) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__2_), .QN(n11639) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12797) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11854) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__16_), .QN(n11694) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__16_), .QN(n11806) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_5__16_), .QN(n11415) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__16_), .QN(n11573) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10520) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12870) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12776) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10927) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__16_), .QN(n12290) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10492) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__16_), .QN(n12261) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__16_), .QN(n12585) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__16_), .QN(n12570) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12441) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12751) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__16_), .QN(n10942) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10493) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__16_), .QN(n12137) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__16_), .QN(n11693) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__16_), .QN(n10767) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12440) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__16_), .QN(n10705) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12869) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12798) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__16_), .QN(n11578) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__16_), .QN(n11757) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__16_), .QN(n10751) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__16_), .QN(n11692) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12439) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12403) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__15_), .QN(n12796) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11853) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12741) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12436) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10504) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__15_), .QN(n12276) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__15_), .QN(n12082) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12868) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12750) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12041) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12437) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10904) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10905) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__15_), .QN(n10688) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__15_), .QN(n12279) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12731) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12435) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10253) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10396) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12952) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12024) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__15_), .QN(n11000) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12867) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__15_), .QN(n12637) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12866) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__15_), .QN(n11414) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12438) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__15_), .QN(n12080) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__15_), .QN(n11372) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10846) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12865) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__15_), .QN(n11596) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12795) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12228) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11845) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12401) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10315) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__14_), .QN(n10699) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__14_), .QN(n10998) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12864) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12775) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10519) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12402) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10902) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10903) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__14_), .QN(n10687) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__14_), .QN(n10334) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12730) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12434) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10866) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10395) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12944) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10856) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__14_), .QN(n10999) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12863) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__14_), .QN(n12636) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12862) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__14_), .QN(n11413) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11887) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__14_), .QN(n10976) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__14_), .QN(n11371) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10380) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12861) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__14_), .QN(n11595) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__13_), .QN(n12794) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11852) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12740) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12431) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10314) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__13_), .QN(n10698) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__13_), .QN(n10996) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12860) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12749) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10518) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12432) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10900) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10901) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__13_), .QN(n10686) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__13_), .QN(n10333) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12729) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12430) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10252) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10394) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12948) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10855) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__13_), .QN(n10997) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12859) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__13_), .QN(n12635) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12858) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__13_), .QN(n11412) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12433) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__13_), .QN(n10975) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__13_), .QN(n11370) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10379) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12857) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__13_), .QN(n11594) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__16_), .QN(n12651) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10415) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__16_), .QN(n10735) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__16_), .QN(n11380) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10278) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__16_), .QN(n12674) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__16_), .QN(n11260) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__16_), .QN(n11294) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__16_), .QN(n10657) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10478) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__16_), .QN(n10595) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__16_), .QN(n12698) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__16_), .QN(n11200) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__16_), .QN(n11447) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__16_), .QN(n11159) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__16_), .QN(n11032) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12337) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12366) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__16_), .QN(n11604) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__16_), .QN(n12247) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__16_), .QN(n11230) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__16_), .QN(n10625) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10216) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__16_), .QN(n11011) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10447) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__16_), .QN(n10576) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__16_), .QN(n11022) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12367) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__16_), .QN(n11324) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__16_), .QN(n11122) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__16_), .QN(n11656) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__16_), .QN(n11624) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12793) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12227) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11844) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12399) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10313) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__12_), .QN(n10697) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__12_), .QN(n10994) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12856) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12774) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10517) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12400) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10898) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10899) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__12_), .QN(n10685) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__12_), .QN(n10332) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12728) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12429) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10865) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10393) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12943) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10854) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__12_), .QN(n10995) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12855) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__12_), .QN(n12634) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12854) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__12_), .QN(n11411) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12773) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__12_), .QN(n10974) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__12_), .QN(n11369) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10378) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12853) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__12_), .QN(n11593) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12792) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12226) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11842) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12394) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10308) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__7_), .QN(n10696) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__7_), .QN(n10992) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12852) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12771) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10512) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12395) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10887) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10888) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__7_), .QN(n10680) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__7_), .QN(n10331) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12727) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12428) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10864) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10886) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12941) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10849) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__7_), .QN(n10993) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12851) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__7_), .QN(n12633) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12850) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__7_), .QN(n12288) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11885) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__7_), .QN(n10973) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__7_), .QN(n11364) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10373) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12849) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__7_), .QN(n11592) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__7_), .QN(n11744) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10406) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__7_), .QN(n10726) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__7_), .QN(n11401) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10269) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__7_), .QN(n11754) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__7_), .QN(n11251) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__7_), .QN(n11354) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__7_), .QN(n10670) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10469) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__7_), .QN(n10646) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__7_), .QN(n11779) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__7_), .QN(n11191) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__7_), .QN(n11438) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__7_), .QN(n11150) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__7_), .QN(n11829) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12328) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12352) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__7_), .QN(n11614) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__7_), .QN(n12238) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__7_), .QN(n11221) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__7_), .QN(n10616) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10207) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__7_), .QN(n11792) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10438) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__7_), .QN(n10567) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__7_), .QN(n11803) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__7_), .QN(n11689) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__7_), .QN(n11315) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__7_), .QN(n11180) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__7_), .QN(n11678) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__7_), .QN(n11646) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__11_), .QN(n12791) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11851) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12739) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12425) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10312) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__11_), .QN(n10695) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__11_), .QN(n10990) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12848) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12748) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10516) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12426) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10896) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10897) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__11_), .QN(n10684) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__11_), .QN(n10330) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12726) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12424) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10859) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10392) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12947) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10853) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__11_), .QN(n10991) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12847) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__11_), .QN(n12632) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12846) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__11_), .QN(n11410) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12427) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__11_), .QN(n10972) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__11_), .QN(n11368) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10377) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12845) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__11_), .QN(n11591) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__11_), .QN(n12646) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10410) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__11_), .QN(n10730) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__11_), .QN(n11375) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10273) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__11_), .QN(n12669) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__11_), .QN(n11255) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__11_), .QN(n11289) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__11_), .QN(n10652) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10473) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__11_), .QN(n10590) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__11_), .QN(n12693) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__11_), .QN(n11195) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__11_), .QN(n11442) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__11_), .QN(n11154) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__11_), .QN(n11027) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12332) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12356) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__11_), .QN(n11599) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__11_), .QN(n12242) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__11_), .QN(n11225) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__11_), .QN(n10620) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10211) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__11_), .QN(n11006) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10442) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__11_), .QN(n10571) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__11_), .QN(n11017) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12357) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__11_), .QN(n11319) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__11_), .QN(n11117) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__11_), .QN(n11651) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__11_), .QN(n11619) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__10_), .QN(n12790) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11850) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12738) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12421) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10311) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__10_), .QN(n10694) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__10_), .QN(n10988) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12844) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12747) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10515) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12422) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10894) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10895) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__10_), .QN(n10683) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__10_), .QN(n10329) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12725) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12420) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10858) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10391) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12946) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10852) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__10_), .QN(n10989) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12843) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__10_), .QN(n12631) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12842) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__10_), .QN(n11409) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12423) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__10_), .QN(n10971) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__10_), .QN(n11367) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10376) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12841) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__10_), .QN(n11590) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__10_), .QN(n12645) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10409) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__10_), .QN(n10729) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__10_), .QN(n11374) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10272) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__10_), .QN(n12668) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__10_), .QN(n11254) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__10_), .QN(n11357) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__10_), .QN(n10651) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10472) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__10_), .QN(n10649) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__10_), .QN(n12692) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__10_), .QN(n11194) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__10_), .QN(n11441) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__10_), .QN(n11153) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__10_), .QN(n11822) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12331) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12355) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__10_), .QN(n11598) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__10_), .QN(n12241) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__10_), .QN(n11224) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__10_), .QN(n10619) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10210) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__10_), .QN(n11785) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10441) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__10_), .QN(n10570) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__10_), .QN(n11796) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__10_), .QN(n11682) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__10_), .QN(n11318) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__10_), .QN(n11183) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__10_), .QN(n11650) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__10_), .QN(n11618) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12789) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12225) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11843) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12396) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10309) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__8_), .QN(n10693) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__8_), .QN(n10986) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12840) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12772) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10513) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12397) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10890) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10891) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__8_), .QN(n10681) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__8_), .QN(n10328) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12724) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12419) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10863) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10889) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12942) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10850) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__8_), .QN(n10987) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12839) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__8_), .QN(n12630) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12838) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__8_), .QN(n12289) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11886) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__8_), .QN(n10970) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__8_), .QN(n11365) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10374) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12837) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__8_), .QN(n11589) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__8_), .QN(n11745) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10407) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__8_), .QN(n10727) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__8_), .QN(n11402) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10270) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__8_), .QN(n11755) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__8_), .QN(n11252) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__8_), .QN(n11355) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__8_), .QN(n10671) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10470) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__8_), .QN(n10647) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__8_), .QN(n11780) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__8_), .QN(n11192) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__8_), .QN(n11439) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__8_), .QN(n11151) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__8_), .QN(n11830) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12329) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12353) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__8_), .QN(n11615) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__8_), .QN(n12239) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__8_), .QN(n11222) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__8_), .QN(n10617) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10208) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__8_), .QN(n11793) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10439) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__8_), .QN(n10568) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__8_), .QN(n11804) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__8_), .QN(n11690) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__8_), .QN(n11316) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__8_), .QN(n11181) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__8_), .QN(n11679) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__8_), .QN(n11647) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__6_), .QN(n12788) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11849) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12737) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12416) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10307) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__6_), .QN(n10692) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__6_), .QN(n10984) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12836) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12746) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10511) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12417) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10884) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10885) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__6_), .QN(n10679) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__6_), .QN(n10327) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12723) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12415) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10857) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10883) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12945) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10848) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__6_), .QN(n10985) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12835) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__6_), .QN(n12629) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12834) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__6_), .QN(n12287) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12418) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__6_), .QN(n10969) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__6_), .QN(n11363) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10372) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12833) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__6_), .QN(n11588) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12787) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11848) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11841) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12392) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10306) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__5_), .QN(n10691) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__5_), .QN(n10982) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12832) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12770) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10510) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12393) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10881) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10882) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__5_), .QN(n10678) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__5_), .QN(n10326) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12722) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12414) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10862) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10880) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12940) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10385) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__5_), .QN(n10983) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12831) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__5_), .QN(n12628) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12830) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__5_), .QN(n12286) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11884) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__5_), .QN(n10968) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__5_), .QN(n11362) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10250) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12829) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__5_), .QN(n11587) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__5_), .QN(n11742) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10404) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__5_), .QN(n10724) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__5_), .QN(n11399) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10267) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__5_), .QN(n11752) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__5_), .QN(n11249) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__5_), .QN(n11352) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__5_), .QN(n10668) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10467) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__5_), .QN(n10644) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__5_), .QN(n11777) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__5_), .QN(n11189) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__5_), .QN(n11436) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__5_), .QN(n11148) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__5_), .QN(n11827) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12326) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12350) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__5_), .QN(n11612) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__5_), .QN(n12236) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__5_), .QN(n11219) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__5_), .QN(n10614) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10205) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__5_), .QN(n11790) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10436) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__5_), .QN(n10565) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__5_), .QN(n11801) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__5_), .QN(n11687) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__5_), .QN(n11313) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__5_), .QN(n11178) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__5_), .QN(n11676) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__5_), .QN(n11644) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__6_), .QN(n11743) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10405) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__6_), .QN(n10725) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__6_), .QN(n11400) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10268) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__6_), .QN(n11753) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__6_), .QN(n11250) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__6_), .QN(n11353) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__6_), .QN(n10669) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10468) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__6_), .QN(n10645) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__6_), .QN(n11778) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__6_), .QN(n11190) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__6_), .QN(n11437) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__6_), .QN(n11149) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__6_), .QN(n11828) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12327) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12351) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__6_), .QN(n11613) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__6_), .QN(n12237) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__6_), .QN(n11220) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__6_), .QN(n10615) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10206) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__6_), .QN(n11791) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10437) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__6_), .QN(n10566) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__6_), .QN(n11802) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__6_), .QN(n11688) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__6_), .QN(n11314) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__6_), .QN(n11179) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__6_), .QN(n11677) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__6_), .QN(n11645) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__12_), .QN(n12647) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10411) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__12_), .QN(n10731) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__12_), .QN(n11376) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10274) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__12_), .QN(n12670) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__12_), .QN(n11256) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__12_), .QN(n11290) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__12_), .QN(n10653) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10474) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__12_), .QN(n10591) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__12_), .QN(n12694) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__12_), .QN(n11196) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__12_), .QN(n11443) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__12_), .QN(n11155) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__12_), .QN(n11028) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12333) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12358) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__12_), .QN(n11600) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__12_), .QN(n12243) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__12_), .QN(n11226) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__12_), .QN(n10621) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10212) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__12_), .QN(n11007) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10443) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__12_), .QN(n10572) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__12_), .QN(n11018) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12359) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__12_), .QN(n11320) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__12_), .QN(n11118) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__12_), .QN(n11652) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__12_), .QN(n11620) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__9_), .QN(n11746) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10408) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__9_), .QN(n10728) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__9_), .QN(n11403) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10271) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__9_), .QN(n11756) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__9_), .QN(n11253) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__9_), .QN(n11356) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__9_), .QN(n10672) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10471) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__9_), .QN(n10648) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__9_), .QN(n11781) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__9_), .QN(n11193) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__9_), .QN(n11440) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__9_), .QN(n11152) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__9_), .QN(n11831) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12330) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12354) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__9_), .QN(n11616) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__9_), .QN(n12240) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__9_), .QN(n11223) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__9_), .QN(n10618) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10209) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__9_), .QN(n11794) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10440) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__9_), .QN(n10569) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__9_), .QN(n11805) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__9_), .QN(n11691) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__9_), .QN(n11317) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__9_), .QN(n11182) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__9_), .QN(n11680) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__9_), .QN(n11648) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__17_), .QN(n12652) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10416) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__17_), .QN(n10736) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__17_), .QN(n11381) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10279) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__17_), .QN(n12675) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__17_), .QN(n11261) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__17_), .QN(n11295) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__17_), .QN(n10658) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10479) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__17_), .QN(n10596) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__17_), .QN(n12699) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__17_), .QN(n11201) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__17_), .QN(n11448) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__17_), .QN(n11160) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__17_), .QN(n11033) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12338) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12368) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__17_), .QN(n11605) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__17_), .QN(n12248) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__17_), .QN(n11231) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__17_), .QN(n10626) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10217) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__17_), .QN(n11012) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10448) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__17_), .QN(n10577) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__17_), .QN(n11023) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12369) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__17_), .QN(n11325) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__17_), .QN(n11123) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__17_), .QN(n11657) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__17_), .QN(n11625) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12786) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11847) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11838) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12382) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10301) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__0_), .QN(n10690) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__0_), .QN(n10958) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12828) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12767) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10505) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12383) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10870) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10871) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__0_), .QN(n10673) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__0_), .QN(n10325) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12721) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12413) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10861) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10869) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12937) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10371) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__0_), .QN(n10959) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12827) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__0_), .QN(n12627) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12826) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__0_), .QN(n12285) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11881) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__0_), .QN(n10949) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__0_), .QN(n11338) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10245) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12825) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__0_), .QN(n11586) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__4_), .QN(n11741) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10403) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__4_), .QN(n10723) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__4_), .QN(n11398) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10266) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__4_), .QN(n11751) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__4_), .QN(n11248) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__4_), .QN(n11351) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__4_), .QN(n10667) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10466) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__4_), .QN(n10643) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__4_), .QN(n11776) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__4_), .QN(n11188) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__4_), .QN(n11435) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__4_), .QN(n11147) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__4_), .QN(n11826) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12325) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12349) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__4_), .QN(n11611) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__4_), .QN(n12235) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__4_), .QN(n11218) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__4_), .QN(n10613) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10204) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__4_), .QN(n11789) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10435) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__4_), .QN(n10564) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__4_), .QN(n11800) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__4_), .QN(n11686) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__4_), .QN(n11312) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__4_), .QN(n11177) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__4_), .QN(n11675) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__4_), .QN(n11643) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__20_), .QN(n12656) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10419) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__20_), .QN(n12283) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__20_), .QN(n11384) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10912) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__20_), .QN(n12679) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__20_), .QN(n12260) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__20_), .QN(n12273) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__20_), .QN(n10661) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10917) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__20_), .QN(n11140) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__20_), .QN(n12703) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__20_), .QN(n12255) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__20_), .QN(n12297) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__20_), .QN(n12252) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__20_), .QN(n12112) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12341) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12374) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__20_), .QN(n12617) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__20_), .QN(n12605) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__20_), .QN(n12257) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__20_), .QN(n11142) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10261) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__20_), .QN(n12090) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10915) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__20_), .QN(n11138) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__20_), .QN(n12101) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12375) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__20_), .QN(n12281) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__20_), .QN(n12222) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__20_), .QN(n11661) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__20_), .QN(n11629) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__21_), .QN(n12657) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10420) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__21_), .QN(n10738) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__21_), .QN(n11385) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10281) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__21_), .QN(n12680) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__21_), .QN(n11263) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__21_), .QN(n11297) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__21_), .QN(n10662) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10481) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__21_), .QN(n10598) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__21_), .QN(n12704) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__21_), .QN(n11203) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__21_), .QN(n11450) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__21_), .QN(n11162) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__21_), .QN(n12113) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12342) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12376) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__21_), .QN(n12618) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__21_), .QN(n12606) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__21_), .QN(n11233) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__21_), .QN(n10628) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10219) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__21_), .QN(n12091) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10450) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__21_), .QN(n10579) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__21_), .QN(n12102) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12377) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__21_), .QN(n11327) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__21_), .QN(n11125) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__21_), .QN(n11662) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__21_), .QN(n11630) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__22_), .QN(n12658) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10421) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__22_), .QN(n10739) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__22_), .QN(n11386) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10282) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__22_), .QN(n12681) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__22_), .QN(n11264) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__22_), .QN(n11298) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__22_), .QN(n10663) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10482) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__22_), .QN(n10599) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__22_), .QN(n12705) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__22_), .QN(n11204) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__22_), .QN(n11451) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__22_), .QN(n11163) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__22_), .QN(n12114) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12343) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12378) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__22_), .QN(n12619) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__22_), .QN(n12607) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__22_), .QN(n11234) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__22_), .QN(n10629) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10220) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__22_), .QN(n12092) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10451) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__22_), .QN(n10580) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__22_), .QN(n12103) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12379) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__22_), .QN(n11328) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__22_), .QN(n11126) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__22_), .QN(n11663) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__22_), .QN(n11631) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__19_), .QN(n12654) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10418) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__19_), .QN(n12282) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__19_), .QN(n11383) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10911) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__19_), .QN(n12677) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__19_), .QN(n12259) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__19_), .QN(n12272) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__19_), .QN(n10660) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10916) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__19_), .QN(n11139) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__19_), .QN(n12701) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__19_), .QN(n12254) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__19_), .QN(n12296) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__19_), .QN(n12251) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__19_), .QN(n12111) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12340) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12372) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__19_), .QN(n12615) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__19_), .QN(n12603) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__19_), .QN(n12256) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__19_), .QN(n11141) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10260) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__19_), .QN(n12089) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10914) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__19_), .QN(n11137) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__19_), .QN(n12100) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12373) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__19_), .QN(n12280) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__19_), .QN(n12221) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__19_), .QN(n11659) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__19_), .QN(n11627) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__23_), .QN(n12659) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10422) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__23_), .QN(n10740) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__23_), .QN(n11387) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10283) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__23_), .QN(n12682) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__23_), .QN(n11265) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__23_), .QN(n11299) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__23_), .QN(n10664) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10483) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__23_), .QN(n10600) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__23_), .QN(n12706) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__23_), .QN(n11205) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__23_), .QN(n11452) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__23_), .QN(n11164) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__23_), .QN(n12115) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12344) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12380) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__23_), .QN(n12620) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__23_), .QN(n12608) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__23_), .QN(n11235) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__23_), .QN(n10630) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10221) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__23_), .QN(n12093) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10452) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__23_), .QN(n10581) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__23_), .QN(n12104) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12381) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__23_), .QN(n11329) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__23_), .QN(n11127) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__23_), .QN(n11664) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__23_), .QN(n11632) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__24_), .QN(n12660) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10423) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__24_), .QN(n11339) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__24_), .QN(n11388) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10284) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__24_), .QN(n12683) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__24_), .QN(n11266) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__24_), .QN(n11300) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__24_), .QN(n11281) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10484) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__24_), .QN(n10601) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__24_), .QN(n12707) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__24_), .QN(n11206) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__24_), .QN(n11453) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__24_), .QN(n11165) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__24_), .QN(n12116) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11479) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11487) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__24_), .QN(n12621) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__24_), .QN(n12609) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__24_), .QN(n11236) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__24_), .QN(n10631) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10222) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__24_), .QN(n12094) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10453) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__24_), .QN(n10582) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__24_), .QN(n12105) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12073) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__24_), .QN(n11330) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__24_), .QN(n11128) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__24_), .QN(n11665) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__24_), .QN(n11633) );
  NAND2_X2 U1315 ( .A1(DMEM_BUS_IN[15]), .A2(net231221), .ZN(n1236) );
  NAND2_X2 U1318 ( .A1(DMEM_BUS_IN[14]), .A2(net231221), .ZN(n1238) );
  NAND2_X2 U1321 ( .A1(DMEM_BUS_IN[13]), .A2(net231263), .ZN(n1240) );
  NAND2_X2 U1324 ( .A1(DMEM_BUS_IN[12]), .A2(net231221), .ZN(n1242) );
  NAND2_X2 U1327 ( .A1(DMEM_BUS_IN[11]), .A2(net231221), .ZN(n1244) );
  NAND2_X2 U1331 ( .A1(DMEM_BUS_IN[10]), .A2(net231221), .ZN(n1248) );
  NAND2_X2 U1334 ( .A1(DMEM_BUS_IN[9]), .A2(net231221), .ZN(n1250) );
  NAND2_X2 U1337 ( .A1(DMEM_BUS_IN[8]), .A2(net231221), .ZN(n1252) );
  NAND2_X2 U1340 ( .A1(DMEM_BUS_IN[7]), .A2(net231221), .ZN(n1254) );
  NAND2_X2 U1343 ( .A1(DMEM_BUS_IN[6]), .A2(net231221), .ZN(n1256) );
  NAND2_X2 U1346 ( .A1(DMEM_BUS_IN[5]), .A2(net231221), .ZN(n1258) );
  NAND2_X2 U1349 ( .A1(DMEM_BUS_IN[4]), .A2(net231221), .ZN(n1260) );
  NAND2_X2 U1352 ( .A1(DMEM_BUS_IN[3]), .A2(net231221), .ZN(n1262) );
  NAND2_X2 U1355 ( .A1(DMEM_BUS_IN[2]), .A2(net231221), .ZN(n1264) );
  NAND2_X2 U1358 ( .A1(DMEM_BUS_IN[1]), .A2(net231221), .ZN(n1266) );
  NAND2_X2 U1362 ( .A1(DMEM_BUS_IN[0]), .A2(net231221), .ZN(n1270) );
  AOI22_X2 U1365 ( .A1(MEM_WB_OUT[68]), .A2(net231307), .B1(net231233), .B2(
        DMEM_BUS_OUT[31]), .ZN(n1271) );
  AOI22_X2 U1376 ( .A1(MEM_WB_OUT[59]), .A2(net231307), .B1(net231233), .B2(
        DMEM_BUS_OUT[22]), .ZN(n1290) );
  AOI22_X2 U1378 ( .A1(MEM_WB_OUT[58]), .A2(net231309), .B1(net231233), .B2(
        DMEM_BUS_OUT[21]), .ZN(n1291) );
  AOI22_X2 U1380 ( .A1(MEM_WB_OUT[57]), .A2(net231309), .B1(net231233), .B2(
        DMEM_BUS_OUT[20]), .ZN(n1292) );
  AOI22_X2 U1382 ( .A1(MEM_WB_OUT[56]), .A2(net231309), .B1(net231233), .B2(
        DMEM_BUS_OUT[19]), .ZN(n1293) );
  AOI22_X2 U1384 ( .A1(MEM_WB_OUT[55]), .A2(net231309), .B1(net231233), .B2(
        DMEM_BUS_OUT[18]), .ZN(n1294) );
  AOI22_X2 U1386 ( .A1(MEM_WB_OUT[54]), .A2(net231309), .B1(net231233), .B2(
        DMEM_BUS_OUT[17]), .ZN(n1295) );
  AOI22_X2 U1389 ( .A1(MEM_WB_OUT[52]), .A2(net231309), .B1(net231233), .B2(
        DMEM_BUS_OUT[15]), .ZN(n1298) );
  AOI22_X2 U1392 ( .A1(MEM_WB_OUT[50]), .A2(net231309), .B1(net231233), .B2(
        DMEM_BUS_OUT[13]), .ZN(n1301) );
  AOI22_X2 U1396 ( .A1(MEM_WB_OUT[48]), .A2(net231309), .B1(net231233), .B2(
        DMEM_BUS_OUT[11]), .ZN(n1306) );
  AOI22_X2 U1398 ( .A1(MEM_WB_OUT[47]), .A2(net231309), .B1(net231233), .B2(
        DMEM_BUS_OUT[10]), .ZN(n1307) );
  AOI22_X2 U1400 ( .A1(MEM_WB_OUT[46]), .A2(net231309), .B1(net231233), .B2(
        DMEM_BUS_OUT[9]), .ZN(n1308) );
  AOI22_X2 U1404 ( .A1(MEM_WB_OUT[43]), .A2(net231309), .B1(net231233), .B2(
        DMEM_BUS_OUT[6]), .ZN(n1313) );
  AOI22_X2 U1407 ( .A1(MEM_WB_OUT[41]), .A2(net231309), .B1(net231233), .B2(
        DMEM_BUS_OUT[4]), .ZN(n1316) );
  AOI22_X2 U1409 ( .A1(MEM_WB_OUT[40]), .A2(net231309), .B1(net231233), .B2(
        DMEM_BUS_OUT[3]), .ZN(n1317) );
  AOI22_X2 U1412 ( .A1(MEM_WB_OUT[39]), .A2(net231309), .B1(net231233), .B2(
        DMEM_BUS_OUT[2]), .ZN(n1320) );
  OAI22_X2 U1413 ( .A1(n12180), .A2(net231263), .B1(net231313), .B2(n10826), 
        .ZN(n7335) );
  OAI22_X2 U1414 ( .A1(n12040), .A2(net231263), .B1(net231313), .B2(n10825), 
        .ZN(n7755) );
  OAI22_X2 U1415 ( .A1(n19320), .A2(net231263), .B1(net231313), .B2(n19319), 
        .ZN(n7874) );
  OAI22_X2 U1416 ( .A1(n19317), .A2(net231261), .B1(net231313), .B2(n19316), 
        .ZN(n7882) );
  OAI22_X2 U1417 ( .A1(n19315), .A2(net231263), .B1(net231313), .B2(n19314), 
        .ZN(n7885) );
  OAI22_X2 U1420 ( .A1(n19311), .A2(net231261), .B1(net231313), .B2(n19310), 
        .ZN(n7891) );
  OAI22_X2 U1422 ( .A1(n12538), .A2(net231263), .B1(net231313), .B2(n11109), 
        .ZN(n7830) );
  OAI22_X2 U1424 ( .A1(n12537), .A2(net231263), .B1(net231313), .B2(n11108), 
        .ZN(n7740) );
  OAI22_X2 U1427 ( .A1(n12499), .A2(net231263), .B1(net231313), .B2(n11115), 
        .ZN(n7725) );
  AOI22_X2 U1430 ( .A1(MEM_WB_OUT[28]), .A2(net231309), .B1(net231233), .B2(
        MEM_WB_REG_MEM_WB_REG_N152), .ZN(n1338) );
  OAI22_X2 U1431 ( .A1(n12224), .A2(net231263), .B1(net231313), .B2(n11107), 
        .ZN(n7681) );
  OAI22_X2 U1433 ( .A1(n12536), .A2(net231263), .B1(net231313), .B2(n11114), 
        .ZN(n7673) );
  OAI22_X2 U1435 ( .A1(n11136), .A2(net231263), .B1(net231313), .B2(n12308), 
        .ZN(n7664) );
  AOI22_X2 U1438 ( .A1(MEM_WB_OUT[24]), .A2(net231309), .B1(net231235), .B2(
        MEM_WB_REG_MEM_WB_REG_N156), .ZN(n1345) );
  OAI22_X2 U1439 ( .A1(n12535), .A2(net231263), .B1(net231313), .B2(n11106), 
        .ZN(n7639) );
  AOI22_X2 U1442 ( .A1(MEM_WB_OUT[22]), .A2(net231309), .B1(net231233), .B2(
        MEM_WB_REG_MEM_WB_REG_N158), .ZN(n1348) );
  OAI22_X2 U1443 ( .A1(n12547), .A2(net231263), .B1(net231315), .B2(n11105), 
        .ZN(n7603) );
  AOI22_X2 U1446 ( .A1(MEM_WB_OUT[20]), .A2(net231309), .B1(net231235), .B2(
        MEM_WB_REG_MEM_WB_REG_N160), .ZN(n1351) );
  OAI22_X2 U1448 ( .A1(n12546), .A2(net231263), .B1(net231313), .B2(n11113), 
        .ZN(n7571) );
  OAI22_X2 U1450 ( .A1(n12545), .A2(net231251), .B1(net231315), .B2(n11104), 
        .ZN(n7563) );
  AOI22_X2 U1453 ( .A1(MEM_WB_OUT[17]), .A2(net231309), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N163), .ZN(n1358) );
  OAI22_X2 U1454 ( .A1(net231247), .A2(n13875), .B1(net231315), .B2(n12204), 
        .ZN(n7758) );
  OAI22_X2 U1455 ( .A1(net231239), .A2(n10365), .B1(net231315), .B2(n12203), 
        .ZN(n7850) );
  OAI22_X2 U1456 ( .A1(net231239), .A2(n10196), .B1(net231315), .B2(n12176), 
        .ZN(n7760) );
  OAI22_X2 U1457 ( .A1(net231239), .A2(n10195), .B1(net231315), .B2(n12175), 
        .ZN(n7734) );
  OAI22_X2 U1458 ( .A1(net231239), .A2(n10194), .B1(net231315), .B2(n12174), 
        .ZN(n7719) );
  OAI22_X2 U1459 ( .A1(net231239), .A2(n10193), .B1(net231315), .B2(n12173), 
        .ZN(n7648) );
  OAI22_X2 U1460 ( .A1(net231237), .A2(n10192), .B1(net231315), .B2(n12172), 
        .ZN(n7707) );
  OAI22_X2 U1461 ( .A1(net231239), .A2(n10191), .B1(net231315), .B2(n12171), 
        .ZN(n7701) );
  OAI22_X2 U1462 ( .A1(net231237), .A2(n10190), .B1(net231315), .B2(n12299), 
        .ZN(n7713) );
  OAI22_X2 U1463 ( .A1(n12223), .A2(net231263), .B1(net231311), .B2(n11103), 
        .ZN(n7471) );
  OAI22_X2 U1465 ( .A1(net231237), .A2(n10189), .B1(net231317), .B2(n12170), 
        .ZN(n7297) );
  OAI22_X2 U1466 ( .A1(net231237), .A2(n10188), .B1(net231317), .B2(n12169), 
        .ZN(n7301) );
  OAI22_X2 U1467 ( .A1(net231237), .A2(n10187), .B1(net231317), .B2(n12168), 
        .ZN(n7309) );
  OAI22_X2 U1468 ( .A1(net231237), .A2(n10186), .B1(net231317), .B2(n12167), 
        .ZN(n7313) );
  OAI22_X2 U1469 ( .A1(net231237), .A2(n10239), .B1(net231317), .B2(n12166), 
        .ZN(n7318) );
  OAI22_X2 U1470 ( .A1(net231237), .A2(n10238), .B1(net231317), .B2(n12165), 
        .ZN(n7305) );
  OAI22_X2 U1471 ( .A1(net231237), .A2(n10185), .B1(net231317), .B2(n12164), 
        .ZN(n7749) );
  OAI22_X2 U1472 ( .A1(net231237), .A2(n10184), .B1(net231317), .B2(n12163), 
        .ZN(n7339) );
  OAI22_X2 U1473 ( .A1(net231237), .A2(n10183), .B1(net231317), .B2(n12162), 
        .ZN(n7438) );
  OAI22_X2 U1474 ( .A1(net231237), .A2(n10182), .B1(net231317), .B2(n12161), 
        .ZN(n7629) );
  OAI22_X2 U1476 ( .A1(net231237), .A2(n10181), .B1(net231317), .B2(n12160), 
        .ZN(n7612) );
  OAI22_X2 U1477 ( .A1(net231235), .A2(n10180), .B1(net231317), .B2(n12159), 
        .ZN(n7595) );
  OAI22_X2 U1478 ( .A1(net231237), .A2(n10179), .B1(net231317), .B2(n12158), 
        .ZN(n7349) );
  OAI22_X2 U1479 ( .A1(net231235), .A2(n10178), .B1(net231317), .B2(n12157), 
        .ZN(n7396) );
  OAI22_X2 U1480 ( .A1(net231235), .A2(n10177), .B1(net231317), .B2(n12156), 
        .ZN(n7386) );
  OAI22_X2 U1481 ( .A1(net231235), .A2(n10176), .B1(net231317), .B2(n12155), 
        .ZN(n7344) );
  OAI22_X2 U1482 ( .A1(net231235), .A2(n10175), .B1(net231315), .B2(n12154), 
        .ZN(n7377) );
  OAI22_X2 U1483 ( .A1(net231235), .A2(n10174), .B1(net231315), .B2(n12153), 
        .ZN(n7406) );
  OAI22_X2 U1484 ( .A1(net231235), .A2(n10173), .B1(net231315), .B2(n12152), 
        .ZN(n7355) );
  OAI22_X2 U1485 ( .A1(net231235), .A2(n10172), .B1(net231315), .B2(n12151), 
        .ZN(n7361) );
  OAI22_X2 U1487 ( .A1(net231237), .A2(n10171), .B1(net231315), .B2(n12150), 
        .ZN(n7323) );
  OAI22_X2 U1488 ( .A1(net231235), .A2(n10170), .B1(net231315), .B2(n12149), 
        .ZN(n7589) );
  OAI22_X2 U1489 ( .A1(net231235), .A2(n10169), .B1(net231315), .B2(n12148), 
        .ZN(n7480) );
  OAI22_X2 U1490 ( .A1(net231235), .A2(n10237), .B1(net231315), .B2(n12147), 
        .ZN(n7533) );
  OAI22_X2 U1491 ( .A1(net231235), .A2(n10168), .B1(net231315), .B2(n12178), 
        .ZN(n7753) );
  AOI22_X2 U1493 ( .A1(net231297), .A2(MEM_WB_OUT[144]), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N35), .ZN(n1433) );
  AOI22_X2 U1495 ( .A1(net231315), .A2(MEM_WB_OUT[143]), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N36), .ZN(n1434) );
  AOI22_X2 U1497 ( .A1(net231315), .A2(MEM_WB_OUT[142]), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N37), .ZN(n1435) );
  AOI22_X2 U1499 ( .A1(net231315), .A2(MEM_WB_OUT[141]), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N38), .ZN(n1436) );
  AOI22_X2 U1501 ( .A1(net231315), .A2(MEM_WB_OUT[140]), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N39), .ZN(n1437) );
  AOI22_X2 U1504 ( .A1(net231315), .A2(MEM_WB_OUT[139]), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N40), .ZN(n1440) );
  AOI22_X2 U1506 ( .A1(net231315), .A2(MEM_WB_OUT[138]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N41), .ZN(n1441) );
  AOI22_X2 U1508 ( .A1(net231315), .A2(MEM_WB_OUT[137]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N42), .ZN(n1442) );
  AOI22_X2 U1510 ( .A1(net231297), .A2(MEM_WB_OUT[136]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N43), .ZN(n1443) );
  AOI22_X2 U1512 ( .A1(net231297), .A2(MEM_WB_OUT[135]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N44), .ZN(n1444) );
  AOI22_X2 U1514 ( .A1(net231315), .A2(MEM_WB_OUT[134]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N45), .ZN(n1445) );
  AOI22_X2 U1516 ( .A1(net231315), .A2(MEM_WB_OUT[133]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N46), .ZN(n1446) );
  AOI22_X2 U1518 ( .A1(net231297), .A2(MEM_WB_OUT[132]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N47), .ZN(n1447) );
  AOI22_X2 U1520 ( .A1(net231315), .A2(MEM_WB_OUT[131]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N48), .ZN(n1448) );
  AOI22_X2 U1522 ( .A1(net231297), .A2(MEM_WB_OUT[130]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N49), .ZN(n1449) );
  AOI22_X2 U1525 ( .A1(net231297), .A2(MEM_WB_OUT[129]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N50), .ZN(n1452) );
  AOI22_X2 U1527 ( .A1(net231297), .A2(MEM_WB_OUT[128]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N51), .ZN(n1453) );
  AOI22_X2 U1529 ( .A1(net231297), .A2(MEM_WB_OUT[127]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N52), .ZN(n1454) );
  AOI22_X2 U1531 ( .A1(net231297), .A2(MEM_WB_OUT[126]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N53), .ZN(n1455) );
  AOI22_X2 U1533 ( .A1(net231297), .A2(MEM_WB_OUT[125]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N54), .ZN(n1456) );
  AOI22_X2 U1535 ( .A1(net231297), .A2(MEM_WB_OUT[124]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N55), .ZN(n1457) );
  AOI22_X2 U1537 ( .A1(net231315), .A2(MEM_WB_OUT[123]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N56), .ZN(n1458) );
  AOI22_X2 U1539 ( .A1(net231297), .A2(MEM_WB_OUT[122]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N57), .ZN(n1459) );
  AOI22_X2 U1541 ( .A1(net231297), .A2(MEM_WB_OUT[121]), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N58), .ZN(n1460) );
  AOI22_X2 U1543 ( .A1(net231315), .A2(MEM_WB_OUT[120]), .B1(net231231), .B2(
        MEM_WB_REG_MEM_WB_REG_N59), .ZN(n1461) );
  AOI22_X2 U1546 ( .A1(net231315), .A2(MEM_WB_OUT[119]), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N60), .ZN(n1464) );
  AOI22_X2 U1548 ( .A1(net231301), .A2(MEM_WB_OUT[118]), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N61), .ZN(n1465) );
  AOI22_X2 U1550 ( .A1(net231297), .A2(MEM_WB_OUT[117]), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N62), .ZN(n1466) );
  AOI22_X2 U1552 ( .A1(net231315), .A2(MEM_WB_OUT[116]), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N63), .ZN(n1467) );
  AOI22_X2 U1554 ( .A1(net231297), .A2(MEM_WB_OUT[115]), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N64), .ZN(n1468) );
  AOI22_X2 U1556 ( .A1(net231315), .A2(MEM_WB_OUT[114]), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N65), .ZN(n1469) );
  AOI22_X2 U1558 ( .A1(net231297), .A2(MEM_WB_OUT[113]), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N66), .ZN(n1470) );
  OAI22_X2 U1559 ( .A1(net231239), .A2(n10947), .B1(net231313), .B2(n12202), 
        .ZN(n7916) );
  OAI22_X2 U1560 ( .A1(net231239), .A2(n10817), .B1(net231313), .B2(n12201), 
        .ZN(n7922) );
  OAI22_X2 U1561 ( .A1(net231239), .A2(n10353), .B1(net231313), .B2(n12200), 
        .ZN(n7928) );
  OAI22_X2 U1563 ( .A1(net231239), .A2(n10802), .B1(net231313), .B2(n12199), 
        .ZN(n7934) );
  OAI22_X2 U1564 ( .A1(net231239), .A2(n10845), .B1(net231313), .B2(n12198), 
        .ZN(n7942) );
  AOI22_X2 U1568 ( .A1(MEM_WB_OUT[104]), .A2(net231309), .B1(net231229), .B2(
        MEM_WB_REG_MEM_WB_REG_N75), .ZN(n1487) );
  OAI22_X2 U1574 ( .A1(n12534), .A2(net231259), .B1(net231311), .B2(n11112), 
        .ZN(n7329) );
  NAND2_X2 U1748 ( .A1(IMEM_BUS_IN[4]), .A2(n19164), .ZN(n1719) );
  OAI22_X2 U1828 ( .A1(net231241), .A2(n12218), .B1(n10828), .B2(net230373), 
        .ZN(n7966) );
  OAI22_X2 U1830 ( .A1(net231241), .A2(n12217), .B1(n10360), .B2(net230373), 
        .ZN(n7969) );
  OAI22_X2 U1845 ( .A1(net231241), .A2(n10357), .B1(n12196), .B2(net230373), 
        .ZN(n7507) );
  OAI22_X2 U1868 ( .A1(net231241), .A2(n10366), .B1(n12195), .B2(net230373), 
        .ZN(n7413) );
  OAI22_X2 U1890 ( .A1(net231241), .A2(n10356), .B1(n12194), .B2(net230373), 
        .ZN(n7502) );
  OAI22_X2 U1906 ( .A1(net231241), .A2(n12550), .B1(net231311), .B2(n1830), 
        .ZN(n7827) );
  NOR4_X2 U1907 ( .A1(n1831), .A2(n1832), .A3(n1833), .A4(n1834), .ZN(n1830)
         );
  OAI221_X2 U1908 ( .B1(n10251), .B2(n13744), .C1(n10689), .C2(n13742), .A(
        n1837), .ZN(n1834) );
  AOI22_X2 U1909 ( .A1(n13187), .A2(REG_FILE_reg_out_29__31_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__31_), .ZN(n1837) );
  OAI221_X2 U1911 ( .B1(n10847), .B2(n13740), .C1(n10461), .C2(n13738), .A(
        n1842), .ZN(n1833) );
  NAND4_X2 U1921 ( .A1(n1858), .A2(n1859), .A3(n1860), .A4(n1861), .ZN(n1831)
         );
  AOI221_X2 U1929 ( .B1(n19154), .B2(REG_FILE_reg_out_26__31_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__31_), .A(n1875), .ZN(n1859) );
  AOI221_X2 U1932 ( .B1(n13495), .B2(REG_FILE_reg_out_13__31_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__31_), .A(n1880), .ZN(n1858) );
  OAI22_X2 U1933 ( .A1(n12025), .A2(n13178), .B1(n10530), .B2(n13732), .ZN(
        n1880) );
  OAI22_X2 U1935 ( .A1(net231241), .A2(n12549), .B1(net231311), .B2(n1884), 
        .ZN(n7736) );
  NOR4_X2 U1936 ( .A1(n1885), .A2(n1886), .A3(n1887), .A4(n1888), .ZN(n1884)
         );
  OAI221_X2 U1937 ( .B1(n10300), .B2(n13745), .C1(n11895), .C2(n13742), .A(
        n1889), .ZN(n1888) );
  AOI22_X2 U1938 ( .A1(n13187), .A2(REG_FILE_reg_out_29__30_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__30_), .ZN(n1889) );
  OAI221_X2 U1940 ( .B1(n10926), .B2(n13740), .C1(n10749), .C2(n13739), .A(
        n1890), .ZN(n1887) );
  NAND4_X2 U1950 ( .A1(n1895), .A2(n1896), .A3(n1897), .A4(n1898), .ZN(n1885)
         );
  AOI221_X2 U1958 ( .B1(n19154), .B2(REG_FILE_reg_out_26__30_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__30_), .A(n1901), .ZN(n1896) );
  AOI221_X2 U1961 ( .B1(n13495), .B2(REG_FILE_reg_out_13__30_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__30_), .A(n1902), .ZN(n1895) );
  OAI22_X2 U1962 ( .A1(n12049), .A2(n13178), .B1(n10529), .B2(n13732), .ZN(
        n1902) );
  OAI22_X2 U1964 ( .A1(net231241), .A2(n12301), .B1(net231311), .B2(n1904), 
        .ZN(n7721) );
  NOR4_X2 U1965 ( .A1(n1905), .A2(n1906), .A3(n1907), .A4(n1908), .ZN(n1904)
         );
  OAI221_X2 U1966 ( .B1(n10299), .B2(n13744), .C1(n11894), .C2(n13742), .A(
        n1909), .ZN(n1908) );
  AOI22_X2 U1967 ( .A1(n13187), .A2(REG_FILE_reg_out_29__29_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__29_), .ZN(n1909) );
  OAI221_X2 U1969 ( .B1(n10925), .B2(n13740), .C1(n10748), .C2(n13738), .A(
        n1910), .ZN(n1907) );
  NAND4_X2 U1979 ( .A1(n1915), .A2(n1916), .A3(n1917), .A4(n1918), .ZN(n1905)
         );
  AOI221_X2 U1987 ( .B1(n19154), .B2(REG_FILE_reg_out_26__29_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__29_), .A(n1921), .ZN(n1916) );
  AOI221_X2 U1990 ( .B1(n13495), .B2(REG_FILE_reg_out_13__29_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__29_), .A(n1922), .ZN(n1915) );
  OAI22_X2 U1991 ( .A1(n12048), .A2(n13178), .B1(n10528), .B2(n13732), .ZN(
        n1922) );
  OAI22_X2 U1993 ( .A1(net231241), .A2(n12231), .B1(net231311), .B2(n1924), 
        .ZN(n7686) );
  NOR4_X2 U1994 ( .A1(n1925), .A2(n1926), .A3(n1927), .A4(n1928), .ZN(n1924)
         );
  OAI221_X2 U1995 ( .B1(n10298), .B2(n13745), .C1(n11893), .C2(n13742), .A(
        n1929), .ZN(n1928) );
  AOI22_X2 U1996 ( .A1(n13187), .A2(REG_FILE_reg_out_29__28_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__28_), .ZN(n1929) );
  OAI221_X2 U1998 ( .B1(n10924), .B2(n13740), .C1(n10747), .C2(n13739), .A(
        n1930), .ZN(n1927) );
  NAND4_X2 U2008 ( .A1(n1935), .A2(n1936), .A3(n1937), .A4(n1938), .ZN(n1925)
         );
  AOI221_X2 U2016 ( .B1(n19154), .B2(REG_FILE_reg_out_26__28_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__28_), .A(n1941), .ZN(n1936) );
  AOI221_X2 U2019 ( .B1(n13495), .B2(REG_FILE_reg_out_13__28_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__28_), .A(n1942), .ZN(n1935) );
  OAI22_X2 U2020 ( .A1(n12047), .A2(n13178), .B1(n10527), .B2(n13732), .ZN(
        n1942) );
  OAI22_X2 U2022 ( .A1(net231241), .A2(n10355), .B1(n12193), .B2(net230373), 
        .ZN(n7497) );
  OAI22_X2 U2024 ( .A1(net231241), .A2(n12230), .B1(net231311), .B2(n1945), 
        .ZN(n7677) );
  NOR4_X2 U2025 ( .A1(n1946), .A2(n1947), .A3(n1948), .A4(n1949), .ZN(n1945)
         );
  OAI221_X2 U2026 ( .B1(n10297), .B2(n13745), .C1(n11892), .C2(n13742), .A(
        n1950), .ZN(n1949) );
  AOI22_X2 U2027 ( .A1(n13187), .A2(REG_FILE_reg_out_29__27_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__27_), .ZN(n1950) );
  OAI221_X2 U2029 ( .B1(n10923), .B2(n13740), .C1(n10746), .C2(n13738), .A(
        n1951), .ZN(n1948) );
  NAND4_X2 U2039 ( .A1(n1956), .A2(n1957), .A3(n1958), .A4(n1959), .ZN(n1946)
         );
  AOI221_X2 U2047 ( .B1(n19154), .B2(REG_FILE_reg_out_26__27_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__27_), .A(n1962), .ZN(n1957) );
  AOI221_X2 U2050 ( .B1(n13495), .B2(REG_FILE_reg_out_13__27_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__27_), .A(n1963), .ZN(n1956) );
  OAI22_X2 U2051 ( .A1(n12046), .A2(n13178), .B1(n10526), .B2(n13732), .ZN(
        n1963) );
  OAI22_X2 U2053 ( .A1(net231241), .A2(n12525), .B1(net231311), .B2(n1965), 
        .ZN(n7669) );
  NOR4_X2 U2054 ( .A1(n1966), .A2(n1967), .A3(n1968), .A4(n1969), .ZN(n1965)
         );
  OAI221_X2 U2055 ( .B1(n10296), .B2(n13745), .C1(n11891), .C2(n13742), .A(
        n1970), .ZN(n1969) );
  AOI22_X2 U2056 ( .A1(n13187), .A2(REG_FILE_reg_out_29__26_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__26_), .ZN(n1970) );
  OAI221_X2 U2058 ( .B1(n10922), .B2(n13740), .C1(n10745), .C2(n13739), .A(
        n1971), .ZN(n1968) );
  NAND4_X2 U2068 ( .A1(n1976), .A2(n1977), .A3(n1978), .A4(n1979), .ZN(n1966)
         );
  AOI221_X2 U2076 ( .B1(n19154), .B2(REG_FILE_reg_out_26__26_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__26_), .A(n1982), .ZN(n1977) );
  AOI221_X2 U2079 ( .B1(n13495), .B2(REG_FILE_reg_out_13__26_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__26_), .A(n1983), .ZN(n1976) );
  OAI22_X2 U2080 ( .A1(n12045), .A2(n13178), .B1(n10525), .B2(n13732), .ZN(
        n1983) );
  OAI22_X2 U2082 ( .A1(net231241), .A2(n12524), .B1(net231311), .B2(n1985), 
        .ZN(n7660) );
  NOR4_X2 U2083 ( .A1(n1986), .A2(n1987), .A3(n1988), .A4(n1989), .ZN(n1985)
         );
  OAI221_X2 U2084 ( .B1(n10295), .B2(n13745), .C1(n11890), .C2(n13742), .A(
        n1990), .ZN(n1989) );
  AOI22_X2 U2085 ( .A1(n13187), .A2(REG_FILE_reg_out_29__25_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__25_), .ZN(n1990) );
  OAI221_X2 U2087 ( .B1(n10921), .B2(n13740), .C1(n10744), .C2(n13738), .A(
        n1991), .ZN(n1988) );
  NAND4_X2 U2097 ( .A1(n1996), .A2(n1997), .A3(n1998), .A4(n1999), .ZN(n1986)
         );
  AOI221_X2 U2105 ( .B1(n19154), .B2(REG_FILE_reg_out_26__25_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__25_), .A(n2002), .ZN(n1997) );
  AOI221_X2 U2108 ( .B1(n13495), .B2(REG_FILE_reg_out_13__25_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__25_), .A(n2003), .ZN(n1996) );
  OAI22_X2 U2109 ( .A1(n12044), .A2(n13178), .B1(n10524), .B2(n13732), .ZN(
        n2003) );
  OAI22_X2 U2111 ( .A1(net231241), .A2(n12548), .B1(net231311), .B2(n2005), 
        .ZN(n7651) );
  NOR4_X2 U2112 ( .A1(n2006), .A2(n2007), .A3(n2008), .A4(n2009), .ZN(n2005)
         );
  OAI221_X2 U2113 ( .B1(n10294), .B2(n13745), .C1(n11889), .C2(n13742), .A(
        n2010), .ZN(n2009) );
  AOI22_X2 U2114 ( .A1(n13187), .A2(REG_FILE_reg_out_29__24_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__24_), .ZN(n2010) );
  OAI221_X2 U2116 ( .B1(n10920), .B2(n13740), .C1(n10743), .C2(n13739), .A(
        n2011), .ZN(n2008) );
  NAND4_X2 U2126 ( .A1(n2016), .A2(n2017), .A3(n2018), .A4(n2019), .ZN(n2006)
         );
  AOI221_X2 U2134 ( .B1(n19154), .B2(REG_FILE_reg_out_26__24_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__24_), .A(n2022), .ZN(n2017) );
  AOI221_X2 U2137 ( .B1(n13495), .B2(REG_FILE_reg_out_13__24_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__24_), .A(n2023), .ZN(n2016) );
  OAI22_X2 U2138 ( .A1(n12043), .A2(n13178), .B1(n10523), .B2(n13732), .ZN(
        n2023) );
  OAI22_X2 U2140 ( .A1(net231241), .A2(n12211), .B1(net231311), .B2(n2025), 
        .ZN(n7635) );
  NOR4_X2 U2141 ( .A1(n2026), .A2(n2027), .A3(n2028), .A4(n2029), .ZN(n2025)
         );
  OAI221_X2 U2142 ( .B1(n10293), .B2(n13745), .C1(n11888), .C2(n13742), .A(
        n2030), .ZN(n2029) );
  AOI22_X2 U2143 ( .A1(n13187), .A2(REG_FILE_reg_out_29__23_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__23_), .ZN(n2030) );
  OAI221_X2 U2145 ( .B1(n10919), .B2(n13740), .C1(n10742), .C2(n13739), .A(
        n2031), .ZN(n2028) );
  NAND4_X2 U2155 ( .A1(n2036), .A2(n2037), .A3(n2038), .A4(n2039), .ZN(n2026)
         );
  AOI221_X2 U2163 ( .B1(n19154), .B2(REG_FILE_reg_out_26__23_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__23_), .A(n2042), .ZN(n2037) );
  AOI221_X2 U2166 ( .B1(n13495), .B2(REG_FILE_reg_out_13__23_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__23_), .A(n2043), .ZN(n2036) );
  OAI22_X2 U2167 ( .A1(n12042), .A2(n13178), .B1(n10522), .B2(n13732), .ZN(
        n2043) );
  OAI221_X2 U2171 ( .B1(n10292), .B2(n13744), .C1(n12815), .C2(n13742), .A(
        n2050), .ZN(n2049) );
  AOI22_X2 U2172 ( .A1(n13187), .A2(REG_FILE_reg_out_29__22_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__22_), .ZN(n2050) );
  OAI221_X2 U2174 ( .B1(n10918), .B2(n13740), .C1(n10741), .C2(n13739), .A(
        n2051), .ZN(n2048) );
  NAND4_X2 U2184 ( .A1(n2056), .A2(n2057), .A3(n2058), .A4(n2059), .ZN(n2046)
         );
  AOI221_X2 U2192 ( .B1(n19154), .B2(REG_FILE_reg_out_26__22_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__22_), .A(n2062), .ZN(n2057) );
  AOI221_X2 U2195 ( .B1(n13495), .B2(REG_FILE_reg_out_13__22_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__22_), .A(n2063), .ZN(n2056) );
  OAI22_X2 U2196 ( .A1(n10321), .A2(n13178), .B1(n10521), .B2(n13732), .ZN(
        n2063) );
  OAI221_X2 U2199 ( .B1(n10503), .B2(n13744), .C1(n12813), .C2(n13742), .A(
        n2070), .ZN(n2069) );
  AOI22_X2 U2200 ( .A1(n13187), .A2(REG_FILE_reg_out_29__21_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__21_), .ZN(n2070) );
  OAI221_X2 U2202 ( .B1(n10502), .B2(n13740), .C1(n11420), .C2(n13739), .A(
        n2071), .ZN(n2068) );
  NAND4_X2 U2212 ( .A1(n2076), .A2(n2077), .A3(n2078), .A4(n2079), .ZN(n2066)
         );
  AOI221_X2 U2220 ( .B1(n19154), .B2(REG_FILE_reg_out_26__21_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__21_), .A(n2082), .ZN(n2077) );
  AOI221_X2 U2223 ( .B1(n13495), .B2(REG_FILE_reg_out_13__21_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__21_), .A(n2083), .ZN(n2076) );
  OAI22_X2 U2224 ( .A1(n10320), .A2(n13178), .B1(n10932), .B2(n13732), .ZN(
        n2083) );
  OAI221_X2 U2227 ( .B1(n10501), .B2(n13744), .C1(n12811), .C2(n13742), .A(
        n2090), .ZN(n2089) );
  AOI22_X2 U2228 ( .A1(n13187), .A2(REG_FILE_reg_out_29__20_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__20_), .ZN(n2090) );
  OAI221_X2 U2230 ( .B1(n10500), .B2(n13741), .C1(n11419), .C2(n13738), .A(
        n2091), .ZN(n2088) );
  NAND4_X2 U2240 ( .A1(n2096), .A2(n2097), .A3(n2098), .A4(n2099), .ZN(n2086)
         );
  AOI221_X2 U2248 ( .B1(n19154), .B2(REG_FILE_reg_out_26__20_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__20_), .A(n2102), .ZN(n2097) );
  AOI221_X2 U2251 ( .B1(n13496), .B2(REG_FILE_reg_out_13__20_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__20_), .A(n2103), .ZN(n2096) );
  OAI22_X2 U2252 ( .A1(n10319), .A2(n13178), .B1(n10931), .B2(n13733), .ZN(
        n2103) );
  OAI221_X2 U2255 ( .B1(n10499), .B2(n13744), .C1(n12809), .C2(n13742), .A(
        n2110), .ZN(n2109) );
  AOI22_X2 U2256 ( .A1(n13187), .A2(REG_FILE_reg_out_29__19_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__19_), .ZN(n2110) );
  OAI221_X2 U2258 ( .B1(n10498), .B2(n13741), .C1(n11418), .C2(n13738), .A(
        n2111), .ZN(n2108) );
  NAND4_X2 U2268 ( .A1(n2116), .A2(n2117), .A3(n2118), .A4(n2119), .ZN(n2106)
         );
  AOI221_X2 U2277 ( .B1(n19154), .B2(REG_FILE_reg_out_26__19_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__19_), .A(n2122), .ZN(n2117) );
  AOI221_X2 U2280 ( .B1(n13496), .B2(REG_FILE_reg_out_13__19_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__19_), .A(n2123), .ZN(n2116) );
  OAI22_X2 U2281 ( .A1(n10318), .A2(n13178), .B1(n10930), .B2(n13733), .ZN(
        n2123) );
  OAI221_X2 U2284 ( .B1(n10497), .B2(n13744), .C1(n12807), .C2(n13742), .A(
        n2130), .ZN(n2129) );
  AOI22_X2 U2285 ( .A1(n13187), .A2(REG_FILE_reg_out_29__18_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__18_), .ZN(n2130) );
  OAI221_X2 U2287 ( .B1(n10496), .B2(n13741), .C1(n11417), .C2(n13738), .A(
        n2131), .ZN(n2128) );
  NAND4_X2 U2297 ( .A1(n2136), .A2(n2137), .A3(n2138), .A4(n2139), .ZN(n2126)
         );
  AOI221_X2 U2306 ( .B1(n19154), .B2(REG_FILE_reg_out_26__18_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__18_), .A(n2142), .ZN(n2137) );
  AOI221_X2 U2309 ( .B1(n13496), .B2(REG_FILE_reg_out_13__18_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__18_), .A(n2143), .ZN(n2136) );
  OAI22_X2 U2310 ( .A1(n10317), .A2(n13178), .B1(n10929), .B2(n13733), .ZN(
        n2143) );
  OAI22_X2 U2311 ( .A1(net231241), .A2(n11914), .B1(n19327), .B2(net230373), 
        .ZN(n7553) );
  OAI221_X2 U2315 ( .B1(n10495), .B2(n13744), .C1(n12803), .C2(n13742), .A(
        n2151), .ZN(n2150) );
  AOI22_X2 U2316 ( .A1(n13187), .A2(REG_FILE_reg_out_29__17_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__17_), .ZN(n2151) );
  OAI221_X2 U2318 ( .B1(n10494), .B2(n13741), .C1(n11416), .C2(n13738), .A(
        n2152), .ZN(n2149) );
  NAND4_X2 U2328 ( .A1(n2157), .A2(n2158), .A3(n2159), .A4(n2160), .ZN(n2147)
         );
  AOI221_X2 U2337 ( .B1(n19154), .B2(REG_FILE_reg_out_26__17_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__17_), .A(n2163), .ZN(n2158) );
  AOI221_X2 U2340 ( .B1(n13496), .B2(REG_FILE_reg_out_13__17_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__17_), .A(n2164), .ZN(n2157) );
  OAI22_X2 U2341 ( .A1(n10316), .A2(n13178), .B1(n10928), .B2(n13733), .ZN(
        n2164) );
  OAI22_X2 U2342 ( .A1(net231243), .A2(n12131), .B1(net231311), .B2(n2166), 
        .ZN(n7470) );
  NOR4_X2 U2343 ( .A1(n2167), .A2(n2168), .A3(n2169), .A4(n2170), .ZN(n2166)
         );
  OAI221_X2 U2344 ( .B1(n10493), .B2(n13744), .C1(n12798), .C2(n13742), .A(
        n2171), .ZN(n2170) );
  AOI22_X2 U2345 ( .A1(n13187), .A2(REG_FILE_reg_out_29__16_), .B1(n10354), 
        .B2(REG_FILE_reg_out_6__16_), .ZN(n2171) );
  OAI221_X2 U2347 ( .B1(n10492), .B2(n13741), .C1(n11415), .C2(n13738), .A(
        n2172), .ZN(n2169) );
  NAND4_X2 U2357 ( .A1(n2177), .A2(n2178), .A3(n2179), .A4(n2180), .ZN(n2167)
         );
  AOI221_X2 U2369 ( .B1(n19154), .B2(REG_FILE_reg_out_26__16_), .C1(n19155), 
        .C2(REG_FILE_reg_out_25__16_), .A(n2185), .ZN(n2178) );
  AOI221_X2 U2374 ( .B1(n13496), .B2(REG_FILE_reg_out_13__16_), .C1(n19160), 
        .C2(REG_FILE_reg_out_27__16_), .A(n2188), .ZN(n2177) );
  OAI22_X2 U2375 ( .A1(n10520), .A2(n13178), .B1(n10927), .B2(n13733), .ZN(
        n2188) );
  OAI221_X2 U2380 ( .B1(n11372), .B2(n13735), .C1(n10688), .C2(n13182), .A(
        n2196), .ZN(n2195) );
  OAI221_X2 U2383 ( .B1(n10846), .B2(n13730), .C1(n12024), .C2(n13727), .A(
        n2198), .ZN(n2194) );
  NAND2_X2 U2385 ( .A1(n2201), .A2(n2202), .ZN(n2193) );
  AOI221_X2 U2386 ( .B1(n19157), .B2(REG_FILE_reg_out_19__15_), .C1(n13496), 
        .C2(REG_FILE_reg_out_13__15_), .A(n2204), .ZN(n2202) );
  AOI221_X2 U2390 ( .B1(n19159), .B2(REG_FILE_reg_out_3__15_), .C1(n13499), 
        .C2(REG_FILE_reg_out_4__15_), .A(n2206), .ZN(n2201) );
  OAI22_X2 U2391 ( .A1(n12041), .A2(n13733), .B1(n10905), .B2(n13176), .ZN(
        n2206) );
  OAI22_X2 U2394 ( .A1(n10504), .A2(n13738), .B1(n10904), .B2(n13741), .ZN(
        n2211) );
  OAI22_X2 U2396 ( .A1(n11414), .A2(n13742), .B1(n10396), .B2(n13744), .ZN(
        n2212) );
  OAI22_X2 U2405 ( .A1(net231243), .A2(n12210), .B1(net231311), .B2(n2216), 
        .ZN(n7453) );
  NOR4_X2 U2406 ( .A1(n2217), .A2(n2218), .A3(n2219), .A4(n2220), .ZN(n2216)
         );
  OAI221_X2 U2407 ( .B1(n11371), .B2(n13735), .C1(n10687), .C2(n13182), .A(
        n2221), .ZN(n2220) );
  OAI221_X2 U2410 ( .B1(n10380), .B2(n13730), .C1(n10856), .C2(n13727), .A(
        n2222), .ZN(n2219) );
  NAND2_X2 U2412 ( .A1(n2223), .A2(n2224), .ZN(n2218) );
  AOI221_X2 U2413 ( .B1(n19157), .B2(REG_FILE_reg_out_19__14_), .C1(n13496), 
        .C2(REG_FILE_reg_out_13__14_), .A(n2225), .ZN(n2224) );
  AOI221_X2 U2417 ( .B1(n19159), .B2(REG_FILE_reg_out_3__14_), .C1(n13499), 
        .C2(REG_FILE_reg_out_4__14_), .A(n2226), .ZN(n2223) );
  OAI22_X2 U2418 ( .A1(n10519), .A2(n13733), .B1(n10903), .B2(n13176), .ZN(
        n2226) );
  OAI22_X2 U2421 ( .A1(n10315), .A2(n13738), .B1(n10902), .B2(n13741), .ZN(
        n2231) );
  OAI22_X2 U2423 ( .A1(n11413), .A2(n13743), .B1(n10395), .B2(n13744), .ZN(
        n2232) );
  OAI221_X2 U2435 ( .B1(n11370), .B2(n13735), .C1(n10686), .C2(n13182), .A(
        n2241), .ZN(n2240) );
  OAI221_X2 U2438 ( .B1(n10379), .B2(n13730), .C1(n10855), .C2(n13727), .A(
        n2242), .ZN(n2239) );
  NAND2_X2 U2440 ( .A1(n2243), .A2(n2244), .ZN(n2238) );
  AOI221_X2 U2441 ( .B1(n19157), .B2(REG_FILE_reg_out_19__13_), .C1(n13496), 
        .C2(REG_FILE_reg_out_13__13_), .A(n2245), .ZN(n2244) );
  AOI221_X2 U2445 ( .B1(n19159), .B2(REG_FILE_reg_out_3__13_), .C1(n13499), 
        .C2(REG_FILE_reg_out_4__13_), .A(n2246), .ZN(n2243) );
  OAI22_X2 U2446 ( .A1(n10518), .A2(n13733), .B1(n10901), .B2(n13176), .ZN(
        n2246) );
  OAI22_X2 U2449 ( .A1(n10314), .A2(n13738), .B1(n10900), .B2(n13741), .ZN(
        n2251) );
  OAI22_X2 U2451 ( .A1(n11412), .A2(n13742), .B1(n10394), .B2(n13744), .ZN(
        n2252) );
  OAI22_X2 U2460 ( .A1(net231243), .A2(n12209), .B1(net231311), .B2(n2256), 
        .ZN(n7428) );
  NOR4_X2 U2461 ( .A1(n2257), .A2(n2258), .A3(n2259), .A4(n2260), .ZN(n2256)
         );
  OAI221_X2 U2462 ( .B1(n11369), .B2(n13735), .C1(n10685), .C2(n13182), .A(
        n2261), .ZN(n2260) );
  OAI221_X2 U2465 ( .B1(n10378), .B2(n13730), .C1(n10854), .C2(n13727), .A(
        n2262), .ZN(n2259) );
  NAND2_X2 U2467 ( .A1(n2263), .A2(n2264), .ZN(n2258) );
  AOI221_X2 U2468 ( .B1(n19157), .B2(REG_FILE_reg_out_19__12_), .C1(n13496), 
        .C2(REG_FILE_reg_out_13__12_), .A(n2265), .ZN(n2264) );
  AOI221_X2 U2472 ( .B1(n19159), .B2(REG_FILE_reg_out_3__12_), .C1(n13499), 
        .C2(REG_FILE_reg_out_4__12_), .A(n2266), .ZN(n2263) );
  OAI22_X2 U2473 ( .A1(n10517), .A2(n13733), .B1(n10899), .B2(n13176), .ZN(
        n2266) );
  OAI22_X2 U2476 ( .A1(n10313), .A2(n13738), .B1(n10898), .B2(n13741), .ZN(
        n2271) );
  OAI22_X2 U2478 ( .A1(n11411), .A2(n13743), .B1(n10393), .B2(n13744), .ZN(
        n2272) );
  OAI221_X2 U2490 ( .B1(n11368), .B2(n13735), .C1(n10684), .C2(n13182), .A(
        n2281), .ZN(n2280) );
  OAI221_X2 U2493 ( .B1(n10377), .B2(n13730), .C1(n10853), .C2(n13727), .A(
        n2282), .ZN(n2279) );
  NAND2_X2 U2495 ( .A1(n2283), .A2(n2284), .ZN(n2278) );
  AOI221_X2 U2496 ( .B1(n19157), .B2(REG_FILE_reg_out_19__11_), .C1(n13496), 
        .C2(REG_FILE_reg_out_13__11_), .A(n2285), .ZN(n2284) );
  AOI221_X2 U2500 ( .B1(n19159), .B2(REG_FILE_reg_out_3__11_), .C1(n13499), 
        .C2(REG_FILE_reg_out_4__11_), .A(n2286), .ZN(n2283) );
  OAI22_X2 U2501 ( .A1(n10516), .A2(n13733), .B1(n10897), .B2(n13176), .ZN(
        n2286) );
  OAI22_X2 U2504 ( .A1(n10312), .A2(n13738), .B1(n10896), .B2(n13741), .ZN(
        n2291) );
  OAI22_X2 U2506 ( .A1(n11410), .A2(n13742), .B1(n10392), .B2(n13744), .ZN(
        n2292) );
  OAI221_X2 U2517 ( .B1(n11367), .B2(n13735), .C1(n10683), .C2(n13182), .A(
        n2301), .ZN(n2300) );
  OAI221_X2 U2520 ( .B1(n10376), .B2(n13730), .C1(n10852), .C2(n13727), .A(
        n2302), .ZN(n2299) );
  NAND2_X2 U2522 ( .A1(n2303), .A2(n2304), .ZN(n2298) );
  AOI221_X2 U2523 ( .B1(n19157), .B2(REG_FILE_reg_out_19__10_), .C1(n13496), 
        .C2(REG_FILE_reg_out_13__10_), .A(n2305), .ZN(n2304) );
  AOI221_X2 U2527 ( .B1(n19159), .B2(REG_FILE_reg_out_3__10_), .C1(n13499), 
        .C2(REG_FILE_reg_out_4__10_), .A(n2306), .ZN(n2303) );
  OAI22_X2 U2528 ( .A1(n10515), .A2(n13733), .B1(n10895), .B2(n13176), .ZN(
        n2306) );
  OAI22_X2 U2531 ( .A1(n10311), .A2(n13738), .B1(n10894), .B2(n13741), .ZN(
        n2311) );
  OAI22_X2 U2533 ( .A1(n11409), .A2(n13742), .B1(n10391), .B2(n13744), .ZN(
        n2312) );
  OAI221_X2 U2544 ( .B1(n11366), .B2(n13735), .C1(n10682), .C2(n13182), .A(
        n2321), .ZN(n2320) );
  OAI221_X2 U2547 ( .B1(n10375), .B2(n13730), .C1(n10851), .C2(n13727), .A(
        n2322), .ZN(n2319) );
  NAND2_X2 U2549 ( .A1(n2323), .A2(n2324), .ZN(n2318) );
  AOI221_X2 U2550 ( .B1(n19157), .B2(REG_FILE_reg_out_19__9_), .C1(n13496), 
        .C2(REG_FILE_reg_out_13__9_), .A(n2325), .ZN(n2324) );
  AOI221_X2 U2554 ( .B1(n19159), .B2(REG_FILE_reg_out_3__9_), .C1(n13499), 
        .C2(REG_FILE_reg_out_4__9_), .A(n2326), .ZN(n2323) );
  OAI22_X2 U2555 ( .A1(n10514), .A2(n13732), .B1(n10893), .B2(n13176), .ZN(
        n2326) );
  OAI22_X2 U2558 ( .A1(n10310), .A2(n13738), .B1(n10892), .B2(n13741), .ZN(
        n2331) );
  OAI22_X2 U2560 ( .A1(n11408), .A2(n13742), .B1(n10390), .B2(n13744), .ZN(
        n2332) );
  OAI22_X2 U2569 ( .A1(net231243), .A2(n12208), .B1(net231311), .B2(n2336), 
        .ZN(n7381) );
  NOR4_X2 U2570 ( .A1(n2337), .A2(n2338), .A3(n2339), .A4(n2340), .ZN(n2336)
         );
  OAI221_X2 U2571 ( .B1(n11365), .B2(n13735), .C1(n10681), .C2(n13182), .A(
        n2341), .ZN(n2340) );
  OAI221_X2 U2574 ( .B1(n10374), .B2(n13730), .C1(n10850), .C2(n13727), .A(
        n2342), .ZN(n2339) );
  NAND2_X2 U2576 ( .A1(n2343), .A2(n2344), .ZN(n2338) );
  AOI221_X2 U2577 ( .B1(n19157), .B2(REG_FILE_reg_out_19__8_), .C1(n13496), 
        .C2(REG_FILE_reg_out_13__8_), .A(n2345), .ZN(n2344) );
  AOI221_X2 U2581 ( .B1(n19159), .B2(REG_FILE_reg_out_3__8_), .C1(n13499), 
        .C2(REG_FILE_reg_out_4__8_), .A(n2346), .ZN(n2343) );
  OAI22_X2 U2582 ( .A1(n10513), .A2(n13732), .B1(n10891), .B2(n13176), .ZN(
        n2346) );
  OAI22_X2 U2585 ( .A1(n10309), .A2(n13739), .B1(n10890), .B2(n13740), .ZN(
        n2351) );
  OAI22_X2 U2587 ( .A1(n12289), .A2(n13743), .B1(n10889), .B2(n13745), .ZN(
        n2352) );
  OAI22_X2 U2597 ( .A1(net231243), .A2(n10364), .B1(n12305), .B2(net230373), 
        .ZN(n7492) );
  OAI22_X2 U2599 ( .A1(net231243), .A2(n12179), .B1(net231311), .B2(n2357), 
        .ZN(n7410) );
  NOR4_X2 U2600 ( .A1(n2358), .A2(n2359), .A3(n2360), .A4(n2361), .ZN(n2357)
         );
  OAI221_X2 U2601 ( .B1(n11364), .B2(n13735), .C1(n10680), .C2(n13182), .A(
        n2362), .ZN(n2361) );
  OAI221_X2 U2604 ( .B1(n10373), .B2(n13730), .C1(n10849), .C2(n13727), .A(
        n2363), .ZN(n2360) );
  NAND2_X2 U2606 ( .A1(n2364), .A2(n2365), .ZN(n2359) );
  AOI221_X2 U2607 ( .B1(n19157), .B2(REG_FILE_reg_out_19__7_), .C1(n13495), 
        .C2(REG_FILE_reg_out_13__7_), .A(n2366), .ZN(n2365) );
  AOI221_X2 U2611 ( .B1(n19159), .B2(REG_FILE_reg_out_3__7_), .C1(n13499), 
        .C2(REG_FILE_reg_out_4__7_), .A(n2367), .ZN(n2364) );
  OAI22_X2 U2612 ( .A1(n10512), .A2(n13733), .B1(n10888), .B2(n13176), .ZN(
        n2367) );
  OAI22_X2 U2615 ( .A1(n10308), .A2(n13739), .B1(n10887), .B2(n13741), .ZN(
        n2372) );
  OAI22_X2 U2617 ( .A1(n12288), .A2(n13743), .B1(n10886), .B2(n13745), .ZN(
        n2373) );
  OAI221_X2 U2629 ( .B1(n11363), .B2(n13735), .C1(n10679), .C2(n13182), .A(
        n2382), .ZN(n2381) );
  OAI221_X2 U2632 ( .B1(n10372), .B2(n13730), .C1(n10848), .C2(n13727), .A(
        n2383), .ZN(n2380) );
  NAND2_X2 U2634 ( .A1(n2384), .A2(n2385), .ZN(n2379) );
  AOI221_X2 U2635 ( .B1(n19157), .B2(REG_FILE_reg_out_19__6_), .C1(n13496), 
        .C2(REG_FILE_reg_out_13__6_), .A(n2386), .ZN(n2385) );
  AOI221_X2 U2639 ( .B1(n19159), .B2(REG_FILE_reg_out_3__6_), .C1(n13499), 
        .C2(REG_FILE_reg_out_4__6_), .A(n2387), .ZN(n2384) );
  OAI22_X2 U2640 ( .A1(n10511), .A2(n13733), .B1(n10885), .B2(n13176), .ZN(
        n2387) );
  OAI22_X2 U2643 ( .A1(n10307), .A2(n13739), .B1(n10884), .B2(n13741), .ZN(
        n2392) );
  OAI22_X2 U2645 ( .A1(n12287), .A2(n13743), .B1(n10883), .B2(n13745), .ZN(
        n2393) );
  OAI22_X2 U2654 ( .A1(net231243), .A2(n12207), .B1(net231311), .B2(n2397), 
        .ZN(n7365) );
  NOR4_X2 U2655 ( .A1(n2398), .A2(n2399), .A3(n2400), .A4(n2401), .ZN(n2397)
         );
  OAI221_X2 U2656 ( .B1(n11362), .B2(n13735), .C1(n10678), .C2(n13182), .A(
        n2402), .ZN(n2401) );
  OAI221_X2 U2659 ( .B1(n10250), .B2(n13730), .C1(n10385), .C2(n13727), .A(
        n2403), .ZN(n2400) );
  NAND2_X2 U2661 ( .A1(n2404), .A2(n2405), .ZN(n2399) );
  AOI221_X2 U2662 ( .B1(n19157), .B2(REG_FILE_reg_out_19__5_), .C1(n13496), 
        .C2(REG_FILE_reg_out_13__5_), .A(n2406), .ZN(n2405) );
  AOI221_X2 U2666 ( .B1(n19159), .B2(REG_FILE_reg_out_3__5_), .C1(n13499), 
        .C2(REG_FILE_reg_out_4__5_), .A(n2407), .ZN(n2404) );
  OAI22_X2 U2667 ( .A1(n10510), .A2(n13732), .B1(n10882), .B2(n13176), .ZN(
        n2407) );
  OAI22_X2 U2670 ( .A1(n10306), .A2(n13739), .B1(n10881), .B2(n13740), .ZN(
        n2412) );
  OAI22_X2 U2672 ( .A1(n12286), .A2(n13743), .B1(n10880), .B2(n13745), .ZN(
        n2413) );
  OAI221_X2 U2684 ( .B1(n11361), .B2(n13735), .C1(n10677), .C2(n13182), .A(
        n2422), .ZN(n2421) );
  OAI221_X2 U2687 ( .B1(n10249), .B2(n13730), .C1(n10384), .C2(n13727), .A(
        n2423), .ZN(n2420) );
  NAND2_X2 U2689 ( .A1(n2424), .A2(n2425), .ZN(n2419) );
  AOI221_X2 U2690 ( .B1(n19157), .B2(REG_FILE_reg_out_19__4_), .C1(n13495), 
        .C2(REG_FILE_reg_out_13__4_), .A(n2426), .ZN(n2425) );
  AOI221_X2 U2694 ( .B1(n19159), .B2(REG_FILE_reg_out_3__4_), .C1(n13499), 
        .C2(REG_FILE_reg_out_4__4_), .A(n2427), .ZN(n2424) );
  OAI22_X2 U2695 ( .A1(n10509), .A2(n13732), .B1(n10879), .B2(n13176), .ZN(
        n2427) );
  OAI22_X2 U2698 ( .A1(n10305), .A2(n13739), .B1(n10878), .B2(n13740), .ZN(
        n2432) );
  OAI22_X2 U2700 ( .A1(n11407), .A2(n13743), .B1(n10389), .B2(n13745), .ZN(
        n2433) );
  OAI221_X2 U2711 ( .B1(n11360), .B2(n13735), .C1(n10676), .C2(n13182), .A(
        n2442), .ZN(n2441) );
  OAI221_X2 U2714 ( .B1(n10248), .B2(n13730), .C1(n10383), .C2(n13727), .A(
        n2443), .ZN(n2440) );
  NAND2_X2 U2716 ( .A1(n2444), .A2(n2445), .ZN(n2439) );
  AOI221_X2 U2717 ( .B1(n19157), .B2(REG_FILE_reg_out_19__3_), .C1(n13495), 
        .C2(REG_FILE_reg_out_13__3_), .A(n2446), .ZN(n2445) );
  AOI221_X2 U2721 ( .B1(n19159), .B2(REG_FILE_reg_out_3__3_), .C1(n13498), 
        .C2(REG_FILE_reg_out_4__3_), .A(n2447), .ZN(n2444) );
  OAI22_X2 U2722 ( .A1(n10508), .A2(n13733), .B1(n10877), .B2(n13176), .ZN(
        n2447) );
  OAI22_X2 U2725 ( .A1(n10304), .A2(n13739), .B1(n10876), .B2(n13741), .ZN(
        n2452) );
  OAI22_X2 U2727 ( .A1(n11406), .A2(n13743), .B1(n10388), .B2(n13745), .ZN(
        n2453) );
  OAI22_X2 U2736 ( .A1(net231243), .A2(n12541), .B1(net231311), .B2(n2457), 
        .ZN(n7484) );
  NOR4_X2 U2737 ( .A1(n2458), .A2(n2459), .A3(n2460), .A4(n2461), .ZN(n2457)
         );
  OAI221_X2 U2738 ( .B1(n11359), .B2(n13735), .C1(n10675), .C2(n13182), .A(
        n2462), .ZN(n2461) );
  OAI221_X2 U2741 ( .B1(n10247), .B2(n13730), .C1(n10382), .C2(n13727), .A(
        n2463), .ZN(n2460) );
  NAND2_X2 U2743 ( .A1(n2464), .A2(n2465), .ZN(n2459) );
  AOI221_X2 U2744 ( .B1(n19157), .B2(REG_FILE_reg_out_19__2_), .C1(n13495), 
        .C2(REG_FILE_reg_out_13__2_), .A(n2466), .ZN(n2465) );
  AOI221_X2 U2748 ( .B1(n19159), .B2(REG_FILE_reg_out_3__2_), .C1(n13498), 
        .C2(REG_FILE_reg_out_4__2_), .A(n2467), .ZN(n2464) );
  OAI22_X2 U2749 ( .A1(n10507), .A2(n13733), .B1(n10875), .B2(n13176), .ZN(
        n2467) );
  OAI22_X2 U2752 ( .A1(n10303), .A2(n13739), .B1(n10874), .B2(n13741), .ZN(
        n2472) );
  OAI22_X2 U2754 ( .A1(n11405), .A2(n13743), .B1(n10387), .B2(n13745), .ZN(
        n2473) );
  OAI22_X2 U2763 ( .A1(net231243), .A2(n12206), .B1(net231311), .B2(n2477), 
        .ZN(n7537) );
  NOR4_X2 U2764 ( .A1(n2478), .A2(n2479), .A3(n2480), .A4(n2481), .ZN(n2477)
         );
  OAI221_X2 U2765 ( .B1(n11358), .B2(n13735), .C1(n10674), .C2(n13182), .A(
        n2482), .ZN(n2481) );
  OAI221_X2 U2768 ( .B1(n10246), .B2(n13730), .C1(n10381), .C2(n13727), .A(
        n2483), .ZN(n2480) );
  NAND2_X2 U2770 ( .A1(n2484), .A2(n2485), .ZN(n2479) );
  AOI221_X2 U2771 ( .B1(n19157), .B2(REG_FILE_reg_out_19__1_), .C1(n13496), 
        .C2(REG_FILE_reg_out_13__1_), .A(n2486), .ZN(n2485) );
  AOI221_X2 U2775 ( .B1(n19159), .B2(REG_FILE_reg_out_3__1_), .C1(n13498), 
        .C2(REG_FILE_reg_out_4__1_), .A(n2487), .ZN(n2484) );
  OAI22_X2 U2776 ( .A1(n10506), .A2(n13732), .B1(n10873), .B2(n13176), .ZN(
        n2487) );
  OAI22_X2 U2779 ( .A1(n10302), .A2(n13739), .B1(n10872), .B2(n13740), .ZN(
        n2492) );
  OAI22_X2 U2781 ( .A1(n11404), .A2(n13743), .B1(n10386), .B2(n13745), .ZN(
        n2493) );
  OAI22_X2 U2791 ( .A1(net231243), .A2(n12229), .B1(net231311), .B2(n2497), 
        .ZN(n7328) );
  NOR4_X2 U2792 ( .A1(n2498), .A2(n2499), .A3(n2500), .A4(n2501), .ZN(n2497)
         );
  OAI221_X2 U2793 ( .B1(n11338), .B2(n13735), .C1(n10673), .C2(n13182), .A(
        n2502), .ZN(n2501) );
  OAI221_X2 U2801 ( .B1(n10245), .B2(n13730), .C1(n10371), .C2(n13727), .A(
        n2509), .ZN(n2500) );
  NAND2_X2 U2810 ( .A1(n2513), .A2(n2514), .ZN(n2499) );
  AOI221_X2 U2811 ( .B1(n19157), .B2(REG_FILE_reg_out_19__0_), .C1(n13495), 
        .C2(REG_FILE_reg_out_13__0_), .A(n2515), .ZN(n2514) );
  AOI221_X2 U2820 ( .B1(n19159), .B2(REG_FILE_reg_out_3__0_), .C1(n13498), 
        .C2(REG_FILE_reg_out_4__0_), .A(n2517), .ZN(n2513) );
  OAI22_X2 U2821 ( .A1(n10505), .A2(n13733), .B1(n10871), .B2(n13176), .ZN(
        n2517) );
  OAI22_X2 U2829 ( .A1(n10301), .A2(n13739), .B1(n10870), .B2(n13740), .ZN(
        n2522) );
  OAI22_X2 U2835 ( .A1(n12285), .A2(n13743), .B1(n10869), .B2(n13745), .ZN(
        n2524) );
  AND2_X2 U2855 ( .A1(n2531), .A2(n2528), .ZN(n2508) );
  OAI22_X2 U2872 ( .A1(net231243), .A2(n10358), .B1(n12304), .B2(net230373), 
        .ZN(n7545) );
  OAI22_X2 U2874 ( .A1(net231243), .A2(net137343), .B1(n12310), .B2(net230373), 
        .ZN(n7727) );
  OAI22_X2 U2876 ( .A1(net231243), .A2(net137317), .B1(n12192), .B2(net230373), 
        .ZN(n7692) );
  OAI22_X2 U2888 ( .A1(net231243), .A2(net137303), .B1(n12191), .B2(net230373), 
        .ZN(n7675) );
  NAND4_X2 U2892 ( .A1(n2565), .A2(n2566), .A3(n2567), .A4(n2568), .ZN(n7292)
         );
  NOR4_X2 U2893 ( .A1(n2569), .A2(n2570), .A3(n2571), .A4(n2572), .ZN(n2568)
         );
  OAI221_X2 U2894 ( .B1(n13725), .B2(n11172), .C1(n13722), .C2(n10589), .A(
        n2577), .ZN(n2572) );
  AOI22_X2 U2895 ( .A1(FP_REG_FILE_reg_out_27__31_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__31_), .B2(n13503), .ZN(n2577) );
  OAI221_X2 U2896 ( .B1(n13721), .B2(n10229), .C1(n13718), .C2(n11135), .A(
        n2584), .ZN(n2571) );
  AOI22_X2 U2897 ( .A1(FP_REG_FILE_reg_out_2__31_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__31_), .B2(n13508), .ZN(n2584) );
  OAI221_X2 U2900 ( .B1(n13716), .B2(n11213), .C1(n13714), .C2(n10608), .A(
        n2598), .ZN(n2569) );
  OAI221_X2 U2903 ( .B1(n13713), .B2(n10291), .C1(n13710), .C2(n10430), .A(
        n2608), .ZN(n2603) );
  AOI22_X2 U2904 ( .A1(FP_REG_FILE_reg_out_9__31_), .A2(n13511), .B1(
        ID_EXEC_OUT[267]), .B2(net231307), .ZN(n2608) );
  AOI221_X2 U2907 ( .B1(FP_REG_FILE_reg_out_28__31_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__31_), .C2(n13514), .A(n2619), .ZN(n2566) );
  OAI22_X2 U2908 ( .A1(n13707), .A2(n10491), .B1(n13704), .B2(n11337), .ZN(
        n2619) );
  AOI221_X2 U2909 ( .B1(FP_REG_FILE_reg_out_29__31_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__31_), .C2(n13518), .A(n2626), .ZN(n2565) );
  OAI22_X2 U2910 ( .A1(n13703), .A2(n10460), .B1(n13700), .B2(n11460), .ZN(
        n2626) );
  NAND4_X2 U2911 ( .A1(n2631), .A2(n2632), .A3(n2633), .A4(n2634), .ZN(n7732)
         );
  NOR4_X2 U2912 ( .A1(n2635), .A2(n2636), .A3(n2637), .A4(n2638), .ZN(n2634)
         );
  OAI221_X2 U2913 ( .B1(n13724), .B2(n11171), .C1(n13722), .C2(n10588), .A(
        n2641), .ZN(n2638) );
  AOI22_X2 U2914 ( .A1(FP_REG_FILE_reg_out_27__30_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__30_), .B2(n13503), .ZN(n2641) );
  OAI221_X2 U2915 ( .B1(n13720), .B2(n10228), .C1(n13718), .C2(n11134), .A(
        n2644), .ZN(n2637) );
  AOI22_X2 U2916 ( .A1(FP_REG_FILE_reg_out_2__30_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__30_), .B2(n13508), .ZN(n2644) );
  OAI221_X2 U2919 ( .B1(n13717), .B2(n11212), .C1(n13714), .C2(n10607), .A(
        n2650), .ZN(n2635) );
  OAI221_X2 U2922 ( .B1(n13712), .B2(n10290), .C1(n13710), .C2(n10429), .A(
        n2655), .ZN(n2652) );
  AOI22_X2 U2923 ( .A1(FP_REG_FILE_reg_out_9__30_), .A2(n13512), .B1(
        ID_EXEC_OUT[266]), .B2(net231305), .ZN(n2655) );
  AOI221_X2 U2926 ( .B1(FP_REG_FILE_reg_out_28__30_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__30_), .C2(n13514), .A(n2659), .ZN(n2632) );
  OAI22_X2 U2927 ( .A1(n13706), .A2(n10490), .B1(n13704), .B2(n11336), .ZN(
        n2659) );
  AOI221_X2 U2928 ( .B1(FP_REG_FILE_reg_out_29__30_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__30_), .C2(n13518), .A(n2662), .ZN(n2631) );
  OAI22_X2 U2929 ( .A1(n13702), .A2(n10459), .B1(n13700), .B2(n11459), .ZN(
        n2662) );
  NAND4_X2 U2930 ( .A1(n2665), .A2(n2666), .A3(n2667), .A4(n2668), .ZN(n7717)
         );
  NOR4_X2 U2931 ( .A1(n2669), .A2(n2670), .A3(n2671), .A4(n2672), .ZN(n2668)
         );
  OAI221_X2 U2932 ( .B1(n13725), .B2(n11170), .C1(n13722), .C2(n10587), .A(
        n2675), .ZN(n2672) );
  AOI22_X2 U2933 ( .A1(FP_REG_FILE_reg_out_27__29_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__29_), .B2(n13503), .ZN(n2675) );
  OAI221_X2 U2934 ( .B1(n13721), .B2(n10227), .C1(n13718), .C2(n11133), .A(
        n2678), .ZN(n2671) );
  AOI22_X2 U2935 ( .A1(FP_REG_FILE_reg_out_2__29_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__29_), .B2(n13508), .ZN(n2678) );
  OAI221_X2 U2938 ( .B1(n13716), .B2(n11211), .C1(n13714), .C2(n10606), .A(
        n2684), .ZN(n2669) );
  OAI221_X2 U2941 ( .B1(n13713), .B2(n10289), .C1(n13710), .C2(n10428), .A(
        n2689), .ZN(n2686) );
  AOI22_X2 U2942 ( .A1(FP_REG_FILE_reg_out_9__29_), .A2(n13511), .B1(
        ID_EXEC_OUT[265]), .B2(net231307), .ZN(n2689) );
  AOI221_X2 U2945 ( .B1(FP_REG_FILE_reg_out_28__29_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__29_), .C2(n13514), .A(n2693), .ZN(n2666) );
  OAI22_X2 U2946 ( .A1(n13707), .A2(n10489), .B1(n13704), .B2(n11335), .ZN(
        n2693) );
  AOI221_X2 U2947 ( .B1(FP_REG_FILE_reg_out_29__29_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__29_), .C2(n13518), .A(n2696), .ZN(n2665) );
  OAI22_X2 U2948 ( .A1(n13703), .A2(n10458), .B1(n13700), .B2(n11458), .ZN(
        n2696) );
  NAND4_X2 U2949 ( .A1(n2699), .A2(n2700), .A3(n2701), .A4(n2702), .ZN(n7646)
         );
  NOR4_X2 U2950 ( .A1(n2703), .A2(n2704), .A3(n2705), .A4(n2706), .ZN(n2702)
         );
  OAI221_X2 U2951 ( .B1(n13724), .B2(n11169), .C1(n13722), .C2(n10586), .A(
        n2709), .ZN(n2706) );
  AOI22_X2 U2952 ( .A1(FP_REG_FILE_reg_out_27__28_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__28_), .B2(n13503), .ZN(n2709) );
  OAI221_X2 U2953 ( .B1(n13720), .B2(n10226), .C1(n13718), .C2(n11132), .A(
        n2712), .ZN(n2705) );
  AOI22_X2 U2954 ( .A1(FP_REG_FILE_reg_out_2__28_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__28_), .B2(n13508), .ZN(n2712) );
  OAI221_X2 U2957 ( .B1(n13717), .B2(n11210), .C1(n13714), .C2(n10605), .A(
        n2718), .ZN(n2703) );
  OAI221_X2 U2960 ( .B1(n13712), .B2(n10288), .C1(n13710), .C2(n10427), .A(
        n2723), .ZN(n2720) );
  AOI22_X2 U2961 ( .A1(FP_REG_FILE_reg_out_9__28_), .A2(n13512), .B1(
        ID_EXEC_OUT[264]), .B2(net231305), .ZN(n2723) );
  AOI221_X2 U2964 ( .B1(FP_REG_FILE_reg_out_28__28_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__28_), .C2(n13514), .A(n2727), .ZN(n2700) );
  OAI22_X2 U2965 ( .A1(n13706), .A2(n10488), .B1(n13704), .B2(n11334), .ZN(
        n2727) );
  AOI221_X2 U2966 ( .B1(FP_REG_FILE_reg_out_29__28_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__28_), .C2(n13518), .A(n2730), .ZN(n2699) );
  OAI22_X2 U2967 ( .A1(n13702), .A2(n10457), .B1(n13700), .B2(n11457), .ZN(
        n2730) );
  NAND4_X2 U2968 ( .A1(n2733), .A2(n2734), .A3(n2735), .A4(n2736), .ZN(n7705)
         );
  NOR4_X2 U2969 ( .A1(n2737), .A2(n2738), .A3(n2739), .A4(n2740), .ZN(n2736)
         );
  OAI221_X2 U2970 ( .B1(n13725), .B2(n11168), .C1(n13722), .C2(n10585), .A(
        n2743), .ZN(n2740) );
  AOI22_X2 U2971 ( .A1(FP_REG_FILE_reg_out_27__27_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__27_), .B2(n13503), .ZN(n2743) );
  OAI221_X2 U2972 ( .B1(n13721), .B2(n10225), .C1(n13718), .C2(n11131), .A(
        n2746), .ZN(n2739) );
  AOI22_X2 U2973 ( .A1(FP_REG_FILE_reg_out_2__27_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__27_), .B2(n13508), .ZN(n2746) );
  OAI221_X2 U2976 ( .B1(n13716), .B2(n11209), .C1(n13714), .C2(n10604), .A(
        n2752), .ZN(n2737) );
  OAI221_X2 U2979 ( .B1(n13713), .B2(n10287), .C1(n13710), .C2(n10426), .A(
        n2757), .ZN(n2754) );
  AOI22_X2 U2980 ( .A1(FP_REG_FILE_reg_out_9__27_), .A2(n13511), .B1(
        ID_EXEC_OUT[263]), .B2(net231307), .ZN(n2757) );
  AOI221_X2 U2983 ( .B1(FP_REG_FILE_reg_out_28__27_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__27_), .C2(n13514), .A(n2761), .ZN(n2734) );
  OAI22_X2 U2984 ( .A1(n13707), .A2(n10487), .B1(n13704), .B2(n11333), .ZN(
        n2761) );
  AOI221_X2 U2985 ( .B1(FP_REG_FILE_reg_out_29__27_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__27_), .C2(n13518), .A(n2764), .ZN(n2733) );
  OAI22_X2 U2986 ( .A1(n13703), .A2(n10456), .B1(n13700), .B2(n11456), .ZN(
        n2764) );
  NAND4_X2 U2987 ( .A1(n2767), .A2(n2768), .A3(n2769), .A4(n2770), .ZN(n7699)
         );
  NOR4_X2 U2988 ( .A1(n2771), .A2(n2772), .A3(n2773), .A4(n2774), .ZN(n2770)
         );
  OAI221_X2 U2989 ( .B1(n13724), .B2(n11167), .C1(n13722), .C2(n10584), .A(
        n2777), .ZN(n2774) );
  AOI22_X2 U2990 ( .A1(FP_REG_FILE_reg_out_27__26_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__26_), .B2(n13503), .ZN(n2777) );
  OAI221_X2 U2991 ( .B1(n13720), .B2(n10224), .C1(n13718), .C2(n11130), .A(
        n2780), .ZN(n2773) );
  AOI22_X2 U2992 ( .A1(FP_REG_FILE_reg_out_2__26_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__26_), .B2(n13508), .ZN(n2780) );
  OAI221_X2 U2995 ( .B1(n13717), .B2(n11208), .C1(n13714), .C2(n10603), .A(
        n2786), .ZN(n2771) );
  OAI221_X2 U2998 ( .B1(n13712), .B2(n10286), .C1(n13710), .C2(n10425), .A(
        n2791), .ZN(n2788) );
  AOI22_X2 U2999 ( .A1(FP_REG_FILE_reg_out_9__26_), .A2(n13512), .B1(
        ID_EXEC_OUT[262]), .B2(net231305), .ZN(n2791) );
  AOI221_X2 U3002 ( .B1(FP_REG_FILE_reg_out_28__26_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__26_), .C2(n13514), .A(n2795), .ZN(n2768) );
  OAI22_X2 U3003 ( .A1(n13706), .A2(n10486), .B1(n13704), .B2(n11332), .ZN(
        n2795) );
  AOI221_X2 U3004 ( .B1(FP_REG_FILE_reg_out_29__26_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__26_), .C2(n13518), .A(n2798), .ZN(n2767) );
  OAI22_X2 U3005 ( .A1(n13702), .A2(n10455), .B1(n13700), .B2(n11455), .ZN(
        n2798) );
  NAND4_X2 U3006 ( .A1(n2801), .A2(n2802), .A3(n2803), .A4(n2804), .ZN(n7711)
         );
  NOR4_X2 U3007 ( .A1(n2805), .A2(n2806), .A3(n2807), .A4(n2808), .ZN(n2804)
         );
  OAI221_X2 U3008 ( .B1(n13725), .B2(n11166), .C1(n13722), .C2(n10583), .A(
        n2811), .ZN(n2808) );
  AOI22_X2 U3009 ( .A1(FP_REG_FILE_reg_out_27__25_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__25_), .B2(n13503), .ZN(n2811) );
  OAI221_X2 U3010 ( .B1(n13721), .B2(n10223), .C1(n13718), .C2(n11129), .A(
        n2814), .ZN(n2807) );
  AOI22_X2 U3011 ( .A1(FP_REG_FILE_reg_out_2__25_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__25_), .B2(n13508), .ZN(n2814) );
  OAI221_X2 U3014 ( .B1(n13716), .B2(n11207), .C1(n13714), .C2(n10602), .A(
        n2820), .ZN(n2805) );
  OAI221_X2 U3017 ( .B1(n13713), .B2(n10285), .C1(n13710), .C2(n10424), .A(
        n2825), .ZN(n2822) );
  AOI22_X2 U3018 ( .A1(FP_REG_FILE_reg_out_9__25_), .A2(n13511), .B1(
        ID_EXEC_OUT[261]), .B2(net231307), .ZN(n2825) );
  AOI221_X2 U3021 ( .B1(FP_REG_FILE_reg_out_28__25_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__25_), .C2(n13514), .A(n2829), .ZN(n2802) );
  OAI22_X2 U3022 ( .A1(n13707), .A2(n10485), .B1(n13704), .B2(n11331), .ZN(
        n2829) );
  AOI221_X2 U3023 ( .B1(FP_REG_FILE_reg_out_29__25_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__25_), .C2(n13518), .A(n2832), .ZN(n2801) );
  OAI22_X2 U3024 ( .A1(n13703), .A2(n10454), .B1(n13700), .B2(n11454), .ZN(
        n2832) );
  NAND4_X2 U3025 ( .A1(n2835), .A2(n2836), .A3(n2837), .A4(n2838), .ZN(n7295)
         );
  NOR4_X2 U3026 ( .A1(n2839), .A2(n2840), .A3(n2841), .A4(n2842), .ZN(n2838)
         );
  OAI221_X2 U3027 ( .B1(n13724), .B2(n11165), .C1(n13722), .C2(n10582), .A(
        n2845), .ZN(n2842) );
  AOI22_X2 U3028 ( .A1(FP_REG_FILE_reg_out_27__24_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__24_), .B2(n13503), .ZN(n2845) );
  OAI221_X2 U3029 ( .B1(n13720), .B2(n10222), .C1(n13718), .C2(n11128), .A(
        n2848), .ZN(n2841) );
  AOI22_X2 U3030 ( .A1(FP_REG_FILE_reg_out_2__24_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__24_), .B2(n13508), .ZN(n2848) );
  OAI221_X2 U3033 ( .B1(n13717), .B2(n11206), .C1(n13714), .C2(n10601), .A(
        n2854), .ZN(n2839) );
  OAI221_X2 U3036 ( .B1(n13712), .B2(n10284), .C1(n13710), .C2(n10423), .A(
        n2859), .ZN(n2856) );
  AOI22_X2 U3037 ( .A1(FP_REG_FILE_reg_out_9__24_), .A2(n13512), .B1(
        ID_EXEC_OUT[260]), .B2(net231305), .ZN(n2859) );
  AOI221_X2 U3040 ( .B1(FP_REG_FILE_reg_out_28__24_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__24_), .C2(n13514), .A(n2863), .ZN(n2836) );
  OAI22_X2 U3041 ( .A1(n13706), .A2(n10484), .B1(n13704), .B2(n11330), .ZN(
        n2863) );
  AOI221_X2 U3042 ( .B1(FP_REG_FILE_reg_out_29__24_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__24_), .C2(n13518), .A(n2866), .ZN(n2835) );
  OAI22_X2 U3043 ( .A1(n13702), .A2(n10453), .B1(n13700), .B2(n11453), .ZN(
        n2866) );
  NAND4_X2 U3046 ( .A1(n2870), .A2(n2871), .A3(n2872), .A4(n2873), .ZN(n7299)
         );
  NOR4_X2 U3047 ( .A1(n2874), .A2(n2875), .A3(n2876), .A4(n2877), .ZN(n2873)
         );
  OAI221_X2 U3048 ( .B1(n13725), .B2(n11164), .C1(n13722), .C2(n10581), .A(
        n2880), .ZN(n2877) );
  AOI22_X2 U3049 ( .A1(FP_REG_FILE_reg_out_27__23_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__23_), .B2(n13503), .ZN(n2880) );
  OAI221_X2 U3050 ( .B1(n13721), .B2(n10221), .C1(n13718), .C2(n11127), .A(
        n2883), .ZN(n2876) );
  AOI22_X2 U3051 ( .A1(FP_REG_FILE_reg_out_2__23_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__23_), .B2(n13508), .ZN(n2883) );
  OAI221_X2 U3054 ( .B1(n13716), .B2(n11205), .C1(n13714), .C2(n10600), .A(
        n2889), .ZN(n2874) );
  OAI221_X2 U3057 ( .B1(n13713), .B2(n10283), .C1(n13710), .C2(n10422), .A(
        n2894), .ZN(n2891) );
  AOI22_X2 U3058 ( .A1(FP_REG_FILE_reg_out_9__23_), .A2(n13511), .B1(
        ID_EXEC_OUT[259]), .B2(net231307), .ZN(n2894) );
  AOI221_X2 U3061 ( .B1(FP_REG_FILE_reg_out_28__23_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__23_), .C2(n13514), .A(n2898), .ZN(n2871) );
  OAI22_X2 U3062 ( .A1(n13707), .A2(n10483), .B1(n13704), .B2(n11329), .ZN(
        n2898) );
  AOI221_X2 U3063 ( .B1(FP_REG_FILE_reg_out_29__23_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__23_), .C2(n13518), .A(n2901), .ZN(n2870) );
  OAI22_X2 U3064 ( .A1(n13703), .A2(n10452), .B1(n13700), .B2(n11452), .ZN(
        n2901) );
  NAND4_X2 U3065 ( .A1(n2904), .A2(n2905), .A3(n2906), .A4(n2907), .ZN(n7307)
         );
  NOR4_X2 U3066 ( .A1(n2908), .A2(n2909), .A3(n2910), .A4(n2911), .ZN(n2907)
         );
  OAI221_X2 U3067 ( .B1(n13724), .B2(n11163), .C1(n13722), .C2(n10580), .A(
        n2914), .ZN(n2911) );
  AOI22_X2 U3068 ( .A1(FP_REG_FILE_reg_out_27__22_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__22_), .B2(n13503), .ZN(n2914) );
  OAI221_X2 U3069 ( .B1(n13720), .B2(n10220), .C1(n13718), .C2(n11126), .A(
        n2917), .ZN(n2910) );
  AOI22_X2 U3070 ( .A1(FP_REG_FILE_reg_out_2__22_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__22_), .B2(n13508), .ZN(n2917) );
  OAI221_X2 U3073 ( .B1(n13717), .B2(n11204), .C1(n13714), .C2(n10599), .A(
        n2923), .ZN(n2908) );
  OAI221_X2 U3076 ( .B1(n13712), .B2(n10282), .C1(n13710), .C2(n10421), .A(
        n2928), .ZN(n2925) );
  AOI22_X2 U3077 ( .A1(FP_REG_FILE_reg_out_9__22_), .A2(n13512), .B1(
        ID_EXEC_OUT[258]), .B2(net231305), .ZN(n2928) );
  AOI221_X2 U3080 ( .B1(FP_REG_FILE_reg_out_28__22_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__22_), .C2(n13514), .A(n2932), .ZN(n2905) );
  OAI22_X2 U3081 ( .A1(n13706), .A2(n10482), .B1(n13704), .B2(n11328), .ZN(
        n2932) );
  AOI221_X2 U3082 ( .B1(FP_REG_FILE_reg_out_29__22_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__22_), .C2(n13518), .A(n2935), .ZN(n2904) );
  OAI22_X2 U3083 ( .A1(n13702), .A2(n10451), .B1(n13700), .B2(n11451), .ZN(
        n2935) );
  NAND4_X2 U3084 ( .A1(n2938), .A2(n2939), .A3(n2940), .A4(n2941), .ZN(n7311)
         );
  NOR4_X2 U3085 ( .A1(n2942), .A2(n2943), .A3(n2944), .A4(n2945), .ZN(n2941)
         );
  OAI221_X2 U3086 ( .B1(n13725), .B2(n11162), .C1(n13722), .C2(n10579), .A(
        n2948), .ZN(n2945) );
  AOI22_X2 U3087 ( .A1(FP_REG_FILE_reg_out_27__21_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__21_), .B2(n13502), .ZN(n2948) );
  OAI221_X2 U3088 ( .B1(n13721), .B2(n10219), .C1(n13718), .C2(n11125), .A(
        n2951), .ZN(n2944) );
  AOI22_X2 U3089 ( .A1(FP_REG_FILE_reg_out_2__21_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__21_), .B2(n13508), .ZN(n2951) );
  OAI221_X2 U3092 ( .B1(n13717), .B2(n11203), .C1(n13714), .C2(n10598), .A(
        n2957), .ZN(n2942) );
  OAI221_X2 U3095 ( .B1(n13713), .B2(n10281), .C1(n13710), .C2(n10420), .A(
        n2962), .ZN(n2959) );
  AOI22_X2 U3096 ( .A1(FP_REG_FILE_reg_out_9__21_), .A2(n13512), .B1(
        ID_EXEC_OUT[257]), .B2(net231307), .ZN(n2962) );
  AOI221_X2 U3099 ( .B1(FP_REG_FILE_reg_out_28__21_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__21_), .C2(n13514), .A(n2966), .ZN(n2939) );
  OAI22_X2 U3100 ( .A1(n13707), .A2(n10481), .B1(n13704), .B2(n11327), .ZN(
        n2966) );
  AOI221_X2 U3101 ( .B1(FP_REG_FILE_reg_out_29__21_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__21_), .C2(n13518), .A(n2969), .ZN(n2938) );
  OAI22_X2 U3102 ( .A1(n13703), .A2(n10450), .B1(n13700), .B2(n11450), .ZN(
        n2969) );
  NAND4_X2 U3103 ( .A1(n2972), .A2(n2973), .A3(n2974), .A4(n2975), .ZN(n7316)
         );
  NOR4_X2 U3104 ( .A1(n2976), .A2(n2977), .A3(n2978), .A4(n2979), .ZN(n2975)
         );
  OAI221_X2 U3105 ( .B1(n13724), .B2(n12252), .C1(n13723), .C2(n11138), .A(
        n2982), .ZN(n2979) );
  AOI22_X2 U3106 ( .A1(FP_REG_FILE_reg_out_27__20_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__20_), .B2(n13502), .ZN(n2982) );
  OAI221_X2 U3107 ( .B1(n13720), .B2(n10261), .C1(n13719), .C2(n12222), .A(
        n2985), .ZN(n2978) );
  AOI22_X2 U3108 ( .A1(FP_REG_FILE_reg_out_2__20_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__20_), .B2(n13507), .ZN(n2985) );
  OAI221_X2 U3111 ( .B1(n13716), .B2(n12255), .C1(n13715), .C2(n11140), .A(
        n2991), .ZN(n2976) );
  OAI221_X2 U3114 ( .B1(n13712), .B2(n10912), .C1(n13711), .C2(n10419), .A(
        n2996), .ZN(n2993) );
  AOI22_X2 U3115 ( .A1(FP_REG_FILE_reg_out_9__20_), .A2(n13512), .B1(
        ID_EXEC_OUT[256]), .B2(net231305), .ZN(n2996) );
  AOI221_X2 U3118 ( .B1(FP_REG_FILE_reg_out_28__20_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__20_), .C2(n13513), .A(n3000), .ZN(n2973) );
  OAI22_X2 U3119 ( .A1(n13706), .A2(n10917), .B1(n13705), .B2(n12281), .ZN(
        n3000) );
  AOI221_X2 U3120 ( .B1(FP_REG_FILE_reg_out_29__20_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__20_), .C2(n13517), .A(n3003), .ZN(n2972) );
  OAI22_X2 U3121 ( .A1(n13702), .A2(n10915), .B1(n13701), .B2(n12297), .ZN(
        n3003) );
  NAND4_X2 U3122 ( .A1(n3006), .A2(n3007), .A3(n3008), .A4(n3009), .ZN(n7303)
         );
  NOR4_X2 U3123 ( .A1(n3010), .A2(n3011), .A3(n3012), .A4(n3013), .ZN(n3009)
         );
  OAI221_X2 U3124 ( .B1(n13724), .B2(n12251), .C1(n13723), .C2(n11137), .A(
        n3016), .ZN(n3013) );
  AOI22_X2 U3125 ( .A1(FP_REG_FILE_reg_out_27__19_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__19_), .B2(n13502), .ZN(n3016) );
  OAI221_X2 U3126 ( .B1(n13720), .B2(n10260), .C1(n13719), .C2(n12221), .A(
        n3019), .ZN(n3012) );
  AOI22_X2 U3127 ( .A1(FP_REG_FILE_reg_out_2__19_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__19_), .B2(n13508), .ZN(n3019) );
  OAI221_X2 U3130 ( .B1(n13716), .B2(n12254), .C1(n13715), .C2(n11139), .A(
        n3025), .ZN(n3010) );
  OAI221_X2 U3133 ( .B1(n13712), .B2(n10911), .C1(n13711), .C2(n10418), .A(
        n3030), .ZN(n3027) );
  AOI22_X2 U3134 ( .A1(FP_REG_FILE_reg_out_9__19_), .A2(n13512), .B1(
        ID_EXEC_OUT[255]), .B2(net231307), .ZN(n3030) );
  AOI221_X2 U3137 ( .B1(FP_REG_FILE_reg_out_28__19_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__19_), .C2(n13514), .A(n3034), .ZN(n3007) );
  OAI22_X2 U3138 ( .A1(n13706), .A2(n10916), .B1(n13705), .B2(n12280), .ZN(
        n3034) );
  AOI221_X2 U3139 ( .B1(FP_REG_FILE_reg_out_29__19_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__19_), .C2(n13518), .A(n3037), .ZN(n3006) );
  OAI22_X2 U3140 ( .A1(n13702), .A2(n10914), .B1(n13701), .B2(n12296), .ZN(
        n3037) );
  NAND4_X2 U3141 ( .A1(n3040), .A2(n3041), .A3(n3042), .A4(n3043), .ZN(n7747)
         );
  NOR4_X2 U3142 ( .A1(n3044), .A2(n3045), .A3(n3046), .A4(n3047), .ZN(n3043)
         );
  OAI221_X2 U3143 ( .B1(n13724), .B2(n11161), .C1(n13723), .C2(n10578), .A(
        n3050), .ZN(n3047) );
  AOI22_X2 U3144 ( .A1(FP_REG_FILE_reg_out_27__18_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__18_), .B2(n13502), .ZN(n3050) );
  OAI221_X2 U3145 ( .B1(n13720), .B2(n10218), .C1(n13719), .C2(n11124), .A(
        n3053), .ZN(n3046) );
  AOI22_X2 U3146 ( .A1(FP_REG_FILE_reg_out_2__18_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__18_), .B2(n13507), .ZN(n3053) );
  OAI221_X2 U3149 ( .B1(n13716), .B2(n11202), .C1(n13715), .C2(n10597), .A(
        n3059), .ZN(n3044) );
  OAI221_X2 U3152 ( .B1(n13712), .B2(n10280), .C1(n13711), .C2(n10417), .A(
        n3064), .ZN(n3061) );
  AOI22_X2 U3153 ( .A1(FP_REG_FILE_reg_out_9__18_), .A2(n13512), .B1(
        ID_EXEC_OUT[254]), .B2(net231305), .ZN(n3064) );
  AOI221_X2 U3156 ( .B1(FP_REG_FILE_reg_out_28__18_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__18_), .C2(n13513), .A(n3068), .ZN(n3041) );
  OAI22_X2 U3157 ( .A1(n13706), .A2(n10480), .B1(n13705), .B2(n11326), .ZN(
        n3068) );
  AOI221_X2 U3158 ( .B1(FP_REG_FILE_reg_out_29__18_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__18_), .C2(n13517), .A(n3071), .ZN(n3040) );
  OAI22_X2 U3159 ( .A1(n13702), .A2(n10449), .B1(n13701), .B2(n11449), .ZN(
        n3071) );
  NAND4_X2 U3160 ( .A1(n3074), .A2(n3075), .A3(n3076), .A4(n3077), .ZN(n7337)
         );
  NOR4_X2 U3161 ( .A1(n3078), .A2(n3079), .A3(n3080), .A4(n3081), .ZN(n3077)
         );
  OAI221_X2 U3162 ( .B1(n13724), .B2(n11160), .C1(n13723), .C2(n10577), .A(
        n3084), .ZN(n3081) );
  AOI22_X2 U3163 ( .A1(FP_REG_FILE_reg_out_27__17_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__17_), .B2(n13502), .ZN(n3084) );
  OAI221_X2 U3164 ( .B1(n13720), .B2(n10217), .C1(n13719), .C2(n11123), .A(
        n3087), .ZN(n3080) );
  AOI22_X2 U3165 ( .A1(FP_REG_FILE_reg_out_2__17_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__17_), .B2(n13508), .ZN(n3087) );
  OAI221_X2 U3168 ( .B1(n13716), .B2(n11201), .C1(n13715), .C2(n10596), .A(
        n3093), .ZN(n3078) );
  OAI221_X2 U3171 ( .B1(n13712), .B2(n10279), .C1(n13711), .C2(n10416), .A(
        n3098), .ZN(n3095) );
  AOI22_X2 U3172 ( .A1(FP_REG_FILE_reg_out_9__17_), .A2(n13512), .B1(
        ID_EXEC_OUT[253]), .B2(net231305), .ZN(n3098) );
  AOI221_X2 U3175 ( .B1(FP_REG_FILE_reg_out_28__17_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__17_), .C2(n13514), .A(n3102), .ZN(n3075) );
  OAI22_X2 U3176 ( .A1(n13706), .A2(n10479), .B1(n13705), .B2(n11325), .ZN(
        n3102) );
  AOI221_X2 U3177 ( .B1(FP_REG_FILE_reg_out_29__17_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__17_), .C2(n13518), .A(n3105), .ZN(n3074) );
  OAI22_X2 U3178 ( .A1(n13702), .A2(n10448), .B1(n13701), .B2(n11448), .ZN(
        n3105) );
  NAND4_X2 U3179 ( .A1(n3108), .A2(n3109), .A3(n3110), .A4(n3111), .ZN(n7436)
         );
  NOR4_X2 U3180 ( .A1(n3112), .A2(n3113), .A3(n3114), .A4(n3115), .ZN(n3111)
         );
  OAI221_X2 U3181 ( .B1(n13724), .B2(n11159), .C1(n13723), .C2(n10576), .A(
        n3118), .ZN(n3115) );
  AOI22_X2 U3182 ( .A1(FP_REG_FILE_reg_out_27__16_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__16_), .B2(n13502), .ZN(n3118) );
  OAI221_X2 U3183 ( .B1(n13720), .B2(n10216), .C1(n13719), .C2(n11122), .A(
        n3121), .ZN(n3114) );
  AOI22_X2 U3184 ( .A1(FP_REG_FILE_reg_out_2__16_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__16_), .B2(n13507), .ZN(n3121) );
  OAI221_X2 U3187 ( .B1(n13716), .B2(n11200), .C1(n13715), .C2(n10595), .A(
        n3127), .ZN(n3112) );
  OAI221_X2 U3190 ( .B1(n13712), .B2(n10278), .C1(n13711), .C2(n10415), .A(
        n3132), .ZN(n3129) );
  AOI22_X2 U3191 ( .A1(FP_REG_FILE_reg_out_9__16_), .A2(n13512), .B1(
        ID_EXEC_OUT[252]), .B2(net231307), .ZN(n3132) );
  AOI221_X2 U3194 ( .B1(FP_REG_FILE_reg_out_28__16_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__16_), .C2(n13513), .A(n3136), .ZN(n3109) );
  OAI22_X2 U3195 ( .A1(n13706), .A2(n10478), .B1(n13705), .B2(n11324), .ZN(
        n3136) );
  AOI221_X2 U3196 ( .B1(FP_REG_FILE_reg_out_29__16_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__16_), .C2(n13517), .A(n3139), .ZN(n3108) );
  OAI22_X2 U3197 ( .A1(n13702), .A2(n10447), .B1(n13701), .B2(n11447), .ZN(
        n3139) );
  NAND4_X2 U3198 ( .A1(n3142), .A2(n3143), .A3(n3144), .A4(n3145), .ZN(n7627)
         );
  NOR4_X2 U3199 ( .A1(n3146), .A2(n3147), .A3(n3148), .A4(n3149), .ZN(n3145)
         );
  OAI221_X2 U3200 ( .B1(n13724), .B2(n11158), .C1(n13723), .C2(n10575), .A(
        n3152), .ZN(n3149) );
  AOI22_X2 U3201 ( .A1(FP_REG_FILE_reg_out_27__15_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__15_), .B2(n13502), .ZN(n3152) );
  OAI221_X2 U3202 ( .B1(n13720), .B2(n10215), .C1(n13719), .C2(n11121), .A(
        n3155), .ZN(n3148) );
  AOI22_X2 U3203 ( .A1(FP_REG_FILE_reg_out_2__15_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__15_), .B2(n13508), .ZN(n3155) );
  OAI221_X2 U3206 ( .B1(n13716), .B2(n11199), .C1(n13715), .C2(n10594), .A(
        n3161), .ZN(n3146) );
  OAI221_X2 U3209 ( .B1(n13712), .B2(n10277), .C1(n13711), .C2(n10414), .A(
        n3166), .ZN(n3163) );
  AOI22_X2 U3210 ( .A1(FP_REG_FILE_reg_out_9__15_), .A2(n13512), .B1(
        ID_EXEC_OUT[251]), .B2(net231307), .ZN(n3166) );
  AOI221_X2 U3213 ( .B1(FP_REG_FILE_reg_out_28__15_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__15_), .C2(n13514), .A(n3170), .ZN(n3143) );
  OAI22_X2 U3214 ( .A1(n13706), .A2(n10477), .B1(n13705), .B2(n11323), .ZN(
        n3170) );
  AOI221_X2 U3215 ( .B1(FP_REG_FILE_reg_out_29__15_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__15_), .C2(n13518), .A(n3173), .ZN(n3142) );
  OAI22_X2 U3216 ( .A1(n13702), .A2(n10446), .B1(n13701), .B2(n11446), .ZN(
        n3173) );
  NAND4_X2 U3217 ( .A1(n3176), .A2(n3177), .A3(n3178), .A4(n3179), .ZN(n7610)
         );
  NOR4_X2 U3218 ( .A1(n3180), .A2(n3181), .A3(n3182), .A4(n3183), .ZN(n3179)
         );
  OAI221_X2 U3219 ( .B1(n13724), .B2(n11157), .C1(n13723), .C2(n10574), .A(
        n3186), .ZN(n3183) );
  AOI22_X2 U3220 ( .A1(FP_REG_FILE_reg_out_27__14_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__14_), .B2(n13502), .ZN(n3186) );
  OAI221_X2 U3221 ( .B1(n13720), .B2(n10214), .C1(n13719), .C2(n11120), .A(
        n3189), .ZN(n3182) );
  AOI22_X2 U3222 ( .A1(FP_REG_FILE_reg_out_2__14_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__14_), .B2(n13507), .ZN(n3189) );
  OAI221_X2 U3225 ( .B1(n13716), .B2(n11198), .C1(n13715), .C2(n10593), .A(
        n3195), .ZN(n3180) );
  OAI221_X2 U3228 ( .B1(n13712), .B2(n10276), .C1(n13711), .C2(n10413), .A(
        n3200), .ZN(n3197) );
  AOI22_X2 U3229 ( .A1(FP_REG_FILE_reg_out_9__14_), .A2(n13512), .B1(
        ID_EXEC_OUT[250]), .B2(net231305), .ZN(n3200) );
  AOI221_X2 U3232 ( .B1(FP_REG_FILE_reg_out_28__14_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__14_), .C2(n13513), .A(n3204), .ZN(n3177) );
  OAI22_X2 U3233 ( .A1(n13706), .A2(n10476), .B1(n13705), .B2(n11322), .ZN(
        n3204) );
  AOI221_X2 U3234 ( .B1(FP_REG_FILE_reg_out_29__14_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__14_), .C2(n13517), .A(n3207), .ZN(n3176) );
  OAI22_X2 U3235 ( .A1(n13702), .A2(n10445), .B1(n13701), .B2(n11445), .ZN(
        n3207) );
  AOI22_X2 U3237 ( .A1(net231315), .A2(nextPC_ex_out[24]), .B1(IF_ID_OUT[24]), 
        .B2(net230393), .ZN(n3210) );
  NAND4_X2 U3238 ( .A1(n3211), .A2(n3212), .A3(n3213), .A4(n3214), .ZN(n7593)
         );
  NOR4_X2 U3239 ( .A1(n3215), .A2(n3216), .A3(n3217), .A4(n3218), .ZN(n3214)
         );
  OAI221_X2 U3240 ( .B1(n13724), .B2(n11156), .C1(n13723), .C2(n10573), .A(
        n3221), .ZN(n3218) );
  AOI22_X2 U3241 ( .A1(FP_REG_FILE_reg_out_27__13_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__13_), .B2(n13502), .ZN(n3221) );
  OAI221_X2 U3242 ( .B1(n13720), .B2(n10213), .C1(n13719), .C2(n11119), .A(
        n3224), .ZN(n3217) );
  AOI22_X2 U3243 ( .A1(FP_REG_FILE_reg_out_2__13_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__13_), .B2(n13508), .ZN(n3224) );
  OAI221_X2 U3246 ( .B1(n13716), .B2(n11197), .C1(n13715), .C2(n10592), .A(
        n3230), .ZN(n3215) );
  OAI221_X2 U3249 ( .B1(n13712), .B2(n10275), .C1(n13711), .C2(n10412), .A(
        n3235), .ZN(n3232) );
  AOI22_X2 U3250 ( .A1(FP_REG_FILE_reg_out_9__13_), .A2(n13512), .B1(
        ID_EXEC_OUT[249]), .B2(net231305), .ZN(n3235) );
  AOI221_X2 U3253 ( .B1(FP_REG_FILE_reg_out_28__13_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__13_), .C2(n13514), .A(n3239), .ZN(n3212) );
  OAI22_X2 U3254 ( .A1(n13706), .A2(n10475), .B1(n13705), .B2(n11321), .ZN(
        n3239) );
  AOI221_X2 U3255 ( .B1(FP_REG_FILE_reg_out_29__13_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__13_), .C2(n13518), .A(n3242), .ZN(n3211) );
  OAI22_X2 U3256 ( .A1(n13702), .A2(n10444), .B1(n13701), .B2(n11444), .ZN(
        n3242) );
  NAND4_X2 U3257 ( .A1(n3245), .A2(n3246), .A3(n3247), .A4(n3248), .ZN(n7347)
         );
  NOR4_X2 U3258 ( .A1(n3249), .A2(n3250), .A3(n3251), .A4(n3252), .ZN(n3248)
         );
  OAI221_X2 U3259 ( .B1(n13724), .B2(n11155), .C1(n13723), .C2(n10572), .A(
        n3255), .ZN(n3252) );
  AOI22_X2 U3260 ( .A1(FP_REG_FILE_reg_out_27__12_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__12_), .B2(n13502), .ZN(n3255) );
  OAI221_X2 U3261 ( .B1(n13720), .B2(n10212), .C1(n13719), .C2(n11118), .A(
        n3258), .ZN(n3251) );
  AOI22_X2 U3262 ( .A1(FP_REG_FILE_reg_out_2__12_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__12_), .B2(n13507), .ZN(n3258) );
  OAI221_X2 U3265 ( .B1(n13716), .B2(n11196), .C1(n13715), .C2(n10591), .A(
        n3264), .ZN(n3249) );
  OAI221_X2 U3268 ( .B1(n13712), .B2(n10274), .C1(n13711), .C2(n10411), .A(
        n3269), .ZN(n3266) );
  AOI22_X2 U3269 ( .A1(FP_REG_FILE_reg_out_9__12_), .A2(n13512), .B1(
        ID_EXEC_OUT[248]), .B2(net231307), .ZN(n3269) );
  AOI221_X2 U3272 ( .B1(FP_REG_FILE_reg_out_28__12_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__12_), .C2(n13513), .A(n3273), .ZN(n3246) );
  OAI22_X2 U3273 ( .A1(n13706), .A2(n10474), .B1(n13705), .B2(n11320), .ZN(
        n3273) );
  AOI221_X2 U3274 ( .B1(FP_REG_FILE_reg_out_29__12_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__12_), .C2(n13517), .A(n3276), .ZN(n3245) );
  OAI22_X2 U3275 ( .A1(n13702), .A2(n10443), .B1(n13701), .B2(n11443), .ZN(
        n3276) );
  NAND4_X2 U3276 ( .A1(n3279), .A2(n3280), .A3(n3281), .A4(n3282), .ZN(n7394)
         );
  NOR4_X2 U3277 ( .A1(n3283), .A2(n3284), .A3(n3285), .A4(n3286), .ZN(n3282)
         );
  OAI221_X2 U3278 ( .B1(n13724), .B2(n11154), .C1(n13723), .C2(n10571), .A(
        n3289), .ZN(n3286) );
  AOI22_X2 U3279 ( .A1(FP_REG_FILE_reg_out_27__11_), .A2(n13506), .B1(
        FP_REG_FILE_reg_out_3__11_), .B2(n13502), .ZN(n3289) );
  OAI221_X2 U3280 ( .B1(n13720), .B2(n10211), .C1(n13719), .C2(n11117), .A(
        n3292), .ZN(n3285) );
  AOI22_X2 U3281 ( .A1(FP_REG_FILE_reg_out_2__11_), .A2(n13510), .B1(
        FP_REG_FILE_reg_out_19__11_), .B2(n13508), .ZN(n3292) );
  OAI221_X2 U3284 ( .B1(n13716), .B2(n11195), .C1(n13715), .C2(n10590), .A(
        n3298), .ZN(n3283) );
  OAI221_X2 U3287 ( .B1(n13712), .B2(n10273), .C1(n13711), .C2(n10410), .A(
        n3303), .ZN(n3300) );
  AOI22_X2 U3288 ( .A1(FP_REG_FILE_reg_out_9__11_), .A2(n13512), .B1(
        ID_EXEC_OUT[247]), .B2(net231305), .ZN(n3303) );
  AOI221_X2 U3291 ( .B1(FP_REG_FILE_reg_out_28__11_), .B2(n13516), .C1(
        FP_REG_FILE_reg_out_4__11_), .C2(n13514), .A(n3307), .ZN(n3280) );
  OAI22_X2 U3292 ( .A1(n13706), .A2(n10473), .B1(n13705), .B2(n11319), .ZN(
        n3307) );
  AOI221_X2 U3293 ( .B1(FP_REG_FILE_reg_out_29__11_), .B2(n13520), .C1(
        FP_REG_FILE_reg_out_5__11_), .C2(n13518), .A(n3310), .ZN(n3279) );
  OAI22_X2 U3294 ( .A1(n13702), .A2(n10442), .B1(n13701), .B2(n11442), .ZN(
        n3310) );
  NAND4_X2 U3295 ( .A1(n3313), .A2(n3314), .A3(n3315), .A4(n3316), .ZN(n7384)
         );
  NOR4_X2 U3296 ( .A1(n3317), .A2(n3318), .A3(n3319), .A4(n3320), .ZN(n3316)
         );
  OAI221_X2 U3297 ( .B1(n13724), .B2(n11153), .C1(n13723), .C2(n10570), .A(
        n3323), .ZN(n3320) );
  AOI22_X2 U3298 ( .A1(FP_REG_FILE_reg_out_27__10_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__10_), .B2(n13501), .ZN(n3323) );
  OAI221_X2 U3299 ( .B1(n13720), .B2(n10210), .C1(n13719), .C2(n11183), .A(
        n3326), .ZN(n3319) );
  AOI22_X2 U3300 ( .A1(FP_REG_FILE_reg_out_2__10_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__10_), .B2(n13507), .ZN(n3326) );
  OAI221_X2 U3303 ( .B1(n13716), .B2(n11194), .C1(n13715), .C2(n10649), .A(
        n3332), .ZN(n3317) );
  OAI221_X2 U3306 ( .B1(n13712), .B2(n10272), .C1(n13711), .C2(n10409), .A(
        n3337), .ZN(n3334) );
  AOI22_X2 U3307 ( .A1(FP_REG_FILE_reg_out_9__10_), .A2(n13511), .B1(
        ID_EXEC_OUT[246]), .B2(net231307), .ZN(n3337) );
  AOI221_X2 U3310 ( .B1(FP_REG_FILE_reg_out_28__10_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__10_), .C2(n13513), .A(n3341), .ZN(n3314) );
  OAI22_X2 U3311 ( .A1(n13706), .A2(n10472), .B1(n13705), .B2(n11318), .ZN(
        n3341) );
  AOI221_X2 U3312 ( .B1(FP_REG_FILE_reg_out_29__10_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__10_), .C2(n13517), .A(n3344), .ZN(n3313) );
  OAI22_X2 U3313 ( .A1(n13702), .A2(n10441), .B1(n13701), .B2(n11441), .ZN(
        n3344) );
  NAND4_X2 U3314 ( .A1(n3347), .A2(n3348), .A3(n3349), .A4(n3350), .ZN(n7342)
         );
  NOR4_X2 U3315 ( .A1(n3351), .A2(n3352), .A3(n3353), .A4(n3354), .ZN(n3350)
         );
  OAI221_X2 U3316 ( .B1(n13725), .B2(n11152), .C1(n13723), .C2(n10569), .A(
        n3357), .ZN(n3354) );
  AOI22_X2 U3317 ( .A1(FP_REG_FILE_reg_out_27__9_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__9_), .B2(n13501), .ZN(n3357) );
  OAI221_X2 U3318 ( .B1(n13721), .B2(n10209), .C1(n13719), .C2(n11182), .A(
        n3360), .ZN(n3353) );
  AOI22_X2 U3319 ( .A1(FP_REG_FILE_reg_out_2__9_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__9_), .B2(n13507), .ZN(n3360) );
  OAI221_X2 U3322 ( .B1(n13717), .B2(n11193), .C1(n13715), .C2(n10648), .A(
        n3366), .ZN(n3351) );
  OAI221_X2 U3325 ( .B1(n13713), .B2(n10271), .C1(n13711), .C2(n10408), .A(
        n3371), .ZN(n3368) );
  AOI22_X2 U3326 ( .A1(FP_REG_FILE_reg_out_9__9_), .A2(n13511), .B1(
        ID_EXEC_OUT[245]), .B2(net231305), .ZN(n3371) );
  AOI221_X2 U3329 ( .B1(FP_REG_FILE_reg_out_28__9_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__9_), .C2(n13513), .A(n3375), .ZN(n3348) );
  OAI22_X2 U3330 ( .A1(n13707), .A2(n10471), .B1(n13705), .B2(n11317), .ZN(
        n3375) );
  AOI221_X2 U3331 ( .B1(FP_REG_FILE_reg_out_29__9_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__9_), .C2(n13517), .A(n3378), .ZN(n3347) );
  OAI22_X2 U3332 ( .A1(n13703), .A2(n10440), .B1(n13701), .B2(n11440), .ZN(
        n3378) );
  NAND4_X2 U3333 ( .A1(n3381), .A2(n3382), .A3(n3383), .A4(n3384), .ZN(n7375)
         );
  NOR4_X2 U3334 ( .A1(n3385), .A2(n3386), .A3(n3387), .A4(n3388), .ZN(n3384)
         );
  OAI221_X2 U3335 ( .B1(n13725), .B2(n11151), .C1(n13722), .C2(n10568), .A(
        n3391), .ZN(n3388) );
  AOI22_X2 U3336 ( .A1(FP_REG_FILE_reg_out_27__8_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__8_), .B2(n13501), .ZN(n3391) );
  OAI221_X2 U3337 ( .B1(n13721), .B2(n10208), .C1(n13718), .C2(n11181), .A(
        n3394), .ZN(n3387) );
  AOI22_X2 U3338 ( .A1(FP_REG_FILE_reg_out_2__8_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__8_), .B2(n13507), .ZN(n3394) );
  OAI221_X2 U3341 ( .B1(n13717), .B2(n11192), .C1(n13714), .C2(n10647), .A(
        n3400), .ZN(n3385) );
  OAI221_X2 U3344 ( .B1(n13713), .B2(n10270), .C1(n13710), .C2(n10407), .A(
        n3405), .ZN(n3402) );
  AOI22_X2 U3345 ( .A1(FP_REG_FILE_reg_out_9__8_), .A2(n13511), .B1(
        ID_EXEC_OUT[244]), .B2(net231307), .ZN(n3405) );
  AOI221_X2 U3348 ( .B1(FP_REG_FILE_reg_out_28__8_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__8_), .C2(n13513), .A(n3409), .ZN(n3382) );
  OAI22_X2 U3349 ( .A1(n13707), .A2(n10470), .B1(n13704), .B2(n11316), .ZN(
        n3409) );
  AOI221_X2 U3350 ( .B1(FP_REG_FILE_reg_out_29__8_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__8_), .C2(n13517), .A(n3412), .ZN(n3381) );
  OAI22_X2 U3351 ( .A1(n13703), .A2(n10439), .B1(n13700), .B2(n11439), .ZN(
        n3412) );
  NAND4_X2 U3352 ( .A1(n3415), .A2(n3416), .A3(n3417), .A4(n3418), .ZN(n7404)
         );
  NOR4_X2 U3353 ( .A1(n3419), .A2(n3420), .A3(n3421), .A4(n3422), .ZN(n3418)
         );
  OAI221_X2 U3354 ( .B1(n13725), .B2(n11150), .C1(n13723), .C2(n10567), .A(
        n3425), .ZN(n3422) );
  AOI22_X2 U3355 ( .A1(FP_REG_FILE_reg_out_27__7_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__7_), .B2(n13501), .ZN(n3425) );
  OAI221_X2 U3356 ( .B1(n13721), .B2(n10207), .C1(n13719), .C2(n11180), .A(
        n3428), .ZN(n3421) );
  AOI22_X2 U3357 ( .A1(FP_REG_FILE_reg_out_2__7_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__7_), .B2(n13507), .ZN(n3428) );
  OAI221_X2 U3360 ( .B1(n13717), .B2(n11191), .C1(n13715), .C2(n10646), .A(
        n3434), .ZN(n3419) );
  OAI221_X2 U3363 ( .B1(n13713), .B2(n10269), .C1(n13711), .C2(n10406), .A(
        n3439), .ZN(n3436) );
  AOI22_X2 U3364 ( .A1(FP_REG_FILE_reg_out_9__7_), .A2(n13511), .B1(
        ID_EXEC_OUT[243]), .B2(net231305), .ZN(n3439) );
  AOI221_X2 U3367 ( .B1(FP_REG_FILE_reg_out_28__7_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__7_), .C2(n13513), .A(n3443), .ZN(n3416) );
  OAI22_X2 U3368 ( .A1(n13707), .A2(n10469), .B1(n13705), .B2(n11315), .ZN(
        n3443) );
  AOI221_X2 U3369 ( .B1(FP_REG_FILE_reg_out_29__7_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__7_), .C2(n13517), .A(n3446), .ZN(n3415) );
  OAI22_X2 U3370 ( .A1(n13703), .A2(n10438), .B1(n13701), .B2(n11438), .ZN(
        n3446) );
  NAND4_X2 U3371 ( .A1(n3449), .A2(n3450), .A3(n3451), .A4(n3452), .ZN(n7353)
         );
  NOR4_X2 U3372 ( .A1(n3453), .A2(n3454), .A3(n3455), .A4(n3456), .ZN(n3452)
         );
  OAI221_X2 U3373 ( .B1(n13725), .B2(n11149), .C1(n13722), .C2(n10566), .A(
        n3459), .ZN(n3456) );
  AOI22_X2 U3374 ( .A1(FP_REG_FILE_reg_out_27__6_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__6_), .B2(n13501), .ZN(n3459) );
  OAI221_X2 U3375 ( .B1(n13721), .B2(n10206), .C1(n13718), .C2(n11179), .A(
        n3462), .ZN(n3455) );
  AOI22_X2 U3376 ( .A1(FP_REG_FILE_reg_out_2__6_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__6_), .B2(n13507), .ZN(n3462) );
  OAI221_X2 U3379 ( .B1(n13717), .B2(n11190), .C1(n13714), .C2(n10645), .A(
        n3468), .ZN(n3453) );
  OAI221_X2 U3382 ( .B1(n13713), .B2(n10268), .C1(n13710), .C2(n10405), .A(
        n3473), .ZN(n3470) );
  AOI22_X2 U3383 ( .A1(FP_REG_FILE_reg_out_9__6_), .A2(n13511), .B1(
        ID_EXEC_OUT[242]), .B2(net231305), .ZN(n3473) );
  AOI221_X2 U3386 ( .B1(FP_REG_FILE_reg_out_28__6_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__6_), .C2(n13513), .A(n3477), .ZN(n3450) );
  OAI22_X2 U3387 ( .A1(n13707), .A2(n10468), .B1(n13704), .B2(n11314), .ZN(
        n3477) );
  AOI221_X2 U3388 ( .B1(FP_REG_FILE_reg_out_29__6_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__6_), .C2(n13517), .A(n3480), .ZN(n3449) );
  OAI22_X2 U3389 ( .A1(n13703), .A2(n10437), .B1(n13700), .B2(n11437), .ZN(
        n3480) );
  NAND4_X2 U3390 ( .A1(n3483), .A2(n3484), .A3(n3485), .A4(n3486), .ZN(n7359)
         );
  NOR4_X2 U3391 ( .A1(n3487), .A2(n3488), .A3(n3489), .A4(n3490), .ZN(n3486)
         );
  OAI221_X2 U3392 ( .B1(n13725), .B2(n11148), .C1(n13723), .C2(n10565), .A(
        n3493), .ZN(n3490) );
  AOI22_X2 U3393 ( .A1(FP_REG_FILE_reg_out_27__5_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__5_), .B2(n13501), .ZN(n3493) );
  OAI221_X2 U3394 ( .B1(n13721), .B2(n10205), .C1(n13719), .C2(n11178), .A(
        n3496), .ZN(n3489) );
  AOI22_X2 U3395 ( .A1(FP_REG_FILE_reg_out_2__5_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__5_), .B2(n13507), .ZN(n3496) );
  OAI221_X2 U3398 ( .B1(n13717), .B2(n11189), .C1(n13715), .C2(n10644), .A(
        n3502), .ZN(n3487) );
  OAI221_X2 U3401 ( .B1(n13713), .B2(n10267), .C1(n13711), .C2(n10404), .A(
        n3507), .ZN(n3504) );
  AOI22_X2 U3402 ( .A1(FP_REG_FILE_reg_out_9__5_), .A2(n13511), .B1(
        ID_EXEC_OUT[241]), .B2(net231305), .ZN(n3507) );
  AOI221_X2 U3405 ( .B1(FP_REG_FILE_reg_out_28__5_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__5_), .C2(n13513), .A(n3511), .ZN(n3484) );
  OAI22_X2 U3406 ( .A1(n13707), .A2(n10467), .B1(n13705), .B2(n11313), .ZN(
        n3511) );
  AOI221_X2 U3407 ( .B1(FP_REG_FILE_reg_out_29__5_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__5_), .C2(n13517), .A(n3514), .ZN(n3483) );
  OAI22_X2 U3408 ( .A1(n13703), .A2(n10436), .B1(n13701), .B2(n11436), .ZN(
        n3514) );
  NAND4_X2 U3409 ( .A1(n3517), .A2(n3518), .A3(n3519), .A4(n3520), .ZN(n7321)
         );
  NOR4_X2 U3410 ( .A1(n3521), .A2(n3522), .A3(n3523), .A4(n3524), .ZN(n3520)
         );
  OAI221_X2 U3411 ( .B1(n13725), .B2(n11147), .C1(n13722), .C2(n10564), .A(
        n3527), .ZN(n3524) );
  AOI22_X2 U3412 ( .A1(FP_REG_FILE_reg_out_27__4_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__4_), .B2(n13501), .ZN(n3527) );
  OAI221_X2 U3413 ( .B1(n13721), .B2(n10204), .C1(n13718), .C2(n11177), .A(
        n3530), .ZN(n3523) );
  AOI22_X2 U3414 ( .A1(FP_REG_FILE_reg_out_2__4_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__4_), .B2(n13507), .ZN(n3530) );
  OAI221_X2 U3417 ( .B1(n13717), .B2(n11188), .C1(n13714), .C2(n10643), .A(
        n3536), .ZN(n3521) );
  OAI221_X2 U3420 ( .B1(n13713), .B2(n10266), .C1(n13710), .C2(n10403), .A(
        n3541), .ZN(n3538) );
  AOI22_X2 U3421 ( .A1(FP_REG_FILE_reg_out_9__4_), .A2(n13511), .B1(
        ID_EXEC_OUT[240]), .B2(net231307), .ZN(n3541) );
  AOI221_X2 U3424 ( .B1(FP_REG_FILE_reg_out_28__4_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__4_), .C2(n13513), .A(n3545), .ZN(n3518) );
  OAI22_X2 U3425 ( .A1(n13707), .A2(n10466), .B1(n13704), .B2(n11312), .ZN(
        n3545) );
  AOI221_X2 U3426 ( .B1(FP_REG_FILE_reg_out_29__4_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__4_), .C2(n13517), .A(n3548), .ZN(n3517) );
  OAI22_X2 U3427 ( .A1(n13703), .A2(n10435), .B1(n13700), .B2(n11435), .ZN(
        n3548) );
  NAND4_X2 U3430 ( .A1(n3552), .A2(n3553), .A3(n3554), .A4(n3555), .ZN(n7587)
         );
  NOR4_X2 U3431 ( .A1(n3556), .A2(n3557), .A3(n3558), .A4(n3559), .ZN(n3555)
         );
  OAI221_X2 U3432 ( .B1(n13725), .B2(n11146), .C1(n13723), .C2(n10563), .A(
        n3562), .ZN(n3559) );
  AOI22_X2 U3433 ( .A1(FP_REG_FILE_reg_out_27__3_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__3_), .B2(n13501), .ZN(n3562) );
  OAI221_X2 U3434 ( .B1(n13721), .B2(n10203), .C1(n13719), .C2(n11176), .A(
        n3565), .ZN(n3558) );
  AOI22_X2 U3435 ( .A1(FP_REG_FILE_reg_out_2__3_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__3_), .B2(n13507), .ZN(n3565) );
  OAI221_X2 U3438 ( .B1(n13717), .B2(n11187), .C1(n13715), .C2(n10642), .A(
        n3571), .ZN(n3556) );
  OAI221_X2 U3441 ( .B1(n13713), .B2(n10265), .C1(n13711), .C2(n10402), .A(
        n3576), .ZN(n3573) );
  AOI22_X2 U3442 ( .A1(FP_REG_FILE_reg_out_9__3_), .A2(n13511), .B1(
        ID_EXEC_OUT[239]), .B2(net231305), .ZN(n3576) );
  AOI221_X2 U3445 ( .B1(FP_REG_FILE_reg_out_28__3_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__3_), .C2(n13513), .A(n3580), .ZN(n3553) );
  OAI22_X2 U3446 ( .A1(n13707), .A2(n10465), .B1(n13705), .B2(n11311), .ZN(
        n3580) );
  AOI221_X2 U3447 ( .B1(FP_REG_FILE_reg_out_29__3_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__3_), .C2(n13517), .A(n3583), .ZN(n3552) );
  OAI22_X2 U3448 ( .A1(n13703), .A2(n10434), .B1(n13701), .B2(n11434), .ZN(
        n3583) );
  NAND4_X2 U3449 ( .A1(n3586), .A2(n3587), .A3(n3588), .A4(n3589), .ZN(n7478)
         );
  NOR4_X2 U3450 ( .A1(n3590), .A2(n3591), .A3(n3592), .A4(n3593), .ZN(n3589)
         );
  OAI221_X2 U3451 ( .B1(n13725), .B2(n11145), .C1(n13722), .C2(n10562), .A(
        n3596), .ZN(n3593) );
  AOI22_X2 U3452 ( .A1(FP_REG_FILE_reg_out_27__2_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__2_), .B2(n13501), .ZN(n3596) );
  OAI221_X2 U3453 ( .B1(n13721), .B2(n10202), .C1(n13718), .C2(n11175), .A(
        n3599), .ZN(n3592) );
  AOI22_X2 U3454 ( .A1(FP_REG_FILE_reg_out_2__2_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__2_), .B2(n13507), .ZN(n3599) );
  OAI221_X2 U3457 ( .B1(n13717), .B2(n11186), .C1(n13714), .C2(n10641), .A(
        n3605), .ZN(n3590) );
  OAI221_X2 U3460 ( .B1(n13713), .B2(n10264), .C1(n13710), .C2(n10401), .A(
        n3610), .ZN(n3607) );
  AOI22_X2 U3461 ( .A1(FP_REG_FILE_reg_out_9__2_), .A2(n13511), .B1(
        ID_EXEC_OUT[238]), .B2(net231307), .ZN(n3610) );
  AOI221_X2 U3464 ( .B1(FP_REG_FILE_reg_out_28__2_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__2_), .C2(n13513), .A(n3614), .ZN(n3587) );
  OAI22_X2 U3465 ( .A1(n13707), .A2(n10464), .B1(n13704), .B2(n11310), .ZN(
        n3614) );
  AOI221_X2 U3466 ( .B1(FP_REG_FILE_reg_out_29__2_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__2_), .C2(n13517), .A(n3617), .ZN(n3586) );
  OAI22_X2 U3467 ( .A1(n13703), .A2(n10433), .B1(n13700), .B2(n11433), .ZN(
        n3617) );
  NAND4_X2 U3468 ( .A1(n3620), .A2(n3621), .A3(n3622), .A4(n3623), .ZN(n7531)
         );
  NOR4_X2 U3469 ( .A1(n3624), .A2(n3625), .A3(n3626), .A4(n3627), .ZN(n3623)
         );
  OAI221_X2 U3470 ( .B1(n13725), .B2(n11144), .C1(n13723), .C2(n10561), .A(
        n3630), .ZN(n3627) );
  AOI22_X2 U3471 ( .A1(FP_REG_FILE_reg_out_27__1_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__1_), .B2(n13501), .ZN(n3630) );
  OAI221_X2 U3472 ( .B1(n13721), .B2(n10201), .C1(n13719), .C2(n11174), .A(
        n3633), .ZN(n3626) );
  AOI22_X2 U3473 ( .A1(FP_REG_FILE_reg_out_2__1_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__1_), .B2(n13507), .ZN(n3633) );
  OAI221_X2 U3476 ( .B1(n13717), .B2(n11185), .C1(n13715), .C2(n10640), .A(
        n3639), .ZN(n3624) );
  OAI221_X2 U3479 ( .B1(n13713), .B2(n10399), .C1(n13711), .C2(n10913), .A(
        n3644), .ZN(n3641) );
  AOI22_X2 U3480 ( .A1(FP_REG_FILE_reg_out_9__1_), .A2(n13511), .B1(
        ID_EXEC_OUT[237]), .B2(net231305), .ZN(n3644) );
  AOI221_X2 U3483 ( .B1(FP_REG_FILE_reg_out_28__1_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__1_), .C2(n13513), .A(n3648), .ZN(n3621) );
  OAI22_X2 U3484 ( .A1(n13707), .A2(n10463), .B1(n13705), .B2(n11309), .ZN(
        n3648) );
  AOI221_X2 U3485 ( .B1(FP_REG_FILE_reg_out_29__1_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__1_), .C2(n13517), .A(n3651), .ZN(n3620) );
  OAI22_X2 U3486 ( .A1(n13703), .A2(n10432), .B1(n13701), .B2(n11432), .ZN(
        n3651) );
  NAND4_X2 U3487 ( .A1(n3654), .A2(n3655), .A3(n3656), .A4(n3657), .ZN(n7293)
         );
  NOR4_X2 U3488 ( .A1(n3658), .A2(n3659), .A3(n3660), .A4(n3661), .ZN(n3657)
         );
  OAI221_X2 U3489 ( .B1(n13725), .B2(n11143), .C1(n13722), .C2(n10560), .A(
        n3664), .ZN(n3661) );
  AOI22_X2 U3490 ( .A1(FP_REG_FILE_reg_out_27__0_), .A2(n13505), .B1(
        FP_REG_FILE_reg_out_3__0_), .B2(n13501), .ZN(n3664) );
  OAI221_X2 U3495 ( .B1(n13721), .B2(n10200), .C1(n13718), .C2(n11173), .A(
        n3674), .ZN(n3660) );
  AOI22_X2 U3496 ( .A1(FP_REG_FILE_reg_out_2__0_), .A2(n13509), .B1(
        FP_REG_FILE_reg_out_19__0_), .B2(n13507), .ZN(n3674) );
  OAI221_X2 U3508 ( .B1(n13717), .B2(n11184), .C1(n13714), .C2(n10639), .A(
        n3684), .ZN(n3658) );
  OAI221_X2 U3516 ( .B1(n13713), .B2(n10263), .C1(n13710), .C2(n10400), .A(
        n3689), .ZN(n3686) );
  AOI22_X2 U3517 ( .A1(FP_REG_FILE_reg_out_9__0_), .A2(n13511), .B1(
        ID_EXEC_OUT[236]), .B2(net231305), .ZN(n3689) );
  AOI221_X2 U3527 ( .B1(FP_REG_FILE_reg_out_28__0_), .B2(n13515), .C1(
        FP_REG_FILE_reg_out_4__0_), .C2(n13513), .A(n3695), .ZN(n3655) );
  OAI22_X2 U3528 ( .A1(n13707), .A2(n10462), .B1(n13704), .B2(n11308), .ZN(
        n3695) );
  AOI221_X2 U3534 ( .B1(FP_REG_FILE_reg_out_29__0_), .B2(n13519), .C1(
        FP_REG_FILE_reg_out_5__0_), .C2(n13517), .A(n3699), .ZN(n3654) );
  OAI22_X2 U3535 ( .A1(n13703), .A2(n10431), .B1(n13700), .B2(n11431), .ZN(
        n3699) );
  NAND4_X2 U3546 ( .A1(n3704), .A2(n3705), .A3(n3706), .A4(n3707), .ZN(n8020)
         );
  NOR4_X2 U3547 ( .A1(n3708), .A2(n3709), .A3(n3710), .A4(n3711), .ZN(n3707)
         );
  OAI221_X2 U3548 ( .B1(n10460), .B2(n13698), .C1(n10229), .C2(n13697), .A(
        n3714), .ZN(n3711) );
  AOI22_X2 U3549 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__31_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__31_), .ZN(n3714) );
  OAI221_X2 U3550 ( .B1(n10491), .B2(n13694), .C1(n11307), .C2(n13693), .A(
        n3720), .ZN(n3710) );
  AOI22_X2 U3551 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__31_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__31_), .ZN(n3720) );
  OAI221_X2 U3557 ( .B1(n10291), .B2(n13690), .C1(n11243), .C2(n13689), .A(
        n3743), .ZN(n3739) );
  OAI221_X2 U3559 ( .B1(n10638), .B2(n13686), .C1(n11273), .C2(n13685), .A(
        n3750), .ZN(n3738) );
  AOI22_X2 U3560 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__31_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__31_), .ZN(n3750) );
  AOI221_X2 U3561 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__31_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__31_), .A(n3755), .ZN(n3705) );
  OAI22_X2 U3562 ( .A1(n11495), .A2(n13682), .B1(n11346), .B2(n13681), .ZN(
        n3755) );
  NAND4_X2 U3565 ( .A1(n3765), .A2(n3766), .A3(n3767), .A4(n3768), .ZN(n7733)
         );
  NOR4_X2 U3566 ( .A1(n3769), .A2(n3770), .A3(n3771), .A4(n3772), .ZN(n3768)
         );
  OAI221_X2 U3567 ( .B1(n10459), .B2(n13698), .C1(n10228), .C2(n13696), .A(
        n3773), .ZN(n3772) );
  AOI22_X2 U3568 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__30_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__30_), .ZN(n3773) );
  OAI221_X2 U3569 ( .B1(n10490), .B2(n13694), .C1(n11306), .C2(n13692), .A(
        n3775), .ZN(n3771) );
  AOI22_X2 U3570 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__30_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__30_), .ZN(n3775) );
  OAI221_X2 U3576 ( .B1(n10290), .B2(n13690), .C1(n11242), .C2(n13688), .A(
        n3785), .ZN(n3783) );
  OAI221_X2 U3578 ( .B1(n10637), .B2(n13686), .C1(n11272), .C2(n13684), .A(
        n3788), .ZN(n3782) );
  AOI22_X2 U3579 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__30_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__30_), .ZN(n3788) );
  AOI221_X2 U3580 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__30_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__30_), .A(n3789), .ZN(n3766) );
  OAI22_X2 U3581 ( .A1(n11493), .A2(n13682), .B1(n11345), .B2(n13680), .ZN(
        n3789) );
  NAND4_X2 U3584 ( .A1(n3794), .A2(n3795), .A3(n3796), .A4(n3797), .ZN(n7718)
         );
  NOR4_X2 U3585 ( .A1(n3798), .A2(n3799), .A3(n3800), .A4(n3801), .ZN(n3797)
         );
  OAI221_X2 U3586 ( .B1(n10458), .B2(n13698), .C1(n10227), .C2(n13697), .A(
        n3802), .ZN(n3801) );
  AOI22_X2 U3587 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__29_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__29_), .ZN(n3802) );
  OAI221_X2 U3588 ( .B1(n10489), .B2(n13694), .C1(n11305), .C2(n13693), .A(
        n3804), .ZN(n3800) );
  AOI22_X2 U3589 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__29_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__29_), .ZN(n3804) );
  OAI221_X2 U3595 ( .B1(n10289), .B2(n13690), .C1(n11241), .C2(n13689), .A(
        n3814), .ZN(n3812) );
  OAI221_X2 U3597 ( .B1(n10636), .B2(n13686), .C1(n11271), .C2(n13685), .A(
        n3817), .ZN(n3811) );
  AOI22_X2 U3598 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__29_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__29_), .ZN(n3817) );
  AOI221_X2 U3599 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__29_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__29_), .A(n3818), .ZN(n3795) );
  OAI22_X2 U3600 ( .A1(n11492), .A2(n13682), .B1(n11344), .B2(n13681), .ZN(
        n3818) );
  NAND4_X2 U3603 ( .A1(n3823), .A2(n3824), .A3(n3825), .A4(n3826), .ZN(n7647)
         );
  NOR4_X2 U3604 ( .A1(n3827), .A2(n3828), .A3(n3829), .A4(n3830), .ZN(n3826)
         );
  OAI221_X2 U3605 ( .B1(n10457), .B2(n13698), .C1(n10226), .C2(n13696), .A(
        n3831), .ZN(n3830) );
  AOI22_X2 U3606 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__28_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__28_), .ZN(n3831) );
  OAI221_X2 U3607 ( .B1(n10488), .B2(n13694), .C1(n11304), .C2(n13692), .A(
        n3833), .ZN(n3829) );
  AOI22_X2 U3608 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__28_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__28_), .ZN(n3833) );
  OAI221_X2 U3614 ( .B1(n10288), .B2(n13690), .C1(n11240), .C2(n13688), .A(
        n3843), .ZN(n3841) );
  OAI221_X2 U3616 ( .B1(n10635), .B2(n13686), .C1(n11270), .C2(n13684), .A(
        n3846), .ZN(n3840) );
  AOI22_X2 U3617 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__28_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__28_), .ZN(n3846) );
  AOI221_X2 U3618 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__28_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__28_), .A(n3847), .ZN(n3824) );
  OAI22_X2 U3619 ( .A1(n11491), .A2(n13682), .B1(n11343), .B2(n13680), .ZN(
        n3847) );
  NAND4_X2 U3622 ( .A1(n3852), .A2(n3853), .A3(n3854), .A4(n3855), .ZN(n7706)
         );
  NOR4_X2 U3623 ( .A1(n3856), .A2(n3857), .A3(n3858), .A4(n3859), .ZN(n3855)
         );
  OAI221_X2 U3624 ( .B1(n10456), .B2(n13698), .C1(n10225), .C2(n13697), .A(
        n3860), .ZN(n3859) );
  AOI22_X2 U3625 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__27_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__27_), .ZN(n3860) );
  OAI221_X2 U3626 ( .B1(n10487), .B2(n13694), .C1(n11303), .C2(n13693), .A(
        n3862), .ZN(n3858) );
  AOI22_X2 U3627 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__27_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__27_), .ZN(n3862) );
  OAI221_X2 U3633 ( .B1(n10287), .B2(n13690), .C1(n11239), .C2(n13689), .A(
        n3872), .ZN(n3870) );
  OAI221_X2 U3635 ( .B1(n10634), .B2(n13686), .C1(n11269), .C2(n13685), .A(
        n3875), .ZN(n3869) );
  AOI22_X2 U3636 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__27_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__27_), .ZN(n3875) );
  AOI221_X2 U3637 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__27_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__27_), .A(n3876), .ZN(n3853) );
  OAI22_X2 U3638 ( .A1(n11490), .A2(n13682), .B1(n11342), .B2(n13681), .ZN(
        n3876) );
  NAND4_X2 U3641 ( .A1(n3881), .A2(n3882), .A3(n3883), .A4(n3884), .ZN(n7700)
         );
  NOR4_X2 U3642 ( .A1(n3885), .A2(n3886), .A3(n3887), .A4(n3888), .ZN(n3884)
         );
  OAI221_X2 U3643 ( .B1(n10455), .B2(n13698), .C1(n10224), .C2(n13696), .A(
        n3889), .ZN(n3888) );
  AOI22_X2 U3644 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__26_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__26_), .ZN(n3889) );
  OAI221_X2 U3645 ( .B1(n10486), .B2(n13694), .C1(n11302), .C2(n13692), .A(
        n3891), .ZN(n3887) );
  AOI22_X2 U3646 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__26_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__26_), .ZN(n3891) );
  OAI221_X2 U3652 ( .B1(n10286), .B2(n13690), .C1(n11238), .C2(n13688), .A(
        n3901), .ZN(n3899) );
  OAI221_X2 U3654 ( .B1(n10633), .B2(n13686), .C1(n11268), .C2(n13684), .A(
        n3904), .ZN(n3898) );
  AOI22_X2 U3655 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__26_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__26_), .ZN(n3904) );
  AOI221_X2 U3656 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__26_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__26_), .A(n3905), .ZN(n3882) );
  OAI22_X2 U3657 ( .A1(n11489), .A2(n13682), .B1(n11341), .B2(n13680), .ZN(
        n3905) );
  OAI22_X2 U3660 ( .A1(net231245), .A2(n10810), .B1(n19324), .B2(net230373), 
        .ZN(n7622) );
  NAND4_X2 U3663 ( .A1(n3911), .A2(n3912), .A3(n3913), .A4(n3914), .ZN(n7712)
         );
  NOR4_X2 U3664 ( .A1(n3915), .A2(n3916), .A3(n3917), .A4(n3918), .ZN(n3914)
         );
  OAI221_X2 U3665 ( .B1(n10454), .B2(n13698), .C1(n10223), .C2(n13697), .A(
        n3919), .ZN(n3918) );
  AOI22_X2 U3666 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__25_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__25_), .ZN(n3919) );
  OAI221_X2 U3667 ( .B1(n10485), .B2(n13694), .C1(n11301), .C2(n13693), .A(
        n3921), .ZN(n3917) );
  AOI22_X2 U3668 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__25_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__25_), .ZN(n3921) );
  OAI221_X2 U3674 ( .B1(n10285), .B2(n13690), .C1(n11237), .C2(n13689), .A(
        n3931), .ZN(n3929) );
  OAI221_X2 U3676 ( .B1(n10632), .B2(n13686), .C1(n11267), .C2(n13685), .A(
        n3934), .ZN(n3928) );
  AOI22_X2 U3677 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__25_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__25_), .ZN(n3934) );
  AOI221_X2 U3678 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__25_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__25_), .A(n3935), .ZN(n3912) );
  OAI22_X2 U3679 ( .A1(n11488), .A2(n13682), .B1(n11340), .B2(n13681), .ZN(
        n3935) );
  NAND4_X2 U3682 ( .A1(n3940), .A2(n3941), .A3(n3942), .A4(n3943), .ZN(n7296)
         );
  NOR4_X2 U3683 ( .A1(n3944), .A2(n3945), .A3(n3946), .A4(n3947), .ZN(n3943)
         );
  OAI221_X2 U3684 ( .B1(n10453), .B2(n13698), .C1(n10222), .C2(n13696), .A(
        n3948), .ZN(n3947) );
  AOI22_X2 U3685 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__24_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__24_), .ZN(n3948) );
  OAI221_X2 U3686 ( .B1(n10484), .B2(n13694), .C1(n11300), .C2(n13692), .A(
        n3950), .ZN(n3946) );
  AOI22_X2 U3687 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__24_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__24_), .ZN(n3950) );
  OAI221_X2 U3693 ( .B1(n10284), .B2(n13690), .C1(n11236), .C2(n13688), .A(
        n3960), .ZN(n3958) );
  OAI221_X2 U3695 ( .B1(n10631), .B2(n13686), .C1(n11266), .C2(n13684), .A(
        n3963), .ZN(n3957) );
  AOI22_X2 U3696 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__24_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__24_), .ZN(n3963) );
  AOI221_X2 U3697 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__24_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__24_), .A(n3964), .ZN(n3941) );
  OAI22_X2 U3698 ( .A1(n11487), .A2(n13682), .B1(n11339), .B2(n13680), .ZN(
        n3964) );
  NAND4_X2 U3701 ( .A1(n3969), .A2(n3970), .A3(n3971), .A4(n3972), .ZN(n7300)
         );
  NOR4_X2 U3702 ( .A1(n3973), .A2(n3974), .A3(n3975), .A4(n3976), .ZN(n3972)
         );
  OAI221_X2 U3703 ( .B1(n10452), .B2(n13698), .C1(n10221), .C2(n13697), .A(
        n3977), .ZN(n3976) );
  AOI22_X2 U3704 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__23_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__23_), .ZN(n3977) );
  OAI221_X2 U3705 ( .B1(n10483), .B2(n13694), .C1(n11299), .C2(n13693), .A(
        n3979), .ZN(n3975) );
  AOI22_X2 U3706 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__23_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__23_), .ZN(n3979) );
  OAI221_X2 U3712 ( .B1(n10283), .B2(n13690), .C1(n11235), .C2(n13689), .A(
        n3989), .ZN(n3987) );
  OAI221_X2 U3714 ( .B1(n10630), .B2(n13686), .C1(n11265), .C2(n13685), .A(
        n3992), .ZN(n3986) );
  AOI22_X2 U3715 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__23_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__23_), .ZN(n3992) );
  AOI221_X2 U3716 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__23_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__23_), .A(n3993), .ZN(n3970) );
  OAI22_X2 U3717 ( .A1(n12380), .A2(n13682), .B1(n10740), .B2(n13681), .ZN(
        n3993) );
  NAND4_X2 U3720 ( .A1(n3998), .A2(n3999), .A3(n4000), .A4(n4001), .ZN(n7308)
         );
  NOR4_X2 U3721 ( .A1(n4002), .A2(n4003), .A3(n4004), .A4(n4005), .ZN(n4001)
         );
  OAI221_X2 U3722 ( .B1(n10451), .B2(n13698), .C1(n10220), .C2(n13696), .A(
        n4006), .ZN(n4005) );
  AOI22_X2 U3723 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__22_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__22_), .ZN(n4006) );
  OAI221_X2 U3724 ( .B1(n10482), .B2(n13694), .C1(n11298), .C2(n13692), .A(
        n4008), .ZN(n4004) );
  AOI22_X2 U3725 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__22_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__22_), .ZN(n4008) );
  OAI221_X2 U3731 ( .B1(n10282), .B2(n13690), .C1(n11234), .C2(n13688), .A(
        n4018), .ZN(n4016) );
  OAI221_X2 U3733 ( .B1(n10629), .B2(n13686), .C1(n11264), .C2(n13684), .A(
        n4021), .ZN(n4015) );
  AOI22_X2 U3734 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__22_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__22_), .ZN(n4021) );
  AOI221_X2 U3735 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__22_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__22_), .A(n4022), .ZN(n3999) );
  OAI22_X2 U3736 ( .A1(n12378), .A2(n13682), .B1(n10739), .B2(n13680), .ZN(
        n4022) );
  NAND4_X2 U3739 ( .A1(n4027), .A2(n4028), .A3(n4029), .A4(n4030), .ZN(n7312)
         );
  NOR4_X2 U3740 ( .A1(n4031), .A2(n4032), .A3(n4033), .A4(n4034), .ZN(n4030)
         );
  OAI221_X2 U3741 ( .B1(n10450), .B2(n13698), .C1(n10219), .C2(n13697), .A(
        n4035), .ZN(n4034) );
  AOI22_X2 U3742 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__21_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__21_), .ZN(n4035) );
  OAI221_X2 U3743 ( .B1(n10481), .B2(n13694), .C1(n11297), .C2(n13693), .A(
        n4037), .ZN(n4033) );
  AOI22_X2 U3744 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__21_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__21_), .ZN(n4037) );
  OAI221_X2 U3750 ( .B1(n10281), .B2(n13690), .C1(n11233), .C2(n13689), .A(
        n4047), .ZN(n4045) );
  OAI221_X2 U3752 ( .B1(n10628), .B2(n13686), .C1(n11263), .C2(n13685), .A(
        n4050), .ZN(n4044) );
  AOI22_X2 U3753 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__21_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__21_), .ZN(n4050) );
  AOI221_X2 U3754 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__21_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__21_), .A(n4051), .ZN(n4028) );
  OAI22_X2 U3755 ( .A1(n12376), .A2(n13682), .B1(n10738), .B2(n13681), .ZN(
        n4051) );
  NAND4_X2 U3758 ( .A1(n4056), .A2(n4057), .A3(n4058), .A4(n4059), .ZN(n7317)
         );
  NOR4_X2 U3759 ( .A1(n4060), .A2(n4061), .A3(n4062), .A4(n4063), .ZN(n4059)
         );
  OAI221_X2 U3760 ( .B1(n10915), .B2(n13699), .C1(n10261), .C2(n13696), .A(
        n4064), .ZN(n4063) );
  AOI22_X2 U3761 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__20_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__20_), .ZN(n4064) );
  OAI221_X2 U3762 ( .B1(n10917), .B2(n13695), .C1(n12273), .C2(n13692), .A(
        n4066), .ZN(n4062) );
  AOI22_X2 U3763 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__20_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__20_), .ZN(n4066) );
  OAI221_X2 U3769 ( .B1(n10912), .B2(n13691), .C1(n12257), .C2(n13688), .A(
        n4076), .ZN(n4074) );
  OAI221_X2 U3771 ( .B1(n11142), .B2(n13687), .C1(n12260), .C2(n13684), .A(
        n4079), .ZN(n4073) );
  AOI22_X2 U3772 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__20_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__20_), .ZN(n4079) );
  AOI221_X2 U3773 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__20_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__20_), .A(n4080), .ZN(n4057) );
  OAI22_X2 U3774 ( .A1(n12374), .A2(n13683), .B1(n12283), .B2(n13680), .ZN(
        n4080) );
  NAND4_X2 U3777 ( .A1(n4085), .A2(n4086), .A3(n4087), .A4(n4088), .ZN(n7304)
         );
  NOR4_X2 U3778 ( .A1(n4089), .A2(n4090), .A3(n4091), .A4(n4092), .ZN(n4088)
         );
  OAI221_X2 U3779 ( .B1(n10914), .B2(n13699), .C1(n10260), .C2(n13696), .A(
        n4093), .ZN(n4092) );
  AOI22_X2 U3780 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__19_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__19_), .ZN(n4093) );
  OAI221_X2 U3781 ( .B1(n10916), .B2(n13695), .C1(n12272), .C2(n13692), .A(
        n4095), .ZN(n4091) );
  AOI22_X2 U3782 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__19_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__19_), .ZN(n4095) );
  OAI221_X2 U3788 ( .B1(n10911), .B2(n13691), .C1(n12256), .C2(n13688), .A(
        n4105), .ZN(n4103) );
  OAI221_X2 U3790 ( .B1(n11141), .B2(n13687), .C1(n12259), .C2(n13684), .A(
        n4108), .ZN(n4102) );
  AOI22_X2 U3791 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__19_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__19_), .ZN(n4108) );
  AOI221_X2 U3792 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__19_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__19_), .A(n4109), .ZN(n4086) );
  OAI22_X2 U3793 ( .A1(n12372), .A2(n13683), .B1(n12282), .B2(n13680), .ZN(
        n4109) );
  NAND4_X2 U3796 ( .A1(n4114), .A2(n4115), .A3(n4116), .A4(n4117), .ZN(n7748)
         );
  NOR4_X2 U3797 ( .A1(n4118), .A2(n4119), .A3(n4120), .A4(n4121), .ZN(n4117)
         );
  OAI221_X2 U3798 ( .B1(n10449), .B2(n13699), .C1(n10218), .C2(n13696), .A(
        n4122), .ZN(n4121) );
  AOI22_X2 U3799 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__18_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__18_), .ZN(n4122) );
  OAI221_X2 U3800 ( .B1(n10480), .B2(n13695), .C1(n11296), .C2(n13692), .A(
        n4124), .ZN(n4120) );
  AOI22_X2 U3801 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__18_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__18_), .ZN(n4124) );
  OAI221_X2 U3807 ( .B1(n10280), .B2(n13691), .C1(n11232), .C2(n13688), .A(
        n4134), .ZN(n4132) );
  OAI221_X2 U3809 ( .B1(n10627), .B2(n13687), .C1(n11262), .C2(n13684), .A(
        n4137), .ZN(n4131) );
  AOI22_X2 U3810 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__18_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__18_), .ZN(n4137) );
  AOI221_X2 U3811 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__18_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__18_), .A(n4138), .ZN(n4115) );
  OAI22_X2 U3812 ( .A1(n12370), .A2(n13683), .B1(n10737), .B2(n13680), .ZN(
        n4138) );
  NAND4_X2 U3815 ( .A1(n4143), .A2(n4144), .A3(n4145), .A4(n4146), .ZN(n7338)
         );
  NOR4_X2 U3816 ( .A1(n4147), .A2(n4148), .A3(n4149), .A4(n4150), .ZN(n4146)
         );
  OAI221_X2 U3817 ( .B1(n10448), .B2(n13699), .C1(n10217), .C2(n13696), .A(
        n4151), .ZN(n4150) );
  AOI22_X2 U3818 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__17_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__17_), .ZN(n4151) );
  OAI221_X2 U3819 ( .B1(n10479), .B2(n13695), .C1(n11295), .C2(n13692), .A(
        n4153), .ZN(n4149) );
  AOI22_X2 U3820 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__17_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__17_), .ZN(n4153) );
  OAI221_X2 U3826 ( .B1(n10279), .B2(n13691), .C1(n11231), .C2(n13688), .A(
        n4163), .ZN(n4161) );
  OAI221_X2 U3828 ( .B1(n10626), .B2(n13687), .C1(n11261), .C2(n13684), .A(
        n4166), .ZN(n4160) );
  AOI22_X2 U3829 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__17_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__17_), .ZN(n4166) );
  AOI221_X2 U3830 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__17_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__17_), .A(n4167), .ZN(n4144) );
  OAI22_X2 U3831 ( .A1(n12368), .A2(n13683), .B1(n10736), .B2(n13680), .ZN(
        n4167) );
  NAND4_X2 U3834 ( .A1(n4172), .A2(n4173), .A3(n4174), .A4(n4175), .ZN(n7437)
         );
  NOR4_X2 U3835 ( .A1(n4176), .A2(n4177), .A3(n4178), .A4(n4179), .ZN(n4175)
         );
  OAI221_X2 U3836 ( .B1(n10447), .B2(n13699), .C1(n10216), .C2(n13696), .A(
        n4180), .ZN(n4179) );
  AOI22_X2 U3837 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__16_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__16_), .ZN(n4180) );
  OAI221_X2 U3838 ( .B1(n10478), .B2(n13695), .C1(n11294), .C2(n13692), .A(
        n4182), .ZN(n4178) );
  AOI22_X2 U3839 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__16_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__16_), .ZN(n4182) );
  OAI221_X2 U3845 ( .B1(n10278), .B2(n13691), .C1(n11230), .C2(n13688), .A(
        n4192), .ZN(n4190) );
  OAI221_X2 U3847 ( .B1(n10625), .B2(n13687), .C1(n11260), .C2(n13684), .A(
        n4195), .ZN(n4189) );
  AOI22_X2 U3848 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__16_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__16_), .ZN(n4195) );
  AOI221_X2 U3849 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__16_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__16_), .A(n4196), .ZN(n4173) );
  OAI22_X2 U3850 ( .A1(n12366), .A2(n13683), .B1(n10735), .B2(n13680), .ZN(
        n4196) );
  NAND4_X2 U3855 ( .A1(n4202), .A2(n4203), .A3(n4204), .A4(n4205), .ZN(n7628)
         );
  NOR4_X2 U3856 ( .A1(n4206), .A2(n4207), .A3(n4208), .A4(n4209), .ZN(n4205)
         );
  OAI221_X2 U3857 ( .B1(n10446), .B2(n13699), .C1(n10215), .C2(n13696), .A(
        n4210), .ZN(n4209) );
  AOI22_X2 U3858 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__15_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__15_), .ZN(n4210) );
  OAI221_X2 U3859 ( .B1(n10477), .B2(n13695), .C1(n11293), .C2(n13692), .A(
        n4212), .ZN(n4208) );
  AOI22_X2 U3860 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__15_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__15_), .ZN(n4212) );
  OAI221_X2 U3866 ( .B1(n10277), .B2(n13691), .C1(n11229), .C2(n13688), .A(
        n4222), .ZN(n4220) );
  OAI221_X2 U3868 ( .B1(n10624), .B2(n13687), .C1(n11259), .C2(n13684), .A(
        n4225), .ZN(n4219) );
  AOI22_X2 U3869 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__15_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__15_), .ZN(n4225) );
  AOI221_X2 U3870 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__15_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__15_), .A(n4226), .ZN(n4203) );
  OAI22_X2 U3871 ( .A1(n12364), .A2(n13683), .B1(n10734), .B2(n13680), .ZN(
        n4226) );
  NAND4_X2 U3874 ( .A1(n4231), .A2(n4232), .A3(n4233), .A4(n4234), .ZN(n7611)
         );
  NOR4_X2 U3875 ( .A1(n4235), .A2(n4236), .A3(n4237), .A4(n4238), .ZN(n4234)
         );
  OAI221_X2 U3876 ( .B1(n10445), .B2(n13699), .C1(n10214), .C2(n13696), .A(
        n4239), .ZN(n4238) );
  AOI22_X2 U3877 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__14_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__14_), .ZN(n4239) );
  OAI221_X2 U3878 ( .B1(n10476), .B2(n13695), .C1(n11292), .C2(n13692), .A(
        n4241), .ZN(n4237) );
  AOI22_X2 U3879 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__14_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__14_), .ZN(n4241) );
  OAI221_X2 U3885 ( .B1(n10276), .B2(n13691), .C1(n11228), .C2(n13688), .A(
        n4251), .ZN(n4249) );
  OAI221_X2 U3887 ( .B1(n10623), .B2(n13687), .C1(n11258), .C2(n13684), .A(
        n4254), .ZN(n4248) );
  AOI22_X2 U3888 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__14_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__14_), .ZN(n4254) );
  AOI221_X2 U3889 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__14_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__14_), .A(n4255), .ZN(n4232) );
  OAI22_X2 U3890 ( .A1(n12362), .A2(n13683), .B1(n10733), .B2(n13680), .ZN(
        n4255) );
  NAND4_X2 U3893 ( .A1(n4260), .A2(n4261), .A3(n4262), .A4(n4263), .ZN(n7594)
         );
  NOR4_X2 U3894 ( .A1(n4264), .A2(n4265), .A3(n4266), .A4(n4267), .ZN(n4263)
         );
  OAI221_X2 U3895 ( .B1(n10444), .B2(n13699), .C1(n10213), .C2(n13696), .A(
        n4268), .ZN(n4267) );
  AOI22_X2 U3896 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__13_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__13_), .ZN(n4268) );
  OAI221_X2 U3897 ( .B1(n10475), .B2(n13695), .C1(n11291), .C2(n13692), .A(
        n4270), .ZN(n4266) );
  AOI22_X2 U3898 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__13_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__13_), .ZN(n4270) );
  OAI221_X2 U3904 ( .B1(n10275), .B2(n13691), .C1(n11227), .C2(n13688), .A(
        n4280), .ZN(n4278) );
  OAI221_X2 U3906 ( .B1(n10622), .B2(n13687), .C1(n11257), .C2(n13684), .A(
        n4283), .ZN(n4277) );
  AOI22_X2 U3907 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__13_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__13_), .ZN(n4283) );
  AOI221_X2 U3908 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__13_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__13_), .A(n4284), .ZN(n4261) );
  OAI22_X2 U3909 ( .A1(n12360), .A2(n13683), .B1(n10732), .B2(n13680), .ZN(
        n4284) );
  NAND4_X2 U3912 ( .A1(n4289), .A2(n4290), .A3(n4291), .A4(n4292), .ZN(n7348)
         );
  NOR4_X2 U3913 ( .A1(n4293), .A2(n4294), .A3(n4295), .A4(n4296), .ZN(n4292)
         );
  OAI221_X2 U3914 ( .B1(n10443), .B2(n13699), .C1(n10212), .C2(n13696), .A(
        n4297), .ZN(n4296) );
  AOI22_X2 U3915 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__12_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__12_), .ZN(n4297) );
  OAI221_X2 U3916 ( .B1(n10474), .B2(n13695), .C1(n11290), .C2(n13692), .A(
        n4299), .ZN(n4295) );
  AOI22_X2 U3917 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__12_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__12_), .ZN(n4299) );
  OAI221_X2 U3923 ( .B1(n10274), .B2(n13691), .C1(n11226), .C2(n13688), .A(
        n4309), .ZN(n4307) );
  OAI221_X2 U3925 ( .B1(n10621), .B2(n13687), .C1(n11256), .C2(n13684), .A(
        n4312), .ZN(n4306) );
  AOI22_X2 U3926 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__12_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__12_), .ZN(n4312) );
  AOI221_X2 U3927 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__12_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__12_), .A(n4313), .ZN(n4290) );
  OAI22_X2 U3928 ( .A1(n12358), .A2(n13683), .B1(n10731), .B2(n13680), .ZN(
        n4313) );
  NAND4_X2 U3931 ( .A1(n4318), .A2(n4319), .A3(n4320), .A4(n4321), .ZN(n7395)
         );
  NOR4_X2 U3932 ( .A1(n4322), .A2(n4323), .A3(n4324), .A4(n4325), .ZN(n4321)
         );
  OAI221_X2 U3933 ( .B1(n10442), .B2(n13699), .C1(n10211), .C2(n13696), .A(
        n4326), .ZN(n4325) );
  AOI22_X2 U3934 ( .A1(n13524), .A2(FP_REG_FILE_reg_out_20__11_), .B1(n13522), 
        .B2(FP_REG_FILE_reg_out_19__11_), .ZN(n4326) );
  OAI221_X2 U3935 ( .B1(n10473), .B2(n13695), .C1(n11289), .C2(n13692), .A(
        n4328), .ZN(n4324) );
  AOI22_X2 U3936 ( .A1(n13528), .A2(FP_REG_FILE_reg_out_15__11_), .B1(n13526), 
        .B2(FP_REG_FILE_reg_out_18__11_), .ZN(n4328) );
  OAI221_X2 U3942 ( .B1(n10273), .B2(n13691), .C1(n11225), .C2(n13688), .A(
        n4338), .ZN(n4336) );
  OAI221_X2 U3944 ( .B1(n10620), .B2(n13687), .C1(n11255), .C2(n13684), .A(
        n4341), .ZN(n4335) );
  AOI22_X2 U3945 ( .A1(n13532), .A2(FP_REG_FILE_reg_out_29__11_), .B1(n13530), 
        .B2(FP_REG_FILE_reg_out_30__11_), .ZN(n4341) );
  AOI221_X2 U3946 ( .B1(n13536), .B2(FP_REG_FILE_reg_out_9__11_), .C1(n13534), 
        .C2(FP_REG_FILE_reg_out_4__11_), .A(n4342), .ZN(n4319) );
  OAI22_X2 U3947 ( .A1(n12356), .A2(n13683), .B1(n10730), .B2(n13680), .ZN(
        n4342) );
  NAND4_X2 U3950 ( .A1(n4347), .A2(n4348), .A3(n4349), .A4(n4350), .ZN(n7385)
         );
  NOR4_X2 U3951 ( .A1(n4351), .A2(n4352), .A3(n4353), .A4(n4354), .ZN(n4350)
         );
  OAI221_X2 U3952 ( .B1(n10441), .B2(n13699), .C1(n10210), .C2(n13696), .A(
        n4355), .ZN(n4354) );
  AOI22_X2 U3953 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__10_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__10_), .ZN(n4355) );
  OAI221_X2 U3954 ( .B1(n10472), .B2(n13695), .C1(n11357), .C2(n13692), .A(
        n4357), .ZN(n4353) );
  AOI22_X2 U3955 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__10_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__10_), .ZN(n4357) );
  OAI221_X2 U3961 ( .B1(n10272), .B2(n13691), .C1(n11224), .C2(n13688), .A(
        n4367), .ZN(n4365) );
  OAI221_X2 U3963 ( .B1(n10619), .B2(n13687), .C1(n11254), .C2(n13684), .A(
        n4370), .ZN(n4364) );
  AOI22_X2 U3964 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__10_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__10_), .ZN(n4370) );
  AOI221_X2 U3965 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__10_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__10_), .A(n4371), .ZN(n4348) );
  OAI22_X2 U3966 ( .A1(n12355), .A2(n13683), .B1(n10729), .B2(n13680), .ZN(
        n4371) );
  NAND4_X2 U3969 ( .A1(n4376), .A2(n4377), .A3(n4378), .A4(n4379), .ZN(n7343)
         );
  NOR4_X2 U3970 ( .A1(n4380), .A2(n4381), .A3(n4382), .A4(n4383), .ZN(n4379)
         );
  OAI221_X2 U3971 ( .B1(n10440), .B2(n13699), .C1(n10209), .C2(n13697), .A(
        n4384), .ZN(n4383) );
  AOI22_X2 U3972 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__9_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__9_), .ZN(n4384) );
  OAI221_X2 U3973 ( .B1(n10471), .B2(n13695), .C1(n11356), .C2(n13693), .A(
        n4386), .ZN(n4382) );
  AOI22_X2 U3974 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__9_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__9_), .ZN(n4386) );
  OAI221_X2 U3980 ( .B1(n10271), .B2(n13691), .C1(n11223), .C2(n13689), .A(
        n4396), .ZN(n4394) );
  OAI221_X2 U3982 ( .B1(n10618), .B2(n13687), .C1(n11253), .C2(n13685), .A(
        n4399), .ZN(n4393) );
  AOI22_X2 U3983 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__9_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__9_), .ZN(n4399) );
  AOI221_X2 U3984 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__9_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__9_), .A(n4400), .ZN(n4377) );
  OAI22_X2 U3985 ( .A1(n12354), .A2(n13683), .B1(n10728), .B2(n13681), .ZN(
        n4400) );
  NAND4_X2 U3988 ( .A1(n4405), .A2(n4406), .A3(n4407), .A4(n4408), .ZN(n7376)
         );
  NOR4_X2 U3989 ( .A1(n4409), .A2(n4410), .A3(n4411), .A4(n4412), .ZN(n4408)
         );
  OAI221_X2 U3990 ( .B1(n10439), .B2(n13698), .C1(n10208), .C2(n13697), .A(
        n4413), .ZN(n4412) );
  AOI22_X2 U3991 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__8_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__8_), .ZN(n4413) );
  OAI221_X2 U3992 ( .B1(n10470), .B2(n13694), .C1(n11355), .C2(n13693), .A(
        n4415), .ZN(n4411) );
  AOI22_X2 U3993 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__8_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__8_), .ZN(n4415) );
  OAI221_X2 U3999 ( .B1(n10270), .B2(n13690), .C1(n11222), .C2(n13689), .A(
        n4425), .ZN(n4423) );
  OAI221_X2 U4001 ( .B1(n10617), .B2(n13686), .C1(n11252), .C2(n13685), .A(
        n4428), .ZN(n4422) );
  AOI22_X2 U4002 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__8_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__8_), .ZN(n4428) );
  AOI221_X2 U4003 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__8_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__8_), .A(n4429), .ZN(n4406) );
  OAI22_X2 U4004 ( .A1(n12353), .A2(n13682), .B1(n10727), .B2(n13681), .ZN(
        n4429) );
  NAND4_X2 U4007 ( .A1(n4434), .A2(n4435), .A3(n4436), .A4(n4437), .ZN(n7405)
         );
  NOR4_X2 U4008 ( .A1(n4438), .A2(n4439), .A3(n4440), .A4(n4441), .ZN(n4437)
         );
  OAI221_X2 U4009 ( .B1(n10438), .B2(n13699), .C1(n10207), .C2(n13697), .A(
        n4442), .ZN(n4441) );
  AOI22_X2 U4010 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__7_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__7_), .ZN(n4442) );
  OAI221_X2 U4011 ( .B1(n10469), .B2(n13695), .C1(n11354), .C2(n13693), .A(
        n4444), .ZN(n4440) );
  AOI22_X2 U4012 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__7_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__7_), .ZN(n4444) );
  OAI221_X2 U4018 ( .B1(n10269), .B2(n13691), .C1(n11221), .C2(n13689), .A(
        n4454), .ZN(n4452) );
  OAI221_X2 U4020 ( .B1(n10616), .B2(n13687), .C1(n11251), .C2(n13685), .A(
        n4457), .ZN(n4451) );
  AOI22_X2 U4021 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__7_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__7_), .ZN(n4457) );
  AOI221_X2 U4022 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__7_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__7_), .A(n4458), .ZN(n4435) );
  OAI22_X2 U4023 ( .A1(n12352), .A2(n13683), .B1(n10726), .B2(n13681), .ZN(
        n4458) );
  NAND4_X2 U4026 ( .A1(n4463), .A2(n4464), .A3(n4465), .A4(n4466), .ZN(n7354)
         );
  NOR4_X2 U4027 ( .A1(n4467), .A2(n4468), .A3(n4469), .A4(n4470), .ZN(n4466)
         );
  OAI221_X2 U4028 ( .B1(n10437), .B2(n13698), .C1(n10206), .C2(n13697), .A(
        n4471), .ZN(n4470) );
  AOI22_X2 U4029 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__6_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__6_), .ZN(n4471) );
  OAI221_X2 U4030 ( .B1(n10468), .B2(n13694), .C1(n11353), .C2(n13693), .A(
        n4473), .ZN(n4469) );
  AOI22_X2 U4031 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__6_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__6_), .ZN(n4473) );
  OAI221_X2 U4037 ( .B1(n10268), .B2(n13690), .C1(n11220), .C2(n13689), .A(
        n4483), .ZN(n4481) );
  OAI221_X2 U4039 ( .B1(n10615), .B2(n13686), .C1(n11250), .C2(n13685), .A(
        n4486), .ZN(n4480) );
  AOI22_X2 U4040 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__6_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__6_), .ZN(n4486) );
  AOI221_X2 U4041 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__6_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__6_), .A(n4487), .ZN(n4464) );
  OAI22_X2 U4042 ( .A1(n12351), .A2(n13682), .B1(n10725), .B2(n13681), .ZN(
        n4487) );
  OAI22_X2 U4045 ( .A1(net231245), .A2(n11927), .B1(n19326), .B2(net230373), 
        .ZN(n7582) );
  NAND4_X2 U4047 ( .A1(n4493), .A2(n4494), .A3(n4495), .A4(n4496), .ZN(n7360)
         );
  NOR4_X2 U4048 ( .A1(n4497), .A2(n4498), .A3(n4499), .A4(n4500), .ZN(n4496)
         );
  OAI221_X2 U4049 ( .B1(n10436), .B2(n13699), .C1(n10205), .C2(n13697), .A(
        n4501), .ZN(n4500) );
  AOI22_X2 U4050 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__5_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__5_), .ZN(n4501) );
  OAI221_X2 U4051 ( .B1(n10467), .B2(n13695), .C1(n11352), .C2(n13693), .A(
        n4503), .ZN(n4499) );
  AOI22_X2 U4052 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__5_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__5_), .ZN(n4503) );
  OAI221_X2 U4058 ( .B1(n10267), .B2(n13691), .C1(n11219), .C2(n13689), .A(
        n4513), .ZN(n4511) );
  OAI221_X2 U4060 ( .B1(n10614), .B2(n13687), .C1(n11249), .C2(n13685), .A(
        n4516), .ZN(n4510) );
  AOI22_X2 U4061 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__5_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__5_), .ZN(n4516) );
  AOI221_X2 U4062 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__5_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__5_), .A(n4517), .ZN(n4494) );
  OAI22_X2 U4063 ( .A1(n12350), .A2(n13683), .B1(n10724), .B2(n13681), .ZN(
        n4517) );
  NAND4_X2 U4066 ( .A1(n4522), .A2(n4523), .A3(n4524), .A4(n4525), .ZN(n7322)
         );
  NOR4_X2 U4067 ( .A1(n4526), .A2(n4527), .A3(n4528), .A4(n4529), .ZN(n4525)
         );
  OAI221_X2 U4068 ( .B1(n10435), .B2(n13698), .C1(n10204), .C2(n13697), .A(
        n4530), .ZN(n4529) );
  AOI22_X2 U4069 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__4_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__4_), .ZN(n4530) );
  OAI221_X2 U4070 ( .B1(n10466), .B2(n13694), .C1(n11351), .C2(n13693), .A(
        n4532), .ZN(n4528) );
  AOI22_X2 U4071 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__4_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__4_), .ZN(n4532) );
  OAI221_X2 U4077 ( .B1(n10266), .B2(n13690), .C1(n11218), .C2(n13689), .A(
        n4542), .ZN(n4540) );
  OAI221_X2 U4079 ( .B1(n10613), .B2(n13686), .C1(n11248), .C2(n13685), .A(
        n4545), .ZN(n4539) );
  AOI22_X2 U4080 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__4_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__4_), .ZN(n4545) );
  AOI221_X2 U4081 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__4_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__4_), .A(n4546), .ZN(n4523) );
  OAI22_X2 U4082 ( .A1(n12349), .A2(n13682), .B1(n10723), .B2(n13681), .ZN(
        n4546) );
  NAND4_X2 U4085 ( .A1(n4551), .A2(n4552), .A3(n4553), .A4(n4554), .ZN(n7588)
         );
  NOR4_X2 U4086 ( .A1(n4555), .A2(n4556), .A3(n4557), .A4(n4558), .ZN(n4554)
         );
  OAI221_X2 U4087 ( .B1(n10434), .B2(n13699), .C1(n10203), .C2(n13697), .A(
        n4559), .ZN(n4558) );
  AOI22_X2 U4088 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__3_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__3_), .ZN(n4559) );
  OAI221_X2 U4089 ( .B1(n10465), .B2(n13695), .C1(n11350), .C2(n13693), .A(
        n4561), .ZN(n4557) );
  AOI22_X2 U4090 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__3_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__3_), .ZN(n4561) );
  OAI221_X2 U4096 ( .B1(n10265), .B2(n13691), .C1(n11217), .C2(n13689), .A(
        n4571), .ZN(n4569) );
  OAI221_X2 U4098 ( .B1(n10612), .B2(n13687), .C1(n11247), .C2(n13685), .A(
        n4574), .ZN(n4568) );
  AOI22_X2 U4099 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__3_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__3_), .ZN(n4574) );
  AOI221_X2 U4100 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__3_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__3_), .A(n4575), .ZN(n4552) );
  OAI22_X2 U4101 ( .A1(n12348), .A2(n13683), .B1(n10722), .B2(n13681), .ZN(
        n4575) );
  NAND4_X2 U4104 ( .A1(n4580), .A2(n4581), .A3(n4582), .A4(n4583), .ZN(n7479)
         );
  NOR4_X2 U4105 ( .A1(n4584), .A2(n4585), .A3(n4586), .A4(n4587), .ZN(n4583)
         );
  OAI221_X2 U4106 ( .B1(n10433), .B2(n13698), .C1(n10202), .C2(n13697), .A(
        n4588), .ZN(n4587) );
  AOI22_X2 U4107 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__2_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__2_), .ZN(n4588) );
  OAI221_X2 U4108 ( .B1(n10464), .B2(n13694), .C1(n11349), .C2(n13693), .A(
        n4590), .ZN(n4586) );
  AOI22_X2 U4109 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__2_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__2_), .ZN(n4590) );
  OAI221_X2 U4115 ( .B1(n10264), .B2(n13690), .C1(n11216), .C2(n13689), .A(
        n4600), .ZN(n4598) );
  OAI221_X2 U4117 ( .B1(n10611), .B2(n13686), .C1(n11246), .C2(n13685), .A(
        n4603), .ZN(n4597) );
  AOI22_X2 U4118 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__2_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__2_), .ZN(n4603) );
  AOI221_X2 U4119 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__2_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__2_), .A(n4604), .ZN(n4581) );
  OAI22_X2 U4120 ( .A1(n12347), .A2(n13682), .B1(n10721), .B2(n13681), .ZN(
        n4604) );
  NAND4_X2 U4123 ( .A1(n4609), .A2(n4610), .A3(n4611), .A4(n4612), .ZN(n7532)
         );
  NOR4_X2 U4124 ( .A1(n4613), .A2(n4614), .A3(n4615), .A4(n4616), .ZN(n4612)
         );
  OAI221_X2 U4125 ( .B1(n10432), .B2(n13699), .C1(n10201), .C2(n13697), .A(
        n4617), .ZN(n4616) );
  AOI22_X2 U4126 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__1_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__1_), .ZN(n4617) );
  OAI221_X2 U4127 ( .B1(n10463), .B2(n13695), .C1(n11348), .C2(n13693), .A(
        n4619), .ZN(n4615) );
  AOI22_X2 U4128 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__1_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__1_), .ZN(n4619) );
  OAI221_X2 U4134 ( .B1(n10399), .B2(n13691), .C1(n11215), .C2(n13689), .A(
        n4629), .ZN(n4627) );
  OAI221_X2 U4136 ( .B1(n10610), .B2(n13687), .C1(n11245), .C2(n13685), .A(
        n4632), .ZN(n4626) );
  AOI22_X2 U4137 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__1_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__1_), .ZN(n4632) );
  AOI221_X2 U4138 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__1_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__1_), .A(n4633), .ZN(n4610) );
  OAI22_X2 U4139 ( .A1(n12346), .A2(n13683), .B1(n10720), .B2(n13681), .ZN(
        n4633) );
  NAND4_X2 U4142 ( .A1(n4638), .A2(n4639), .A3(n4640), .A4(n4641), .ZN(n7757)
         );
  NOR4_X2 U4143 ( .A1(n4642), .A2(n4643), .A3(n4644), .A4(n4645), .ZN(n4641)
         );
  OAI221_X2 U4144 ( .B1(n10431), .B2(n13698), .C1(n10200), .C2(n13697), .A(
        n4646), .ZN(n4645) );
  AOI22_X2 U4145 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_20__0_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_19__0_), .ZN(n4646) );
  OAI221_X2 U4150 ( .B1(n10462), .B2(n13694), .C1(n11347), .C2(n13693), .A(
        n4650), .ZN(n4644) );
  AOI22_X2 U4151 ( .A1(n13527), .A2(FP_REG_FILE_reg_out_15__0_), .B1(n13525), 
        .B2(FP_REG_FILE_reg_out_18__0_), .ZN(n4650) );
  OAI221_X2 U4170 ( .B1(n10263), .B2(n13690), .C1(n11214), .C2(n13689), .A(
        n4662), .ZN(n4660) );
  OAI221_X2 U4179 ( .B1(n10609), .B2(n13686), .C1(n11244), .C2(n13685), .A(
        n4665), .ZN(n4659) );
  AOI22_X2 U4180 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_29__0_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_30__0_), .ZN(n4665) );
  AOI221_X2 U4187 ( .B1(n13535), .B2(FP_REG_FILE_reg_out_9__0_), .C1(n13533), 
        .C2(FP_REG_FILE_reg_out_4__0_), .A(n4666), .ZN(n4639) );
  OAI22_X2 U4188 ( .A1(n12345), .A2(n13682), .B1(n10719), .B2(n13681), .ZN(
        n4666) );
  OAI22_X2 U4213 ( .A1(net231245), .A2(n10362), .B1(n12303), .B2(net230373), 
        .ZN(n7540) );
  OAI22_X2 U4215 ( .A1(net231245), .A2(n10242), .B1(n12190), .B2(net230379), 
        .ZN(n7573) );
  OAI22_X2 U5688 ( .A1(net231245), .A2(n11955), .B1(n12189), .B2(net230379), 
        .ZN(n7464) );
  OAI22_X2 U5694 ( .A1(net231245), .A2(n11913), .B1(n5482), .B2(net230379), 
        .ZN(n7841) );
  OAI22_X2 U5701 ( .A1(net231245), .A2(n11915), .B1(n5499), .B2(net230379), 
        .ZN(n7842) );
  OAI22_X2 U5714 ( .A1(net231245), .A2(n10236), .B1(n5518), .B2(net230379), 
        .ZN(n7843) );
  XOR2_X2 U5753 ( .A(n10838), .B(ID_STAGE_imm16_aluA[28]), .Z(n5546) );
  OAI22_X2 U5787 ( .A1(net231245), .A2(n10948), .B1(n12555), .B2(n4685), .ZN(
        n7898) );
  OAI22_X2 U5789 ( .A1(net231245), .A2(n12197), .B1(net230381), .B2(n5558), 
        .ZN(n7881) );
  OAI22_X2 U5851 ( .A1(net231247), .A2(n11921), .B1(n12188), .B2(net230379), 
        .ZN(n7431) );
  AOI22_X2 U5854 ( .A1(net231301), .A2(EXEC_STAGE_imm16_32[23]), .B1(
        ID_STAGE_imm16_aluA[23]), .B2(net230393), .ZN(n5595) );
  AOI22_X2 U5857 ( .A1(net231301), .A2(EXEC_STAGE_imm16_32[21]), .B1(
        ID_STAGE_imm16_aluA[21]), .B2(net230393), .ZN(n5597) );
  OAI22_X2 U5881 ( .A1(net231247), .A2(net137569), .B1(n12300), .B2(net230379), 
        .ZN(n7990) );
  AOI22_X2 U5887 ( .A1(net231301), .A2(EXEC_STAGE_imm26_32[23]), .B1(
        ID_STAGE_imm16_aluA[23]), .B2(net230393), .ZN(n5612) );
  AOI22_X2 U5891 ( .A1(net231301), .A2(EXEC_STAGE_imm26_32[21]), .B1(
        ID_STAGE_imm16_aluA[21]), .B2(net230393), .ZN(n5614) );
  OAI22_X2 U5894 ( .A1(net231247), .A2(n11919), .B1(n19331), .B2(net230379), 
        .ZN(n7418) );
  NAND2_X2 U5899 ( .A1(net230393), .A2(ID_STAGE_imm16_aluA[18]), .ZN(n2559) );
  OAI22_X2 U5915 ( .A1(net231247), .A2(n12216), .B1(n11922), .B2(net230379), 
        .ZN(n7836) );
  OAI22_X2 U5918 ( .A1(net231247), .A2(n12215), .B1(n10824), .B2(net230379), 
        .ZN(n7838) );
  OAI22_X2 U5924 ( .A1(net231247), .A2(n10243), .B1(n15638), .B2(net230379), 
        .ZN(n7331) );
  OAI22_X2 U5926 ( .A1(n10176), .A2(n13678), .B1(n11746), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5928 ( .A1(n10175), .A2(n13678), .B1(n11745), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5930 ( .A1(n10174), .A2(n13678), .B1(n11744), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5932 ( .A1(n10173), .A2(n13678), .B1(n11743), .B2(n5630), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5934 ( .A1(n10172), .A2(n13678), .B1(n11742), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5936 ( .A1(n10171), .A2(n13678), .B1(n11741), .B2(n5630), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5938 ( .A1(n10170), .A2(n13678), .B1(n11740), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5940 ( .A1(n10196), .A2(n13678), .B1(n11739), .B2(n5630), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5942 ( .A1(n10195), .A2(n13678), .B1(n11738), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5944 ( .A1(n10169), .A2(n13678), .B1(n11737), .B2(n5630), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5946 ( .A1(n10194), .A2(n13678), .B1(n12665), .B2(n5630), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5948 ( .A1(n10193), .A2(n13679), .B1(n12664), .B2(n5630), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5950 ( .A1(n10192), .A2(n13679), .B1(n12663), .B2(n5630), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5952 ( .A1(n10191), .A2(n13679), .B1(n12662), .B2(n5630), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5954 ( .A1(n10190), .A2(n13679), .B1(n12661), .B2(n5630), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5956 ( .A1(n10189), .A2(n13679), .B1(n12660), .B2(n5630), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5958 ( .A1(n10188), .A2(n13679), .B1(n12659), .B2(n5630), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5960 ( .A1(n10187), .A2(n13679), .B1(n12658), .B2(n5630), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5962 ( .A1(n10186), .A2(n13679), .B1(n12657), .B2(n5630), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5964 ( .A1(n10239), .A2(n13679), .B1(n12656), .B2(n5630), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5966 ( .A1(n10237), .A2(n13679), .B1(n12655), .B2(n5630), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5968 ( .A1(n10238), .A2(n13679), .B1(n12654), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5970 ( .A1(n10185), .A2(n13679), .B1(n12653), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5972 ( .A1(n10184), .A2(n13678), .B1(n12652), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5974 ( .A1(n10183), .A2(n13679), .B1(n12651), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5976 ( .A1(n10182), .A2(n13678), .B1(n12650), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5978 ( .A1(n10181), .A2(n13679), .B1(n12649), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5980 ( .A1(n10180), .A2(n13678), .B1(n12648), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5982 ( .A1(n10179), .A2(n13679), .B1(n12647), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5984 ( .A1(n10178), .A2(n13678), .B1(n12646), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5986 ( .A1(n10177), .A2(n13679), .B1(n12645), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5988 ( .A1(n10168), .A2(n13678), .B1(n12644), .B2(n13676), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5992 ( .A1(n10176), .A2(n13674), .B1(n10408), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5994 ( .A1(n10175), .A2(n13674), .B1(n10407), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5996 ( .A1(n10174), .A2(n13674), .B1(n10406), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U5998 ( .A1(n10173), .A2(n13674), .B1(n10405), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6000 ( .A1(n10172), .A2(n13674), .B1(n10404), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6002 ( .A1(n10171), .A2(n13674), .B1(n10403), .B2(n5667), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6004 ( .A1(n10170), .A2(n13674), .B1(n10402), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6006 ( .A1(n10196), .A2(n13674), .B1(n10430), .B2(n5667), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6008 ( .A1(n10195), .A2(n13674), .B1(n10429), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6010 ( .A1(n10169), .A2(n13674), .B1(n10401), .B2(n5667), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6012 ( .A1(n10194), .A2(n13674), .B1(n10428), .B2(n5667), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6014 ( .A1(n10193), .A2(n13675), .B1(n10427), .B2(n5667), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6016 ( .A1(n10192), .A2(n13675), .B1(n10426), .B2(n5667), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6018 ( .A1(n10191), .A2(n13675), .B1(n10425), .B2(n5667), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6020 ( .A1(n10190), .A2(n13675), .B1(n10424), .B2(n5667), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6022 ( .A1(n10189), .A2(n13675), .B1(n10423), .B2(n5667), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6024 ( .A1(n10188), .A2(n13675), .B1(n10422), .B2(n5667), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6026 ( .A1(n10187), .A2(n13675), .B1(n10421), .B2(n5667), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6028 ( .A1(n10186), .A2(n13675), .B1(n10420), .B2(n5667), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6030 ( .A1(n10239), .A2(n13675), .B1(n10419), .B2(n5667), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6032 ( .A1(n10237), .A2(n13675), .B1(n10913), .B2(n5667), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6034 ( .A1(n10238), .A2(n13675), .B1(n10418), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6036 ( .A1(n10185), .A2(n13675), .B1(n10417), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6038 ( .A1(n10184), .A2(n13674), .B1(n10416), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6040 ( .A1(n10183), .A2(n13675), .B1(n10415), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6042 ( .A1(n10182), .A2(n13674), .B1(n10414), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6044 ( .A1(n10181), .A2(n13675), .B1(n10413), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6046 ( .A1(n10180), .A2(n13674), .B1(n10412), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6048 ( .A1(n10179), .A2(n13675), .B1(n10411), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6050 ( .A1(n10178), .A2(n13674), .B1(n10410), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6052 ( .A1(n10177), .A2(n13675), .B1(n10409), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6054 ( .A1(n10168), .A2(n13674), .B1(n10400), .B2(n13672), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6058 ( .A1(n10176), .A2(n13670), .B1(n10728), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6060 ( .A1(n10175), .A2(n13670), .B1(n10727), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6062 ( .A1(n10174), .A2(n13670), .B1(n10726), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6064 ( .A1(n10173), .A2(n13670), .B1(n10725), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6066 ( .A1(n10172), .A2(n13670), .B1(n10724), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6068 ( .A1(n10171), .A2(n13670), .B1(n10723), .B2(n5673), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6070 ( .A1(n10170), .A2(n13670), .B1(n10722), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6072 ( .A1(n10196), .A2(n13670), .B1(n11346), .B2(n5673), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6074 ( .A1(n10195), .A2(n13670), .B1(n11345), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6076 ( .A1(n10169), .A2(n13670), .B1(n10721), .B2(n5673), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6078 ( .A1(n10194), .A2(n13670), .B1(n11344), .B2(n5673), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6080 ( .A1(n10193), .A2(n13671), .B1(n11343), .B2(n5673), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6082 ( .A1(n10192), .A2(n13671), .B1(n11342), .B2(n5673), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6084 ( .A1(n10191), .A2(n13671), .B1(n11341), .B2(n5673), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6086 ( .A1(n10190), .A2(n13671), .B1(n11340), .B2(n5673), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6088 ( .A1(n10189), .A2(n13671), .B1(n11339), .B2(n5673), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6090 ( .A1(n10188), .A2(n13671), .B1(n10740), .B2(n5673), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6092 ( .A1(n10187), .A2(n13671), .B1(n10739), .B2(n5673), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6094 ( .A1(n10186), .A2(n13671), .B1(n10738), .B2(n5673), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6096 ( .A1(n10239), .A2(n13671), .B1(n12283), .B2(n5673), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6098 ( .A1(n10237), .A2(n13671), .B1(n10720), .B2(n5673), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6100 ( .A1(n10238), .A2(n13671), .B1(n12282), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6102 ( .A1(n10185), .A2(n13671), .B1(n10737), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6104 ( .A1(n10184), .A2(n13670), .B1(n10736), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6106 ( .A1(n10183), .A2(n13671), .B1(n10735), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6108 ( .A1(n10182), .A2(n13670), .B1(n10734), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6110 ( .A1(n10181), .A2(n13671), .B1(n10733), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6112 ( .A1(n10180), .A2(n13670), .B1(n10732), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6114 ( .A1(n10179), .A2(n13671), .B1(n10731), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6116 ( .A1(n10178), .A2(n13670), .B1(n10730), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6118 ( .A1(n10177), .A2(n13671), .B1(n10729), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6120 ( .A1(n10168), .A2(n13670), .B1(n10719), .B2(n13668), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6124 ( .A1(n10176), .A2(n13666), .B1(n11403), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6126 ( .A1(n10175), .A2(n13666), .B1(n11402), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6128 ( .A1(n10174), .A2(n13666), .B1(n11401), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6130 ( .A1(n10173), .A2(n13666), .B1(n11400), .B2(n5675), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6132 ( .A1(n10172), .A2(n13666), .B1(n11399), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6134 ( .A1(n10171), .A2(n13666), .B1(n11398), .B2(n5675), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6136 ( .A1(n10170), .A2(n13666), .B1(n11397), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6138 ( .A1(n10196), .A2(n13666), .B1(n11396), .B2(n5675), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6140 ( .A1(n10195), .A2(n13666), .B1(n11395), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6142 ( .A1(n10169), .A2(n13666), .B1(n11394), .B2(n5675), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6144 ( .A1(n10194), .A2(n13666), .B1(n11393), .B2(n5675), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6146 ( .A1(n10193), .A2(n13667), .B1(n11392), .B2(n5675), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6148 ( .A1(n10192), .A2(n13667), .B1(n11391), .B2(n5675), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6150 ( .A1(n10191), .A2(n13667), .B1(n11390), .B2(n5675), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6152 ( .A1(n10190), .A2(n13667), .B1(n11389), .B2(n5675), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6154 ( .A1(n10189), .A2(n13667), .B1(n11388), .B2(n5675), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6156 ( .A1(n10188), .A2(n13667), .B1(n11387), .B2(n5675), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6158 ( .A1(n10187), .A2(n13667), .B1(n11386), .B2(n5675), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6160 ( .A1(n10186), .A2(n13667), .B1(n11385), .B2(n5675), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6162 ( .A1(n10239), .A2(n13667), .B1(n11384), .B2(n5675), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6164 ( .A1(n10237), .A2(n13667), .B1(n12284), .B2(n5675), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6166 ( .A1(n10238), .A2(n13667), .B1(n11383), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6168 ( .A1(n10185), .A2(n13667), .B1(n11382), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6170 ( .A1(n10184), .A2(n13666), .B1(n11381), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6172 ( .A1(n10183), .A2(n13667), .B1(n11380), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6174 ( .A1(n10182), .A2(n13666), .B1(n11379), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6176 ( .A1(n10181), .A2(n13667), .B1(n11378), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6178 ( .A1(n10180), .A2(n13666), .B1(n11377), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6180 ( .A1(n10179), .A2(n13667), .B1(n11376), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6182 ( .A1(n10178), .A2(n13666), .B1(n11375), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6184 ( .A1(n10177), .A2(n13667), .B1(n11374), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6186 ( .A1(n10168), .A2(n13666), .B1(n11373), .B2(n13664), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6190 ( .A1(n10176), .A2(n13662), .B1(n10271), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6192 ( .A1(n10175), .A2(n13662), .B1(n10270), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6194 ( .A1(n10174), .A2(n13662), .B1(n10269), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6196 ( .A1(n10173), .A2(n13662), .B1(n10268), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6198 ( .A1(n10172), .A2(n13662), .B1(n10267), .B2(n5679), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6200 ( .A1(n10171), .A2(n13662), .B1(n10266), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6202 ( .A1(n10170), .A2(n13662), .B1(n10265), .B2(n5679), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6204 ( .A1(n10196), .A2(n13662), .B1(n10291), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6206 ( .A1(n10195), .A2(n13662), .B1(n10290), .B2(n5679), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6208 ( .A1(n10169), .A2(n13662), .B1(n10264), .B2(n5679), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6210 ( .A1(n10194), .A2(n13662), .B1(n10289), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6212 ( .A1(n10193), .A2(n13663), .B1(n10288), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6214 ( .A1(n10192), .A2(n13663), .B1(n10287), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6216 ( .A1(n10191), .A2(n13663), .B1(n10286), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6218 ( .A1(n10190), .A2(n13663), .B1(n10285), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6220 ( .A1(n10189), .A2(n13663), .B1(n10284), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6222 ( .A1(n10188), .A2(n13663), .B1(n10283), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6224 ( .A1(n10187), .A2(n13663), .B1(n10282), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6226 ( .A1(n10186), .A2(n13663), .B1(n10281), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6228 ( .A1(n10239), .A2(n13663), .B1(n10912), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6230 ( .A1(n10237), .A2(n13663), .B1(n10399), .B2(n13660), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6232 ( .A1(n10238), .A2(n13663), .B1(n10911), .B2(n5679), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6234 ( .A1(n10185), .A2(n13663), .B1(n10280), .B2(n5679), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6236 ( .A1(n10184), .A2(n13662), .B1(n10279), .B2(n5679), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6238 ( .A1(n10183), .A2(n13663), .B1(n10278), .B2(n5679), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6240 ( .A1(n10182), .A2(n13662), .B1(n10277), .B2(n5679), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6242 ( .A1(n10181), .A2(n13663), .B1(n10276), .B2(n5679), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6244 ( .A1(n10180), .A2(n13662), .B1(n10275), .B2(n5679), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6246 ( .A1(n10179), .A2(n13663), .B1(n10274), .B2(n5679), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6248 ( .A1(n10178), .A2(n13662), .B1(n10273), .B2(n5679), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6250 ( .A1(n10177), .A2(n13663), .B1(n10272), .B2(n5679), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6252 ( .A1(n10168), .A2(n13662), .B1(n10263), .B2(n5679), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6256 ( .A1(n10176), .A2(n13658), .B1(n11756), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6258 ( .A1(n10175), .A2(n13658), .B1(n11755), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6260 ( .A1(n10174), .A2(n13658), .B1(n11754), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6262 ( .A1(n10173), .A2(n13658), .B1(n11753), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6264 ( .A1(n10172), .A2(n13658), .B1(n11752), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6266 ( .A1(n10171), .A2(n13658), .B1(n11751), .B2(n5684), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6268 ( .A1(n10170), .A2(n13658), .B1(n11750), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6270 ( .A1(n10196), .A2(n13658), .B1(n11749), .B2(n5684), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6272 ( .A1(n10195), .A2(n13658), .B1(n11748), .B2(n5684), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6274 ( .A1(n10169), .A2(n13658), .B1(n11747), .B2(n5684), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6276 ( .A1(n10194), .A2(n13658), .B1(n12688), .B2(n5684), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6278 ( .A1(n10193), .A2(n13659), .B1(n12687), .B2(n5684), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6280 ( .A1(n10192), .A2(n13659), .B1(n12686), .B2(n5684), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6282 ( .A1(n10191), .A2(n13659), .B1(n12685), .B2(n5684), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6284 ( .A1(n10190), .A2(n13659), .B1(n12684), .B2(n5684), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6286 ( .A1(n10189), .A2(n13659), .B1(n12683), .B2(n5684), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6288 ( .A1(n10188), .A2(n13659), .B1(n12682), .B2(n5684), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6290 ( .A1(n10187), .A2(n13659), .B1(n12681), .B2(n5684), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6292 ( .A1(n10186), .A2(n13659), .B1(n12680), .B2(n5684), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6294 ( .A1(n10239), .A2(n13659), .B1(n12679), .B2(n5684), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6296 ( .A1(n10237), .A2(n13659), .B1(n12678), .B2(n5684), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6298 ( .A1(n10238), .A2(n13659), .B1(n12677), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6300 ( .A1(n10185), .A2(n13659), .B1(n12676), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6302 ( .A1(n10184), .A2(n13658), .B1(n12675), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6304 ( .A1(n10183), .A2(n13659), .B1(n12674), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6306 ( .A1(n10182), .A2(n13658), .B1(n12673), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6308 ( .A1(n10181), .A2(n13659), .B1(n12672), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6310 ( .A1(n10180), .A2(n13658), .B1(n12671), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6312 ( .A1(n10179), .A2(n13659), .B1(n12670), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6314 ( .A1(n10178), .A2(n13658), .B1(n12669), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6316 ( .A1(n10177), .A2(n13659), .B1(n12668), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6318 ( .A1(n10168), .A2(n13658), .B1(n12667), .B2(n13656), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6322 ( .A1(n10176), .A2(n13654), .B1(n11253), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6324 ( .A1(n10175), .A2(n13654), .B1(n11252), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6326 ( .A1(n10174), .A2(n13654), .B1(n11251), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6328 ( .A1(n10173), .A2(n13654), .B1(n11250), .B2(n5717), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6330 ( .A1(n10172), .A2(n13654), .B1(n11249), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6332 ( .A1(n10171), .A2(n13654), .B1(n11248), .B2(n5717), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6334 ( .A1(n10170), .A2(n13654), .B1(n11247), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6336 ( .A1(n10196), .A2(n13654), .B1(n11273), .B2(n5717), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6338 ( .A1(n10195), .A2(n13654), .B1(n11272), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6340 ( .A1(n10169), .A2(n13654), .B1(n11246), .B2(n5717), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6342 ( .A1(n10194), .A2(n13654), .B1(n11271), .B2(n5717), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6344 ( .A1(n10193), .A2(n13655), .B1(n11270), .B2(n5717), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6346 ( .A1(n10192), .A2(n13655), .B1(n11269), .B2(n5717), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6348 ( .A1(n10191), .A2(n13655), .B1(n11268), .B2(n5717), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6350 ( .A1(n10190), .A2(n13655), .B1(n11267), .B2(n5717), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6352 ( .A1(n10189), .A2(n13655), .B1(n11266), .B2(n5717), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6354 ( .A1(n10188), .A2(n13655), .B1(n11265), .B2(n5717), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6356 ( .A1(n10187), .A2(n13655), .B1(n11264), .B2(n5717), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6358 ( .A1(n10186), .A2(n13655), .B1(n11263), .B2(n5717), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6360 ( .A1(n10239), .A2(n13655), .B1(n12260), .B2(n5717), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6362 ( .A1(n10237), .A2(n13655), .B1(n11245), .B2(n5717), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6364 ( .A1(n10238), .A2(n13655), .B1(n12259), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6366 ( .A1(n10185), .A2(n13655), .B1(n11262), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6368 ( .A1(n10184), .A2(n13654), .B1(n11261), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6370 ( .A1(n10183), .A2(n13655), .B1(n11260), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6372 ( .A1(n10182), .A2(n13654), .B1(n11259), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6374 ( .A1(n10181), .A2(n13655), .B1(n11258), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6376 ( .A1(n10180), .A2(n13654), .B1(n11257), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6378 ( .A1(n10179), .A2(n13655), .B1(n11256), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6380 ( .A1(n10178), .A2(n13654), .B1(n11255), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6382 ( .A1(n10177), .A2(n13655), .B1(n11254), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6384 ( .A1(n10168), .A2(n13654), .B1(n11244), .B2(n13652), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6388 ( .A1(n10176), .A2(n13650), .B1(n11356), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6390 ( .A1(n10175), .A2(n13650), .B1(n11355), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6392 ( .A1(n10174), .A2(n13650), .B1(n11354), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6394 ( .A1(n10173), .A2(n13650), .B1(n11353), .B2(n5721), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6396 ( .A1(n10172), .A2(n13650), .B1(n11352), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6398 ( .A1(n10171), .A2(n13650), .B1(n11351), .B2(n5721), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6400 ( .A1(n10170), .A2(n13650), .B1(n11350), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6402 ( .A1(n10196), .A2(n13650), .B1(n11307), .B2(n5721), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6404 ( .A1(n10195), .A2(n13650), .B1(n11306), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6406 ( .A1(n10169), .A2(n13650), .B1(n11349), .B2(n5721), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6408 ( .A1(n10194), .A2(n13650), .B1(n11305), .B2(n5721), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6410 ( .A1(n10193), .A2(n13651), .B1(n11304), .B2(n5721), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6412 ( .A1(n10192), .A2(n13651), .B1(n11303), .B2(n5721), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6414 ( .A1(n10191), .A2(n13651), .B1(n11302), .B2(n5721), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6416 ( .A1(n10190), .A2(n13651), .B1(n11301), .B2(n5721), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6418 ( .A1(n10189), .A2(n13651), .B1(n11300), .B2(n5721), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6420 ( .A1(n10188), .A2(n13651), .B1(n11299), .B2(n5721), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6422 ( .A1(n10187), .A2(n13651), .B1(n11298), .B2(n5721), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6424 ( .A1(n10186), .A2(n13651), .B1(n11297), .B2(n5721), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6426 ( .A1(n10239), .A2(n13651), .B1(n12273), .B2(n5721), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6428 ( .A1(n10237), .A2(n13651), .B1(n11348), .B2(n5721), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6430 ( .A1(n10238), .A2(n13651), .B1(n12272), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6432 ( .A1(n10185), .A2(n13651), .B1(n11296), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6434 ( .A1(n10184), .A2(n13650), .B1(n11295), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6436 ( .A1(n10183), .A2(n13651), .B1(n11294), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6438 ( .A1(n10182), .A2(n13650), .B1(n11293), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6440 ( .A1(n10181), .A2(n13651), .B1(n11292), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6442 ( .A1(n10180), .A2(n13650), .B1(n11291), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6444 ( .A1(n10179), .A2(n13651), .B1(n11290), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6446 ( .A1(n10178), .A2(n13650), .B1(n11289), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6448 ( .A1(n10177), .A2(n13651), .B1(n11357), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6450 ( .A1(n10168), .A2(n13650), .B1(n11347), .B2(n13648), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6454 ( .A1(n10176), .A2(n13646), .B1(n10672), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6456 ( .A1(n10175), .A2(n13646), .B1(n10671), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6458 ( .A1(n10174), .A2(n13646), .B1(n10670), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6460 ( .A1(n10173), .A2(n13646), .B1(n10669), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6462 ( .A1(n10172), .A2(n13646), .B1(n10668), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6464 ( .A1(n10171), .A2(n13646), .B1(n10667), .B2(n5723), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6466 ( .A1(n10170), .A2(n13646), .B1(n10666), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6468 ( .A1(n10196), .A2(n13646), .B1(n11288), .B2(n5723), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6470 ( .A1(n10195), .A2(n13646), .B1(n11287), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6472 ( .A1(n10169), .A2(n13646), .B1(n10665), .B2(n5723), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6474 ( .A1(n10194), .A2(n13646), .B1(n11286), .B2(n5723), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6476 ( .A1(n10193), .A2(n13647), .B1(n11285), .B2(n5723), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6478 ( .A1(n10192), .A2(n13647), .B1(n11284), .B2(n5723), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6480 ( .A1(n10191), .A2(n13647), .B1(n11283), .B2(n5723), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6482 ( .A1(n10190), .A2(n13647), .B1(n11282), .B2(n5723), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6484 ( .A1(n10189), .A2(n13647), .B1(n11281), .B2(n5723), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6486 ( .A1(n10188), .A2(n13647), .B1(n10664), .B2(n5723), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6488 ( .A1(n10187), .A2(n13647), .B1(n10663), .B2(n5723), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6490 ( .A1(n10186), .A2(n13647), .B1(n10662), .B2(n5723), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6492 ( .A1(n10239), .A2(n13647), .B1(n10661), .B2(n5723), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6494 ( .A1(n10237), .A2(n13647), .B1(n12271), .B2(n5723), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6496 ( .A1(n10238), .A2(n13647), .B1(n10660), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6498 ( .A1(n10185), .A2(n13647), .B1(n10659), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6500 ( .A1(n10184), .A2(n13646), .B1(n10658), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6502 ( .A1(n10183), .A2(n13647), .B1(n10657), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6504 ( .A1(n10182), .A2(n13646), .B1(n10656), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6506 ( .A1(n10181), .A2(n13647), .B1(n10655), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6508 ( .A1(n10180), .A2(n13646), .B1(n10654), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6510 ( .A1(n10179), .A2(n13647), .B1(n10653), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6512 ( .A1(n10178), .A2(n13646), .B1(n10652), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6514 ( .A1(n10177), .A2(n13647), .B1(n10651), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6516 ( .A1(n10168), .A2(n13646), .B1(n10650), .B2(n13644), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6520 ( .A1(n10176), .A2(n13642), .B1(n10471), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6522 ( .A1(n10175), .A2(n13642), .B1(n10470), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6524 ( .A1(n10174), .A2(n13642), .B1(n10469), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6526 ( .A1(n10173), .A2(n13642), .B1(n10468), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6528 ( .A1(n10172), .A2(n13642), .B1(n10467), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6530 ( .A1(n10171), .A2(n13642), .B1(n10466), .B2(n5727), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6532 ( .A1(n10170), .A2(n13642), .B1(n10465), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6534 ( .A1(n10196), .A2(n13642), .B1(n10491), .B2(n5727), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6536 ( .A1(n10195), .A2(n13642), .B1(n10490), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6538 ( .A1(n10169), .A2(n13642), .B1(n10464), .B2(n5727), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6540 ( .A1(n10194), .A2(n13642), .B1(n10489), .B2(n5727), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6542 ( .A1(n10193), .A2(n13643), .B1(n10488), .B2(n5727), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6544 ( .A1(n10192), .A2(n13643), .B1(n10487), .B2(n5727), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6546 ( .A1(n10191), .A2(n13643), .B1(n10486), .B2(n5727), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6548 ( .A1(n10190), .A2(n13643), .B1(n10485), .B2(n5727), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6550 ( .A1(n10189), .A2(n13643), .B1(n10484), .B2(n5727), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6552 ( .A1(n10188), .A2(n13643), .B1(n10483), .B2(n5727), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6554 ( .A1(n10187), .A2(n13643), .B1(n10482), .B2(n5727), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6556 ( .A1(n10186), .A2(n13643), .B1(n10481), .B2(n5727), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6558 ( .A1(n10239), .A2(n13643), .B1(n10917), .B2(n5727), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6560 ( .A1(n10237), .A2(n13643), .B1(n10463), .B2(n5727), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6562 ( .A1(n10238), .A2(n13643), .B1(n10916), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6564 ( .A1(n10185), .A2(n13643), .B1(n10480), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6566 ( .A1(n10184), .A2(n13642), .B1(n10479), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6568 ( .A1(n10183), .A2(n13643), .B1(n10478), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6570 ( .A1(n10182), .A2(n13642), .B1(n10477), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6572 ( .A1(n10181), .A2(n13643), .B1(n10476), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6574 ( .A1(n10180), .A2(n13642), .B1(n10475), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6576 ( .A1(n10179), .A2(n13643), .B1(n10474), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6578 ( .A1(n10178), .A2(n13642), .B1(n10473), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6580 ( .A1(n10177), .A2(n13643), .B1(n10472), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6582 ( .A1(n10168), .A2(n13642), .B1(n10462), .B2(n13640), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6586 ( .A1(n10176), .A2(n13638), .B1(n10648), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6588 ( .A1(n10175), .A2(n13638), .B1(n10647), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6590 ( .A1(n10174), .A2(n13638), .B1(n10646), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6592 ( .A1(n10173), .A2(n13638), .B1(n10645), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6594 ( .A1(n10172), .A2(n13638), .B1(n10644), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6596 ( .A1(n10171), .A2(n13638), .B1(n10643), .B2(n5729), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6598 ( .A1(n10170), .A2(n13638), .B1(n10642), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6600 ( .A1(n10196), .A2(n13638), .B1(n10608), .B2(n5729), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6602 ( .A1(n10195), .A2(n13638), .B1(n10607), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6604 ( .A1(n10169), .A2(n13638), .B1(n10641), .B2(n5729), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6606 ( .A1(n10194), .A2(n13638), .B1(n10606), .B2(n5729), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6608 ( .A1(n10193), .A2(n13639), .B1(n10605), .B2(n5729), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6610 ( .A1(n10192), .A2(n13639), .B1(n10604), .B2(n5729), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6612 ( .A1(n10191), .A2(n13639), .B1(n10603), .B2(n5729), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6614 ( .A1(n10190), .A2(n13639), .B1(n10602), .B2(n5729), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6616 ( .A1(n10189), .A2(n13639), .B1(n10601), .B2(n5729), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6618 ( .A1(n10188), .A2(n13639), .B1(n10600), .B2(n5729), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6620 ( .A1(n10187), .A2(n13639), .B1(n10599), .B2(n5729), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6622 ( .A1(n10186), .A2(n13639), .B1(n10598), .B2(n5729), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6624 ( .A1(n10239), .A2(n13639), .B1(n11140), .B2(n5729), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6626 ( .A1(n10237), .A2(n13639), .B1(n10640), .B2(n5729), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6628 ( .A1(n10238), .A2(n13639), .B1(n11139), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6630 ( .A1(n10185), .A2(n13639), .B1(n10597), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6632 ( .A1(n10184), .A2(n13638), .B1(n10596), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6634 ( .A1(n10183), .A2(n13639), .B1(n10595), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6636 ( .A1(n10182), .A2(n13638), .B1(n10594), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6638 ( .A1(n10181), .A2(n13639), .B1(n10593), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6640 ( .A1(n10180), .A2(n13638), .B1(n10592), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6642 ( .A1(n10179), .A2(n13639), .B1(n10591), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6644 ( .A1(n10178), .A2(n13638), .B1(n10590), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6646 ( .A1(n10177), .A2(n13639), .B1(n10649), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6648 ( .A1(n10168), .A2(n13638), .B1(n10639), .B2(n13636), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6652 ( .A1(n10176), .A2(n13634), .B1(n11781), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6654 ( .A1(n10175), .A2(n13634), .B1(n11780), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6656 ( .A1(n10174), .A2(n13634), .B1(n11779), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6658 ( .A1(n10173), .A2(n13634), .B1(n11778), .B2(n5732), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6660 ( .A1(n10172), .A2(n13634), .B1(n11777), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6662 ( .A1(n10171), .A2(n13634), .B1(n11776), .B2(n5732), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6664 ( .A1(n10170), .A2(n13634), .B1(n11775), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6666 ( .A1(n10196), .A2(n13634), .B1(n11774), .B2(n5732), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6668 ( .A1(n10195), .A2(n13634), .B1(n11773), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6670 ( .A1(n10169), .A2(n13634), .B1(n11772), .B2(n5732), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6672 ( .A1(n10194), .A2(n13634), .B1(n12712), .B2(n5732), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6674 ( .A1(n10193), .A2(n13635), .B1(n12711), .B2(n5732), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6676 ( .A1(n10192), .A2(n13635), .B1(n12710), .B2(n5732), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6678 ( .A1(n10191), .A2(n13635), .B1(n12709), .B2(n5732), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6680 ( .A1(n10190), .A2(n13635), .B1(n12708), .B2(n5732), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6682 ( .A1(n10189), .A2(n13635), .B1(n12707), .B2(n5732), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6684 ( .A1(n10188), .A2(n13635), .B1(n12706), .B2(n5732), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6686 ( .A1(n10187), .A2(n13635), .B1(n12705), .B2(n5732), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6688 ( .A1(n10186), .A2(n13635), .B1(n12704), .B2(n5732), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6690 ( .A1(n10239), .A2(n13635), .B1(n12703), .B2(n5732), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6692 ( .A1(n10237), .A2(n13635), .B1(n12702), .B2(n5732), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6694 ( .A1(n10238), .A2(n13635), .B1(n12701), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6696 ( .A1(n10185), .A2(n13635), .B1(n12700), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6698 ( .A1(n10184), .A2(n13634), .B1(n12699), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6700 ( .A1(n10183), .A2(n13635), .B1(n12698), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6702 ( .A1(n10182), .A2(n13634), .B1(n12697), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6704 ( .A1(n10181), .A2(n13635), .B1(n12696), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6706 ( .A1(n10180), .A2(n13634), .B1(n12695), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6708 ( .A1(n10179), .A2(n13635), .B1(n12694), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6710 ( .A1(n10178), .A2(n13634), .B1(n12693), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6712 ( .A1(n10177), .A2(n13635), .B1(n12692), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6714 ( .A1(n10168), .A2(n13634), .B1(n12691), .B2(n13632), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6718 ( .A1(n10176), .A2(n13630), .B1(n11193), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6720 ( .A1(n10175), .A2(n13630), .B1(n11192), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6722 ( .A1(n10174), .A2(n13630), .B1(n11191), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6724 ( .A1(n10173), .A2(n13630), .B1(n11190), .B2(n5767), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6726 ( .A1(n10172), .A2(n13630), .B1(n11189), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6728 ( .A1(n10171), .A2(n13630), .B1(n11188), .B2(n5767), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6730 ( .A1(n10170), .A2(n13630), .B1(n11187), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6732 ( .A1(n10196), .A2(n13630), .B1(n11213), .B2(n5767), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6734 ( .A1(n10195), .A2(n13630), .B1(n11212), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6736 ( .A1(n10169), .A2(n13630), .B1(n11186), .B2(n5767), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6738 ( .A1(n10194), .A2(n13630), .B1(n11211), .B2(n5767), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6740 ( .A1(n10193), .A2(n13631), .B1(n11210), .B2(n5767), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6742 ( .A1(n10192), .A2(n13631), .B1(n11209), .B2(n5767), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6744 ( .A1(n10191), .A2(n13631), .B1(n11208), .B2(n5767), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6746 ( .A1(n10190), .A2(n13631), .B1(n11207), .B2(n5767), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6748 ( .A1(n10189), .A2(n13631), .B1(n11206), .B2(n5767), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6750 ( .A1(n10188), .A2(n13631), .B1(n11205), .B2(n5767), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6752 ( .A1(n10187), .A2(n13631), .B1(n11204), .B2(n5767), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6754 ( .A1(n10186), .A2(n13631), .B1(n11203), .B2(n5767), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6756 ( .A1(n10239), .A2(n13631), .B1(n12255), .B2(n5767), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6758 ( .A1(n10237), .A2(n13631), .B1(n11185), .B2(n5767), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6760 ( .A1(n10238), .A2(n13631), .B1(n12254), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6762 ( .A1(n10185), .A2(n13631), .B1(n11202), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6764 ( .A1(n10184), .A2(n13630), .B1(n11201), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6766 ( .A1(n10183), .A2(n13631), .B1(n11200), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6768 ( .A1(n10182), .A2(n13630), .B1(n11199), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6770 ( .A1(n10181), .A2(n13631), .B1(n11198), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6772 ( .A1(n10180), .A2(n13630), .B1(n11197), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6774 ( .A1(n10179), .A2(n13631), .B1(n11196), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6776 ( .A1(n10178), .A2(n13630), .B1(n11195), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6778 ( .A1(n10177), .A2(n13631), .B1(n11194), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6780 ( .A1(n10168), .A2(n13630), .B1(n11184), .B2(n13628), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6784 ( .A1(n10176), .A2(n13626), .B1(n11440), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6786 ( .A1(n10175), .A2(n13626), .B1(n11439), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6788 ( .A1(n10174), .A2(n13626), .B1(n11438), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6790 ( .A1(n10173), .A2(n13626), .B1(n11437), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6792 ( .A1(n10172), .A2(n13626), .B1(n11436), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6794 ( .A1(n10171), .A2(n13626), .B1(n11435), .B2(n5769), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6796 ( .A1(n10170), .A2(n13626), .B1(n11434), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6798 ( .A1(n10196), .A2(n13626), .B1(n11460), .B2(n5769), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6800 ( .A1(n10195), .A2(n13626), .B1(n11459), .B2(n5769), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6802 ( .A1(n10169), .A2(n13626), .B1(n11433), .B2(n5769), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6804 ( .A1(n10194), .A2(n13626), .B1(n11458), .B2(n5769), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6806 ( .A1(n10193), .A2(n13627), .B1(n11457), .B2(n5769), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6808 ( .A1(n10192), .A2(n13627), .B1(n11456), .B2(n5769), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6810 ( .A1(n10191), .A2(n13627), .B1(n11455), .B2(n5769), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6812 ( .A1(n10190), .A2(n13627), .B1(n11454), .B2(n5769), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6814 ( .A1(n10189), .A2(n13627), .B1(n11453), .B2(n5769), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6816 ( .A1(n10188), .A2(n13627), .B1(n11452), .B2(n5769), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6818 ( .A1(n10187), .A2(n13627), .B1(n11451), .B2(n5769), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6820 ( .A1(n10186), .A2(n13627), .B1(n11450), .B2(n5769), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6822 ( .A1(n10239), .A2(n13627), .B1(n12297), .B2(n5769), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6824 ( .A1(n10237), .A2(n13627), .B1(n11432), .B2(n5769), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6826 ( .A1(n10238), .A2(n13627), .B1(n12296), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6828 ( .A1(n10185), .A2(n13627), .B1(n11449), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6830 ( .A1(n10184), .A2(n13626), .B1(n11448), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6832 ( .A1(n10183), .A2(n13627), .B1(n11447), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6834 ( .A1(n10182), .A2(n13626), .B1(n11446), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6836 ( .A1(n10181), .A2(n13627), .B1(n11445), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6838 ( .A1(n10180), .A2(n13626), .B1(n11444), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6840 ( .A1(n10179), .A2(n13627), .B1(n11443), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6842 ( .A1(n10178), .A2(n13626), .B1(n11442), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6844 ( .A1(n10177), .A2(n13627), .B1(n11441), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6846 ( .A1(n10168), .A2(n13626), .B1(n11431), .B2(n13624), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6850 ( .A1(n10176), .A2(n13622), .B1(n11152), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6852 ( .A1(n10175), .A2(n13622), .B1(n11151), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6854 ( .A1(n10174), .A2(n13622), .B1(n11150), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6856 ( .A1(n10173), .A2(n13622), .B1(n11149), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6858 ( .A1(n10172), .A2(n13622), .B1(n11148), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6860 ( .A1(n10171), .A2(n13622), .B1(n11147), .B2(n5773), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6862 ( .A1(n10170), .A2(n13622), .B1(n11146), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6864 ( .A1(n10196), .A2(n13622), .B1(n11172), .B2(n5773), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6866 ( .A1(n10195), .A2(n13622), .B1(n11171), .B2(n5773), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6868 ( .A1(n10169), .A2(n13622), .B1(n11145), .B2(n5773), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6870 ( .A1(n10194), .A2(n13622), .B1(n11170), .B2(n5773), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6872 ( .A1(n10193), .A2(n13623), .B1(n11169), .B2(n5773), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6874 ( .A1(n10192), .A2(n13623), .B1(n11168), .B2(n5773), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6876 ( .A1(n10191), .A2(n13623), .B1(n11167), .B2(n5773), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6878 ( .A1(n10190), .A2(n13623), .B1(n11166), .B2(n5773), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6880 ( .A1(n10189), .A2(n13623), .B1(n11165), .B2(n5773), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6882 ( .A1(n10188), .A2(n13623), .B1(n11164), .B2(n5773), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6884 ( .A1(n10187), .A2(n13623), .B1(n11163), .B2(n5773), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6886 ( .A1(n10186), .A2(n13623), .B1(n11162), .B2(n5773), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6888 ( .A1(n10239), .A2(n13623), .B1(n12252), .B2(n5773), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6890 ( .A1(n10237), .A2(n13623), .B1(n11144), .B2(n5773), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6892 ( .A1(n10238), .A2(n13623), .B1(n12251), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6894 ( .A1(n10185), .A2(n13623), .B1(n11161), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6896 ( .A1(n10184), .A2(n13622), .B1(n11160), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6898 ( .A1(n10183), .A2(n13623), .B1(n11159), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6900 ( .A1(n10182), .A2(n13622), .B1(n11158), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6902 ( .A1(n10181), .A2(n13623), .B1(n11157), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6904 ( .A1(n10180), .A2(n13622), .B1(n11156), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6906 ( .A1(n10179), .A2(n13623), .B1(n11155), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6908 ( .A1(n10178), .A2(n13622), .B1(n11154), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6910 ( .A1(n10177), .A2(n13623), .B1(n11153), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6912 ( .A1(n10168), .A2(n13622), .B1(n11143), .B2(n13620), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6918 ( .A1(n10176), .A2(n13618), .B1(n11831), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6921 ( .A1(n10175), .A2(n13618), .B1(n11830), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6924 ( .A1(n10174), .A2(n13618), .B1(n11829), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6927 ( .A1(n10173), .A2(n13618), .B1(n11828), .B2(n5776), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6930 ( .A1(n10172), .A2(n13618), .B1(n11827), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6933 ( .A1(n10171), .A2(n13618), .B1(n11826), .B2(n5776), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6936 ( .A1(n10170), .A2(n13618), .B1(n11825), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6939 ( .A1(n10196), .A2(n13618), .B1(n11036), .B2(n5776), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6942 ( .A1(n10195), .A2(n13618), .B1(n11035), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6945 ( .A1(n10169), .A2(n13618), .B1(n11824), .B2(n5776), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6948 ( .A1(n10194), .A2(n13618), .B1(n12121), .B2(n5776), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6951 ( .A1(n10193), .A2(n13619), .B1(n12120), .B2(n5776), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6954 ( .A1(n10192), .A2(n13619), .B1(n12119), .B2(n5776), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6957 ( .A1(n10191), .A2(n13619), .B1(n12118), .B2(n5776), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6960 ( .A1(n10190), .A2(n13619), .B1(n12117), .B2(n5776), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6963 ( .A1(n10189), .A2(n13619), .B1(n12116), .B2(n5776), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6966 ( .A1(n10188), .A2(n13619), .B1(n12115), .B2(n5776), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6969 ( .A1(n10187), .A2(n13619), .B1(n12114), .B2(n5776), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6972 ( .A1(n10186), .A2(n13619), .B1(n12113), .B2(n5776), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6975 ( .A1(n10239), .A2(n13619), .B1(n12112), .B2(n5776), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6978 ( .A1(n10237), .A2(n13619), .B1(n11823), .B2(n5776), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6981 ( .A1(n10238), .A2(n13619), .B1(n12111), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6984 ( .A1(n10185), .A2(n13619), .B1(n11034), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6987 ( .A1(n10184), .A2(n13618), .B1(n11033), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6990 ( .A1(n10183), .A2(n13619), .B1(n11032), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6993 ( .A1(n10182), .A2(n13618), .B1(n11031), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6996 ( .A1(n10181), .A2(n13619), .B1(n11030), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6999 ( .A1(n10180), .A2(n13618), .B1(n11029), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7002 ( .A1(n10179), .A2(n13619), .B1(n11028), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7005 ( .A1(n10178), .A2(n13618), .B1(n11027), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7008 ( .A1(n10177), .A2(n13619), .B1(n11822), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7011 ( .A1(n10168), .A2(n13618), .B1(n11821), .B2(n13616), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U7017 ( .A1(n12978), .A2(n10947), .ZN(n5774) );
  OAI22_X2 U7020 ( .A1(n12330), .A2(n13614), .B1(n13612), .B2(n5779), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7022 ( .A1(n12329), .A2(n5777), .B1(n13612), .B2(n5780), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7024 ( .A1(n12328), .A2(n13614), .B1(n13612), .B2(n5781), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7026 ( .A1(n12327), .A2(n5777), .B1(n13612), .B2(n5782), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7028 ( .A1(n12326), .A2(n13614), .B1(n13612), .B2(n5783), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7030 ( .A1(n12325), .A2(n5777), .B1(n13612), .B2(n5784), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7032 ( .A1(n12324), .A2(n13614), .B1(n13612), .B2(n5785), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7034 ( .A1(n11486), .A2(n5777), .B1(n13612), .B2(n5786), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7036 ( .A1(n11485), .A2(n13614), .B1(n13612), .B2(n5787), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7038 ( .A1(n12323), .A2(n5777), .B1(n13612), .B2(n5788), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7040 ( .A1(n11484), .A2(n5777), .B1(n13612), .B2(n5789), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7042 ( .A1(n11483), .A2(n5777), .B1(n13613), .B2(n5790), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7044 ( .A1(n11482), .A2(n5777), .B1(n13613), .B2(n5791), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7046 ( .A1(n11481), .A2(n5777), .B1(n13613), .B2(n5792), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7048 ( .A1(n11480), .A2(n5777), .B1(n13613), .B2(n5793), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7050 ( .A1(n11479), .A2(n5777), .B1(n13613), .B2(n5794), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7052 ( .A1(n12344), .A2(n5777), .B1(n13613), .B2(n5795), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7054 ( .A1(n12343), .A2(n13614), .B1(n13613), .B2(n5796), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7056 ( .A1(n12342), .A2(n5777), .B1(n13613), .B2(n5797), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7058 ( .A1(n12341), .A2(n5777), .B1(n13613), .B2(n5798), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7060 ( .A1(n12322), .A2(n5777), .B1(n13613), .B2(n5799), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7062 ( .A1(n12340), .A2(n13614), .B1(n13613), .B2(n5800), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7064 ( .A1(n12339), .A2(n13614), .B1(n13613), .B2(n5801), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7066 ( .A1(n12338), .A2(n13614), .B1(n13612), .B2(n5802), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7068 ( .A1(n12337), .A2(n13614), .B1(n13613), .B2(n5803), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7070 ( .A1(n12336), .A2(n13614), .B1(n13612), .B2(n5804), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7072 ( .A1(n12335), .A2(n13614), .B1(n13613), .B2(n5805), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7074 ( .A1(n12334), .A2(n13614), .B1(n13612), .B2(n5806), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7076 ( .A1(n12333), .A2(n13614), .B1(n13613), .B2(n5807), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7078 ( .A1(n12332), .A2(n13614), .B1(n13612), .B2(n5808), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7080 ( .A1(n12331), .A2(n13614), .B1(n13613), .B2(n5809), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7082 ( .A1(n12321), .A2(n13614), .B1(n13612), .B2(n5810), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7086 ( .A1(n12354), .A2(n13610), .B1(n5779), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7088 ( .A1(n12353), .A2(n5813), .B1(n5780), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7090 ( .A1(n12352), .A2(n13610), .B1(n5781), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7092 ( .A1(n12351), .A2(n5813), .B1(n5782), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7094 ( .A1(n12350), .A2(n13610), .B1(n5783), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7096 ( .A1(n12349), .A2(n5813), .B1(n5784), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7098 ( .A1(n12348), .A2(n13610), .B1(n5785), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7100 ( .A1(n11495), .A2(n5813), .B1(n5786), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7102 ( .A1(n11493), .A2(n13610), .B1(n5787), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7104 ( .A1(n12347), .A2(n5813), .B1(n5788), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7106 ( .A1(n11492), .A2(n5813), .B1(n5789), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7108 ( .A1(n11491), .A2(n5813), .B1(n5790), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7110 ( .A1(n11490), .A2(n5813), .B1(n5791), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7112 ( .A1(n11489), .A2(n5813), .B1(n5792), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7114 ( .A1(n11488), .A2(n5813), .B1(n5793), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7116 ( .A1(n11487), .A2(n5813), .B1(n5794), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7118 ( .A1(n12380), .A2(n5813), .B1(n5795), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7120 ( .A1(n12378), .A2(n13610), .B1(n5796), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7122 ( .A1(n12376), .A2(n5813), .B1(n5797), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7124 ( .A1(n12374), .A2(n5813), .B1(n5798), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7126 ( .A1(n12346), .A2(n5813), .B1(n5799), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7128 ( .A1(n12372), .A2(n13610), .B1(n5800), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7130 ( .A1(n12370), .A2(n13610), .B1(n5801), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7132 ( .A1(n12368), .A2(n13610), .B1(n5802), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7134 ( .A1(n12366), .A2(n13610), .B1(n5803), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7136 ( .A1(n12364), .A2(n13610), .B1(n5804), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7138 ( .A1(n12362), .A2(n13610), .B1(n5805), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7140 ( .A1(n12360), .A2(n13610), .B1(n5806), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7142 ( .A1(n12358), .A2(n13610), .B1(n5807), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7144 ( .A1(n12356), .A2(n13610), .B1(n5808), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7146 ( .A1(n12355), .A2(n13610), .B1(n5809), .B2(n13609), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7148 ( .A1(n12345), .A2(n13610), .B1(n5810), .B2(n13608), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7152 ( .A1(n11616), .A2(n13606), .B1(n5779), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7154 ( .A1(n11615), .A2(n5818), .B1(n5780), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7156 ( .A1(n11614), .A2(n13606), .B1(n5781), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7158 ( .A1(n11613), .A2(n5818), .B1(n5782), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7160 ( .A1(n11612), .A2(n13606), .B1(n5783), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7162 ( .A1(n11611), .A2(n5818), .B1(n5784), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7164 ( .A1(n11610), .A2(n13606), .B1(n5785), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7166 ( .A1(n11609), .A2(n5818), .B1(n5786), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7168 ( .A1(n11608), .A2(n13606), .B1(n5787), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7170 ( .A1(n11607), .A2(n5818), .B1(n5788), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7172 ( .A1(n12626), .A2(n5818), .B1(n5789), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7174 ( .A1(n12625), .A2(n5818), .B1(n5790), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7176 ( .A1(n12624), .A2(n5818), .B1(n5791), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7178 ( .A1(n12623), .A2(n5818), .B1(n5792), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7180 ( .A1(n12622), .A2(n5818), .B1(n5793), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7182 ( .A1(n12621), .A2(n5818), .B1(n5794), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7184 ( .A1(n12620), .A2(n5818), .B1(n5795), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7186 ( .A1(n12619), .A2(n13606), .B1(n5796), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7188 ( .A1(n12618), .A2(n5818), .B1(n5797), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7190 ( .A1(n12617), .A2(n5818), .B1(n5798), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7192 ( .A1(n12616), .A2(n5818), .B1(n5799), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7194 ( .A1(n12615), .A2(n13606), .B1(n5800), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7196 ( .A1(n11606), .A2(n13606), .B1(n5801), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7198 ( .A1(n11605), .A2(n13606), .B1(n5802), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7200 ( .A1(n11604), .A2(n13606), .B1(n5803), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7202 ( .A1(n11603), .A2(n13606), .B1(n5804), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7204 ( .A1(n11602), .A2(n13606), .B1(n5805), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7206 ( .A1(n11601), .A2(n13606), .B1(n5806), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7208 ( .A1(n11600), .A2(n13606), .B1(n5807), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7210 ( .A1(n11599), .A2(n13606), .B1(n5808), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7212 ( .A1(n11598), .A2(n13606), .B1(n5809), .B2(n13605), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7214 ( .A1(n11597), .A2(n13606), .B1(n5810), .B2(n13604), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7220 ( .A1(n12240), .A2(n13602), .B1(n5779), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7222 ( .A1(n12239), .A2(n5853), .B1(n5780), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7224 ( .A1(n12238), .A2(n13602), .B1(n5781), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7226 ( .A1(n12237), .A2(n5853), .B1(n5782), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7228 ( .A1(n12236), .A2(n13602), .B1(n5783), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7230 ( .A1(n12235), .A2(n5853), .B1(n5784), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7232 ( .A1(n12234), .A2(n13602), .B1(n5785), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7234 ( .A1(n11585), .A2(n5853), .B1(n5786), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7236 ( .A1(n11584), .A2(n5853), .B1(n5787), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7238 ( .A1(n12233), .A2(n5853), .B1(n5788), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7240 ( .A1(n12614), .A2(n5853), .B1(n5789), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7242 ( .A1(n12613), .A2(n5853), .B1(n5790), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7244 ( .A1(n12612), .A2(n5853), .B1(n5791), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7246 ( .A1(n12611), .A2(n5853), .B1(n5792), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7248 ( .A1(n12610), .A2(n5853), .B1(n5793), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7250 ( .A1(n12609), .A2(n5853), .B1(n5794), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7252 ( .A1(n12608), .A2(n5853), .B1(n5795), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7254 ( .A1(n12607), .A2(n13602), .B1(n5796), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7256 ( .A1(n12606), .A2(n5853), .B1(n5797), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7258 ( .A1(n12605), .A2(n13602), .B1(n5798), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7260 ( .A1(n12604), .A2(n5853), .B1(n5799), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7262 ( .A1(n12603), .A2(n13602), .B1(n5800), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7264 ( .A1(n12249), .A2(n13602), .B1(n5801), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7266 ( .A1(n12248), .A2(n13602), .B1(n5802), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7268 ( .A1(n12247), .A2(n13602), .B1(n5803), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7270 ( .A1(n12246), .A2(n13602), .B1(n5804), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7272 ( .A1(n12245), .A2(n13602), .B1(n5805), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7274 ( .A1(n12244), .A2(n13602), .B1(n5806), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7276 ( .A1(n12243), .A2(n13602), .B1(n5807), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7278 ( .A1(n12242), .A2(n13602), .B1(n5808), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7280 ( .A1(n12241), .A2(n13602), .B1(n5809), .B2(n13601), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7282 ( .A1(n12232), .A2(n13602), .B1(n5810), .B2(n13600), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7286 ( .A1(n11223), .A2(n13598), .B1(n5779), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7288 ( .A1(n11222), .A2(n5886), .B1(n5780), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7290 ( .A1(n11221), .A2(n13598), .B1(n5781), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7292 ( .A1(n11220), .A2(n5886), .B1(n5782), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7294 ( .A1(n11219), .A2(n13598), .B1(n5783), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7296 ( .A1(n11218), .A2(n5886), .B1(n5784), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7298 ( .A1(n11217), .A2(n13598), .B1(n5785), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7300 ( .A1(n11243), .A2(n5886), .B1(n5786), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7302 ( .A1(n11242), .A2(n13598), .B1(n5787), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7304 ( .A1(n11216), .A2(n5886), .B1(n5788), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7306 ( .A1(n11241), .A2(n5886), .B1(n5789), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7308 ( .A1(n11240), .A2(n5886), .B1(n5790), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7310 ( .A1(n11239), .A2(n5886), .B1(n5791), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7312 ( .A1(n11238), .A2(n5886), .B1(n5792), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7314 ( .A1(n11237), .A2(n5886), .B1(n5793), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7316 ( .A1(n11236), .A2(n5886), .B1(n5794), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7318 ( .A1(n11235), .A2(n5886), .B1(n5795), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7320 ( .A1(n11234), .A2(n13598), .B1(n5796), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7322 ( .A1(n11233), .A2(n5886), .B1(n5797), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7324 ( .A1(n12257), .A2(n5886), .B1(n5798), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7326 ( .A1(n11215), .A2(n5886), .B1(n5799), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7328 ( .A1(n12256), .A2(n13598), .B1(n5800), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7330 ( .A1(n11232), .A2(n13598), .B1(n5801), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7332 ( .A1(n11231), .A2(n13598), .B1(n5802), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7334 ( .A1(n11230), .A2(n13598), .B1(n5803), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7336 ( .A1(n11229), .A2(n13598), .B1(n5804), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7338 ( .A1(n11228), .A2(n13598), .B1(n5805), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7340 ( .A1(n11227), .A2(n13598), .B1(n5806), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7342 ( .A1(n11226), .A2(n13598), .B1(n5807), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7344 ( .A1(n11225), .A2(n13598), .B1(n5808), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7346 ( .A1(n11224), .A2(n13598), .B1(n5809), .B2(n13597), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7348 ( .A1(n11214), .A2(n13598), .B1(n5810), .B2(n13596), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7352 ( .A1(n10618), .A2(n13594), .B1(n5779), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7354 ( .A1(n10617), .A2(n5888), .B1(n5780), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7356 ( .A1(n10616), .A2(n13594), .B1(n5781), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7358 ( .A1(n10615), .A2(n5888), .B1(n5782), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7360 ( .A1(n10614), .A2(n13594), .B1(n5783), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7362 ( .A1(n10613), .A2(n5888), .B1(n5784), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7364 ( .A1(n10612), .A2(n13594), .B1(n5785), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7366 ( .A1(n10638), .A2(n5888), .B1(n5786), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7368 ( .A1(n10637), .A2(n13594), .B1(n5787), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7370 ( .A1(n10611), .A2(n5888), .B1(n5788), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7372 ( .A1(n10636), .A2(n5888), .B1(n5789), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7374 ( .A1(n10635), .A2(n5888), .B1(n5790), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7376 ( .A1(n10634), .A2(n5888), .B1(n5791), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7378 ( .A1(n10633), .A2(n5888), .B1(n5792), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7380 ( .A1(n10632), .A2(n5888), .B1(n5793), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7382 ( .A1(n10631), .A2(n5888), .B1(n5794), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7384 ( .A1(n10630), .A2(n5888), .B1(n5795), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7386 ( .A1(n10629), .A2(n13594), .B1(n5796), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7388 ( .A1(n10628), .A2(n5888), .B1(n5797), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7390 ( .A1(n11142), .A2(n5888), .B1(n5798), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7392 ( .A1(n10610), .A2(n5888), .B1(n5799), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7394 ( .A1(n11141), .A2(n13594), .B1(n5800), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7396 ( .A1(n10627), .A2(n13594), .B1(n5801), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7398 ( .A1(n10626), .A2(n13594), .B1(n5802), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7400 ( .A1(n10625), .A2(n13594), .B1(n5803), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7402 ( .A1(n10624), .A2(n13594), .B1(n5804), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7404 ( .A1(n10623), .A2(n13594), .B1(n5805), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7406 ( .A1(n10622), .A2(n13594), .B1(n5806), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7408 ( .A1(n10621), .A2(n13594), .B1(n5807), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7410 ( .A1(n10620), .A2(n13594), .B1(n5808), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7412 ( .A1(n10619), .A2(n13594), .B1(n5809), .B2(n13593), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7414 ( .A1(n10609), .A2(n13594), .B1(n5810), .B2(n13592), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7420 ( .A1(n10209), .A2(n13590), .B1(n5779), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7422 ( .A1(n10208), .A2(n5891), .B1(n5780), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7424 ( .A1(n10207), .A2(n13590), .B1(n5781), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7426 ( .A1(n10206), .A2(n5891), .B1(n5782), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7428 ( .A1(n10205), .A2(n13590), .B1(n5783), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7430 ( .A1(n10204), .A2(n5891), .B1(n5784), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7432 ( .A1(n10203), .A2(n13590), .B1(n5785), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7434 ( .A1(n10229), .A2(n5891), .B1(n5786), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7436 ( .A1(n10228), .A2(n13590), .B1(n5787), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7438 ( .A1(n10202), .A2(n5891), .B1(n5788), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7440 ( .A1(n10227), .A2(n5891), .B1(n5789), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7442 ( .A1(n10226), .A2(n5891), .B1(n5790), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7444 ( .A1(n10225), .A2(n5891), .B1(n5791), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7446 ( .A1(n10224), .A2(n5891), .B1(n5792), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7448 ( .A1(n10223), .A2(n5891), .B1(n5793), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7450 ( .A1(n10222), .A2(n5891), .B1(n5794), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7452 ( .A1(n10221), .A2(n5891), .B1(n5795), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7454 ( .A1(n10220), .A2(n13590), .B1(n5796), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7456 ( .A1(n10219), .A2(n5891), .B1(n5797), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7458 ( .A1(n10261), .A2(n5891), .B1(n5798), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7460 ( .A1(n10201), .A2(n5891), .B1(n5799), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7462 ( .A1(n10260), .A2(n13590), .B1(n5800), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7464 ( .A1(n10218), .A2(n13590), .B1(n5801), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7466 ( .A1(n10217), .A2(n13590), .B1(n5802), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7468 ( .A1(n10216), .A2(n13590), .B1(n5803), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7470 ( .A1(n10215), .A2(n13590), .B1(n5804), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7472 ( .A1(n10214), .A2(n13590), .B1(n5805), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7474 ( .A1(n10213), .A2(n13590), .B1(n5806), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7476 ( .A1(n10212), .A2(n13590), .B1(n5807), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7478 ( .A1(n10211), .A2(n13590), .B1(n5808), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7480 ( .A1(n10210), .A2(n13590), .B1(n5809), .B2(n13589), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7482 ( .A1(n10200), .A2(n13590), .B1(n5810), .B2(n13588), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7486 ( .A1(n11794), .A2(n13586), .B1(n5779), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7488 ( .A1(n11793), .A2(n5893), .B1(n5780), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7490 ( .A1(n11792), .A2(n13586), .B1(n5781), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7492 ( .A1(n11791), .A2(n5893), .B1(n5782), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7494 ( .A1(n11790), .A2(n13586), .B1(n5783), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7496 ( .A1(n11789), .A2(n5893), .B1(n5784), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7498 ( .A1(n11788), .A2(n13586), .B1(n5785), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7500 ( .A1(n11015), .A2(n5893), .B1(n5786), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7502 ( .A1(n11014), .A2(n13586), .B1(n5787), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7504 ( .A1(n11787), .A2(n5893), .B1(n5788), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7506 ( .A1(n12099), .A2(n5893), .B1(n5789), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7508 ( .A1(n12098), .A2(n5893), .B1(n5790), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7510 ( .A1(n12097), .A2(n5893), .B1(n5791), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7512 ( .A1(n12096), .A2(n5893), .B1(n5792), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7514 ( .A1(n12095), .A2(n5893), .B1(n5793), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7516 ( .A1(n12094), .A2(n5893), .B1(n5794), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7518 ( .A1(n12093), .A2(n5893), .B1(n5795), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7520 ( .A1(n12092), .A2(n13586), .B1(n5796), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7522 ( .A1(n12091), .A2(n5893), .B1(n5797), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7524 ( .A1(n12090), .A2(n5893), .B1(n5798), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7526 ( .A1(n11786), .A2(n5893), .B1(n5799), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7528 ( .A1(n12089), .A2(n13586), .B1(n5800), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7530 ( .A1(n11013), .A2(n13586), .B1(n5801), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7532 ( .A1(n11012), .A2(n13586), .B1(n5802), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7534 ( .A1(n11011), .A2(n13586), .B1(n5803), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7536 ( .A1(n11010), .A2(n13586), .B1(n5804), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7538 ( .A1(n11009), .A2(n13586), .B1(n5805), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7540 ( .A1(n11008), .A2(n13586), .B1(n5806), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7542 ( .A1(n11007), .A2(n13586), .B1(n5807), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7544 ( .A1(n11006), .A2(n13586), .B1(n5808), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7546 ( .A1(n11785), .A2(n13586), .B1(n5809), .B2(n13585), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7548 ( .A1(n11784), .A2(n13586), .B1(n5810), .B2(n13584), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7554 ( .A1(n10440), .A2(n13582), .B1(n5779), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7556 ( .A1(n10439), .A2(n5895), .B1(n5780), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7558 ( .A1(n10438), .A2(n13582), .B1(n5781), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7560 ( .A1(n10437), .A2(n5895), .B1(n5782), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7562 ( .A1(n10436), .A2(n13582), .B1(n5783), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7564 ( .A1(n10435), .A2(n5895), .B1(n5784), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7566 ( .A1(n10434), .A2(n13582), .B1(n5785), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7568 ( .A1(n10460), .A2(n5895), .B1(n5786), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7570 ( .A1(n10459), .A2(n13582), .B1(n5787), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7572 ( .A1(n10433), .A2(n5895), .B1(n5788), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7574 ( .A1(n10458), .A2(n5895), .B1(n5789), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7576 ( .A1(n10457), .A2(n5895), .B1(n5790), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7578 ( .A1(n10456), .A2(n5895), .B1(n5791), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7580 ( .A1(n10455), .A2(n5895), .B1(n5792), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7582 ( .A1(n10454), .A2(n5895), .B1(n5793), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7584 ( .A1(n10453), .A2(n5895), .B1(n5794), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7586 ( .A1(n10452), .A2(n5895), .B1(n5795), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7588 ( .A1(n10451), .A2(n13582), .B1(n5796), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7590 ( .A1(n10450), .A2(n5895), .B1(n5797), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7592 ( .A1(n10915), .A2(n5895), .B1(n5798), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7594 ( .A1(n10432), .A2(n5895), .B1(n5799), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7596 ( .A1(n10914), .A2(n13582), .B1(n5800), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7598 ( .A1(n10449), .A2(n13582), .B1(n5801), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7600 ( .A1(n10448), .A2(n13582), .B1(n5802), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7602 ( .A1(n10447), .A2(n13582), .B1(n5803), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7604 ( .A1(n10446), .A2(n13582), .B1(n5804), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7606 ( .A1(n10445), .A2(n13582), .B1(n5805), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7608 ( .A1(n10444), .A2(n13582), .B1(n5806), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7610 ( .A1(n10443), .A2(n13582), .B1(n5807), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7612 ( .A1(n10442), .A2(n13582), .B1(n5808), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7614 ( .A1(n10441), .A2(n13582), .B1(n5809), .B2(n13581), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7616 ( .A1(n10431), .A2(n13582), .B1(n5810), .B2(n13580), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7620 ( .A1(n10569), .A2(n13578), .B1(n5779), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7622 ( .A1(n10568), .A2(n5897), .B1(n5780), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7624 ( .A1(n10567), .A2(n13578), .B1(n5781), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7626 ( .A1(n10566), .A2(n5897), .B1(n5782), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7628 ( .A1(n10565), .A2(n13578), .B1(n5783), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7630 ( .A1(n10564), .A2(n5897), .B1(n5784), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7632 ( .A1(n10563), .A2(n13578), .B1(n5785), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7634 ( .A1(n10589), .A2(n5897), .B1(n5786), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7636 ( .A1(n10588), .A2(n13578), .B1(n5787), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7638 ( .A1(n10562), .A2(n5897), .B1(n5788), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7640 ( .A1(n10587), .A2(n5897), .B1(n5789), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7642 ( .A1(n10586), .A2(n5897), .B1(n5790), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7644 ( .A1(n10585), .A2(n5897), .B1(n5791), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7646 ( .A1(n10584), .A2(n5897), .B1(n5792), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7648 ( .A1(n10583), .A2(n5897), .B1(n5793), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7650 ( .A1(n10582), .A2(n5897), .B1(n5794), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7652 ( .A1(n10581), .A2(n5897), .B1(n5795), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7654 ( .A1(n10580), .A2(n13578), .B1(n5796), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7656 ( .A1(n10579), .A2(n5897), .B1(n5797), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7658 ( .A1(n11138), .A2(n5897), .B1(n5798), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7660 ( .A1(n10561), .A2(n5897), .B1(n5799), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7662 ( .A1(n11137), .A2(n13578), .B1(n5800), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7664 ( .A1(n10578), .A2(n13578), .B1(n5801), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7666 ( .A1(n10577), .A2(n13578), .B1(n5802), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7668 ( .A1(n10576), .A2(n13578), .B1(n5803), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7670 ( .A1(n10575), .A2(n13578), .B1(n5804), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7672 ( .A1(n10574), .A2(n13578), .B1(n5805), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7674 ( .A1(n10573), .A2(n13578), .B1(n5806), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7676 ( .A1(n10572), .A2(n13578), .B1(n5807), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7678 ( .A1(n10571), .A2(n13578), .B1(n5808), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7680 ( .A1(n10570), .A2(n13578), .B1(n5809), .B2(n13577), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7682 ( .A1(n10560), .A2(n13578), .B1(n5810), .B2(n13576), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7688 ( .A1(n11805), .A2(n13574), .B1(n5779), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7690 ( .A1(n11804), .A2(n5899), .B1(n5780), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7692 ( .A1(n11803), .A2(n13574), .B1(n5781), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7694 ( .A1(n11802), .A2(n5899), .B1(n5782), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7696 ( .A1(n11801), .A2(n13574), .B1(n5783), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7698 ( .A1(n11800), .A2(n5899), .B1(n5784), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7700 ( .A1(n11799), .A2(n13574), .B1(n5785), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7702 ( .A1(n11026), .A2(n5899), .B1(n5786), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7704 ( .A1(n11025), .A2(n13574), .B1(n5787), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7706 ( .A1(n11798), .A2(n5899), .B1(n5788), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7708 ( .A1(n12110), .A2(n5899), .B1(n5789), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7710 ( .A1(n12109), .A2(n5899), .B1(n5790), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7712 ( .A1(n12108), .A2(n5899), .B1(n5791), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7714 ( .A1(n12107), .A2(n5899), .B1(n5792), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7716 ( .A1(n12106), .A2(n5899), .B1(n5793), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7718 ( .A1(n12105), .A2(n5899), .B1(n5794), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7720 ( .A1(n12104), .A2(n5899), .B1(n5795), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7722 ( .A1(n12103), .A2(n13574), .B1(n5796), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7724 ( .A1(n12102), .A2(n5899), .B1(n5797), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7726 ( .A1(n12101), .A2(n5899), .B1(n5798), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7728 ( .A1(n11797), .A2(n5899), .B1(n5799), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7730 ( .A1(n12100), .A2(n13574), .B1(n5800), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7732 ( .A1(n11024), .A2(n13574), .B1(n5801), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7734 ( .A1(n11023), .A2(n13574), .B1(n5802), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7736 ( .A1(n11022), .A2(n13574), .B1(n5803), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7738 ( .A1(n11021), .A2(n13574), .B1(n5804), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7740 ( .A1(n11020), .A2(n13574), .B1(n5805), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7742 ( .A1(n11019), .A2(n13574), .B1(n5806), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7744 ( .A1(n11018), .A2(n13574), .B1(n5807), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7746 ( .A1(n11017), .A2(n13574), .B1(n5808), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7748 ( .A1(n11796), .A2(n13574), .B1(n5809), .B2(n13573), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7750 ( .A1(n11795), .A2(n13574), .B1(n5810), .B2(n13572), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7754 ( .A1(n11691), .A2(n13570), .B1(n5779), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7756 ( .A1(n11690), .A2(n5901), .B1(n5780), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7758 ( .A1(n11689), .A2(n13570), .B1(n5781), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7760 ( .A1(n11688), .A2(n5901), .B1(n5782), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7762 ( .A1(n11687), .A2(n13570), .B1(n5783), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7764 ( .A1(n11686), .A2(n5901), .B1(n5784), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7766 ( .A1(n11685), .A2(n13570), .B1(n5785), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7768 ( .A1(n11496), .A2(n5901), .B1(n5786), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7770 ( .A1(n11494), .A2(n13570), .B1(n5787), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7772 ( .A1(n11684), .A2(n5901), .B1(n5788), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7774 ( .A1(n12078), .A2(n5901), .B1(n5789), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7776 ( .A1(n12077), .A2(n5901), .B1(n5790), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7778 ( .A1(n12076), .A2(n5901), .B1(n5791), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7780 ( .A1(n12075), .A2(n5901), .B1(n5792), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7782 ( .A1(n12074), .A2(n5901), .B1(n5793), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7784 ( .A1(n12073), .A2(n5901), .B1(n5794), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7786 ( .A1(n12381), .A2(n5901), .B1(n5795), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7788 ( .A1(n12379), .A2(n13570), .B1(n5796), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7790 ( .A1(n12377), .A2(n5901), .B1(n5797), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7792 ( .A1(n12375), .A2(n5901), .B1(n5798), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7794 ( .A1(n11683), .A2(n5901), .B1(n5799), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7796 ( .A1(n12373), .A2(n13570), .B1(n5800), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7798 ( .A1(n12371), .A2(n13570), .B1(n5801), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7800 ( .A1(n12369), .A2(n13570), .B1(n5802), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7802 ( .A1(n12367), .A2(n13570), .B1(n5803), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7804 ( .A1(n12365), .A2(n13570), .B1(n5804), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7806 ( .A1(n12363), .A2(n13570), .B1(n5805), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7808 ( .A1(n12361), .A2(n13570), .B1(n5806), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7810 ( .A1(n12359), .A2(n13570), .B1(n5807), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7812 ( .A1(n12357), .A2(n13570), .B1(n5808), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7814 ( .A1(n11682), .A2(n13570), .B1(n5809), .B2(n13569), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7816 ( .A1(n11681), .A2(n13570), .B1(n5810), .B2(n13568), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7824 ( .A1(n11317), .A2(n13566), .B1(n5779), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7826 ( .A1(n11316), .A2(n5903), .B1(n5780), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7828 ( .A1(n11315), .A2(n13566), .B1(n5781), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7830 ( .A1(n11314), .A2(n5903), .B1(n5782), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7832 ( .A1(n11313), .A2(n13566), .B1(n5783), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7834 ( .A1(n11312), .A2(n5903), .B1(n5784), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7836 ( .A1(n11311), .A2(n13566), .B1(n5785), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7838 ( .A1(n11337), .A2(n5903), .B1(n5786), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7840 ( .A1(n11336), .A2(n5903), .B1(n5787), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7842 ( .A1(n11310), .A2(n5903), .B1(n5788), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7844 ( .A1(n11335), .A2(n5903), .B1(n5789), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7846 ( .A1(n11334), .A2(n5903), .B1(n5790), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7848 ( .A1(n11333), .A2(n5903), .B1(n5791), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7850 ( .A1(n11332), .A2(n5903), .B1(n5792), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7852 ( .A1(n11331), .A2(n5903), .B1(n5793), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7854 ( .A1(n11330), .A2(n5903), .B1(n5794), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7856 ( .A1(n11329), .A2(n5903), .B1(n5795), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7858 ( .A1(n11328), .A2(n13566), .B1(n5796), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7860 ( .A1(n11327), .A2(n5903), .B1(n5797), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7862 ( .A1(n12281), .A2(n13566), .B1(n5798), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7864 ( .A1(n11309), .A2(n5903), .B1(n5799), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7866 ( .A1(n12280), .A2(n13566), .B1(n5800), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7868 ( .A1(n11326), .A2(n13566), .B1(n5801), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7870 ( .A1(n11325), .A2(n13566), .B1(n5802), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7872 ( .A1(n11324), .A2(n13566), .B1(n5803), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7874 ( .A1(n11323), .A2(n13566), .B1(n5804), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7876 ( .A1(n11322), .A2(n13566), .B1(n5805), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7878 ( .A1(n11321), .A2(n13566), .B1(n5806), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7880 ( .A1(n11320), .A2(n13566), .B1(n5807), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7882 ( .A1(n11319), .A2(n13566), .B1(n5808), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7884 ( .A1(n11318), .A2(n13566), .B1(n5809), .B2(n13565), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7886 ( .A1(n11308), .A2(n13566), .B1(n5810), .B2(n13564), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7890 ( .A1(n11182), .A2(n13562), .B1(n5779), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7892 ( .A1(n11181), .A2(n5905), .B1(n5780), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7894 ( .A1(n11180), .A2(n13562), .B1(n5781), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7896 ( .A1(n11179), .A2(n5905), .B1(n5782), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7898 ( .A1(n11178), .A2(n13562), .B1(n5783), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7900 ( .A1(n11177), .A2(n5905), .B1(n5784), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7902 ( .A1(n11176), .A2(n13562), .B1(n5785), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7904 ( .A1(n11135), .A2(n5905), .B1(n5786), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7906 ( .A1(n11134), .A2(n13562), .B1(n5787), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7908 ( .A1(n11175), .A2(n5905), .B1(n5788), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7910 ( .A1(n11133), .A2(n5905), .B1(n5789), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7912 ( .A1(n11132), .A2(n5905), .B1(n5790), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7914 ( .A1(n11131), .A2(n5905), .B1(n5791), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7916 ( .A1(n11130), .A2(n5905), .B1(n5792), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7918 ( .A1(n11129), .A2(n5905), .B1(n5793), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7920 ( .A1(n11128), .A2(n5905), .B1(n5794), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7922 ( .A1(n11127), .A2(n5905), .B1(n5795), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7924 ( .A1(n11126), .A2(n13562), .B1(n5796), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7926 ( .A1(n11125), .A2(n5905), .B1(n5797), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7928 ( .A1(n12222), .A2(n5905), .B1(n5798), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7930 ( .A1(n11174), .A2(n5905), .B1(n5799), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7932 ( .A1(n12221), .A2(n13562), .B1(n5800), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7934 ( .A1(n11124), .A2(n13562), .B1(n5801), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7936 ( .A1(n11123), .A2(n13562), .B1(n5802), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7938 ( .A1(n11122), .A2(n13562), .B1(n5803), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7940 ( .A1(n11121), .A2(n13562), .B1(n5804), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7942 ( .A1(n11120), .A2(n13562), .B1(n5805), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7944 ( .A1(n11119), .A2(n13562), .B1(n5806), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7946 ( .A1(n11118), .A2(n13562), .B1(n5807), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7948 ( .A1(n11117), .A2(n13562), .B1(n5808), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7950 ( .A1(n11183), .A2(n13562), .B1(n5809), .B2(n13561), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7952 ( .A1(n11173), .A2(n13562), .B1(n5810), .B2(n13560), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7958 ( .A1(n11680), .A2(n13558), .B1(n5779), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7960 ( .A1(n11679), .A2(n5907), .B1(n5780), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7962 ( .A1(n11678), .A2(n13558), .B1(n5781), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7964 ( .A1(n11677), .A2(n5907), .B1(n5782), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7966 ( .A1(n11676), .A2(n13558), .B1(n5783), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7968 ( .A1(n11675), .A2(n5907), .B1(n5784), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7970 ( .A1(n11674), .A2(n13558), .B1(n5785), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7972 ( .A1(n11673), .A2(n5907), .B1(n5786), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7974 ( .A1(n11672), .A2(n13558), .B1(n5787), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7976 ( .A1(n11671), .A2(n5907), .B1(n5788), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7978 ( .A1(n11670), .A2(n5907), .B1(n5789), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7980 ( .A1(n11669), .A2(n5907), .B1(n5790), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7982 ( .A1(n11668), .A2(n5907), .B1(n5791), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7984 ( .A1(n11667), .A2(n5907), .B1(n5792), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7986 ( .A1(n11666), .A2(n5907), .B1(n5793), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7988 ( .A1(n11665), .A2(n5907), .B1(n5794), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7990 ( .A1(n11664), .A2(n5907), .B1(n5795), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7992 ( .A1(n11663), .A2(n13558), .B1(n5796), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7994 ( .A1(n11662), .A2(n5907), .B1(n5797), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7996 ( .A1(n11661), .A2(n5907), .B1(n5798), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7998 ( .A1(n11660), .A2(n5907), .B1(n5799), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8000 ( .A1(n11659), .A2(n13558), .B1(n5800), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8002 ( .A1(n11658), .A2(n13558), .B1(n5801), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8004 ( .A1(n11657), .A2(n13558), .B1(n5802), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8006 ( .A1(n11656), .A2(n13558), .B1(n5803), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8008 ( .A1(n11655), .A2(n13558), .B1(n5804), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8010 ( .A1(n11654), .A2(n13558), .B1(n5805), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8012 ( .A1(n11653), .A2(n13558), .B1(n5806), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8014 ( .A1(n11652), .A2(n13558), .B1(n5807), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8016 ( .A1(n11651), .A2(n13558), .B1(n5808), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8018 ( .A1(n11650), .A2(n13558), .B1(n5809), .B2(n13557), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8020 ( .A1(n11649), .A2(n13558), .B1(n5810), .B2(n13556), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8028 ( .A1(n11648), .A2(n13554), .B1(n5779), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8031 ( .A1(n11647), .A2(n5910), .B1(n5780), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8034 ( .A1(n11646), .A2(n13554), .B1(n5781), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8037 ( .A1(n11645), .A2(n5910), .B1(n5782), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8040 ( .A1(n11644), .A2(n13554), .B1(n5783), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8043 ( .A1(n11643), .A2(n5910), .B1(n5784), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8046 ( .A1(n11642), .A2(n13554), .B1(n5785), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8049 ( .A1(n11641), .A2(n5910), .B1(n5786), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8052 ( .A1(n11640), .A2(n13554), .B1(n5787), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8055 ( .A1(n11639), .A2(n5910), .B1(n5788), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8058 ( .A1(n11638), .A2(n5910), .B1(n5789), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8061 ( .A1(n11637), .A2(n5910), .B1(n5790), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8064 ( .A1(n11636), .A2(n5910), .B1(n5791), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8067 ( .A1(n11635), .A2(n5910), .B1(n5792), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8070 ( .A1(n11634), .A2(n5910), .B1(n5793), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8073 ( .A1(n11633), .A2(n5910), .B1(n5794), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8076 ( .A1(n11632), .A2(n5910), .B1(n5795), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8079 ( .A1(n11631), .A2(n13554), .B1(n5796), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8082 ( .A1(n11630), .A2(n5910), .B1(n5797), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8085 ( .A1(n11629), .A2(n5910), .B1(n5798), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8088 ( .A1(n11628), .A2(n5910), .B1(n5799), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8091 ( .A1(n11627), .A2(n13554), .B1(n5800), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8094 ( .A1(n11626), .A2(n13554), .B1(n5801), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8097 ( .A1(n11625), .A2(n13554), .B1(n5802), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8100 ( .A1(n11624), .A2(n13554), .B1(n5803), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8103 ( .A1(n11623), .A2(n13554), .B1(n5804), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8106 ( .A1(n11622), .A2(n13554), .B1(n5805), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8109 ( .A1(n11621), .A2(n13554), .B1(n5806), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8112 ( .A1(n11620), .A2(n13554), .B1(n5807), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8115 ( .A1(n11619), .A2(n13554), .B1(n5808), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8118 ( .A1(n11618), .A2(n13554), .B1(n5809), .B2(n13553), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8121 ( .A1(n11617), .A2(n13554), .B1(n5810), .B2(n13552), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U8129 ( .A1(MEM_WB_OUT[112]), .A2(n12978), .ZN(n5909) );
  OAI22_X2 U8275 ( .A1(net231247), .A2(n11554), .B1(net230381), .B2(n10357), 
        .ZN(n7506) );
  OAI22_X2 U8445 ( .A1(net231247), .A2(n11553), .B1(net230381), .B2(n10366), 
        .ZN(n7412) );
  OAI22_X2 U8625 ( .A1(net231247), .A2(n11552), .B1(net230381), .B2(n10356), 
        .ZN(n7501) );
  OAI22_X2 U8797 ( .A1(net231247), .A2(n19319), .B1(net230381), .B2(n12184), 
        .ZN(n7875) );
  OAI22_X2 U8800 ( .A1(net231239), .A2(n19316), .B1(net230381), .B2(n12307), 
        .ZN(n7883) );
  OAI22_X2 U8803 ( .A1(net231247), .A2(n19314), .B1(net230381), .B2(n12183), 
        .ZN(n7886) );
  OAI22_X2 U8806 ( .A1(net231247), .A2(n19312), .B1(net230381), .B2(n12306), 
        .ZN(n7889) );
  OAI22_X2 U8809 ( .A1(net231247), .A2(n19310), .B1(net230381), .B2(n12182), 
        .ZN(n7892) );
  OAI22_X2 U8812 ( .A1(net231247), .A2(n11551), .B1(net230381), .B2(n10355), 
        .ZN(n7496) );
  OAI22_X2 U8814 ( .A1(net231245), .A2(n11550), .B1(net230383), .B2(n11914), 
        .ZN(n7552) );
  OAI22_X2 U8816 ( .A1(net231245), .A2(n11549), .B1(net230383), .B2(n10364), 
        .ZN(n7491) );
  OAI22_X2 U8822 ( .A1(net231245), .A2(n11548), .B1(net230383), .B2(n10358), 
        .ZN(n7544) );
  OAI22_X2 U8824 ( .A1(net231245), .A2(n11115), .B1(net230383), .B2(net137343), 
        .ZN(n7726) );
  OAI22_X2 U8826 ( .A1(net231245), .A2(n12523), .B1(net230383), .B2(net137317), 
        .ZN(n7691) );
  OAI22_X2 U8830 ( .A1(net231245), .A2(n11114), .B1(net230383), .B2(net137303), 
        .ZN(n7674) );
  OAI22_X2 U8834 ( .A1(net231243), .A2(n12204), .B1(n10941), .B2(net230379), 
        .ZN(n7759) );
  AOI22_X2 U8837 ( .A1(net231301), .A2(MEM_WB_REG_MEM_WB_REG_N156), .B1(
        net230393), .B2(nextPC_ex_out[24]), .ZN(n6744) );
  OAI22_X2 U8838 ( .A1(net231243), .A2(n12203), .B1(net230383), .B2(n11102), 
        .ZN(n7851) );
  NAND2_X2 U8842 ( .A1(EXEC_STAGE_mul_result_long[63]), .A2(n13551), .ZN(n6746) );
  NAND2_X2 U8845 ( .A1(EXEC_STAGE_mul_result_long[62]), .A2(n13551), .ZN(n6748) );
  NAND2_X2 U8848 ( .A1(EXEC_STAGE_mul_result_long[61]), .A2(n13551), .ZN(n6749) );
  NAND2_X2 U8851 ( .A1(EXEC_STAGE_mul_result_long[60]), .A2(n13551), .ZN(n6750) );
  NAND2_X2 U8854 ( .A1(EXEC_STAGE_mul_result_long[59]), .A2(n13548), .ZN(n6751) );
  NAND2_X2 U8857 ( .A1(EXEC_STAGE_mul_result_long[58]), .A2(n13549), .ZN(n6752) );
  NAND2_X2 U8860 ( .A1(EXEC_STAGE_mul_result_long[57]), .A2(n13550), .ZN(n6753) );
  NAND2_X2 U8863 ( .A1(EXEC_STAGE_mul_result_long[56]), .A2(n13550), .ZN(n6754) );
  NAND2_X2 U8866 ( .A1(EXEC_STAGE_mul_result_long[55]), .A2(n13550), .ZN(n6756) );
  NAND2_X2 U8871 ( .A1(EXEC_STAGE_mul_result_long[54]), .A2(n13550), .ZN(n6757) );
  NAND2_X2 U8874 ( .A1(EXEC_STAGE_mul_result_long[53]), .A2(n13550), .ZN(n6759) );
  NAND2_X2 U8877 ( .A1(EXEC_STAGE_mul_result_long[52]), .A2(n13550), .ZN(n6760) );
  NAND2_X2 U8880 ( .A1(EXEC_STAGE_mul_result_long[51]), .A2(n13550), .ZN(n6761) );
  NAND2_X2 U8883 ( .A1(EXEC_STAGE_mul_result_long[50]), .A2(n13550), .ZN(n6762) );
  NAND2_X2 U8886 ( .A1(EXEC_STAGE_mul_result_long[49]), .A2(n13550), .ZN(n6763) );
  NAND2_X2 U8889 ( .A1(EXEC_STAGE_mul_result_long[48]), .A2(n13550), .ZN(n6764) );
  NAND2_X2 U8892 ( .A1(EXEC_STAGE_mul_result_long[47]), .A2(n13550), .ZN(n6765) );
  NAND2_X2 U8895 ( .A1(EXEC_STAGE_mul_result_long[46]), .A2(n13550), .ZN(n6766) );
  NAND2_X2 U8898 ( .A1(EXEC_STAGE_mul_result_long[45]), .A2(n13551), .ZN(n6768) );
  AOI22_X2 U8901 ( .A1(net231301), .A2(MEM_WB_REG_MEM_WB_REG_N158), .B1(
        net230387), .B2(nextPC_ex_out[22]), .ZN(n6769) );
  NAND2_X2 U8903 ( .A1(EXEC_STAGE_mul_result_long[44]), .A2(n13551), .ZN(n6770) );
  NAND2_X2 U8906 ( .A1(EXEC_STAGE_mul_result_long[43]), .A2(n13551), .ZN(n6771) );
  NAND2_X2 U8909 ( .A1(EXEC_STAGE_mul_result_long[42]), .A2(n13551), .ZN(n6772) );
  NAND2_X2 U8912 ( .A1(EXEC_STAGE_mul_result_long[41]), .A2(n13551), .ZN(n6773) );
  NAND2_X2 U8915 ( .A1(EXEC_STAGE_mul_result_long[40]), .A2(n13551), .ZN(n6774) );
  NAND2_X2 U8918 ( .A1(EXEC_STAGE_mul_result_long[39]), .A2(n13551), .ZN(n6775) );
  NAND2_X2 U8921 ( .A1(EXEC_STAGE_mul_result_long[38]), .A2(n13551), .ZN(n6776) );
  NAND2_X2 U8924 ( .A1(EXEC_STAGE_mul_result_long[37]), .A2(n13551), .ZN(n6777) );
  NAND2_X2 U8927 ( .A1(EXEC_STAGE_mul_result_long[36]), .A2(n13551), .ZN(n6778) );
  NAND2_X2 U8930 ( .A1(EXEC_STAGE_mul_result_long[35]), .A2(n13551), .ZN(n6779) );
  NAND2_X2 U8935 ( .A1(EXEC_STAGE_mul_result_long[34]), .A2(n13551), .ZN(n6780) );
  NAND2_X2 U8938 ( .A1(EXEC_STAGE_mul_result_long[33]), .A2(n13550), .ZN(n6781) );
  NAND2_X2 U8941 ( .A1(EXEC_STAGE_mul_result_long[32]), .A2(n13550), .ZN(n6782) );
  AOI22_X2 U8945 ( .A1(net231301), .A2(MEM_WB_REG_MEM_WB_REG_N35), .B1(n13550), 
        .B2(EXEC_STAGE_mul_result_long[31]), .ZN(n6783) );
  AOI22_X2 U8947 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N36), .B1(n13550), 
        .B2(EXEC_STAGE_mul_result_long[30]), .ZN(n6784) );
  AOI22_X2 U8949 ( .A1(net231301), .A2(MEM_WB_REG_MEM_WB_REG_N37), .B1(n13550), 
        .B2(EXEC_STAGE_mul_result_long[29]), .ZN(n6785) );
  AOI22_X2 U8951 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N38), .B1(n13550), 
        .B2(EXEC_STAGE_mul_result_long[28]), .ZN(n6786) );
  AOI22_X2 U8953 ( .A1(net231301), .A2(MEM_WB_REG_MEM_WB_REG_N39), .B1(n13550), 
        .B2(EXEC_STAGE_mul_result_long[27]), .ZN(n6787) );
  AOI22_X2 U8955 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N40), .B1(n13550), 
        .B2(EXEC_STAGE_mul_result_long[26]), .ZN(n6788) );
  AOI22_X2 U8957 ( .A1(net231301), .A2(MEM_WB_REG_MEM_WB_REG_N41), .B1(n13550), 
        .B2(EXEC_STAGE_mul_result_long[25]), .ZN(n6789) );
  AOI22_X2 U8959 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N160), .B1(
        net230393), .B2(nextPC_ex_out[20]), .ZN(n6790) );
  AOI22_X2 U8961 ( .A1(net231301), .A2(MEM_WB_REG_MEM_WB_REG_N42), .B1(n13550), 
        .B2(EXEC_STAGE_mul_result_long[24]), .ZN(n6791) );
  AOI22_X2 U8963 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N43), .B1(n13550), 
        .B2(EXEC_STAGE_mul_result_long[23]), .ZN(n6792) );
  AOI22_X2 U8965 ( .A1(net231301), .A2(MEM_WB_REG_MEM_WB_REG_N44), .B1(n13550), 
        .B2(EXEC_STAGE_mul_result_long[22]), .ZN(n6793) );
  AOI22_X2 U8967 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N45), .B1(n13549), 
        .B2(EXEC_STAGE_mul_result_long[21]), .ZN(n6794) );
  AOI22_X2 U8969 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N46), .B1(n13549), 
        .B2(EXEC_STAGE_mul_result_long[20]), .ZN(n6795) );
  AOI22_X2 U8971 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N47), .B1(n13549), 
        .B2(EXEC_STAGE_mul_result_long[19]), .ZN(n6796) );
  AOI22_X2 U8973 ( .A1(net231301), .A2(MEM_WB_REG_MEM_WB_REG_N48), .B1(n13549), 
        .B2(EXEC_STAGE_mul_result_long[18]), .ZN(n6797) );
  AOI22_X2 U8975 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N49), .B1(n13549), 
        .B2(EXEC_STAGE_mul_result_long[17]), .ZN(n6798) );
  AOI22_X2 U8977 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N50), .B1(n13549), 
        .B2(EXEC_STAGE_mul_result_long[16]), .ZN(n6799) );
  AOI22_X2 U8979 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N51), .B1(n13549), 
        .B2(EXEC_STAGE_mul_result_long[15]), .ZN(n6800) );
  OAI22_X2 U8980 ( .A1(net231243), .A2(n11547), .B1(net230383), .B2(n10362), 
        .ZN(n7539) );
  OAI22_X2 U8982 ( .A1(net231243), .A2(n11113), .B1(net230383), .B2(n10242), 
        .ZN(n7572) );
  AOI22_X2 U8985 ( .A1(net231301), .A2(MEM_WB_REG_MEM_WB_REG_N52), .B1(n13549), 
        .B2(EXEC_STAGE_mul_result_long[14]), .ZN(n6801) );
  AOI22_X2 U8987 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N53), .B1(n13549), 
        .B2(EXEC_STAGE_mul_result_long[13]), .ZN(n6802) );
  AOI22_X2 U8989 ( .A1(net231301), .A2(MEM_WB_REG_MEM_WB_REG_N54), .B1(n13549), 
        .B2(EXEC_STAGE_mul_result_long[12]), .ZN(n6803) );
  AOI22_X2 U8991 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N55), .B1(n13549), 
        .B2(EXEC_STAGE_mul_result_long[11]), .ZN(n6804) );
  AOI22_X2 U8993 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N56), .B1(n13548), 
        .B2(EXEC_STAGE_mul_result_long[10]), .ZN(n6805) );
  AOI22_X2 U8995 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N57), .B1(n13548), 
        .B2(EXEC_STAGE_mul_result_long[9]), .ZN(n6806) );
  AOI22_X2 U8997 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N58), .B1(n13548), 
        .B2(EXEC_STAGE_mul_result_long[8]), .ZN(n6807) );
  AOI22_X2 U8999 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N59), .B1(n13548), 
        .B2(EXEC_STAGE_mul_result_long[7]), .ZN(n6808) );
  AOI22_X2 U9001 ( .A1(net231301), .A2(MEM_WB_REG_MEM_WB_REG_N60), .B1(n13548), 
        .B2(EXEC_STAGE_mul_result_long[6]), .ZN(n6809) );
  AOI22_X2 U9003 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N61), .B1(n13548), 
        .B2(EXEC_STAGE_mul_result_long[5]), .ZN(n6810) );
  AOI22_X2 U9007 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N62), .B1(n13548), 
        .B2(EXEC_STAGE_mul_result_long[4]), .ZN(n6811) );
  AOI22_X2 U9009 ( .A1(net231305), .A2(MEM_WB_REG_MEM_WB_REG_N63), .B1(n13548), 
        .B2(EXEC_STAGE_mul_result_long[3]), .ZN(n6812) );
  AOI22_X2 U9011 ( .A1(net231303), .A2(MEM_WB_REG_MEM_WB_REG_N64), .B1(n13548), 
        .B2(EXEC_STAGE_mul_result_long[2]), .ZN(n6813) );
  AOI22_X2 U9013 ( .A1(net231305), .A2(MEM_WB_REG_MEM_WB_REG_N65), .B1(n13548), 
        .B2(EXEC_STAGE_mul_result_long[1]), .ZN(n6814) );
  AOI22_X2 U9015 ( .A1(net231301), .A2(MEM_WB_REG_MEM_WB_REG_N66), .B1(n13548), 
        .B2(EXEC_STAGE_mul_result_long[0]), .ZN(n6815) );
  OAI22_X2 U9017 ( .A1(net231241), .A2(n12202), .B1(net230383), .B2(n10939), 
        .ZN(n7917) );
  OAI22_X2 U9020 ( .A1(net231241), .A2(n12201), .B1(net230383), .B2(n10938), 
        .ZN(n7923) );
  OAI22_X2 U9023 ( .A1(net231239), .A2(n12200), .B1(net230383), .B2(n10937), 
        .ZN(n7929) );
  OAI22_X2 U9026 ( .A1(net231239), .A2(n12199), .B1(net230383), .B2(n10936), 
        .ZN(n7935) );
  OAI22_X2 U9029 ( .A1(net231239), .A2(n12198), .B1(net230383), .B2(n10935), 
        .ZN(n7943) );
  OAI22_X2 U9079 ( .A1(net231239), .A2(n11546), .B1(net230383), .B2(n11955), 
        .ZN(n7463) );
  OAI22_X2 U9153 ( .A1(n10157), .A2(net231251), .B1(n6889), .B2(net230379), 
        .ZN(n8018) );
  XOR2_X2 U9155 ( .A(n12212), .B(n6891), .Z(n6890) );
  OAI22_X2 U9215 ( .A1(net231237), .A2(n11545), .B1(net230383), .B2(n11921), 
        .ZN(n7430) );
  OAI22_X2 U9322 ( .A1(net231237), .A2(n11544), .B1(net230381), .B2(n11919), 
        .ZN(n7417) );
  OAI22_X2 U9488 ( .A1(net231237), .A2(n11471), .B1(net230383), .B2(n12052), 
        .ZN(n7845) );
  OAI22_X2 U9491 ( .A1(net231235), .A2(n10781), .B1(net230381), .B2(n11542), 
        .ZN(n7848) );
  OAI22_X2 U9494 ( .A1(net231235), .A2(n12522), .B1(net230383), .B2(n10933), 
        .ZN(n7904) );
  OAI22_X2 U9497 ( .A1(net231235), .A2(n12601), .B1(net230381), .B2(n19318), 
        .ZN(n7835) );
  OAI22_X2 U9502 ( .A1(net231235), .A2(n10860), .B1(net230383), .B2(n12051), 
        .ZN(n7871) );
  OAI22_X2 U9505 ( .A1(net231239), .A2(n11543), .B1(net230383), .B2(n12197), 
        .ZN(n7880) );
  NAND2_X2 U10055 ( .A1(n13218), .A2(n10236), .ZN(n7280) );
  XOR2_X2 U10056 ( .A(n11913), .B(n13218), .Z(n7279) );
  OAI22_X2 U10063 ( .A1(net231249), .A2(n11112), .B1(net230379), .B2(n10243), 
        .ZN(n7330) );
  OR2_X2 U10071 ( .A1(n13544), .A2(n13542), .ZN(EXEC_STAGE_mul_ex_N479) );
  AND2_X2 U10073 ( .A1(EXEC_STAGE_mul_ex_N185), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N476) );
  AND2_X2 U10074 ( .A1(EXEC_STAGE_mul_ex_N184), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N475) );
  AND2_X2 U10075 ( .A1(EXEC_STAGE_mul_ex_N183), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N474) );
  AND2_X2 U10076 ( .A1(EXEC_STAGE_mul_ex_N182), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N473) );
  AND2_X2 U10077 ( .A1(EXEC_STAGE_mul_ex_N181), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N472) );
  AND2_X2 U10078 ( .A1(EXEC_STAGE_mul_ex_N180), .A2(n19191), .ZN(
        EXEC_STAGE_mul_ex_N471) );
  AND2_X2 U10079 ( .A1(EXEC_STAGE_mul_ex_N179), .A2(n19191), .ZN(
        EXEC_STAGE_mul_ex_N470) );
  AND2_X2 U10080 ( .A1(EXEC_STAGE_mul_ex_N178), .A2(n19191), .ZN(
        EXEC_STAGE_mul_ex_N469) );
  AND2_X2 U10081 ( .A1(EXEC_STAGE_mul_ex_N177), .A2(n19191), .ZN(
        EXEC_STAGE_mul_ex_N468) );
  AND2_X2 U10082 ( .A1(EXEC_STAGE_mul_ex_N176), .A2(n19191), .ZN(
        EXEC_STAGE_mul_ex_N467) );
  AND2_X2 U10083 ( .A1(EXEC_STAGE_mul_ex_N175), .A2(n19191), .ZN(
        EXEC_STAGE_mul_ex_N466) );
  AND2_X2 U10084 ( .A1(EXEC_STAGE_mul_ex_N174), .A2(n19191), .ZN(
        EXEC_STAGE_mul_ex_N465) );
  AND2_X2 U10085 ( .A1(EXEC_STAGE_mul_ex_N173), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N464) );
  AND2_X2 U10086 ( .A1(EXEC_STAGE_mul_ex_N172), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N463) );
  AND2_X2 U10087 ( .A1(EXEC_STAGE_mul_ex_N171), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N462) );
  AND2_X2 U10088 ( .A1(EXEC_STAGE_mul_ex_N170), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N461) );
  AND2_X2 U10089 ( .A1(EXEC_STAGE_mul_ex_N169), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N460) );
  AND2_X2 U10090 ( .A1(EXEC_STAGE_mul_ex_N168), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N459) );
  AND2_X2 U10091 ( .A1(EXEC_STAGE_mul_ex_N167), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N458) );
  AND2_X2 U10092 ( .A1(EXEC_STAGE_mul_ex_N166), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N457) );
  AND2_X2 U10093 ( .A1(EXEC_STAGE_mul_ex_N165), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N456) );
  AND2_X2 U10094 ( .A1(EXEC_STAGE_mul_ex_N164), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N455) );
  AND2_X2 U10095 ( .A1(EXEC_STAGE_mul_ex_N163), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N454) );
  AND2_X2 U10096 ( .A1(EXEC_STAGE_mul_ex_N162), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N453) );
  AND2_X2 U10097 ( .A1(EXEC_STAGE_mul_ex_N161), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N452) );
  AND2_X2 U10098 ( .A1(EXEC_STAGE_mul_ex_N160), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N451) );
  AND2_X2 U10099 ( .A1(EXEC_STAGE_mul_ex_N159), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N450) );
  AND2_X2 U10100 ( .A1(EXEC_STAGE_mul_ex_N158), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N449) );
  AND2_X2 U10101 ( .A1(EXEC_STAGE_mul_ex_N157), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N448) );
  AND2_X2 U10102 ( .A1(EXEC_STAGE_mul_ex_N156), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N447) );
  AND2_X2 U10103 ( .A1(EXEC_STAGE_mul_ex_N155), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N446) );
  AND2_X2 U10104 ( .A1(EXEC_STAGE_mul_ex_N154), .A2(n13541), .ZN(
        EXEC_STAGE_mul_ex_N445) );
  NAND2_X2 U10105 ( .A1(n7283), .A2(n7284), .ZN(EXEC_STAGE_mul_ex_N444) );
  AND2_X2 U10106 ( .A1(EXEC_STAGE_mul_ex_N249), .A2(n19189), .ZN(
        EXEC_STAGE_mul_ex_N443) );
  AND2_X2 U10107 ( .A1(EXEC_STAGE_mul_ex_N248), .A2(n13537), .ZN(
        EXEC_STAGE_mul_ex_N442) );
  AND2_X2 U10108 ( .A1(EXEC_STAGE_mul_ex_N247), .A2(n13538), .ZN(
        EXEC_STAGE_mul_ex_N441) );
  AND2_X2 U10109 ( .A1(EXEC_STAGE_mul_ex_N246), .A2(n19189), .ZN(
        EXEC_STAGE_mul_ex_N440) );
  AND2_X2 U10110 ( .A1(EXEC_STAGE_mul_ex_N245), .A2(n13537), .ZN(
        EXEC_STAGE_mul_ex_N439) );
  AND2_X2 U10111 ( .A1(EXEC_STAGE_mul_ex_N244), .A2(n13538), .ZN(
        EXEC_STAGE_mul_ex_N438) );
  AND2_X2 U10112 ( .A1(EXEC_STAGE_mul_ex_N243), .A2(n19189), .ZN(
        EXEC_STAGE_mul_ex_N437) );
  AND2_X2 U10113 ( .A1(EXEC_STAGE_mul_ex_N242), .A2(n19189), .ZN(
        EXEC_STAGE_mul_ex_N436) );
  AND2_X2 U10114 ( .A1(EXEC_STAGE_mul_ex_N241), .A2(n13537), .ZN(
        EXEC_STAGE_mul_ex_N435) );
  AND2_X2 U10115 ( .A1(EXEC_STAGE_mul_ex_N240), .A2(n13538), .ZN(
        EXEC_STAGE_mul_ex_N434) );
  AND2_X2 U10116 ( .A1(EXEC_STAGE_mul_ex_N239), .A2(n13538), .ZN(
        EXEC_STAGE_mul_ex_N433) );
  AND2_X2 U10117 ( .A1(EXEC_STAGE_mul_ex_N238), .A2(n13538), .ZN(
        EXEC_STAGE_mul_ex_N432) );
  AND2_X2 U10118 ( .A1(EXEC_STAGE_mul_ex_N237), .A2(n13538), .ZN(
        EXEC_STAGE_mul_ex_N431) );
  AND2_X2 U10119 ( .A1(EXEC_STAGE_mul_ex_N236), .A2(n13538), .ZN(
        EXEC_STAGE_mul_ex_N430) );
  AND2_X2 U10121 ( .A1(EXEC_STAGE_mul_ex_N235), .A2(n13538), .ZN(
        EXEC_STAGE_mul_ex_N429) );
  AND2_X2 U10122 ( .A1(EXEC_STAGE_mul_ex_N234), .A2(n13538), .ZN(
        EXEC_STAGE_mul_ex_N428) );
  AND2_X2 U10123 ( .A1(EXEC_STAGE_mul_ex_N233), .A2(n13538), .ZN(
        EXEC_STAGE_mul_ex_N427) );
  AND2_X2 U10124 ( .A1(EXEC_STAGE_mul_ex_N232), .A2(n13538), .ZN(
        EXEC_STAGE_mul_ex_N426) );
  AND2_X2 U10125 ( .A1(EXEC_STAGE_mul_ex_N231), .A2(n13538), .ZN(
        EXEC_STAGE_mul_ex_N425) );
  AND2_X2 U10126 ( .A1(EXEC_STAGE_mul_ex_N230), .A2(n13538), .ZN(
        EXEC_STAGE_mul_ex_N424) );
  AND2_X2 U10127 ( .A1(EXEC_STAGE_mul_ex_N229), .A2(n13538), .ZN(
        EXEC_STAGE_mul_ex_N423) );
  AND2_X2 U10128 ( .A1(EXEC_STAGE_mul_ex_N228), .A2(n13537), .ZN(
        EXEC_STAGE_mul_ex_N422) );
  AND2_X2 U10129 ( .A1(EXEC_STAGE_mul_ex_N227), .A2(n13537), .ZN(
        EXEC_STAGE_mul_ex_N421) );
  AND2_X2 U10130 ( .A1(EXEC_STAGE_mul_ex_N226), .A2(n13537), .ZN(
        EXEC_STAGE_mul_ex_N420) );
  AND2_X2 U10131 ( .A1(EXEC_STAGE_mul_ex_N225), .A2(n13537), .ZN(
        EXEC_STAGE_mul_ex_N419) );
  AND2_X2 U10132 ( .A1(EXEC_STAGE_mul_ex_N224), .A2(n13537), .ZN(
        EXEC_STAGE_mul_ex_N418) );
  AND2_X2 U10133 ( .A1(EXEC_STAGE_mul_ex_N223), .A2(n13537), .ZN(
        EXEC_STAGE_mul_ex_N417) );
  AND2_X2 U10134 ( .A1(EXEC_STAGE_mul_ex_N222), .A2(n13537), .ZN(
        EXEC_STAGE_mul_ex_N416) );
  AND2_X2 U10135 ( .A1(EXEC_STAGE_mul_ex_N221), .A2(n13537), .ZN(
        EXEC_STAGE_mul_ex_N415) );
  AND2_X2 U10136 ( .A1(EXEC_STAGE_mul_ex_N220), .A2(n13537), .ZN(
        EXEC_STAGE_mul_ex_N414) );
  AND2_X2 U10137 ( .A1(EXEC_STAGE_mul_ex_N219), .A2(n13537), .ZN(
        EXEC_STAGE_mul_ex_N413) );
  AND2_X2 U10138 ( .A1(EXEC_STAGE_mul_ex_N218), .A2(n13537), .ZN(
        EXEC_STAGE_mul_ex_N412) );
  NAND2_X2 U10140 ( .A1(n7283), .A2(n7286), .ZN(EXEC_STAGE_mul_ex_N411) );
  AND2_X2 U10141 ( .A1(EXEC_STAGE_mul_ex_N119), .A2(n19190), .ZN(
        EXEC_STAGE_mul_ex_N410) );
  AND2_X2 U10142 ( .A1(EXEC_STAGE_mul_ex_N118), .A2(n13539), .ZN(
        EXEC_STAGE_mul_ex_N409) );
  AND2_X2 U10143 ( .A1(EXEC_STAGE_mul_ex_N117), .A2(n13540), .ZN(
        EXEC_STAGE_mul_ex_N408) );
  AND2_X2 U10144 ( .A1(EXEC_STAGE_mul_ex_N116), .A2(n19190), .ZN(
        EXEC_STAGE_mul_ex_N407) );
  AND2_X2 U10145 ( .A1(EXEC_STAGE_mul_ex_N115), .A2(n13539), .ZN(
        EXEC_STAGE_mul_ex_N406) );
  AND2_X2 U10146 ( .A1(EXEC_STAGE_mul_ex_N114), .A2(n13540), .ZN(
        EXEC_STAGE_mul_ex_N405) );
  AND2_X2 U10147 ( .A1(EXEC_STAGE_mul_ex_N113), .A2(n19190), .ZN(
        EXEC_STAGE_mul_ex_N404) );
  AND2_X2 U10148 ( .A1(EXEC_STAGE_mul_ex_N112), .A2(n19190), .ZN(
        EXEC_STAGE_mul_ex_N403) );
  AND2_X2 U10149 ( .A1(EXEC_STAGE_mul_ex_N111), .A2(n13539), .ZN(
        EXEC_STAGE_mul_ex_N402) );
  AND2_X2 U10150 ( .A1(EXEC_STAGE_mul_ex_N110), .A2(n13540), .ZN(
        EXEC_STAGE_mul_ex_N401) );
  AND2_X2 U10151 ( .A1(EXEC_STAGE_mul_ex_N109), .A2(n13540), .ZN(
        EXEC_STAGE_mul_ex_N400) );
  AND2_X2 U10152 ( .A1(EXEC_STAGE_mul_ex_N108), .A2(n13540), .ZN(
        EXEC_STAGE_mul_ex_N399) );
  AND2_X2 U10153 ( .A1(EXEC_STAGE_mul_ex_N107), .A2(n13540), .ZN(
        EXEC_STAGE_mul_ex_N398) );
  AND2_X2 U10154 ( .A1(EXEC_STAGE_mul_ex_N106), .A2(n13540), .ZN(
        EXEC_STAGE_mul_ex_N397) );
  AND2_X2 U10155 ( .A1(EXEC_STAGE_mul_ex_N105), .A2(n13540), .ZN(
        EXEC_STAGE_mul_ex_N396) );
  AND2_X2 U10156 ( .A1(EXEC_STAGE_mul_ex_N104), .A2(n13540), .ZN(
        EXEC_STAGE_mul_ex_N395) );
  AND2_X2 U10157 ( .A1(EXEC_STAGE_mul_ex_N103), .A2(n13540), .ZN(
        EXEC_STAGE_mul_ex_N394) );
  AND2_X2 U10158 ( .A1(EXEC_STAGE_mul_ex_N102), .A2(n13540), .ZN(
        EXEC_STAGE_mul_ex_N393) );
  AND2_X2 U10159 ( .A1(EXEC_STAGE_mul_ex_N101), .A2(n13540), .ZN(
        EXEC_STAGE_mul_ex_N392) );
  AND2_X2 U10160 ( .A1(EXEC_STAGE_mul_ex_N100), .A2(n13540), .ZN(
        EXEC_STAGE_mul_ex_N391) );
  AND2_X2 U10161 ( .A1(EXEC_STAGE_mul_ex_N99), .A2(n13540), .ZN(
        EXEC_STAGE_mul_ex_N390) );
  AND2_X2 U10162 ( .A1(EXEC_STAGE_mul_ex_N98), .A2(n13539), .ZN(
        EXEC_STAGE_mul_ex_N389) );
  AND2_X2 U10163 ( .A1(EXEC_STAGE_mul_ex_N97), .A2(n13539), .ZN(
        EXEC_STAGE_mul_ex_N388) );
  AND2_X2 U10164 ( .A1(EXEC_STAGE_mul_ex_N96), .A2(n13539), .ZN(
        EXEC_STAGE_mul_ex_N387) );
  AND2_X2 U10165 ( .A1(EXEC_STAGE_mul_ex_N95), .A2(n13539), .ZN(
        EXEC_STAGE_mul_ex_N386) );
  AND2_X2 U10166 ( .A1(EXEC_STAGE_mul_ex_N94), .A2(n13539), .ZN(
        EXEC_STAGE_mul_ex_N385) );
  AND2_X2 U10167 ( .A1(EXEC_STAGE_mul_ex_N93), .A2(n13539), .ZN(
        EXEC_STAGE_mul_ex_N384) );
  AND2_X2 U10168 ( .A1(EXEC_STAGE_mul_ex_N92), .A2(n13539), .ZN(
        EXEC_STAGE_mul_ex_N383) );
  AND2_X2 U10169 ( .A1(EXEC_STAGE_mul_ex_N91), .A2(n13539), .ZN(
        EXEC_STAGE_mul_ex_N382) );
  AND2_X2 U10170 ( .A1(EXEC_STAGE_mul_ex_N90), .A2(n13539), .ZN(
        EXEC_STAGE_mul_ex_N381) );
  AND2_X2 U10171 ( .A1(EXEC_STAGE_mul_ex_N89), .A2(n13539), .ZN(
        EXEC_STAGE_mul_ex_N380) );
  AND2_X2 U10172 ( .A1(EXEC_STAGE_mul_ex_N88), .A2(n13539), .ZN(
        EXEC_STAGE_mul_ex_N379) );
  NAND2_X2 U10174 ( .A1(n7283), .A2(n7288), .ZN(EXEC_STAGE_mul_ex_N378) );
  NAND2_X2 U10175 ( .A1(n7289), .A2(n10543), .ZN(n7283) );
  NAND2_X2 U10186 ( .A1(EXEC_STAGE_mul_ex_CurrentState_1_), .A2(n7289), .ZN(
        n7284) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_47_ ( .D(n7948), .CK(clk), .RN(n13924), 
        .Q(offset_26_id[9]), .QN(n12984) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_37_ ( .D(n7897), .CK(clk), .RN(n13888), 
        .Q(IF_ID_OUT[37]), .QN(n12020) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_159_ ( .D(n7840), .CK(clk), .RN(n13896), 
        .QN(n11041) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_3_ ( .D(n7492), .CK(clk), .RN(n13919), 
        .Q(nextPC_ex_out[3]), .QN(n10364) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_146_ ( .D(n7902), .CK(clk), .RN(n13897), 
        .Q(net239627), .QN(net233216) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_105_ ( .D(n7847), .CK(clk), .RN(n13887), .QN(n13124) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_193_ ( .D(n7970), .CK(clk), .RN(n13895), 
        .Q(ID_EXEC_OUT[193]), .QN(n13120) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_36_ ( .D(n7874), .CK(clk), .RN(n13929), 
        .Q(destReg_wb_out[4]), .QN(n13140) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_64_ ( .D(n7892), .CK(clk), .RN(
        n13911), .Q(MEM_WB_REG_MEM_WB_REG_N148), .QN(n13121) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_104_ ( .D(n7895), .CK(clk), .RN(
        n13892), .Q(MEM_WB_REG_MEM_WB_REG_N76), .QN(n13099) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_199_ ( .D(n7837), .CK(clk), .RN(n13894), 
        .Q(ID_EXEC_OUT[199]), .QN(n13145) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_67_ ( .D(n7883), .CK(clk), .RN(
        n13899), .Q(MEM_WB_REG_MEM_WB_REG_N145), .QN(n13132) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_192_ ( .D(n7899), .CK(clk), .RN(n13916), 
        .Q(ID_EXEC_OUT[192]), .QN(n13045) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_68_ ( .D(n7875), .CK(clk), .RN(
        n13911), .Q(MEM_WB_REG_MEM_WB_REG_N144), .QN(n13112) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_120_ ( .D(n7973), .CK(clk), .RN(n13906), 
        .Q(EXEC_STAGE_imm26_32[30]), .QN(net239083) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_102_ ( .D(n7870), .CK(clk), .RN(n13925), .Q(RegWrite_wb_out), .QN(n11916) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_101_ ( .D(n7879), .CK(clk), .RN(n13887), .Q(n12568), .QN(n13117) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_30_ ( .D(n7742), .CK(clk), .RN(n13919), 
        .QN(net233233) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_95_ ( .D(n7704), .CK(clk), .RN(
        n13912), .Q(DMEM_BUS_OUT[26]), .QN(n13134) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_198_ ( .D(n7839), .CK(clk), .RN(n13916), 
        .Q(ID_EXEC_OUT[198]), .QN(n13129) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_119_ ( .D(n19292), .CK(clk), .RN(n13905), 
        .Q(EXEC_STAGE_imm26_32[29]), .QN(n13075) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_106_ ( .D(n7844), .CK(clk), .RN(n13925), .QN(n13127) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_32_ ( .D(n7891), .CK(clk), .RN(n13929), 
        .Q(destReg_wb_out[0]), .QN(n13130) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_197_ ( .D(n7958), .CK(clk), .RN(n13895), 
        .Q(ID_EXEC_OUT[197]), .QN(n13135) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_103_ ( .D(n7871), .CK(clk), .RN(
        n13899), .Q(MEM_WB_REG_MEM_WB_REG_N77), .QN(n10860) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_104_ ( .D(n19278), .CK(clk), .RN(
        n13925), .Q(MEM_WB_OUT[104]), .QN(n13108) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_121_ ( .D(n19285), .CK(clk), .RN(n13913), 
        .Q(EXEC_STAGE_imm26_32[31]), .QN(net239370) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_34_ ( .D(n7885), .CK(clk), .RN(n13929), 
        .QN(n13105) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_29_ ( .D(n7727), .CK(clk), .RN(n13919), 
        .Q(nextPC_ex_out[29]), .QN(net239329) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_28_ ( .D(n7692), .CK(clk), .RN(n13892), 
        .Q(nextPC_ex_out[28]), .QN(net239555) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_27_ ( .D(n7683), .CK(clk), .RN(n13919), 
        .Q(nextPC_ex_out[27]), .QN(net239554) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_135_ ( .D(n19293), .CK(clk), .RN(n13897), 
        .Q(EXEC_STAGE_imm16_32[29]), .QN(n13077) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_103_ ( .D(n7894), .CK(clk), .RN(n13887), .Q(MEM_WB_OUT[103]), .QN(n13153) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_134_ ( .D(n7982), .CK(clk), .RN(n13913), 
        .Q(EXEC_STAGE_imm16_32[28]), .QN(n13062) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_196_ ( .D(n7961), .CK(clk), .RN(n13916), 
        .Q(ID_EXEC_OUT[196]), .QN(n13133) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_118_ ( .D(n7981), .CK(clk), .RN(n13913), 
        .Q(EXEC_STAGE_imm26_32[28]), .QN(n13042) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_65_ ( .D(n7889), .CK(clk), .RN(
        n13899), .Q(MEM_WB_REG_MEM_WB_REG_N147), .QN(n13137) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_200_ ( .D(n19280), .CK(clk), .RN(n13916), 
        .Q(ID_EXEC_OUT[200]), .QN(n13054) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_25_ ( .D(n7666), .CK(clk), .RN(n13889), 
        .Q(nextPC_ex_out[25]), .QN(net239756) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_136_ ( .D(n7974), .CK(clk), .RN(n13913), 
        .Q(EXEC_STAGE_imm16_32[30]), .QN(net239035) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_115_ ( .D(n7990), .CK(clk), .RN(n13885), 
        .Q(EXEC_STAGE_imm26_32[25]), .QN(net239806) );
  OAI22_X2 U8137 ( .A1(n11540), .A2(net231253), .B1(net230381), .B2(n11920), 
        .ZN(n7514) );
  OAI22_X2 U1822 ( .A1(net231239), .A2(n11920), .B1(net137185), .B2(net230373), 
        .ZN(n7515) );
  OAI22_X2 U4767 ( .A1(net231245), .A2(n11995), .B1(n12186), .B2(net230373), 
        .ZN(n7526) );
  AOI22_X2 U9033 ( .A1(net231315), .A2(MEM_WB_REG_MEM_WB_REG_N163), .B1(
        net230393), .B2(nextPC_ex_out[17]), .ZN(n6816) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_46_ ( .D(n7951), .CK(clk), .RN(n13888), 
        .Q(offset_26_id[8]), .QN(n12982) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_195_ ( .D(n7964), .CK(clk), .RN(n13895), 
        .Q(ID_EXEC_OUT[195]), .QN(n13122) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_33_ ( .D(n7888), .CK(clk), .RN(n13884), 
        .Q(n10351), .QN(n13059) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_42_ ( .D(n7959), .CK(clk), .RN(n13888), 
        .Q(offset_26_id[4]), .QN(n10368) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_41_ ( .D(n7962), .CK(clk), .RN(n13924), 
        .Q(offset_26_id[3]), .QN(n10844) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[17]), .QN(n12993) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_84_ ( .D(n7632), .CK(clk), .RN(
        n13912), .Q(DMEM_BUS_OUT[15]), .QN(n12130) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_40_ ( .D(n7965), .CK(clk), .RN(n13888), 
        .Q(offset_26_id[2]), .QN(n12026) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[13]), .QN(n12989) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[14]), .QN(n12988) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_93_ ( .D(n7698), .CK(clk), .RN(
        n13912), .Q(DMEM_BUS_OUT[24]) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_61_ ( .D(n7980), .CK(clk), .RN(n13925), 
        .Q(ID_STAGE_imm16_aluA[29]), .QN(n12039) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_39_ ( .D(n7968), .CK(clk), .RN(n13888), 
        .Q(offset_26_id[1]), .QN(n10828) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_98_ ( .D(n7731), .CK(clk), .RN(
        n13892), .Q(DMEM_BUS_OUT[29]), .QN(n12037) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_50_ ( .D(n7933), .CK(clk), .RN(n13924), 
        .Q(ID_STAGE_imm16_aluA[18]), .QN(n11045) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[19]), .QN(n12716) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_51_ ( .D(n7927), .CK(clk), .RN(n13888), 
        .Q(ID_STAGE_imm16_aluA[19]), .QN(n10806) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_49_ ( .D(n7939), .CK(clk), .RN(n13924), 
        .Q(ID_STAGE_imm16_aluA[17]), .QN(n10807) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[20]), .QN(n12567) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_125_ ( .D(n7925), .CK(clk), .RN(n13913), 
        .Q(EXEC_STAGE_imm16_32[19]), .QN(n12565) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_128_ ( .D(n7911), .CK(clk), .RN(n13888), 
        .Q(EXEC_STAGE_imm16_32[22]), .QN(n12564) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_130_ ( .D(n7994), .CK(clk), .RN(n13913), 
        .Q(EXEC_STAGE_imm16_32[24]), .QN(n12563) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_132_ ( .D(n7988), .CK(clk), .RN(n13913), 
        .Q(EXEC_STAGE_imm16_32[26]), .QN(n12562) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_126_ ( .D(n7919), .CK(clk), .RN(n13928), 
        .Q(EXEC_STAGE_imm16_32[20]), .QN(n12561) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[18]), .QN(n12560) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[6]), .QN(n12559) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_127_ ( .D(n19284), .CK(clk), .RN(n13913), 
        .Q(EXEC_STAGE_imm16_32[21]), .QN(n12557) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_129_ ( .D(n19283), .CK(clk), .RN(n13913), 
        .Q(EXEC_STAGE_imm16_32[23]), .QN(n12556) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[15]), .QN(n12554) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_31_ ( .D(n7832), .CK(clk), .RN(n13892), 
        .Q(nextPC_ex_out[31]), .QN(net239557) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[7]), .QN(n12544) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[16]), .QN(n12542) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[24]), .QN(n12319) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[8]), .QN(n12318) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[12]), .QN(n12317) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[9]), .QN(n12315) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[21]), .QN(n12314) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[23]), .QN(n12313) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( .D(n10105), 
        .CK(clk), .Q(IMEM_BUS_OUT[31]), .QN(n12312) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( .D(n10104), 
        .CK(clk), .Q(IMEM_BUS_OUT[30]), .QN(n12311) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_133_ ( .D(n19282), .CK(clk), .RN(n13897), 
        .Q(EXEC_STAGE_imm16_32[27]), .QN(n12258) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_194_ ( .D(n7967), .CK(clk), .RN(n13916), 
        .QN(n13138) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[22]), .QN(n12181) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_73_ ( .D(n8005), .CK(clk), .RN(n13882), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[20]), .QN(n12060) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_60_ ( .D(n7983), .CK(clk), .RN(n13887), 
        .Q(ID_STAGE_imm16_aluA[28]), .QN(n10840) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_52_ ( .D(n7921), .CK(clk), .RN(n13924), 
        .Q(ID_STAGE_imm16_aluA[20]), .QN(n12021) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_23_ ( .D(n7641), .CK(clk), .RN(n13918), 
        .Q(nextPC_ex_out[23]), .QN(n11985) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_53_ ( .D(n7915), .CK(clk), .RN(n13888), 
        .Q(ID_STAGE_imm16_aluA[21]), .QN(n11983) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_15_ ( .D(n7462), .CK(clk), .RN(n13928), 
        .Q(MEM_WB_OUT[15]), .QN(n11980) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_26_ ( .D(n7675), .CK(clk), .RN(n13892), 
        .Q(nextPC_ex_out[26]), .QN(n11962) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_24_ ( .D(n19279), .CK(clk), .RN(n13893), 
        .Q(nextPC_ex_out[24]), .QN(n11950) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_96_ ( .D(n7710), .CK(clk), .RN(
        n13886), .Q(DMEM_BUS_OUT[27]), .QN(n11949) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_97_ ( .D(n7696), .CK(clk), .RN(
        n13913), .Q(DMEM_BUS_OUT[28]), .QN(n11947) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_85_ ( .D(n7477), .CK(clk), .RN(
        n13898), .Q(DMEM_BUS_OUT[16]), .QN(n11938) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_20_ ( .D(n7582), .CK(clk), .RN(n13894), 
        .Q(nextPC_ex_out[20]), .QN(n11927) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_21_ ( .D(n7605), .CK(clk), .RN(n13917), 
        .Q(nextPC_ex_out[21]), .QN(n11918) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_18_ ( .D(n7565), .CK(clk), .RN(n13895), 
        .Q(nextPC_ex_out[18]), .QN(n11917) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_48_ ( .D(n7945), .CK(clk), .RN(n13888), 
        .Q(ID_STAGE_imm16_aluA[16]), .QN(n10816) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_109_ ( .D(n7926), .CK(clk), .RN(n13887), 
        .Q(EXEC_STAGE_imm26_32[19]), .QN(n11568) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_112_ ( .D(n7910), .CK(clk), .RN(n13887), 
        .Q(EXEC_STAGE_imm26_32[22]), .QN(n11567) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_114_ ( .D(n7993), .CK(clk), .RN(n13931), 
        .Q(EXEC_STAGE_imm26_32[24]), .QN(n11566) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_116_ ( .D(n7987), .CK(clk), .RN(n13924), 
        .Q(EXEC_STAGE_imm26_32[26]), .QN(n11565) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_110_ ( .D(n7920), .CK(clk), .RN(n13925), 
        .Q(EXEC_STAGE_imm26_32[20]), .QN(n11564) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_111_ ( .D(n19288), .CK(clk), .RN(n13913), 
        .Q(EXEC_STAGE_imm26_32[21]), .QN(n11559) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_113_ ( .D(n19287), .CK(clk), .RN(n13927), 
        .Q(EXEC_STAGE_imm26_32[23]), .QN(n11558) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_100_ ( .D(n8016), .CK(clk), .RN(n13925), .Q(MEM_WB_OUT[100]), .QN(n11555) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_81_ ( .D(n7867), .CK(clk), .RN(n13931), 
        .QN(n12069) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_82_ ( .D(n7866), .CK(clk), .RN(n13881), 
        .QN(n12070) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_80_ ( .D(n7868), .CK(clk), .RN(n13881), 
        .QN(n12068) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[11]), .QN(n11470) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_83_ ( .D(n7865), .CK(clk), .RN(n13931), 
        .QN(n12071) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_63_ ( .D(n7703), .CK(clk), .RN(n13931), 
        .Q(MEM_WB_OUT[63]), .QN(n11116) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[10]), .QN(n11097) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_76_ ( .D(n8008), .CK(clk), .RN(n13931), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[23]), .QN(n12032) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_75_ ( .D(n8007), .CK(clk), .RN(n13882), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[22]), .QN(n12031) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_117_ ( .D(n19286), .CK(clk), .RN(n13931), 
        .Q(EXEC_STAGE_imm26_32[27]), .QN(n11082) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_77_ ( .D(n8009), .CK(clk), .RN(n13882), 
        .QN(n12066) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_78_ ( .D(n8010), .CK(clk), .RN(n13931), 
        .QN(n12067) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_153_ ( .D(n8017), .CK(clk), .RN(n13897), 
        .Q(EXEC_MEM_IN_250), .QN(n10941) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_60_ ( .D(n7644), .CK(clk), .RN(n13882), 
        .Q(MEM_WB_OUT[60]), .QN(n10940) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_68_ ( .D(n19225), .CK(clk), .RN(n13882), .Q(MEM_WB_OUT[68]), .QN(n10910) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_22_ ( .D(n7622), .CK(clk), .RN(n13915), 
        .Q(nextPC_ex_out[22]), .QN(n10810) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_43_ ( .D(n7956), .CK(clk), .RN(n13924), 
        .Q(offset_26_id[5]), .QN(n10824) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_165_ ( .D(n7318), .CK(clk), .RN(n13928), .Q(MEM_WB_OUT[165]), .QN(n10239) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_164_ ( .D(n7305), .CK(clk), .RN(n13885), .Q(MEM_WB_OUT[164]), .QN(n10238) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_146_ ( .D(n7533), .CK(clk), .RN(n13886), .Q(MEM_WB_OUT[146]), .QN(n10237) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_176_ ( .D(n7760), .CK(clk), .RN(n13928), .Q(MEM_WB_OUT[176]), .QN(n10196) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_175_ ( .D(n7734), .CK(clk), .RN(n13884), .Q(MEM_WB_OUT[175]), .QN(n10195) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_174_ ( .D(n7719), .CK(clk), .RN(n13928), .Q(MEM_WB_OUT[174]), .QN(n10194) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_173_ ( .D(n7648), .CK(clk), .RN(n13885), .Q(MEM_WB_OUT[173]), .QN(n10193) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_172_ ( .D(n7707), .CK(clk), .RN(n13928), .Q(MEM_WB_OUT[172]), .QN(n10192) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_171_ ( .D(n7701), .CK(clk), .RN(n13885), .Q(MEM_WB_OUT[171]), .QN(n10191) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_170_ ( .D(n7713), .CK(clk), .RN(n13928), .Q(MEM_WB_OUT[170]), .QN(n10190) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_169_ ( .D(n7297), .CK(clk), .RN(n13928), .Q(MEM_WB_OUT[169]), .QN(n10189) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_168_ ( .D(n7301), .CK(clk), .RN(n13885), .Q(MEM_WB_OUT[168]), .QN(n10188) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_167_ ( .D(n7309), .CK(clk), .RN(n13928), .Q(MEM_WB_OUT[167]), .QN(n10187) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_166_ ( .D(n7313), .CK(clk), .RN(n13885), .Q(MEM_WB_OUT[166]), .QN(n10186) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_163_ ( .D(n7749), .CK(clk), .RN(n13928), .Q(MEM_WB_OUT[163]), .QN(n10185) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_162_ ( .D(n7339), .CK(clk), .RN(n13885), .Q(MEM_WB_OUT[162]), .QN(n10184) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_161_ ( .D(n7438), .CK(clk), .RN(n13928), .Q(MEM_WB_OUT[161]), .QN(n10183) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_160_ ( .D(n7629), .CK(clk), .RN(n13885), .Q(MEM_WB_OUT[160]), .QN(n10182) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_159_ ( .D(n7612), .CK(clk), .RN(n13885), .Q(MEM_WB_OUT[159]), .QN(n10181) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_158_ ( .D(n7595), .CK(clk), .RN(n13927), .Q(MEM_WB_OUT[158]), .QN(n10180) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_157_ ( .D(n7349), .CK(clk), .RN(n13885), .Q(MEM_WB_OUT[157]), .QN(n10179) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_156_ ( .D(n7396), .CK(clk), .RN(n13927), .Q(MEM_WB_OUT[156]), .QN(n10178) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_155_ ( .D(n7386), .CK(clk), .RN(n13885), .Q(MEM_WB_OUT[155]), .QN(n10177) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_154_ ( .D(n7344), .CK(clk), .RN(n13927), .Q(MEM_WB_OUT[154]), .QN(n10176) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_153_ ( .D(n7377), .CK(clk), .RN(n13885), .Q(MEM_WB_OUT[153]), .QN(n10175) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_152_ ( .D(n7406), .CK(clk), .RN(n13927), .Q(MEM_WB_OUT[152]), .QN(n10174) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_151_ ( .D(n7355), .CK(clk), .RN(n13886), .Q(MEM_WB_OUT[151]), .QN(n10173) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_150_ ( .D(n7361), .CK(clk), .RN(n13927), .Q(MEM_WB_OUT[150]), .QN(n10172) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_149_ ( .D(n7323), .CK(clk), .RN(n13927), .Q(MEM_WB_OUT[149]), .QN(n10171) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_148_ ( .D(n7589), .CK(clk), .RN(n13886), .Q(MEM_WB_OUT[148]), .QN(n10170) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_147_ ( .D(n7480), .CK(clk), .RN(n13927), .Q(MEM_WB_OUT[147]), .QN(n10169) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_145_ ( .D(n7753), .CK(clk), .RN(n13927), .Q(MEM_WB_OUT[145]), .QN(n10168) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_137_ ( .D(n19281), .CK(clk), .RN(n13897), 
        .Q(EXEC_STAGE_imm16_32[31]), .QN(n10110) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_131_ ( .D(n7991), .CK(clk), .RN(n13890), 
        .QN(net239744) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_201_ ( .D(n7950), .CK(clk), .RN(n13894), 
        .Q(ID_EXEC_OUT[201]), .QN(n13053) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_66_ ( .D(n7886), .CK(clk), .RN(
        n13911), .Q(MEM_WB_REG_MEM_WB_REG_N146), .QN(n13113) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_89_ ( .D(n7586), .CK(clk), .RN(
        n13898), .Q(DMEM_BUS_OUT[20]), .QN(n11963) );
  NAND2_X1 U10188 ( .A1(net227068), .A2(net225824), .ZN(n10117) );
  INV_X2 U10190 ( .A(net223742), .ZN(net227247) );
  NOR2_X1 U10191 ( .A1(n10144), .A2(net227186), .ZN(net227225) );
  OAI21_X2 U10192 ( .B1(net227226), .B2(net227247), .A(nextPC_ex_out[24]), 
        .ZN(net227246) );
  INV_X2 U10193 ( .A(net239475), .ZN(net227256) );
  NAND2_X1 U10194 ( .A1(n15530), .A2(net239782), .ZN(n10147) );
  NAND2_X2 U10195 ( .A1(n13111), .A2(net223743), .ZN(n17675) );
  INV_X4 U10196 ( .A(net227247), .ZN(n10107) );
  XNOR2_X2 U10197 ( .A(net233233), .B(net239035), .ZN(n15530) );
  OAI221_X2 U10198 ( .B1(n19350), .B2(net227188), .C1(net239737), .C2(
        net227191), .A(net227192), .ZN(n10108) );
  BUF_X32 U10199 ( .A(net227259), .Z(net239828) );
  INV_X2 U10200 ( .A(net225823), .ZN(net225892) );
  INV_X4 U10202 ( .A(n10110), .ZN(n10111) );
  NAND2_X4 U10203 ( .A1(n10146), .A2(n10147), .ZN(net222980) );
  NAND3_X4 U10204 ( .A1(net223797), .A2(n15544), .A3(n15545), .ZN(n10123) );
  BUF_X32 U10210 ( .A(net224955), .Z(net239674) );
  NAND3_X4 U10211 ( .A1(n15536), .A2(net227216), .A3(net227217), .ZN(n15544)
         );
  INV_X2 U10212 ( .A(net239782), .ZN(net239628) );
  NOR2_X1 U10213 ( .A1(n11995), .A2(net227117), .ZN(net227116) );
  XNOR2_X1 U10214 ( .A(nextPC_ex_out[24]), .B(net223743), .ZN(n18020) );
  XNOR2_X1 U10215 ( .A(nextPC_ex_out[22]), .B(net223985), .ZN(n17830) );
  INV_X4 U10216 ( .A(net233233), .ZN(net233156) );
  INV_X8 U10217 ( .A(n10139), .ZN(net227255) );
  BUF_X32 U10218 ( .A(net239473), .Z(n10116) );
  NAND2_X4 U10219 ( .A1(net239507), .A2(n10355), .ZN(n13029) );
  INV_X4 U10220 ( .A(net239572), .ZN(net227197) );
  AOI21_X2 U10221 ( .B1(n17207), .B2(n17206), .A(n17205), .ZN(n17208) );
  NAND2_X4 U10222 ( .A1(net224403), .A2(nextPC_ex_out[20]), .ZN(net239404) );
  INV_X8 U10223 ( .A(net233142), .ZN(net227262) );
  INV_X4 U10224 ( .A(net233078), .ZN(net227002) );
  BUF_X8 U10225 ( .A(net227081), .Z(net233102) );
  INV_X4 U10227 ( .A(net239597), .ZN(net225527) );
  NAND2_X4 U10228 ( .A1(net239678), .A2(net239718), .ZN(n16618) );
  NAND2_X2 U10229 ( .A1(n13386), .A2(n18862), .ZN(n17540) );
  INV_X32 U10230 ( .A(n13387), .ZN(n13386) );
  INV_X8 U10231 ( .A(n16007), .ZN(n18271) );
  OAI21_X2 U10232 ( .B1(n19354), .B2(n16007), .A(n16064), .ZN(n16877) );
  AOI222_X2 U10233 ( .A1(n17924), .A2(n17923), .B1(n18575), .B2(n18302), .C1(
        n18577), .C2(n18360), .ZN(n17925) );
  NAND2_X4 U10234 ( .A1(n10141), .A2(n10109), .ZN(net225448) );
  INV_X16 U10235 ( .A(net222300), .ZN(net232816) );
  AOI21_X2 U10236 ( .B1(n13492), .B2(n17507), .A(n17506), .ZN(n17555) );
  AOI21_X2 U10237 ( .B1(n13492), .B2(n17888), .A(n17887), .ZN(n17889) );
  NAND2_X4 U10238 ( .A1(n16782), .A2(n16781), .ZN(n18562) );
  NAND2_X2 U10240 ( .A1(n17044), .A2(n13492), .ZN(n17065) );
  NAND3_X4 U10241 ( .A1(n14057), .A2(n14056), .A3(n14055), .ZN(n15686) );
  NOR3_X2 U10242 ( .A1(n13976), .A2(n13975), .A3(n13974), .ZN(n13981) );
  INV_X8 U10243 ( .A(n14091), .ZN(n14098) );
  OAI21_X2 U10244 ( .B1(n17730), .B2(n17729), .A(n17728), .ZN(n17731) );
  OAI21_X2 U10245 ( .B1(n17883), .B2(n17733), .A(n17732), .ZN(n17735) );
  XNOR2_X2 U10246 ( .A(n13120), .B(n13121), .ZN(n13143) );
  INV_X8 U10247 ( .A(n13147), .ZN(n13219) );
  INV_X8 U10248 ( .A(n13153), .ZN(n13073) );
  NAND2_X1 U10249 ( .A1(net231615), .A2(n13151), .ZN(n18748) );
  NAND2_X1 U10250 ( .A1(n13409), .A2(n13151), .ZN(n18685) );
  NAND2_X1 U10251 ( .A1(n10363), .A2(n13151), .ZN(n18460) );
  NAND2_X1 U10252 ( .A1(n18644), .A2(n13151), .ZN(n18265) );
  NAND4_X1 U10253 ( .A1(n19126), .A2(n13151), .A3(ID_EXEC_OUT[156]), .A4(
        n19124), .ZN(n19127) );
  NAND3_X1 U10254 ( .A1(n19107), .A2(n13151), .A3(n19106), .ZN(n19121) );
  INV_X1 U10255 ( .A(n18281), .ZN(n18282) );
  XNOR2_X2 U10256 ( .A(n10125), .B(n16141), .ZN(n16143) );
  OAI21_X2 U10257 ( .B1(n15907), .B2(n15906), .A(n15905), .ZN(n10125) );
  INV_X4 U10259 ( .A(n17979), .ZN(n17836) );
  NOR2_X2 U10260 ( .A1(n14073), .A2(n14074), .ZN(n14076) );
  INV_X2 U10261 ( .A(n17493), .ZN(n15843) );
  OAI21_X2 U10262 ( .B1(n10121), .B2(n17706), .A(n17501), .ZN(n17504) );
  INV_X1 U10263 ( .A(n18930), .ZN(n10118) );
  OAI21_X2 U10264 ( .B1(n18304), .B2(n10120), .A(n10119), .ZN(n17710) );
  INV_X2 U10265 ( .A(n18304), .ZN(n18305) );
  NAND2_X4 U10266 ( .A1(n18304), .A2(n17834), .ZN(n17979) );
  NAND2_X4 U10267 ( .A1(n18396), .A2(n17499), .ZN(n17706) );
  NAND2_X4 U10268 ( .A1(n17896), .A2(n17894), .ZN(n18396) );
  XNOR2_X2 U10269 ( .A(n17838), .B(n12999), .ZN(n17839) );
  NAND2_X1 U10270 ( .A1(n17839), .A2(n13492), .ZN(n17865) );
  NAND2_X2 U10271 ( .A1(net224844), .A2(net239032), .ZN(n17032) );
  AOI21_X4 U10272 ( .B1(n15934), .B2(n15935), .A(n15933), .ZN(n19150) );
  BUF_X32 U10273 ( .A(n17708), .Z(n10119) );
  NAND2_X4 U10274 ( .A1(n13097), .A2(n13096), .ZN(n18684) );
  INV_X1 U10275 ( .A(n19358), .ZN(n10120) );
  INV_X8 U10276 ( .A(n17709), .ZN(n15775) );
  INV_X8 U10278 ( .A(n15777), .ZN(n17708) );
  BUF_X32 U10279 ( .A(n15668), .Z(n10122) );
  INV_X1 U10280 ( .A(ID_EXEC_OUT[198]), .ZN(n18753) );
  NAND2_X1 U10281 ( .A1(net231325), .A2(ID_EXEC_OUT[199]), .ZN(n18751) );
  NAND2_X2 U10282 ( .A1(n16396), .A2(n16395), .ZN(n16536) );
  INV_X1 U10283 ( .A(MEM_WB_REG_MEM_WB_REG_N144), .ZN(n19319) );
  INV_X2 U10284 ( .A(n18588), .ZN(n18620) );
  CLKBUF_X2 U10285 ( .A(net227079), .Z(net239678) );
  INV_X4 U10286 ( .A(net227274), .ZN(n10124) );
  INV_X8 U10287 ( .A(net227274), .ZN(net227261) );
  NAND2_X4 U10288 ( .A1(DMEM_BUS_OUT[23]), .A2(n13484), .ZN(n15763) );
  NAND2_X1 U10289 ( .A1(n17142), .A2(n18890), .ZN(n17143) );
  NAND2_X2 U10291 ( .A1(net239454), .A2(n13080), .ZN(n13082) );
  INV_X32 U10292 ( .A(n13404), .ZN(n13403) );
  INV_X16 U10293 ( .A(n18625), .ZN(n13404) );
  INV_X8 U10294 ( .A(n13073), .ZN(n10126) );
  INV_X1 U10295 ( .A(n18383), .ZN(n10127) );
  INV_X4 U10296 ( .A(n10127), .ZN(n10128) );
  AOI21_X2 U10298 ( .B1(n15561), .B2(n15560), .A(n15559), .ZN(n15581) );
  INV_X16 U10300 ( .A(n13997), .ZN(n15712) );
  NAND3_X2 U10301 ( .A1(n15816), .A2(n15817), .A3(n15818), .ZN(n10129) );
  NAND3_X4 U10303 ( .A1(n15685), .A2(n15684), .A3(n15683), .ZN(n10130) );
  NAND3_X2 U10304 ( .A1(n15685), .A2(n15684), .A3(n15683), .ZN(n18960) );
  NAND2_X2 U10305 ( .A1(ID_EXEC_OUT[91]), .A2(n18625), .ZN(n15685) );
  NAND2_X1 U10306 ( .A1(n13409), .A2(n13163), .ZN(n18019) );
  NAND2_X1 U10307 ( .A1(net231615), .A2(n13163), .ZN(n18241) );
  INV_X2 U10308 ( .A(n13163), .ZN(n18365) );
  AOI22_X1 U10309 ( .A1(n18533), .A2(n16207), .B1(n10843), .B2(n13163), .ZN(
        n18545) );
  NOR2_X2 U10310 ( .A1(n18962), .A2(n18960), .ZN(n13109) );
  NAND2_X2 U10311 ( .A1(n18860), .A2(n10130), .ZN(net222304) );
  INV_X4 U10312 ( .A(n10130), .ZN(n18373) );
  NAND2_X2 U10313 ( .A1(n16879), .A2(n10130), .ZN(n16795) );
  NAND2_X4 U10314 ( .A1(n13068), .A2(n13067), .ZN(n18953) );
  INV_X4 U10316 ( .A(net225198), .ZN(net224837) );
  INV_X2 U10317 ( .A(net225214), .ZN(n10132) );
  INV_X8 U10318 ( .A(net227229), .ZN(n10154) );
  INV_X1 U10319 ( .A(n18961), .ZN(n10133) );
  INV_X8 U10320 ( .A(net227221), .ZN(n13006) );
  INV_X1 U10321 ( .A(n19360), .ZN(n18886) );
  INV_X1 U10322 ( .A(n17137), .ZN(n17138) );
  NAND2_X4 U10325 ( .A1(n16959), .A2(net225198), .ZN(net225196) );
  NAND3_X2 U10326 ( .A1(n17226), .A2(n17227), .A3(n17228), .ZN(n7547) );
  NOR2_X2 U10327 ( .A1(n17225), .A2(n17224), .ZN(n17226) );
  OAI21_X4 U10329 ( .B1(n15578), .B2(n15577), .A(n15576), .ZN(n15579) );
  BUF_X32 U10330 ( .A(net227282), .Z(n10135) );
  BUF_X32 U10332 ( .A(net223442), .Z(n10137) );
  INV_X4 U10333 ( .A(n10158), .ZN(net232881) );
  INV_X2 U10334 ( .A(net232881), .ZN(net227290) );
  AND3_X4 U10335 ( .A1(net227015), .A2(net227009), .A3(net225077), .ZN(n10138)
         );
  BUF_X32 U10336 ( .A(net225780), .Z(net239508) );
  NAND3_X2 U10337 ( .A1(ID_EXEC_OUT[94]), .A2(n13092), .A3(n13098), .ZN(n15703) );
  NAND2_X2 U10338 ( .A1(net227282), .A2(net239805), .ZN(n13018) );
  NAND2_X4 U10339 ( .A1(net233142), .A2(nextPC_ex_out[26]), .ZN(n15533) );
  NAND2_X2 U10340 ( .A1(n18945), .A2(n13163), .ZN(n18950) );
  AOI21_X4 U10341 ( .B1(n18920), .B2(n13061), .A(n18919), .ZN(n19010) );
  NAND4_X2 U10342 ( .A1(net227163), .A2(net227164), .A3(n13035), .A4(n13034), 
        .ZN(n13036) );
  NAND2_X4 U10343 ( .A1(net227199), .A2(net239533), .ZN(n10139) );
  NAND2_X2 U10344 ( .A1(net239533), .A2(net227199), .ZN(net227191) );
  OAI22_X4 U10345 ( .A1(net227180), .A2(net239496), .B1(n13033), .B2(net227148), .ZN(net239082) );
  OAI21_X2 U10346 ( .B1(net227188), .B2(n15534), .A(net227224), .ZN(n15535) );
  INV_X2 U10347 ( .A(n10145), .ZN(n10140) );
  INV_X2 U10348 ( .A(n19136), .ZN(n19132) );
  NAND2_X1 U10349 ( .A1(n18945), .A2(n10130), .ZN(net222300) );
  XNOR2_X1 U10350 ( .A(n10130), .B(n13494), .ZN(n15844) );
  BUF_X32 U10353 ( .A(net227139), .Z(n10142) );
  AND2_X2 U10354 ( .A1(n10140), .A2(net232881), .ZN(n10369) );
  AND2_X2 U10355 ( .A1(net239782), .A2(EXEC_STAGE_imm16_32[16]), .ZN(n10158)
         );
  INV_X1 U10356 ( .A(net239782), .ZN(n10145) );
  BUF_X32 U10357 ( .A(n18445), .Z(n10143) );
  NAND2_X4 U10358 ( .A1(net227282), .A2(net239805), .ZN(net239390) );
  INV_X4 U10359 ( .A(n10144), .ZN(net239761) );
  INV_X4 U10360 ( .A(net223663), .ZN(net233141) );
  NAND2_X4 U10361 ( .A1(net239767), .A2(n10153), .ZN(n13020) );
  INV_X2 U10362 ( .A(net223589), .ZN(n10144) );
  INV_X4 U10363 ( .A(net223589), .ZN(net227226) );
  INV_X4 U10364 ( .A(net233156), .ZN(net222982) );
  NAND2_X1 U10365 ( .A1(n10145), .A2(n15531), .ZN(n10146) );
  INV_X4 U10366 ( .A(net227142), .ZN(net227139) );
  NOR2_X4 U10367 ( .A1(net239527), .A2(net227241), .ZN(net227248) );
  INV_X8 U10368 ( .A(n13004), .ZN(net239477) );
  INV_X4 U10369 ( .A(n13004), .ZN(n13005) );
  NAND2_X2 U10370 ( .A1(net227277), .A2(net227276), .ZN(n18445) );
  INV_X4 U10371 ( .A(net233141), .ZN(n10148) );
  BUF_X32 U10372 ( .A(net225908), .Z(net239598) );
  INV_X4 U10373 ( .A(net233156), .ZN(n10149) );
  INV_X4 U10374 ( .A(net223666), .ZN(n10150) );
  INV_X8 U10375 ( .A(n10150), .ZN(n10151) );
  NAND3_X2 U10376 ( .A1(net227088), .A2(net227089), .A3(net227087), .ZN(
        net239414) );
  NAND2_X1 U10377 ( .A1(net227225), .A2(net223666), .ZN(n15534) );
  NAND2_X2 U10378 ( .A1(n13030), .A2(n13029), .ZN(net225201) );
  NAND2_X4 U10379 ( .A1(n15651), .A2(n12745), .ZN(n13116) );
  NAND2_X1 U10380 ( .A1(net225214), .A2(n10152), .ZN(n13030) );
  AND2_X2 U10381 ( .A1(net225209), .A2(nextPC_ex_out[5]), .ZN(n10152) );
  NAND3_X4 U10382 ( .A1(net227070), .A2(net227069), .A3(n11921), .ZN(net227068) );
  INV_X4 U10383 ( .A(net239744), .ZN(n10153) );
  NAND2_X4 U10384 ( .A1(net227121), .A2(n15551), .ZN(n15552) );
  NAND2_X2 U10385 ( .A1(n15551), .A2(net227121), .ZN(net227106) );
  NAND2_X4 U10386 ( .A1(net225075), .A2(net225076), .ZN(net224844) );
  INV_X8 U10387 ( .A(net239254), .ZN(net227188) );
  AND2_X2 U10388 ( .A1(n10143), .A2(nextPC_ex_out[29]), .ZN(n10155) );
  NAND2_X1 U10389 ( .A1(net227149), .A2(net227150), .ZN(n13032) );
  BUF_X32 U10390 ( .A(net224182), .Z(n10156) );
  NAND3_X2 U10391 ( .A1(net224491), .A2(net239404), .A3(n10242), .ZN(net224661) );
  NAND3_X4 U10392 ( .A1(n15555), .A2(n17197), .A3(net224816), .ZN(n15651) );
  NAND2_X2 U10393 ( .A1(n10138), .A2(n15566), .ZN(n15641) );
  NAND2_X2 U10394 ( .A1(n15642), .A2(n15641), .ZN(n15555) );
  NAND2_X4 U10395 ( .A1(net233242), .A2(n13076), .ZN(net227276) );
  INV_X16 U10396 ( .A(net233242), .ZN(net239767) );
  NAND3_X4 U10397 ( .A1(n10151), .A2(net239254), .A3(net239761), .ZN(net227207) );
  CLKBUF_X3 U10398 ( .A(net227220), .Z(net239825) );
  NAND3_X4 U10399 ( .A1(net225452), .A2(net225453), .A3(nextPC_ex_out[16]), 
        .ZN(net227098) );
  NAND2_X4 U10400 ( .A1(net227008), .A2(net227002), .ZN(n15648) );
  INV_X4 U10401 ( .A(net227014), .ZN(net227052) );
  INV_X4 U10402 ( .A(net233181), .ZN(net239737) );
  NAND2_X4 U10403 ( .A1(n15544), .A2(n15545), .ZN(net227175) );
  NOR2_X2 U10404 ( .A1(net227058), .A2(n12205), .ZN(net239379) );
  INV_X4 U10405 ( .A(net227062), .ZN(net227058) );
  INV_X8 U10406 ( .A(net224708), .ZN(net233106) );
  AOI221_X4 U10407 ( .B1(net233242), .B2(net239083), .C1(net239767), .C2(
        net239221), .A(net222982), .ZN(net239220) );
  NAND3_X4 U10408 ( .A1(n10154), .A2(n10123), .A3(net223985), .ZN(net224174)
         );
  OAI211_X4 U10409 ( .C1(net239380), .C2(net227013), .A(n13026), .B(n11016), 
        .ZN(net224842) );
  INV_X4 U10410 ( .A(n14193), .ZN(n14998) );
  NAND3_X2 U10411 ( .A1(n12026), .A2(n10844), .A3(n10368), .ZN(n14193) );
  INV_X8 U10412 ( .A(n18540), .ZN(n13398) );
  INV_X8 U10414 ( .A(n18340), .ZN(n13391) );
  INV_X16 U10415 ( .A(n13398), .ZN(n13397) );
  NOR2_X2 U10416 ( .A1(n7280), .A2(n11913), .ZN(n15674) );
  NOR2_X2 U10417 ( .A1(n7279), .A2(n10236), .ZN(n15675) );
  INV_X4 U10418 ( .A(n16059), .ZN(n13395) );
  NAND2_X1 U10419 ( .A1(n18756), .A2(ID_STAGE_imm16_aluA[29]), .ZN(n14241) );
  INV_X4 U10420 ( .A(n13437), .ZN(n13434) );
  NAND3_X2 U10421 ( .A1(n12953), .A2(n12982), .A3(n12984), .ZN(n14192) );
  NOR2_X2 U10422 ( .A1(net227071), .A2(n12018), .ZN(net227067) );
  NOR2_X2 U10423 ( .A1(n12018), .A2(n11921), .ZN(net227072) );
  INV_X4 U10424 ( .A(n15336), .ZN(n13283) );
  NAND2_X1 U10425 ( .A1(n2511), .A2(n14998), .ZN(n15336) );
  NAND2_X1 U10426 ( .A1(n14995), .A2(n2511), .ZN(n2184) );
  NAND2_X2 U10427 ( .A1(n18664), .A2(n17868), .ZN(n14151) );
  INV_X4 U10428 ( .A(n13737), .ZN(n13736) );
  INV_X4 U10429 ( .A(n13728), .ZN(n13726) );
  INV_X4 U10430 ( .A(n13731), .ZN(n13729) );
  INV_X4 U10431 ( .A(n18714), .ZN(n13196) );
  NAND2_X2 U10432 ( .A1(n15608), .A2(n15617), .ZN(n18714) );
  NAND2_X2 U10433 ( .A1(n15621), .A2(n15617), .ZN(n18712) );
  NAND2_X1 U10434 ( .A1(n15616), .A2(n15613), .ZN(n18730) );
  INV_X4 U10435 ( .A(n10834), .ZN(n13475) );
  NAND2_X2 U10436 ( .A1(n14288), .A2(n14998), .ZN(n13171) );
  NOR2_X1 U10437 ( .A1(n13218), .A2(ID_EXEC_OUT[157]), .ZN(n15710) );
  NOR2_X1 U10438 ( .A1(n14011), .A2(net222304), .ZN(n15695) );
  NOR2_X2 U10439 ( .A1(n15739), .A2(n16060), .ZN(n15744) );
  NAND2_X2 U10440 ( .A1(n14288), .A2(n14998), .ZN(n13170) );
  INV_X4 U10441 ( .A(n17773), .ZN(n13375) );
  INV_X4 U10442 ( .A(n17772), .ZN(n13372) );
  INV_X4 U10443 ( .A(n17774), .ZN(n13378) );
  INV_X16 U10444 ( .A(n10782), .ZN(n13184) );
  INV_X4 U10445 ( .A(n10805), .ZN(n13458) );
  NOR3_X2 U10446 ( .A1(n19095), .A2(n19094), .A3(n19093), .ZN(n19102) );
  NAND3_X1 U10447 ( .A1(ID_STAGE_imm16_aluA[26]), .A2(n10838), .A3(n13167), 
        .ZN(n14218) );
  NAND3_X2 U10448 ( .A1(nextPC_ex_out[0]), .A2(net224704), .A3(
        nextPC_ex_out[1]), .ZN(n15568) );
  INV_X4 U10449 ( .A(n13283), .ZN(n13282) );
  INV_X4 U10450 ( .A(n13274), .ZN(n13273) );
  NAND3_X2 U10451 ( .A1(n16312), .A2(n16795), .A3(n16311), .ZN(n17747) );
  INV_X4 U10452 ( .A(n13283), .ZN(n13281) );
  NOR2_X2 U10453 ( .A1(net224847), .A2(net224848), .ZN(net224839) );
  INV_X4 U10454 ( .A(n13274), .ZN(n13272) );
  INV_X4 U10455 ( .A(n13271), .ZN(n13269) );
  INV_X4 U10456 ( .A(n13731), .ZN(n13730) );
  INV_X4 U10457 ( .A(net225185), .ZN(net224704) );
  NAND3_X2 U10458 ( .A1(n16029), .A2(n16028), .A3(n16027), .ZN(n16030) );
  NAND3_X2 U10459 ( .A1(n14033), .A2(n14032), .A3(n14031), .ZN(n17382) );
  NAND3_X2 U10460 ( .A1(n14003), .A2(n14002), .A3(n14001), .ZN(n17546) );
  NAND3_X1 U10461 ( .A1(n16302), .A2(n16795), .A3(n16301), .ZN(n17585) );
  INV_X4 U10462 ( .A(n13369), .ZN(n13368) );
  INV_X4 U10463 ( .A(n13208), .ZN(n13209) );
  INV_X4 U10464 ( .A(n18569), .ZN(n17982) );
  INV_X4 U10465 ( .A(n17870), .ZN(n18566) );
  INV_X4 U10466 ( .A(n13366), .ZN(n13365) );
  NAND3_X2 U10467 ( .A1(n14028), .A2(n14027), .A3(n14026), .ZN(n17331) );
  NAND3_X1 U10468 ( .A1(n16391), .A2(n16795), .A3(n16390), .ZN(n17586) );
  INV_X8 U10469 ( .A(n10559), .ZN(n13207) );
  NAND3_X2 U10470 ( .A1(n16525), .A2(n16795), .A3(n16524), .ZN(n17910) );
  NAND2_X2 U10471 ( .A1(n13208), .A2(n13406), .ZN(n18569) );
  INV_X4 U10472 ( .A(n13369), .ZN(n13367) );
  INV_X4 U10473 ( .A(net231353), .ZN(net231331) );
  INV_X8 U10474 ( .A(n13166), .ZN(n13167) );
  INV_X4 U10475 ( .A(net231359), .ZN(net231355) );
  NAND3_X2 U10476 ( .A1(n14260), .A2(n14259), .A3(n14258), .ZN(n18760) );
  NOR2_X2 U10477 ( .A1(n15558), .A2(n15644), .ZN(n15559) );
  INV_X16 U10479 ( .A(n10349), .ZN(n13182) );
  INV_X8 U10480 ( .A(n13737), .ZN(n13735) );
  NAND3_X2 U10481 ( .A1(n17303), .A2(n17302), .A3(n17301), .ZN(n17575) );
  INV_X4 U10482 ( .A(n18451), .ZN(n13212) );
  INV_X4 U10483 ( .A(n18550), .ZN(n13492) );
  INV_X4 U10484 ( .A(n13490), .ZN(n13491) );
  NAND3_X2 U10485 ( .A1(n18669), .A2(n10236), .A3(n15931), .ZN(n18550) );
  NOR2_X2 U10486 ( .A1(ID_EXEC_OUT[157]), .A2(ID_EXEC_OUT[158]), .ZN(n15931)
         );
  NAND2_X2 U10487 ( .A1(n18664), .A2(n17981), .ZN(n14071) );
  INV_X4 U10488 ( .A(n19104), .ZN(n18651) );
  INV_X16 U10489 ( .A(n13162), .ZN(n13163) );
  INV_X4 U10490 ( .A(n13478), .ZN(n13483) );
  INV_X4 U10491 ( .A(n18456), .ZN(n13208) );
  NAND2_X2 U10492 ( .A1(n18669), .A2(n15714), .ZN(n18456) );
  INV_X4 U10493 ( .A(n19110), .ZN(n13490) );
  INV_X8 U10494 ( .A(n13210), .ZN(n13211) );
  INV_X8 U10496 ( .A(n19125), .ZN(n13150) );
  INV_X4 U10497 ( .A(net231277), .ZN(net231243) );
  OAI21_X1 U10498 ( .B1(n18781), .B2(n14220), .A(n14212), .ZN(n14213) );
  INV_X2 U10499 ( .A(n13109), .ZN(n13110) );
  OAI21_X1 U10500 ( .B1(n18925), .B2(n18924), .A(n18975), .ZN(n18974) );
  NAND3_X2 U10501 ( .A1(n18595), .A2(n18606), .A3(n18594), .ZN(n18604) );
  INV_X4 U10502 ( .A(n13437), .ZN(n13436) );
  AOI22_X2 U10503 ( .A1(MEM_WB_OUT[16]), .A2(n13877), .B1(MEM_WB_OUT[85]), 
        .B2(n14102), .ZN(n14108) );
  INV_X16 U10504 ( .A(n13437), .ZN(n13435) );
  NOR2_X1 U10505 ( .A1(n11985), .A2(n10810), .ZN(net227224) );
  NOR3_X2 U10506 ( .A1(n2539), .A2(n2538), .A3(n12053), .ZN(n14978) );
  NOR2_X2 U10507 ( .A1(n14103), .A2(n12067), .ZN(n14038) );
  NAND2_X2 U10508 ( .A1(n13087), .A2(n13088), .ZN(n15502) );
  NAND2_X2 U10509 ( .A1(n13085), .A2(n13086), .ZN(n13088) );
  INV_X4 U10510 ( .A(n13425), .ZN(n13428) );
  NOR2_X2 U10511 ( .A1(n19089), .A2(n18878), .ZN(n19037) );
  NOR2_X2 U10512 ( .A1(n12113), .A2(n13169), .ZN(n14523) );
  NOR2_X2 U10513 ( .A1(n12112), .A2(n13169), .ZN(n14512) );
  NAND3_X2 U10514 ( .A1(net227026), .A2(net224846), .A3(net224845), .ZN(
        net227062) );
  INV_X4 U10515 ( .A(n10827), .ZN(n13421) );
  NAND3_X2 U10517 ( .A1(net224954), .A2(net224955), .A3(net227104), .ZN(
        net227103) );
  NOR2_X2 U10518 ( .A1(n16732), .A2(n16731), .ZN(n16733) );
  NOR2_X2 U10519 ( .A1(n13432), .A2(n12440), .ZN(n16732) );
  NOR2_X2 U10520 ( .A1(n13427), .A2(n12441), .ZN(n16731) );
  NOR2_X2 U10521 ( .A1(n16730), .A2(n16729), .ZN(n16735) );
  NOR2_X2 U10522 ( .A1(n13422), .A2(n12439), .ZN(n16730) );
  NOR2_X2 U10523 ( .A1(n13423), .A2(n12869), .ZN(n16729) );
  NOR2_X2 U10524 ( .A1(n17073), .A2(n17072), .ZN(n17074) );
  NOR2_X2 U10525 ( .A1(n13432), .A2(n12452), .ZN(n17073) );
  NOR2_X2 U10526 ( .A1(n13427), .A2(n12453), .ZN(n17072) );
  NOR2_X2 U10527 ( .A1(n17071), .A2(n17070), .ZN(n17076) );
  NOR2_X2 U10528 ( .A1(n13422), .A2(n12451), .ZN(n17071) );
  NOR2_X2 U10529 ( .A1(n13423), .A2(n12883), .ZN(n17070) );
  INV_X8 U10530 ( .A(n13433), .ZN(n13431) );
  INV_X8 U10531 ( .A(n13433), .ZN(n13432) );
  NOR2_X2 U10532 ( .A1(n17341), .A2(n17340), .ZN(n17346) );
  NOR2_X2 U10533 ( .A1(n13422), .A2(n12459), .ZN(n17341) );
  NOR2_X2 U10534 ( .A1(n13423), .A2(n12893), .ZN(n17340) );
  NOR2_X2 U10535 ( .A1(n17343), .A2(n17342), .ZN(n17344) );
  NOR2_X1 U10536 ( .A1(n13426), .A2(n12461), .ZN(n17342) );
  NOR2_X2 U10537 ( .A1(n13431), .A2(n12460), .ZN(n17343) );
  NOR2_X2 U10538 ( .A1(n17392), .A2(n17391), .ZN(n17397) );
  NOR2_X2 U10539 ( .A1(n13421), .A2(n12462), .ZN(n17392) );
  NOR2_X2 U10540 ( .A1(n13423), .A2(n12895), .ZN(n17391) );
  NOR2_X2 U10541 ( .A1(n17394), .A2(n17393), .ZN(n17395) );
  NOR2_X1 U10542 ( .A1(n13426), .A2(n12464), .ZN(n17393) );
  NOR2_X2 U10543 ( .A1(n13431), .A2(n12463), .ZN(n17394) );
  AOI21_X2 U10544 ( .B1(n13196), .B2(REG_FILE_reg_out_22__20_), .A(n17471), 
        .ZN(n17472) );
  NOR2_X2 U10545 ( .A1(n17470), .A2(n13452), .ZN(n17471) );
  NOR2_X2 U10546 ( .A1(n17447), .A2(n17446), .ZN(n17452) );
  NOR2_X2 U10547 ( .A1(n13421), .A2(n12465), .ZN(n17447) );
  NOR2_X2 U10548 ( .A1(n13423), .A2(n12897), .ZN(n17446) );
  NOR2_X2 U10549 ( .A1(n17449), .A2(n17448), .ZN(n17450) );
  NOR2_X1 U10550 ( .A1(n13426), .A2(n12467), .ZN(n17448) );
  NOR2_X2 U10551 ( .A1(n13431), .A2(n12466), .ZN(n17449) );
  NAND2_X2 U10552 ( .A1(n13111), .A2(net223743), .ZN(n13093) );
  INV_X4 U10553 ( .A(n15474), .ZN(n15398) );
  NAND2_X1 U10554 ( .A1(n15616), .A2(n15610), .ZN(n18700) );
  NAND2_X1 U10555 ( .A1(n15610), .A2(n10241), .ZN(n18701) );
  INV_X4 U10556 ( .A(n10803), .ZN(n13451) );
  INV_X4 U10557 ( .A(n13449), .ZN(n13448) );
  INV_X4 U10558 ( .A(n10805), .ZN(n13459) );
  INV_X4 U10559 ( .A(n13469), .ZN(n13467) );
  INV_X4 U10560 ( .A(n10804), .ZN(n13472) );
  OAI21_X1 U10561 ( .B1(n13485), .B2(n18666), .A(n18654), .ZN(n18655) );
  NOR2_X2 U10562 ( .A1(n18902), .A2(net232817), .ZN(n15694) );
  NOR2_X1 U10563 ( .A1(n18925), .A2(net222304), .ZN(n18633) );
  OAI21_X1 U10564 ( .B1(n15732), .B2(net232817), .A(n17125), .ZN(n15734) );
  INV_X4 U10565 ( .A(n17769), .ZN(n13366) );
  INV_X4 U10566 ( .A(n19158), .ZN(n13500) );
  INV_X4 U10567 ( .A(n19156), .ZN(n13497) );
  INV_X4 U10568 ( .A(n1881), .ZN(n13177) );
  NAND2_X2 U10569 ( .A1(n14982), .A2(n2511), .ZN(n1881) );
  INV_X4 U10570 ( .A(n15327), .ZN(n13179) );
  NAND2_X2 U10571 ( .A1(n14982), .A2(n2503), .ZN(n15327) );
  INV_X8 U10572 ( .A(n13196), .ZN(n13197) );
  INV_X8 U10573 ( .A(n11572), .ZN(n13193) );
  INV_X4 U10574 ( .A(n10803), .ZN(n13450) );
  INV_X4 U10575 ( .A(n13449), .ZN(n13447) );
  INV_X8 U10576 ( .A(n11992), .ZN(n13202) );
  NAND3_X1 U10577 ( .A1(n18854), .A2(n19011), .A3(n18853), .ZN(n18857) );
  NOR2_X2 U10578 ( .A1(n18850), .A2(n19023), .ZN(n18854) );
  NOR3_X2 U10579 ( .A1(n18852), .A2(n18919), .A3(n18881), .ZN(n18853) );
  NAND3_X1 U10580 ( .A1(n19047), .A2(n19076), .A3(n19111), .ZN(n18856) );
  NOR2_X1 U10581 ( .A1(n19105), .A2(n19104), .ZN(n19106) );
  AOI211_X2 U10582 ( .C1(n19118), .C2(n19117), .A(n19116), .B(n19115), .ZN(
        n19119) );
  NOR2_X2 U10583 ( .A1(net231345), .A2(n11990), .ZN(n19116) );
  NOR2_X2 U10584 ( .A1(n19114), .A2(n10815), .ZN(n19115) );
  NAND2_X2 U10585 ( .A1(DMEM_BUS_OUT[28]), .A2(n13484), .ZN(n15680) );
  INV_X4 U10586 ( .A(n13072), .ZN(n14148) );
  NOR2_X2 U10587 ( .A1(n14974), .A2(n14973), .ZN(n14975) );
  NOR2_X2 U10588 ( .A1(n11015), .A2(n14972), .ZN(n14974) );
  NOR3_X2 U10589 ( .A1(n14655), .A2(n14654), .A3(n14653), .ZN(n3684) );
  NOR2_X2 U10590 ( .A1(n13258), .A2(n11649), .ZN(n14655) );
  NOR2_X2 U10591 ( .A1(n13260), .A2(n11681), .ZN(n14653) );
  NOR2_X2 U10592 ( .A1(n14902), .A2(n14901), .ZN(n14903) );
  NOR2_X2 U10593 ( .A1(n12094), .A2(n13173), .ZN(n14902) );
  NOR2_X2 U10594 ( .A1(n14556), .A2(n14555), .ZN(n14557) );
  NOR2_X2 U10595 ( .A1(n12073), .A2(n13171), .ZN(n14555) );
  NOR2_X2 U10596 ( .A1(n14892), .A2(n14891), .ZN(n14893) );
  NOR2_X2 U10597 ( .A1(n12093), .A2(n13172), .ZN(n14892) );
  NOR2_X2 U10598 ( .A1(n14545), .A2(n14544), .ZN(n14546) );
  NOR2_X2 U10599 ( .A1(n12381), .A2(n13170), .ZN(n14544) );
  NOR2_X2 U10600 ( .A1(n14852), .A2(n14851), .ZN(n14853) );
  NOR2_X2 U10601 ( .A1(n12089), .A2(n14972), .ZN(n14852) );
  NOR2_X2 U10602 ( .A1(n14501), .A2(n14500), .ZN(n14502) );
  NOR2_X2 U10603 ( .A1(n12373), .A2(n14633), .ZN(n14500) );
  NOR2_X2 U10604 ( .A1(n14882), .A2(n14881), .ZN(n14883) );
  NOR2_X2 U10605 ( .A1(n12092), .A2(n14972), .ZN(n14882) );
  NOR2_X2 U10606 ( .A1(n14534), .A2(n14533), .ZN(n14535) );
  NOR2_X2 U10607 ( .A1(n12379), .A2(n14633), .ZN(n14533) );
  NOR2_X2 U10608 ( .A1(n14872), .A2(n14871), .ZN(n14873) );
  NOR2_X2 U10609 ( .A1(n12091), .A2(n13173), .ZN(n14872) );
  NOR2_X2 U10610 ( .A1(n14862), .A2(n14861), .ZN(n14863) );
  NOR2_X2 U10611 ( .A1(n12090), .A2(n13172), .ZN(n14862) );
  NOR2_X2 U10612 ( .A1(n13183), .A2(n12382), .ZN(n14989) );
  NOR2_X2 U10613 ( .A1(n13188), .A2(n12383), .ZN(n14992) );
  NOR3_X2 U10614 ( .A1(n15002), .A2(n15001), .A3(n15000), .ZN(n15003) );
  NOR2_X2 U10615 ( .A1(n12825), .A2(n13275), .ZN(n14983) );
  NOR2_X2 U10616 ( .A1(n14832), .A2(n14831), .ZN(n14833) );
  NOR2_X2 U10617 ( .A1(n11012), .A2(n13172), .ZN(n14832) );
  NOR2_X2 U10618 ( .A1(n14479), .A2(n14478), .ZN(n14480) );
  NOR2_X2 U10619 ( .A1(n12369), .A2(n13170), .ZN(n14478) );
  NOR2_X2 U10620 ( .A1(n14782), .A2(n14781), .ZN(n14783) );
  NOR2_X2 U10621 ( .A1(n11007), .A2(n13173), .ZN(n14782) );
  NOR2_X2 U10622 ( .A1(n14424), .A2(n14423), .ZN(n14425) );
  NOR2_X2 U10623 ( .A1(n12359), .A2(n13171), .ZN(n14423) );
  NOR2_X2 U10624 ( .A1(n13183), .A2(n12392), .ZN(n15054) );
  NOR2_X2 U10625 ( .A1(n13188), .A2(n12393), .ZN(n15055) );
  NOR3_X2 U10626 ( .A1(n15060), .A2(n15059), .A3(n15058), .ZN(n15061) );
  NOR2_X2 U10627 ( .A1(n12829), .A2(n13276), .ZN(n15049) );
  NOR2_X2 U10628 ( .A1(n13183), .A2(n12396), .ZN(n15091) );
  NOR2_X2 U10629 ( .A1(n13188), .A2(n12397), .ZN(n15092) );
  NOR3_X2 U10630 ( .A1(n15097), .A2(n15096), .A3(n15095), .ZN(n15098) );
  NOR2_X2 U10631 ( .A1(n12837), .A2(n13276), .ZN(n15086) );
  NOR2_X2 U10632 ( .A1(n11966), .A2(n17870), .ZN(n16298) );
  NOR2_X2 U10633 ( .A1(n14772), .A2(n14771), .ZN(n14773) );
  NOR2_X2 U10634 ( .A1(n11006), .A2(n13172), .ZN(n14772) );
  NOR2_X2 U10635 ( .A1(n14413), .A2(n14412), .ZN(n14414) );
  NOR2_X2 U10636 ( .A1(n12357), .A2(n13170), .ZN(n14412) );
  NOR2_X2 U10637 ( .A1(n13183), .A2(n12394), .ZN(n15075) );
  NOR2_X2 U10638 ( .A1(n13188), .A2(n12395), .ZN(n15076) );
  NOR3_X2 U10639 ( .A1(n15081), .A2(n15080), .A3(n15079), .ZN(n15082) );
  NOR2_X2 U10640 ( .A1(n12849), .A2(n13276), .ZN(n15070) );
  NOR2_X2 U10642 ( .A1(n13183), .A2(n12399), .ZN(n15122) );
  NOR2_X2 U10643 ( .A1(n13188), .A2(n12400), .ZN(n15123) );
  NOR3_X2 U10644 ( .A1(n15128), .A2(n15127), .A3(n15126), .ZN(n15129) );
  NOR2_X2 U10645 ( .A1(n12853), .A2(n13275), .ZN(n15117) );
  NOR2_X2 U10646 ( .A1(n14822), .A2(n14821), .ZN(n14823) );
  NOR2_X2 U10647 ( .A1(n11011), .A2(n14972), .ZN(n14822) );
  NOR2_X2 U10648 ( .A1(n14468), .A2(n14467), .ZN(n14469) );
  NOR2_X2 U10649 ( .A1(n12367), .A2(n14633), .ZN(n14467) );
  NOR2_X2 U10650 ( .A1(n13183), .A2(n12401), .ZN(n15143) );
  NOR2_X2 U10651 ( .A1(n13188), .A2(n12402), .ZN(n15144) );
  NOR3_X2 U10652 ( .A1(n15149), .A2(n15148), .A3(n15147), .ZN(n15150) );
  NOR2_X2 U10653 ( .A1(n12861), .A2(n13275), .ZN(n15138) );
  NOR2_X2 U10654 ( .A1(n12869), .A2(n13273), .ZN(n15159) );
  NOR2_X2 U10655 ( .A1(n13726), .A2(n11693), .ZN(n15160) );
  NOR3_X2 U10656 ( .A1(n15164), .A2(n15163), .A3(n15162), .ZN(n2180) );
  NOR2_X2 U10657 ( .A1(n13282), .A2(n12403), .ZN(n15162) );
  NOR2_X2 U10658 ( .A1(n13729), .A2(n11692), .ZN(n15163) );
  NOR2_X2 U10659 ( .A1(n13183), .A2(n12388), .ZN(n15028) );
  NOR2_X2 U10660 ( .A1(n13188), .A2(n12389), .ZN(n15029) );
  NOR3_X2 U10661 ( .A1(n15034), .A2(n15033), .A3(n15032), .ZN(n15035) );
  NOR2_X2 U10662 ( .A1(n12871), .A2(n13275), .ZN(n15023) );
  AOI21_X1 U10663 ( .B1(n16874), .B2(n16873), .A(n18874), .ZN(n16875) );
  AOI21_X1 U10664 ( .B1(n17982), .B2(n16872), .A(n16871), .ZN(n16874) );
  NOR2_X1 U10665 ( .A1(n13209), .A2(n16870), .ZN(n16871) );
  NOR2_X1 U10666 ( .A1(n19047), .A2(n13491), .ZN(n16893) );
  OAI21_X2 U10667 ( .B1(n19114), .B2(n11943), .A(n16891), .ZN(n16894) );
  OAI21_X1 U10668 ( .B1(EXEC_STAGE_imm26_32[6]), .B2(net227290), .A(net232877), 
        .ZN(net224816) );
  OAI21_X1 U10669 ( .B1(EXEC_STAGE_imm26_32[7]), .B2(net227290), .A(net232877), 
        .ZN(n16969) );
  OAI21_X1 U10670 ( .B1(EXEC_STAGE_imm26_32[8]), .B2(net227290), .A(net232877), 
        .ZN(net225195) );
  NOR2_X2 U10672 ( .A1(n12883), .A2(n13273), .ZN(n15173) );
  NOR2_X2 U10673 ( .A1(n13726), .A2(n11696), .ZN(n15174) );
  NOR3_X2 U10674 ( .A1(n15179), .A2(n15178), .A3(n15177), .ZN(n2160) );
  NOR2_X2 U10675 ( .A1(n13282), .A2(n12404), .ZN(n15177) );
  NOR2_X2 U10676 ( .A1(n13729), .A2(n11695), .ZN(n15178) );
  NAND3_X2 U10677 ( .A1(n14022), .A2(n14021), .A3(n14020), .ZN(n17094) );
  INV_X8 U10678 ( .A(n10801), .ZN(n13181) );
  INV_X4 U10679 ( .A(n13497), .ZN(n13496) );
  INV_X8 U10680 ( .A(n13175), .ZN(n13176) );
  INV_X4 U10681 ( .A(n2189), .ZN(n13175) );
  NAND2_X2 U10682 ( .A1(n14982), .A2(n2506), .ZN(n2189) );
  NOR2_X2 U10683 ( .A1(n13183), .A2(n12385), .ZN(n15012) );
  NOR2_X2 U10684 ( .A1(n13188), .A2(n12386), .ZN(n15013) );
  NOR3_X2 U10685 ( .A1(n15018), .A2(n15017), .A3(n15016), .ZN(n15019) );
  NOR2_X2 U10686 ( .A1(n12885), .A2(n13276), .ZN(n15007) );
  NAND3_X2 U10687 ( .A1(net224704), .A2(nextPC_ex_out[2]), .A3(
        nextPC_ex_out[3]), .ZN(n17201) );
  INV_X8 U10688 ( .A(n10354), .ZN(n13183) );
  INV_X4 U10689 ( .A(n13728), .ZN(n13727) );
  INV_X16 U10690 ( .A(n13489), .ZN(n13487) );
  NOR3_X2 U10691 ( .A1(n15186), .A2(n15185), .A3(n15184), .ZN(n2139) );
  NOR2_X2 U10692 ( .A1(n13282), .A2(n12405), .ZN(n15184) );
  NOR2_X2 U10693 ( .A1(n13729), .A2(n11698), .ZN(n15185) );
  NOR3_X2 U10694 ( .A1(n15182), .A2(n15181), .A3(n15180), .ZN(n2138) );
  NOR2_X2 U10695 ( .A1(n13726), .A2(n11699), .ZN(n15181) );
  NOR2_X2 U10696 ( .A1(n12893), .A2(n13273), .ZN(n15180) );
  INV_X16 U10697 ( .A(n13500), .ZN(n13499) );
  NOR3_X2 U10698 ( .A1(n15193), .A2(n15192), .A3(n15191), .ZN(n2119) );
  NOR2_X2 U10699 ( .A1(n13282), .A2(n12406), .ZN(n15191) );
  NOR2_X2 U10700 ( .A1(n13729), .A2(n11701), .ZN(n15192) );
  NOR3_X2 U10701 ( .A1(n15189), .A2(n15188), .A3(n15187), .ZN(n2118) );
  NOR2_X2 U10702 ( .A1(n13726), .A2(n11702), .ZN(n15188) );
  NOR2_X2 U10703 ( .A1(n12895), .A2(n13273), .ZN(n15187) );
  NOR3_X2 U10704 ( .A1(n15199), .A2(n15198), .A3(n15197), .ZN(n2099) );
  NOR2_X2 U10705 ( .A1(n13282), .A2(n12407), .ZN(n15197) );
  NOR2_X2 U10706 ( .A1(n13729), .A2(n11704), .ZN(n15198) );
  NOR3_X2 U10707 ( .A1(n15196), .A2(n15195), .A3(n15194), .ZN(n2098) );
  NOR2_X2 U10708 ( .A1(n13726), .A2(n11705), .ZN(n15195) );
  NOR2_X2 U10709 ( .A1(n12897), .A2(n13273), .ZN(n15194) );
  NAND3_X2 U10710 ( .A1(n16881), .A2(n16880), .A3(n17305), .ZN(n17565) );
  AOI21_X1 U10711 ( .B1(n18611), .B2(n18601), .A(n18612), .ZN(n15914) );
  NOR2_X2 U10712 ( .A1(n14792), .A2(n14791), .ZN(n14793) );
  NOR2_X2 U10713 ( .A1(n11008), .A2(n14972), .ZN(n14792) );
  NOR2_X2 U10714 ( .A1(n14435), .A2(n14434), .ZN(n14436) );
  NOR2_X2 U10715 ( .A1(n12361), .A2(n14633), .ZN(n14434) );
  NOR3_X2 U10716 ( .A1(n15205), .A2(n15204), .A3(n15203), .ZN(n2079) );
  NOR2_X2 U10717 ( .A1(n13282), .A2(n12408), .ZN(n15203) );
  NOR2_X2 U10718 ( .A1(n13729), .A2(n11707), .ZN(n15204) );
  NOR3_X2 U10719 ( .A1(n15202), .A2(n15201), .A3(n15200), .ZN(n2078) );
  NOR2_X2 U10720 ( .A1(n13726), .A2(n11708), .ZN(n15201) );
  NOR2_X2 U10721 ( .A1(n12899), .A2(n13273), .ZN(n15200) );
  NAND3_X2 U10722 ( .A1(n17658), .A2(n17657), .A3(n17656), .ZN(n17661) );
  AOI21_X2 U10723 ( .B1(n13196), .B2(REG_FILE_reg_out_22__21_), .A(n17655), 
        .ZN(n17656) );
  NOR3_X2 U10724 ( .A1(n17640), .A2(n17639), .A3(n17638), .ZN(n17665) );
  NAND3_X2 U10725 ( .A1(n17637), .A2(n17636), .A3(n17635), .ZN(n17640) );
  NOR3_X2 U10726 ( .A1(n17654), .A2(n17653), .A3(n17652), .ZN(n17663) );
  NAND3_X2 U10727 ( .A1(n14008), .A2(n14007), .A3(n14006), .ZN(n17622) );
  NOR2_X2 U10728 ( .A1(n14802), .A2(n14801), .ZN(n14803) );
  NOR2_X2 U10729 ( .A1(n11009), .A2(n13172), .ZN(n14802) );
  NOR2_X2 U10730 ( .A1(n14446), .A2(n14445), .ZN(n14447) );
  NOR2_X2 U10731 ( .A1(n12363), .A2(n13170), .ZN(n14445) );
  INV_X4 U10732 ( .A(n13363), .ZN(n13361) );
  NOR3_X2 U10733 ( .A1(n15211), .A2(n15210), .A3(n15209), .ZN(n2059) );
  NOR2_X2 U10734 ( .A1(n13282), .A2(n12409), .ZN(n15209) );
  NOR2_X2 U10735 ( .A1(n13729), .A2(n11710), .ZN(n15210) );
  NOR3_X2 U10736 ( .A1(n15208), .A2(n15207), .A3(n15206), .ZN(n2058) );
  NOR2_X2 U10737 ( .A1(n13726), .A2(n11711), .ZN(n15207) );
  NOR2_X2 U10738 ( .A1(n12901), .A2(n13273), .ZN(n15206) );
  NOR3_X2 U10739 ( .A1(n17793), .A2(n17792), .A3(n17791), .ZN(n17819) );
  NAND3_X2 U10740 ( .A1(n17790), .A2(n17789), .A3(n17788), .ZN(n17793) );
  NOR3_X2 U10741 ( .A1(n17815), .A2(n17814), .A3(n17813), .ZN(n17816) );
  NAND3_X2 U10742 ( .A1(n17812), .A2(n17811), .A3(n17810), .ZN(n17815) );
  AOI22_X2 U10743 ( .A1(MEM_WB_OUT[22]), .A2(n13878), .B1(MEM_WB_OUT[91]), 
        .B2(n14102), .ZN(n14016) );
  NOR2_X2 U10744 ( .A1(n14812), .A2(n14811), .ZN(n14813) );
  NOR2_X2 U10745 ( .A1(n11010), .A2(n13173), .ZN(n14812) );
  NOR2_X2 U10746 ( .A1(n14457), .A2(n14456), .ZN(n14458) );
  NOR2_X2 U10747 ( .A1(n12365), .A2(n13171), .ZN(n14456) );
  NAND3_X2 U10748 ( .A1(n15805), .A2(n15804), .A3(n15803), .ZN(n18914) );
  NOR2_X2 U10749 ( .A1(n12903), .A2(n13273), .ZN(n15212) );
  NOR2_X2 U10750 ( .A1(n13726), .A2(n11714), .ZN(n15213) );
  NOR3_X2 U10751 ( .A1(n15217), .A2(n15216), .A3(n15215), .ZN(n2039) );
  NOR2_X2 U10752 ( .A1(n13282), .A2(n12410), .ZN(n15215) );
  NOR2_X2 U10753 ( .A1(n13729), .A2(n11713), .ZN(n15216) );
  NAND3_X2 U10754 ( .A1(n17961), .A2(n17960), .A3(n17959), .ZN(n17964) );
  AOI21_X2 U10755 ( .B1(n13196), .B2(REG_FILE_reg_out_22__23_), .A(n17958), 
        .ZN(n17959) );
  NAND3_X2 U10756 ( .A1(n17939), .A2(n17938), .A3(n17937), .ZN(n17942) );
  NOR2_X2 U10757 ( .A1(n14942), .A2(n14941), .ZN(n14943) );
  NOR2_X2 U10758 ( .A1(n12098), .A2(n14972), .ZN(n14942) );
  NOR2_X2 U10759 ( .A1(n14600), .A2(n14599), .ZN(n14601) );
  NOR2_X2 U10760 ( .A1(n12077), .A2(n14633), .ZN(n14599) );
  INV_X4 U10761 ( .A(n13381), .ZN(n13379) );
  NOR2_X2 U10762 ( .A1(n12905), .A2(n13273), .ZN(n15226) );
  NOR2_X2 U10763 ( .A1(n13726), .A2(n11717), .ZN(n15227) );
  NOR3_X2 U10764 ( .A1(n15231), .A2(n15230), .A3(n15229), .ZN(n2019) );
  NOR2_X2 U10765 ( .A1(n13281), .A2(n11497), .ZN(n15229) );
  NOR2_X2 U10766 ( .A1(n13729), .A2(n11716), .ZN(n15230) );
  NAND3_X2 U10767 ( .A1(n18051), .A2(n18050), .A3(n18049), .ZN(n18054) );
  AOI21_X2 U10768 ( .B1(n13196), .B2(REG_FILE_reg_out_22__24_), .A(n18048), 
        .ZN(n18049) );
  NAND3_X2 U10769 ( .A1(n18029), .A2(n18028), .A3(n18027), .ZN(n18032) );
  NOR2_X2 U10770 ( .A1(n13729), .A2(n11719), .ZN(n15244) );
  NOR2_X2 U10771 ( .A1(n13281), .A2(n11498), .ZN(n15243) );
  NOR3_X2 U10772 ( .A1(n15242), .A2(n15241), .A3(n15240), .ZN(n1998) );
  NOR2_X2 U10773 ( .A1(n13726), .A2(n11720), .ZN(n15241) );
  NOR2_X2 U10774 ( .A1(n12907), .A2(n13272), .ZN(n15240) );
  NAND3_X2 U10775 ( .A1(n18094), .A2(n18093), .A3(n18092), .ZN(n18097) );
  AOI21_X2 U10776 ( .B1(n13196), .B2(REG_FILE_reg_out_22__25_), .A(n18091), 
        .ZN(n18092) );
  NAND3_X2 U10777 ( .A1(n18072), .A2(n18071), .A3(n18070), .ZN(n18075) );
  NOR2_X2 U10778 ( .A1(n13729), .A2(n11722), .ZN(n15259) );
  NOR2_X2 U10779 ( .A1(n13281), .A2(n11499), .ZN(n15258) );
  NOR3_X2 U10780 ( .A1(n15256), .A2(n15255), .A3(n15254), .ZN(n1978) );
  NOR2_X2 U10781 ( .A1(n13726), .A2(n11723), .ZN(n15255) );
  NOR2_X2 U10782 ( .A1(n12909), .A2(n13273), .ZN(n15254) );
  NAND3_X2 U10783 ( .A1(n18139), .A2(n18138), .A3(n18137), .ZN(n18142) );
  AOI21_X2 U10784 ( .B1(n13196), .B2(REG_FILE_reg_out_22__26_), .A(n18136), 
        .ZN(n18137) );
  NAND3_X2 U10785 ( .A1(n18117), .A2(n18116), .A3(n18115), .ZN(n18120) );
  NOR2_X2 U10786 ( .A1(n12911), .A2(n13272), .ZN(n15269) );
  NOR2_X2 U10787 ( .A1(n13726), .A2(n11726), .ZN(n15270) );
  NOR3_X2 U10788 ( .A1(n15274), .A2(n15273), .A3(n15272), .ZN(n1959) );
  NOR2_X2 U10789 ( .A1(n13281), .A2(n11500), .ZN(n15272) );
  NOR2_X2 U10790 ( .A1(n13729), .A2(n11725), .ZN(n15273) );
  NAND3_X2 U10791 ( .A1(n18180), .A2(n18179), .A3(n18178), .ZN(n18183) );
  AOI21_X2 U10792 ( .B1(n13196), .B2(REG_FILE_reg_out_22__27_), .A(n18177), 
        .ZN(n18178) );
  NAND3_X2 U10793 ( .A1(n18158), .A2(n18157), .A3(n18156), .ZN(n18161) );
  NOR2_X2 U10794 ( .A1(n13727), .A2(n11729), .ZN(n15284) );
  NOR2_X2 U10795 ( .A1(n12913), .A2(n13272), .ZN(n15283) );
  NOR3_X2 U10796 ( .A1(n15290), .A2(n15289), .A3(n15288), .ZN(n1938) );
  NOR2_X2 U10797 ( .A1(n13281), .A2(n11501), .ZN(n15288) );
  NOR2_X2 U10798 ( .A1(n13730), .A2(n11728), .ZN(n15289) );
  NAND3_X2 U10799 ( .A1(n18225), .A2(n18224), .A3(n18223), .ZN(n18228) );
  AOI21_X2 U10800 ( .B1(n13196), .B2(REG_FILE_reg_out_22__28_), .A(n18222), 
        .ZN(n18223) );
  NAND3_X2 U10801 ( .A1(n18203), .A2(n18202), .A3(n18201), .ZN(n18206) );
  NOR2_X2 U10802 ( .A1(n14922), .A2(n14921), .ZN(n14923) );
  NOR2_X2 U10803 ( .A1(n12096), .A2(n13172), .ZN(n14922) );
  NOR2_X2 U10804 ( .A1(n14578), .A2(n14577), .ZN(n14579) );
  NOR2_X2 U10805 ( .A1(n12075), .A2(n13170), .ZN(n14577) );
  AOI21_X2 U10806 ( .B1(n13964), .B2(n13963), .A(n13962), .ZN(n13965) );
  NOR2_X2 U10807 ( .A1(n14932), .A2(n14931), .ZN(n14933) );
  NOR2_X2 U10808 ( .A1(n12097), .A2(n13173), .ZN(n14932) );
  NOR2_X2 U10809 ( .A1(n14589), .A2(n14588), .ZN(n14590) );
  NOR2_X2 U10810 ( .A1(n12076), .A2(n13171), .ZN(n14588) );
  NOR2_X2 U10811 ( .A1(n14912), .A2(n14911), .ZN(n14913) );
  NOR2_X2 U10812 ( .A1(n12095), .A2(n14972), .ZN(n14912) );
  NOR2_X2 U10813 ( .A1(n14567), .A2(n14566), .ZN(n14568) );
  NOR2_X2 U10814 ( .A1(n12074), .A2(n14633), .ZN(n14566) );
  NOR2_X2 U10815 ( .A1(n14952), .A2(n14951), .ZN(n14953) );
  NOR2_X2 U10816 ( .A1(n12099), .A2(n13172), .ZN(n14952) );
  NOR2_X2 U10817 ( .A1(n14611), .A2(n14610), .ZN(n14612) );
  NOR2_X2 U10818 ( .A1(n12078), .A2(n13170), .ZN(n14610) );
  NOR2_X2 U10819 ( .A1(n13727), .A2(n11732), .ZN(n15300) );
  NOR2_X2 U10820 ( .A1(n12915), .A2(n13273), .ZN(n15299) );
  NOR3_X2 U10821 ( .A1(n15304), .A2(n15303), .A3(n15302), .ZN(n1918) );
  NOR2_X2 U10822 ( .A1(n13281), .A2(n11502), .ZN(n15302) );
  NOR2_X2 U10823 ( .A1(n13730), .A2(n11731), .ZN(n15303) );
  NAND3_X2 U10824 ( .A1(n18433), .A2(n18432), .A3(n18431), .ZN(n18436) );
  AOI21_X2 U10825 ( .B1(n13196), .B2(REG_FILE_reg_out_22__29_), .A(n18430), 
        .ZN(n18431) );
  NAND3_X2 U10826 ( .A1(n18411), .A2(n18410), .A3(n18409), .ZN(n18414) );
  NOR2_X2 U10827 ( .A1(n14962), .A2(n14961), .ZN(n14963) );
  NOR2_X2 U10828 ( .A1(n11014), .A2(n13173), .ZN(n14962) );
  NOR2_X2 U10829 ( .A1(n14622), .A2(n14621), .ZN(n14623) );
  NOR2_X2 U10830 ( .A1(n11494), .A2(n13171), .ZN(n14621) );
  NOR2_X2 U10831 ( .A1(n13727), .A2(n11735), .ZN(n15314) );
  NOR2_X2 U10832 ( .A1(n12917), .A2(n13272), .ZN(n15313) );
  NOR3_X2 U10833 ( .A1(n15318), .A2(n15317), .A3(n15316), .ZN(n1898) );
  NOR2_X2 U10834 ( .A1(n13281), .A2(n11503), .ZN(n15316) );
  NOR2_X2 U10835 ( .A1(n13730), .A2(n11734), .ZN(n15317) );
  NAND3_X2 U10836 ( .A1(n18514), .A2(n18513), .A3(n18512), .ZN(n18517) );
  AOI21_X2 U10837 ( .B1(n13196), .B2(REG_FILE_reg_out_22__30_), .A(n18511), 
        .ZN(n18512) );
  NAND3_X2 U10838 ( .A1(n18489), .A2(n18488), .A3(n18487), .ZN(n18492) );
  NOR2_X2 U10840 ( .A1(n14842), .A2(n14841), .ZN(n14843) );
  NOR2_X2 U10841 ( .A1(n11013), .A2(n13173), .ZN(n14842) );
  NOR2_X2 U10842 ( .A1(n14490), .A2(n14489), .ZN(n14491) );
  NOR2_X2 U10843 ( .A1(n12371), .A2(n13171), .ZN(n14489) );
  INV_X8 U10844 ( .A(n18664), .ZN(n13408) );
  NAND3_X2 U10845 ( .A1(n16775), .A2(n16795), .A3(n16774), .ZN(n17587) );
  INV_X4 U10846 ( .A(net231353), .ZN(net231335) );
  INV_X4 U10847 ( .A(n13375), .ZN(n13373) );
  INV_X4 U10848 ( .A(n13372), .ZN(n13371) );
  INV_X4 U10849 ( .A(n13366), .ZN(n13364) );
  INV_X8 U10850 ( .A(n13184), .ZN(n19153) );
  INV_X16 U10851 ( .A(n13500), .ZN(n13498) );
  NOR2_X2 U10852 ( .A1(n13727), .A2(n12411), .ZN(n15332) );
  NOR2_X2 U10853 ( .A1(n12919), .A2(n13273), .ZN(n15331) );
  INV_X4 U10854 ( .A(n13497), .ZN(n13495) );
  INV_X4 U10855 ( .A(n13176), .ZN(n19160) );
  INV_X4 U10856 ( .A(n13181), .ZN(n19155) );
  NOR3_X2 U10857 ( .A1(n15339), .A2(n15338), .A3(n15337), .ZN(n1861) );
  NOR2_X2 U10858 ( .A1(n13281), .A2(n12135), .ZN(n15337) );
  NOR2_X2 U10859 ( .A1(n13730), .A2(n12412), .ZN(n15338) );
  INV_X4 U10860 ( .A(n10842), .ZN(n13742) );
  INV_X4 U10861 ( .A(net231339), .ZN(net231273) );
  NOR2_X2 U10862 ( .A1(n14635), .A2(n14634), .ZN(n14636) );
  NOR2_X2 U10863 ( .A1(n11496), .A2(n14633), .ZN(n14634) );
  NAND3_X2 U10864 ( .A1(n14263), .A2(n14262), .A3(n14261), .ZN(n14268) );
  AOI21_X1 U10865 ( .B1(n16812), .B2(n16811), .A(n18885), .ZN(n16813) );
  OAI21_X2 U10866 ( .B1(n19114), .B2(n10813), .A(n16822), .ZN(n16825) );
  NOR2_X2 U10867 ( .A1(net231217), .A2(n11947), .ZN(n18259) );
  OAI21_X1 U10868 ( .B1(n18455), .B2(n18463), .A(n18285), .ZN(n18286) );
  NAND3_X1 U10869 ( .A1(n19107), .A2(n13163), .A3(n18360), .ZN(n18285) );
  NOR2_X1 U10870 ( .A1(n17494), .A2(n18280), .ZN(n18283) );
  NAND3_X2 U10871 ( .A1(n18278), .A2(n18277), .A3(n18276), .ZN(n18367) );
  OAI21_X2 U10872 ( .B1(n18365), .B2(n18463), .A(n18364), .ZN(n18366) );
  NAND3_X1 U10873 ( .A1(n10363), .A2(n18644), .A3(n13159), .ZN(n18364) );
  NOR3_X2 U10874 ( .A1(n18378), .A2(n18377), .A3(n18376), .ZN(n18379) );
  NOR2_X2 U10875 ( .A1(net231217), .A2(n11949), .ZN(n18377) );
  NOR2_X2 U10876 ( .A1(net231217), .A2(n12037), .ZN(n18453) );
  NOR2_X2 U10877 ( .A1(n18463), .A2(n18462), .ZN(n18464) );
  NOR2_X2 U10878 ( .A1(n19114), .A2(n11933), .ZN(n18390) );
  NAND3_X2 U10879 ( .A1(n16315), .A2(n16314), .A3(n16313), .ZN(n16422) );
  NOR2_X1 U10880 ( .A1(n19001), .A2(n13491), .ZN(n16420) );
  OAI21_X2 U10881 ( .B1(n19114), .B2(n11942), .A(n16419), .ZN(n16421) );
  NAND3_X2 U10882 ( .A1(n16394), .A2(n16393), .A3(n16392), .ZN(n16530) );
  OAI21_X2 U10883 ( .B1(n19114), .B2(n11936), .A(n18344), .ZN(n18353) );
  NOR3_X1 U10884 ( .A1(n18325), .A2(n14011), .A3(n13209), .ZN(n18326) );
  NOR2_X2 U10885 ( .A1(n13221), .A2(n12029), .ZN(n18755) );
  NOR2_X2 U10886 ( .A1(n14966), .A2(n14965), .ZN(n14967) );
  NOR2_X2 U10887 ( .A1(n13251), .A2(n11495), .ZN(n14966) );
  NOR2_X2 U10888 ( .A1(n13253), .A2(n11585), .ZN(n14965) );
  NOR2_X2 U10889 ( .A1(n14651), .A2(n14650), .ZN(n14652) );
  NOR2_X2 U10890 ( .A1(n13250), .A2(n12345), .ZN(n14651) );
  NOR2_X2 U10891 ( .A1(n13252), .A2(n12232), .ZN(n14650) );
  NOR2_X2 U10892 ( .A1(n14896), .A2(n14895), .ZN(n14897) );
  NOR2_X2 U10893 ( .A1(n13250), .A2(n11487), .ZN(n14896) );
  NOR2_X2 U10894 ( .A1(n13252), .A2(n12609), .ZN(n14895) );
  NOR2_X2 U10895 ( .A1(n13245), .A2(n11479), .ZN(n14561) );
  NOR2_X2 U10896 ( .A1(net231241), .A2(n10811), .ZN(n14559) );
  NOR2_X2 U10897 ( .A1(n14886), .A2(n14885), .ZN(n14887) );
  NOR2_X2 U10898 ( .A1(n13251), .A2(n12380), .ZN(n14886) );
  NOR2_X2 U10899 ( .A1(n13253), .A2(n12608), .ZN(n14885) );
  NOR2_X2 U10900 ( .A1(n13245), .A2(n12344), .ZN(n14550) );
  NOR2_X2 U10901 ( .A1(net231241), .A2(n11932), .ZN(n14548) );
  NOR2_X2 U10902 ( .A1(n14846), .A2(n14845), .ZN(n14847) );
  NOR2_X2 U10903 ( .A1(n13251), .A2(n12372), .ZN(n14846) );
  NOR2_X2 U10904 ( .A1(n13253), .A2(n12603), .ZN(n14845) );
  NOR2_X2 U10905 ( .A1(n13245), .A2(n12340), .ZN(n14506) );
  NOR2_X2 U10906 ( .A1(net231217), .A2(n11959), .ZN(n14504) );
  NOR2_X2 U10907 ( .A1(n14876), .A2(n14875), .ZN(n14877) );
  NOR2_X2 U10908 ( .A1(n13251), .A2(n12378), .ZN(n14876) );
  NOR2_X2 U10909 ( .A1(n13253), .A2(n12607), .ZN(n14875) );
  NOR2_X2 U10910 ( .A1(n13245), .A2(n12343), .ZN(n14539) );
  NOR2_X2 U10911 ( .A1(net231217), .A2(n10818), .ZN(n14537) );
  NOR2_X2 U10912 ( .A1(n14866), .A2(n14865), .ZN(n14867) );
  NOR2_X2 U10913 ( .A1(n13251), .A2(n12376), .ZN(n14866) );
  NOR2_X2 U10914 ( .A1(n13253), .A2(n12606), .ZN(n14865) );
  NOR2_X2 U10915 ( .A1(n14856), .A2(n14855), .ZN(n14857) );
  NOR2_X2 U10916 ( .A1(n13251), .A2(n12374), .ZN(n14856) );
  NOR2_X2 U10917 ( .A1(n13253), .A2(n12605), .ZN(n14855) );
  NOR2_X2 U10918 ( .A1(n14695), .A2(n14694), .ZN(n14696) );
  NOR2_X2 U10919 ( .A1(n13250), .A2(n12349), .ZN(n14695) );
  NOR2_X2 U10920 ( .A1(n13252), .A2(n12235), .ZN(n14694) );
  NOR2_X2 U10921 ( .A1(n13244), .A2(n12325), .ZN(n14340) );
  NOR2_X2 U10922 ( .A1(net231223), .A2(n11944), .ZN(n14338) );
  NOR2_X2 U10923 ( .A1(n4539), .A2(n4540), .ZN(n4524) );
  NOR2_X2 U10924 ( .A1(nextPC_ex_out[0]), .A2(n15652), .ZN(n15560) );
  NAND3_X2 U10925 ( .A1(n15575), .A2(n15573), .A3(n15572), .ZN(n15577) );
  OAI21_X2 U10926 ( .B1(nextPC_ex_out[0]), .B2(n15647), .A(n15557), .ZN(n15563) );
  AOI21_X2 U10927 ( .B1(n17924), .B2(n16882), .A(n15727), .ZN(n15752) );
  NOR2_X2 U10928 ( .A1(n14826), .A2(n14825), .ZN(n14827) );
  NOR2_X2 U10929 ( .A1(n13251), .A2(n12368), .ZN(n14826) );
  NOR2_X2 U10930 ( .A1(n13253), .A2(n12248), .ZN(n14825) );
  NOR2_X2 U10931 ( .A1(n13245), .A2(n12338), .ZN(n14484) );
  NOR2_X2 U10932 ( .A1(net231223), .A2(n11935), .ZN(n14482) );
  NOR2_X2 U10933 ( .A1(n14745), .A2(n14744), .ZN(n14746) );
  NOR2_X2 U10934 ( .A1(n13250), .A2(n12354), .ZN(n14745) );
  NOR2_X2 U10935 ( .A1(n13252), .A2(n12240), .ZN(n14744) );
  NOR2_X2 U10936 ( .A1(n13244), .A2(n12330), .ZN(n14395) );
  NOR2_X2 U10937 ( .A1(net231223), .A2(n11961), .ZN(n14393) );
  NOR2_X2 U10938 ( .A1(n4393), .A2(n4394), .ZN(n4378) );
  NOR2_X2 U10939 ( .A1(n14776), .A2(n14775), .ZN(n14777) );
  NOR2_X2 U10940 ( .A1(n13251), .A2(n12358), .ZN(n14776) );
  NOR2_X2 U10941 ( .A1(n13253), .A2(n12243), .ZN(n14775) );
  NOR2_X2 U10942 ( .A1(n13245), .A2(n12333), .ZN(n14429) );
  NOR2_X2 U10943 ( .A1(net231243), .A2(n10821), .ZN(n14427) );
  NOR2_X2 U10944 ( .A1(n14715), .A2(n14714), .ZN(n14716) );
  NOR2_X2 U10945 ( .A1(n13250), .A2(n12351), .ZN(n14715) );
  NOR2_X2 U10946 ( .A1(n13252), .A2(n12237), .ZN(n14714) );
  NOR2_X2 U10947 ( .A1(n13244), .A2(n12327), .ZN(n14362) );
  NOR2_X2 U10948 ( .A1(net231223), .A2(n11941), .ZN(n14360) );
  NOR2_X2 U10949 ( .A1(n4480), .A2(n4481), .ZN(n4465) );
  NOR2_X2 U10950 ( .A1(n14705), .A2(n14704), .ZN(n14706) );
  NOR2_X2 U10951 ( .A1(n13250), .A2(n12350), .ZN(n14705) );
  NOR2_X2 U10952 ( .A1(n13252), .A2(n12236), .ZN(n14704) );
  NOR2_X1 U10953 ( .A1(n19040), .A2(n13491), .ZN(n16004) );
  OAI21_X1 U10954 ( .B1(n17316), .B2(n13213), .A(n16036), .ZN(n16037) );
  NOR2_X2 U10955 ( .A1(n16023), .A2(n13207), .ZN(n16038) );
  NOR2_X2 U10956 ( .A1(net231217), .A2(n11967), .ZN(n16006) );
  NOR2_X2 U10957 ( .A1(n15069), .A2(n15068), .ZN(n2382) );
  NOR2_X2 U10958 ( .A1(n12834), .A2(n13272), .ZN(n15069) );
  NOR2_X2 U10959 ( .A1(n12835), .A2(n13269), .ZN(n15068) );
  NOR2_X2 U10960 ( .A1(n13183), .A2(n12416), .ZN(n16129) );
  NOR2_X2 U10961 ( .A1(n13188), .A2(n12417), .ZN(n16127) );
  NOR3_X2 U10962 ( .A1(n16135), .A2(n16134), .A3(n16133), .ZN(n16136) );
  NAND3_X2 U10963 ( .A1(n12526), .A2(n11461), .A3(n16132), .ZN(n16135) );
  AOI21_X1 U10964 ( .B1(n16149), .B2(n16148), .A(n19039), .ZN(n16150) );
  AOI21_X1 U10965 ( .B1(n17982), .B2(n16147), .A(n16146), .ZN(n16149) );
  NOR2_X1 U10966 ( .A1(n13209), .A2(n16145), .ZN(n16146) );
  OAI21_X2 U10967 ( .B1(n13217), .B2(n11941), .A(n16153), .ZN(n16156) );
  NOR2_X1 U10968 ( .A1(n19035), .A2(n13491), .ZN(n16155) );
  NOR2_X2 U10969 ( .A1(n14735), .A2(n14734), .ZN(n14736) );
  NOR2_X2 U10970 ( .A1(n13250), .A2(n12353), .ZN(n14735) );
  NOR2_X2 U10971 ( .A1(n13252), .A2(n12239), .ZN(n14734) );
  NOR2_X2 U10972 ( .A1(n13244), .A2(n12329), .ZN(n14384) );
  NOR2_X2 U10973 ( .A1(net231223), .A2(n10820), .ZN(n14382) );
  NOR2_X2 U10974 ( .A1(n4422), .A2(n4423), .ZN(n4407) );
  NOR2_X2 U10975 ( .A1(n16226), .A2(n13213), .ZN(n16227) );
  NAND3_X2 U10976 ( .A1(n16225), .A2(n16224), .A3(n16223), .ZN(n16228) );
  NOR2_X1 U10977 ( .A1(n19025), .A2(n13491), .ZN(n16216) );
  NOR2_X2 U10978 ( .A1(n14755), .A2(n14754), .ZN(n14756) );
  NOR2_X2 U10979 ( .A1(n13250), .A2(n12355), .ZN(n14755) );
  NOR2_X2 U10980 ( .A1(n13252), .A2(n12241), .ZN(n14754) );
  NOR2_X2 U10981 ( .A1(n13244), .A2(n12331), .ZN(n14407) );
  NOR2_X2 U10982 ( .A1(net231241), .A2(n11958), .ZN(n14405) );
  NOR2_X2 U10983 ( .A1(n4364), .A2(n4365), .ZN(n4349) );
  NOR2_X2 U10984 ( .A1(n15111), .A2(n15110), .ZN(n2301) );
  NOR2_X2 U10985 ( .A1(n12842), .A2(n13272), .ZN(n15111) );
  NOR2_X2 U10986 ( .A1(n12843), .A2(n13269), .ZN(n15110) );
  NOR2_X2 U10987 ( .A1(n13183), .A2(n12421), .ZN(n16278) );
  NOR2_X2 U10988 ( .A1(n13188), .A2(n12422), .ZN(n16276) );
  NOR3_X2 U10989 ( .A1(n16284), .A2(n16283), .A3(n16282), .ZN(n16285) );
  NAND3_X2 U10990 ( .A1(n12527), .A2(n11462), .A3(n16281), .ZN(n16284) );
  NOR2_X2 U10991 ( .A1(n14766), .A2(n14765), .ZN(n14767) );
  NOR2_X2 U10992 ( .A1(n13250), .A2(n12356), .ZN(n14766) );
  NOR2_X2 U10993 ( .A1(n13252), .A2(n12242), .ZN(n14765) );
  NOR2_X2 U10994 ( .A1(n13244), .A2(n12332), .ZN(n14418) );
  NOR2_X2 U10995 ( .A1(net231223), .A2(n11942), .ZN(n14416) );
  NOR2_X2 U10996 ( .A1(n15116), .A2(n15115), .ZN(n2281) );
  NOR2_X2 U10997 ( .A1(n12846), .A2(n13272), .ZN(n15116) );
  NOR2_X2 U10998 ( .A1(n12847), .A2(n13269), .ZN(n15115) );
  NOR2_X2 U10999 ( .A1(n13183), .A2(n12425), .ZN(n16378) );
  NOR2_X2 U11000 ( .A1(n13188), .A2(n12426), .ZN(n16376) );
  NOR3_X2 U11001 ( .A1(n16383), .A2(n16382), .A3(n16381), .ZN(n16384) );
  NAND3_X2 U11002 ( .A1(n12528), .A2(n11463), .A3(n16380), .ZN(n16383) );
  NOR2_X2 U11003 ( .A1(n14725), .A2(n14724), .ZN(n14726) );
  NOR2_X2 U11004 ( .A1(n13250), .A2(n12352), .ZN(n14725) );
  NOR2_X2 U11005 ( .A1(n13252), .A2(n12238), .ZN(n14724) );
  NOR2_X2 U11006 ( .A1(n13244), .A2(n12328), .ZN(n14373) );
  NOR2_X2 U11007 ( .A1(net231243), .A2(n11957), .ZN(n14371) );
  NOR2_X2 U11008 ( .A1(n4451), .A2(n4452), .ZN(n4436) );
  NOR2_X2 U11009 ( .A1(n14816), .A2(n14815), .ZN(n14817) );
  NOR2_X2 U11010 ( .A1(n13251), .A2(n12366), .ZN(n14816) );
  NOR2_X2 U11011 ( .A1(n13253), .A2(n12247), .ZN(n14815) );
  NOR2_X2 U11012 ( .A1(n13245), .A2(n12337), .ZN(n14473) );
  NOR2_X2 U11013 ( .A1(net231217), .A2(n10813), .ZN(n14471) );
  NOR2_X2 U11014 ( .A1(n15137), .A2(n15136), .ZN(n2241) );
  NOR2_X2 U11015 ( .A1(n12858), .A2(n13273), .ZN(n15137) );
  NOR2_X2 U11016 ( .A1(n12859), .A2(n13270), .ZN(n15136) );
  NOR2_X2 U11017 ( .A1(n13183), .A2(n12431), .ZN(n16606) );
  NOR2_X2 U11018 ( .A1(n13188), .A2(n12432), .ZN(n16604) );
  NOR3_X2 U11019 ( .A1(n16611), .A2(n16610), .A3(n16609), .ZN(n16612) );
  NAND3_X2 U11020 ( .A1(n12529), .A2(n11464), .A3(n16608), .ZN(n16611) );
  NOR2_X2 U11021 ( .A1(n15158), .A2(n15157), .ZN(n2196) );
  NOR2_X2 U11022 ( .A1(n12866), .A2(n13273), .ZN(n15158) );
  NOR2_X2 U11023 ( .A1(n12867), .A2(n13270), .ZN(n15157) );
  NOR2_X2 U11024 ( .A1(n13183), .A2(n12436), .ZN(n16710) );
  NOR2_X2 U11025 ( .A1(n13188), .A2(n12437), .ZN(n16708) );
  NOR3_X2 U11026 ( .A1(n16716), .A2(n16715), .A3(n16714), .ZN(n16717) );
  NAND3_X2 U11027 ( .A1(n12530), .A2(n11465), .A3(n16713), .ZN(n16716) );
  INV_X4 U11028 ( .A(n10832), .ZN(n13741) );
  NOR2_X2 U11029 ( .A1(n14675), .A2(n14674), .ZN(n14676) );
  NOR2_X2 U11030 ( .A1(n13250), .A2(n12347), .ZN(n14675) );
  NOR2_X2 U11031 ( .A1(n13252), .A2(n12233), .ZN(n14674) );
  NOR2_X2 U11032 ( .A1(n13244), .A2(n12323), .ZN(n14318) );
  NOR2_X2 U11033 ( .A1(net231223), .A2(n11943), .ZN(n14316) );
  NOR2_X2 U11034 ( .A1(n4597), .A2(n4598), .ZN(n4582) );
  NOR2_X2 U11035 ( .A1(n15043), .A2(n15042), .ZN(n2442) );
  NOR2_X2 U11036 ( .A1(n12876), .A2(n13272), .ZN(n15043) );
  NOR2_X2 U11037 ( .A1(n12877), .A2(n13269), .ZN(n15042) );
  NOR2_X2 U11038 ( .A1(n13183), .A2(n12444), .ZN(n16946) );
  NOR2_X2 U11039 ( .A1(n13188), .A2(n12445), .ZN(n16944) );
  NOR3_X2 U11040 ( .A1(n16951), .A2(n16950), .A3(n16949), .ZN(n16952) );
  NAND3_X2 U11041 ( .A1(n12531), .A2(n11466), .A3(n16948), .ZN(n16951) );
  AOI21_X2 U11042 ( .B1(net224711), .B2(n10356), .A(net225191), .ZN(n16962) );
  OAI21_X2 U11043 ( .B1(n10356), .B2(net224713), .A(net225188), .ZN(n16960) );
  NOR2_X2 U11044 ( .A1(nextPC_ex_out[6]), .A2(net225185), .ZN(net225192) );
  NOR2_X2 U11045 ( .A1(net231225), .A2(n12123), .ZN(n16964) );
  NOR2_X2 U11046 ( .A1(n15106), .A2(n15105), .ZN(n2321) );
  NOR2_X2 U11047 ( .A1(n12880), .A2(n13272), .ZN(n15106) );
  NOR2_X2 U11048 ( .A1(n12881), .A2(n13269), .ZN(n15105) );
  NOR2_X2 U11049 ( .A1(n13183), .A2(n12448), .ZN(n17019) );
  NOR2_X2 U11050 ( .A1(n13188), .A2(n12449), .ZN(n17017) );
  NOR3_X2 U11051 ( .A1(n17025), .A2(n17024), .A3(n17023), .ZN(n17026) );
  NAND3_X2 U11052 ( .A1(n12532), .A2(n11467), .A3(n17022), .ZN(n17025) );
  INV_X4 U11053 ( .A(net231339), .ZN(net231295) );
  OAI21_X1 U11054 ( .B1(EXEC_STAGE_imm26_32[9]), .B2(net227290), .A(net232877), 
        .ZN(net225077) );
  NOR2_X2 U11055 ( .A1(n11977), .A2(n17870), .ZN(n17048) );
  AOI21_X2 U11056 ( .B1(n17040), .B2(n17039), .A(n17038), .ZN(n17043) );
  OAI21_X2 U11057 ( .B1(n19114), .B2(n11935), .A(n17146), .ZN(n17148) );
  NOR2_X2 U11058 ( .A1(n14665), .A2(n14664), .ZN(n14666) );
  NOR2_X2 U11059 ( .A1(n13250), .A2(n12346), .ZN(n14665) );
  NOR2_X2 U11060 ( .A1(n13252), .A2(n12604), .ZN(n14664) );
  NOR2_X2 U11061 ( .A1(n13244), .A2(n12322), .ZN(n14307) );
  NOR2_X2 U11062 ( .A1(net231239), .A2(n11939), .ZN(n14305) );
  NOR2_X2 U11063 ( .A1(n4626), .A2(n4627), .ZN(n4611) );
  NOR2_X2 U11064 ( .A1(nextPC_ex_out[3]), .A2(n10358), .ZN(n17202) );
  NOR2_X2 U11065 ( .A1(net231229), .A2(n12124), .ZN(n17195) );
  NOR2_X2 U11066 ( .A1(n15048), .A2(n15047), .ZN(n2422) );
  NOR2_X2 U11067 ( .A1(n12890), .A2(n13272), .ZN(n15048) );
  NOR2_X2 U11068 ( .A1(n12891), .A2(n13269), .ZN(n15047) );
  NOR2_X2 U11069 ( .A1(n13183), .A2(n12456), .ZN(n17273) );
  NOR2_X2 U11070 ( .A1(n13188), .A2(n12457), .ZN(n17271) );
  NOR3_X2 U11071 ( .A1(n17278), .A2(n17277), .A3(n17276), .ZN(n17279) );
  NAND3_X2 U11072 ( .A1(n12533), .A2(n11468), .A3(n17275), .ZN(n17278) );
  OAI21_X2 U11073 ( .B1(n13217), .B2(n11944), .A(n17319), .ZN(n17321) );
  INV_X4 U11074 ( .A(n13207), .ZN(n18644) );
  NOR2_X1 U11075 ( .A1(n19044), .A2(n13491), .ZN(n17320) );
  OAI21_X2 U11076 ( .B1(n17316), .B2(n13211), .A(n17315), .ZN(n17317) );
  NOR2_X2 U11077 ( .A1(n17574), .A2(n13213), .ZN(n17318) );
  NOR2_X1 U11078 ( .A1(n18990), .A2(n13491), .ZN(n17506) );
  AOI21_X2 U11079 ( .B1(n17549), .B2(n17548), .A(n17547), .ZN(n17550) );
  AOI21_X1 U11080 ( .B1(n17982), .B2(n17546), .A(n17545), .ZN(n17549) );
  NOR2_X2 U11081 ( .A1(net231229), .A2(n11963), .ZN(n17508) );
  NOR2_X2 U11082 ( .A1(n14685), .A2(n14684), .ZN(n14686) );
  NOR2_X2 U11083 ( .A1(n13250), .A2(n12348), .ZN(n14685) );
  NOR2_X2 U11084 ( .A1(n13252), .A2(n12234), .ZN(n14684) );
  NOR2_X2 U11085 ( .A1(n13244), .A2(n12324), .ZN(n14329) );
  NOR2_X2 U11086 ( .A1(net231223), .A2(n11930), .ZN(n14327) );
  NOR2_X2 U11087 ( .A1(n4568), .A2(n4569), .ZN(n4553) );
  AOI21_X1 U11088 ( .B1(ID_EXEC_OUT[207]), .B2(n13216), .A(n17562), .ZN(n17563) );
  NOR2_X2 U11089 ( .A1(net231217), .A2(n11964), .ZN(n17562) );
  NOR2_X2 U11090 ( .A1(n17576), .A2(n13207), .ZN(n17577) );
  NOR2_X2 U11091 ( .A1(n14786), .A2(n14785), .ZN(n14787) );
  NOR2_X2 U11092 ( .A1(n13251), .A2(n12360), .ZN(n14786) );
  NOR2_X2 U11093 ( .A1(n13253), .A2(n12244), .ZN(n14785) );
  NOR2_X2 U11094 ( .A1(n13245), .A2(n12334), .ZN(n14440) );
  NOR2_X2 U11095 ( .A1(net231217), .A2(n11945), .ZN(n14438) );
  AOI211_X2 U11096 ( .C1(n19118), .C2(n17617), .A(n17616), .B(n17615), .ZN(
        n17618) );
  OAI21_X2 U11097 ( .B1(n19114), .B2(n11945), .A(n17614), .ZN(n17616) );
  NOR2_X1 U11098 ( .A1(n18917), .A2(n13491), .ZN(n17615) );
  NOR2_X2 U11099 ( .A1(n13207), .A2(n17689), .ZN(n17690) );
  NOR2_X1 U11100 ( .A1(n18989), .A2(n13491), .ZN(n17713) );
  NOR2_X2 U11101 ( .A1(n14796), .A2(n14795), .ZN(n14797) );
  NOR2_X2 U11102 ( .A1(n13251), .A2(n12362), .ZN(n14796) );
  NOR2_X2 U11103 ( .A1(n13253), .A2(n12245), .ZN(n14795) );
  NOR2_X2 U11104 ( .A1(n13245), .A2(n12335), .ZN(n14451) );
  NOR2_X2 U11105 ( .A1(net231217), .A2(n11940), .ZN(n14449) );
  NOR2_X2 U11106 ( .A1(n19114), .A2(n11940), .ZN(n17762) );
  NOR2_X2 U11107 ( .A1(net231217), .A2(n11968), .ZN(n17763) );
  INV_X4 U11108 ( .A(net231335), .ZN(net231307) );
  NOR2_X2 U11109 ( .A1(n13207), .A2(n17855), .ZN(n17856) );
  NOR2_X2 U11110 ( .A1(n18009), .A2(n13211), .ZN(n17857) );
  NOR2_X1 U11111 ( .A1(n18976), .A2(n13491), .ZN(n17860) );
  NOR2_X2 U11112 ( .A1(n14806), .A2(n14805), .ZN(n14807) );
  NOR2_X2 U11113 ( .A1(n13251), .A2(n12364), .ZN(n14806) );
  NOR2_X2 U11114 ( .A1(n13253), .A2(n12246), .ZN(n14805) );
  NOR2_X2 U11115 ( .A1(n13245), .A2(n12336), .ZN(n14462) );
  NOR2_X2 U11116 ( .A1(net231223), .A2(n10822), .ZN(n14460) );
  OAI21_X2 U11117 ( .B1(net231221), .B2(n11965), .A(n17928), .ZN(n17929) );
  OAI21_X1 U11118 ( .B1(n18009), .B2(n18008), .A(n18007), .ZN(n18010) );
  NOR2_X2 U11119 ( .A1(n19114), .A2(n11932), .ZN(n18012) );
  NOR2_X2 U11120 ( .A1(net231229), .A2(n11969), .ZN(n18013) );
  NOR2_X2 U11121 ( .A1(n14936), .A2(n14935), .ZN(n14937) );
  NOR2_X2 U11122 ( .A1(n13250), .A2(n11491), .ZN(n14936) );
  NOR2_X2 U11123 ( .A1(n13252), .A2(n12613), .ZN(n14935) );
  NOR2_X2 U11124 ( .A1(n13245), .A2(n11483), .ZN(n14605) );
  NOR2_X2 U11125 ( .A1(net231217), .A2(n11981), .ZN(n14603) );
  NOR2_X2 U11126 ( .A1(n14916), .A2(n14915), .ZN(n14917) );
  NOR2_X2 U11127 ( .A1(n13250), .A2(n11489), .ZN(n14916) );
  NOR2_X2 U11128 ( .A1(n13252), .A2(n12611), .ZN(n14915) );
  NOR2_X2 U11129 ( .A1(n13245), .A2(n11481), .ZN(n14583) );
  NOR2_X2 U11130 ( .A1(net231225), .A2(n11936), .ZN(n14581) );
  NOR2_X2 U11131 ( .A1(n14926), .A2(n14925), .ZN(n14927) );
  NOR2_X2 U11132 ( .A1(n13251), .A2(n11490), .ZN(n14926) );
  NOR2_X2 U11133 ( .A1(n13253), .A2(n12612), .ZN(n14925) );
  NOR2_X2 U11134 ( .A1(n13244), .A2(n11482), .ZN(n14594) );
  NOR2_X2 U11135 ( .A1(net231239), .A2(n10819), .ZN(n14592) );
  NOR2_X2 U11136 ( .A1(n14906), .A2(n14905), .ZN(n14907) );
  NOR2_X2 U11137 ( .A1(n13251), .A2(n11488), .ZN(n14906) );
  NOR2_X2 U11138 ( .A1(n13253), .A2(n12610), .ZN(n14905) );
  NOR2_X2 U11139 ( .A1(n13244), .A2(n11480), .ZN(n14572) );
  NOR2_X2 U11140 ( .A1(net231217), .A2(n11933), .ZN(n14570) );
  NOR2_X2 U11141 ( .A1(n14946), .A2(n14945), .ZN(n14947) );
  NOR2_X2 U11142 ( .A1(n13251), .A2(n11492), .ZN(n14946) );
  NOR2_X2 U11143 ( .A1(n13253), .A2(n12614), .ZN(n14945) );
  NOR2_X2 U11144 ( .A1(n13244), .A2(n11484), .ZN(n14616) );
  NOR2_X2 U11145 ( .A1(net231239), .A2(n10823), .ZN(n14614) );
  NOR2_X2 U11146 ( .A1(n14956), .A2(n14955), .ZN(n14957) );
  NOR2_X2 U11147 ( .A1(n13250), .A2(n11493), .ZN(n14956) );
  NOR2_X2 U11148 ( .A1(n13252), .A2(n11584), .ZN(n14955) );
  NOR2_X2 U11149 ( .A1(n13245), .A2(n11485), .ZN(n14627) );
  NOR2_X2 U11150 ( .A1(net231243), .A2(n11937), .ZN(n14625) );
  INV_X4 U11151 ( .A(n10831), .ZN(n13739) );
  INV_X4 U11152 ( .A(net231339), .ZN(net231293) );
  OAI21_X2 U11153 ( .B1(n13217), .B2(n11937), .A(n18546), .ZN(n18553) );
  NOR2_X2 U11154 ( .A1(n18551), .A2(n18550), .ZN(n18552) );
  NAND2_X2 U11155 ( .A1(DMEM_BUS_OUT[30]), .A2(n18927), .ZN(n15702) );
  NOR2_X2 U11156 ( .A1(n14836), .A2(n14835), .ZN(n14837) );
  NOR2_X2 U11157 ( .A1(n13251), .A2(n12370), .ZN(n14836) );
  NOR2_X2 U11158 ( .A1(n13253), .A2(n12249), .ZN(n14835) );
  NOR2_X2 U11159 ( .A1(n13245), .A2(n12339), .ZN(n14495) );
  NOR2_X2 U11160 ( .A1(net231223), .A2(n10814), .ZN(n14493) );
  OAI21_X2 U11161 ( .B1(n19114), .B2(n10814), .A(n18576), .ZN(n18580) );
  NAND4_X2 U11162 ( .A1(n17912), .A2(n17915), .A3(n17913), .A4(n17914), .ZN(
        n18575) );
  OAI21_X2 U11163 ( .B1(n18573), .B2(n13214), .A(n18572), .ZN(n18574) );
  AOI21_X2 U11164 ( .B1(n18675), .B2(DMEM_BUS_OUT[0]), .A(n18674), .ZN(n18676)
         );
  AOI21_X2 U11165 ( .B1(n18673), .B2(n18672), .A(n18671), .ZN(n18674) );
  OAI21_X2 U11166 ( .B1(n18659), .B2(n12035), .A(net231229), .ZN(n18675) );
  NOR2_X2 U11167 ( .A1(n18651), .A2(n18650), .ZN(n18680) );
  NOR3_X1 U11168 ( .A1(n18649), .A2(n19138), .A3(n18648), .ZN(n18650) );
  NOR2_X2 U11170 ( .A1(n13244), .A2(n12321), .ZN(n14296) );
  NOR2_X2 U11171 ( .A1(net231223), .A2(n11960), .ZN(n14294) );
  NOR2_X2 U11172 ( .A1(n4659), .A2(n4660), .ZN(n4640) );
  INV_X4 U11173 ( .A(net231279), .ZN(net231229) );
  INV_X4 U11174 ( .A(net231339), .ZN(net231297) );
  INV_X4 U11175 ( .A(n10832), .ZN(n13740) );
  INV_X4 U11176 ( .A(n10831), .ZN(n13738) );
  OAI21_X2 U11177 ( .B1(n14246), .B2(n14245), .A(n14244), .ZN(n14257) );
  AOI21_X2 U11178 ( .B1(n14236), .B2(n14235), .A(n14234), .ZN(n14248) );
  NOR2_X2 U11179 ( .A1(n14233), .A2(n14232), .ZN(n14234) );
  OAI21_X2 U11180 ( .B1(n14241), .B2(n14240), .A(n12690), .ZN(n18759) );
  NOR2_X2 U11181 ( .A1(n14225), .A2(n14224), .ZN(n14226) );
  OAI21_X1 U11182 ( .B1(n18788), .B2(n18780), .A(IF_ID_OUT[32]), .ZN(n15393)
         );
  NOR2_X2 U11183 ( .A1(n12029), .A2(n12020), .ZN(n5506) );
  INV_X4 U11184 ( .A(net231331), .ZN(net231319) );
  NOR2_X1 U11185 ( .A1(n14209), .A2(n14208), .ZN(n14214) );
  NOR2_X2 U11186 ( .A1(n12134), .A2(n12016), .ZN(n14207) );
  NAND3_X1 U11187 ( .A1(n14238), .A2(n13167), .A3(n11991), .ZN(n18769) );
  OAI21_X2 U11188 ( .B1(offset_26_id[9]), .B2(n15370), .A(n15359), .ZN(n18773)
         );
  NOR2_X1 U11189 ( .A1(n13221), .A2(IF_ID_OUT[35]), .ZN(n18780) );
  NOR2_X2 U11190 ( .A1(n13221), .A2(IF_ID_OUT[36]), .ZN(n14205) );
  INV_X4 U11191 ( .A(net231329), .ZN(net231325) );
  INV_X4 U11192 ( .A(net231279), .ZN(net231235) );
  NOR3_X1 U11193 ( .A1(n14135), .A2(n18872), .A3(n18873), .ZN(n14186) );
  NOR2_X1 U11194 ( .A1(n18559), .A2(n18911), .ZN(n14114) );
  NOR2_X2 U11195 ( .A1(n14025), .A2(n12600), .ZN(n14115) );
  INV_X4 U11196 ( .A(net231273), .ZN(net231251) );
  INV_X8 U11197 ( .A(n11041), .ZN(n13218) );
  NOR2_X2 U11198 ( .A1(n13244), .A2(n11486), .ZN(n14640) );
  NOR2_X2 U11199 ( .A1(net231225), .A2(n10815), .ZN(n14638) );
  AOI222_X1 U11200 ( .A1(DMEM_BUS_OUT[24]), .A2(net231289), .B1(n18292), .B2(
        n18360), .C1(ID_EXEC_OUT[228]), .C2(n13216), .ZN(n18320) );
  OAI21_X2 U11201 ( .B1(n13480), .B2(n18834), .A(n18833), .ZN(n7977) );
  NOR3_X2 U11202 ( .A1(n14528), .A2(n14527), .A3(n14526), .ZN(n4027) );
  NOR2_X2 U11203 ( .A1(n4044), .A2(n4045), .ZN(n4029) );
  NOR3_X2 U11204 ( .A1(n14517), .A2(n14516), .A3(n14515), .ZN(n4056) );
  NOR2_X2 U11205 ( .A1(n4073), .A2(n4074), .ZN(n4058) );
  NOR3_X2 U11206 ( .A1(n14351), .A2(n14350), .A3(n14349), .ZN(n4493) );
  OAI21_X2 U11207 ( .B1(net231245), .B2(n12136), .A(n4685), .ZN(n7900) );
  NOR2_X2 U11208 ( .A1(n18952), .A2(n18951), .ZN(n18955) );
  OAI21_X2 U11209 ( .B1(n13104), .B2(n18941), .A(n18940), .ZN(n18948) );
  NOR2_X1 U11210 ( .A1(n14011), .A2(n18958), .ZN(n18965) );
  NOR2_X1 U11211 ( .A1(n18986), .A2(n18985), .ZN(n18987) );
  NOR2_X1 U11212 ( .A1(n18992), .A2(n18991), .ZN(n18994) );
  NOR2_X2 U11213 ( .A1(n19017), .A2(n19016), .ZN(n19018) );
  NOR2_X2 U11214 ( .A1(IMEM_BUS_IN[3]), .A2(IMEM_BUS_IN[0]), .ZN(n15381) );
  NOR2_X2 U11215 ( .A1(IMEM_BUS_IN[5]), .A2(IMEM_BUS_IN[1]), .ZN(n15380) );
  AOI21_X2 U11216 ( .B1(IMEM_BUS_IN[4]), .B2(n18786), .A(IMEM_BUS_IN[1]), .ZN(
        n15367) );
  NOR2_X2 U11217 ( .A1(IMEM_BUS_IN[3]), .A2(n15366), .ZN(n15368) );
  INV_X8 U11218 ( .A(n18690), .ZN(n13437) );
  INV_X4 U11219 ( .A(n12713), .ZN(n13425) );
  NOR2_X2 U11220 ( .A1(nextPC_ex_out[13]), .A2(nextPC_ex_out[14]), .ZN(
        net227090) );
  NOR2_X2 U11221 ( .A1(nextPC_ex_out[16]), .A2(nextPC_ex_out[17]), .ZN(
        net227104) );
  NOR2_X2 U11222 ( .A1(nextPC_ex_out[18]), .A2(nextPC_ex_out[19]), .ZN(
        net227119) );
  NOR2_X2 U11223 ( .A1(n11920), .A2(net225906), .ZN(net227053) );
  NOR2_X2 U11224 ( .A1(nextPC_ex_out[9]), .A2(nextPC_ex_out[8]), .ZN(net224846) );
  NOR2_X1 U11225 ( .A1(nextPC_ex_out[21]), .A2(net227177), .ZN(net227176) );
  NAND2_X2 U11227 ( .A1(net223444), .A2(nextPC_ex_out[27]), .ZN(net239527) );
  NOR2_X2 U11228 ( .A1(net227243), .A2(net227242), .ZN(net227265) );
  INV_X8 U11229 ( .A(n13429), .ZN(n13426) );
  INV_X4 U11230 ( .A(n13425), .ZN(n13429) );
  NOR3_X2 U11231 ( .A1(n12921), .A2(IMEM_BUS_IN[3]), .A3(n1719), .ZN(n15394)
         );
  INV_X8 U11232 ( .A(n13202), .ZN(n18502) );
  INV_X4 U11233 ( .A(n19161), .ZN(n13504) );
  INV_X4 U11234 ( .A(n10352), .ZN(n13174) );
  OAI21_X1 U11235 ( .B1(n17498), .B2(n17496), .A(n17897), .ZN(n15847) );
  NOR2_X2 U11236 ( .A1(n19092), .A2(net232817), .ZN(n19093) );
  NOR2_X1 U11237 ( .A1(n19089), .A2(net222304), .ZN(n19095) );
  NOR3_X1 U11238 ( .A1(EXEC_MEM_OUT_141), .A2(offset_26_id[0]), .A3(n10828), 
        .ZN(n2531) );
  INV_X4 U11239 ( .A(n14179), .ZN(n13164) );
  NAND2_X2 U11240 ( .A1(n14119), .A2(n14118), .ZN(n14179) );
  INV_X4 U11241 ( .A(n13955), .ZN(n13938) );
  NAND3_X2 U11242 ( .A1(n14047), .A2(n14048), .A3(n14049), .ZN(n15682) );
  AOI22_X2 U11243 ( .A1(MEM_WB_OUT[27]), .A2(n13877), .B1(MEM_WB_OUT[96]), 
        .B2(n14102), .ZN(n14049) );
  NOR2_X2 U11244 ( .A1(n14054), .A2(n14053), .ZN(n14055) );
  NOR2_X2 U11245 ( .A1(n5812), .A2(n13956), .ZN(n5811) );
  NOR2_X2 U11246 ( .A1(n5816), .A2(n13955), .ZN(n5815) );
  NOR2_X2 U11247 ( .A1(n10845), .A2(n10365), .ZN(n5890) );
  NOR2_X2 U11248 ( .A1(n10365), .A2(MEM_WB_OUT[108]), .ZN(n5851) );
  INV_X4 U11249 ( .A(reset), .ZN(n13954) );
  NOR2_X2 U11250 ( .A1(n5662), .A2(n13955), .ZN(n5664) );
  INV_X4 U11251 ( .A(n13955), .ZN(n13936) );
  NOR2_X2 U11252 ( .A1(n19315), .A2(n11916), .ZN(n15354) );
  INV_X4 U11253 ( .A(n13954), .ZN(n13937) );
  NOR2_X2 U11254 ( .A1(n5668), .A2(n13955), .ZN(n5670) );
  NOR2_X2 U11255 ( .A1(n11026), .A2(n13174), .ZN(n14973) );
  NOR2_X2 U11256 ( .A1(n13256), .A2(n11617), .ZN(n14654) );
  NOR2_X2 U11257 ( .A1(n12105), .A2(n13174), .ZN(n14901) );
  NOR2_X2 U11258 ( .A1(n12116), .A2(n13169), .ZN(n14556) );
  NOR2_X2 U11259 ( .A1(n12104), .A2(n13174), .ZN(n14891) );
  NOR2_X2 U11260 ( .A1(n12115), .A2(n13169), .ZN(n14545) );
  NOR2_X2 U11261 ( .A1(n12100), .A2(n13174), .ZN(n14851) );
  NOR2_X2 U11262 ( .A1(n12111), .A2(n13169), .ZN(n14501) );
  NOR2_X2 U11263 ( .A1(n12103), .A2(n13174), .ZN(n14881) );
  NOR2_X2 U11264 ( .A1(n12114), .A2(n13169), .ZN(n14534) );
  NOR2_X2 U11265 ( .A1(n12102), .A2(n13174), .ZN(n14871) );
  NOR2_X2 U11266 ( .A1(n12101), .A2(n13174), .ZN(n14861) );
  NOR2_X2 U11267 ( .A1(nextPC_ex_out[9]), .A2(net224847), .ZN(net227042) );
  NOR2_X2 U11268 ( .A1(n11023), .A2(n13174), .ZN(n14831) );
  NOR2_X2 U11269 ( .A1(n11033), .A2(n13169), .ZN(n14479) );
  NOR2_X2 U11270 ( .A1(n11018), .A2(n13174), .ZN(n14781) );
  NOR2_X2 U11271 ( .A1(n11028), .A2(n13169), .ZN(n14424) );
  NOR2_X2 U11272 ( .A1(n11017), .A2(n13174), .ZN(n14771) );
  NOR2_X2 U11273 ( .A1(n11027), .A2(n13169), .ZN(n14413) );
  NOR2_X2 U11274 ( .A1(n11022), .A2(n13174), .ZN(n14821) );
  NOR2_X2 U11275 ( .A1(n11032), .A2(n13169), .ZN(n14468) );
  OAI21_X2 U11276 ( .B1(EXEC_STAGE_imm26_32[14]), .B2(net227290), .A(net232877), .ZN(net227077) );
  AOI21_X2 U11277 ( .B1(n13196), .B2(REG_FILE_reg_out_22__16_), .A(n16754), 
        .ZN(n16755) );
  NOR2_X2 U11278 ( .A1(n16753), .A2(n13453), .ZN(n16754) );
  INV_X8 U11279 ( .A(n16810), .ZN(n16753) );
  NOR2_X2 U11280 ( .A1(n11995), .A2(n11917), .ZN(n13015) );
  NOR2_X2 U11281 ( .A1(nextPC_ex_out[11]), .A2(nextPC_ex_out[10]), .ZN(n13028)
         );
  INV_X4 U11282 ( .A(n15882), .ZN(n12995) );
  AOI21_X2 U11283 ( .B1(n13196), .B2(REG_FILE_reg_out_22__17_), .A(n17095), 
        .ZN(n17096) );
  NOR2_X2 U11284 ( .A1(n17141), .A2(n13453), .ZN(n17095) );
  NOR3_X2 U11285 ( .A1(n10828), .A2(EXEC_MEM_OUT_141), .A3(n10360), .ZN(n2533)
         );
  NAND2_X2 U11286 ( .A1(n2511), .A2(n14986), .ZN(n1882) );
  AOI21_X2 U11287 ( .B1(n13196), .B2(REG_FILE_reg_out_22__18_), .A(n17364), 
        .ZN(n17365) );
  NOR2_X2 U11288 ( .A1(n18570), .A2(n13453), .ZN(n17364) );
  AOI21_X2 U11289 ( .B1(n13196), .B2(REG_FILE_reg_out_22__19_), .A(n17415), 
        .ZN(n17416) );
  NOR2_X2 U11290 ( .A1(n17905), .A2(n13453), .ZN(n17415) );
  NAND3_X2 U11291 ( .A1(net227164), .A2(n13034), .A3(nextPC_ex_out[21]), .ZN(
        n13038) );
  INV_X4 U11292 ( .A(n13172), .ZN(n14760) );
  INV_X4 U11293 ( .A(n13504), .ZN(n13501) );
  NOR2_X2 U11294 ( .A1(n11019), .A2(n13174), .ZN(n14791) );
  NOR2_X2 U11295 ( .A1(n11029), .A2(n13169), .ZN(n14435) );
  NOR2_X2 U11296 ( .A1(n15860), .A2(n15859), .ZN(n15861) );
  NOR2_X2 U11297 ( .A1(n17681), .A2(n13452), .ZN(n17655) );
  NOR2_X2 U11298 ( .A1(n17632), .A2(n17631), .ZN(n17637) );
  NOR2_X2 U11299 ( .A1(n13421), .A2(n12468), .ZN(n17632) );
  NOR2_X2 U11300 ( .A1(n13424), .A2(n12899), .ZN(n17631) );
  NOR2_X2 U11301 ( .A1(n17634), .A2(n17633), .ZN(n17635) );
  NOR2_X2 U11302 ( .A1(n13426), .A2(n12470), .ZN(n17633) );
  NOR2_X2 U11303 ( .A1(n13431), .A2(n12469), .ZN(n17634) );
  NOR2_X2 U11304 ( .A1(n11020), .A2(n13174), .ZN(n14801) );
  NOR2_X2 U11305 ( .A1(n11030), .A2(n13169), .ZN(n14446) );
  NOR2_X2 U11306 ( .A1(n17785), .A2(n17784), .ZN(n17790) );
  NOR2_X2 U11307 ( .A1(n13421), .A2(n12471), .ZN(n17785) );
  NOR2_X2 U11308 ( .A1(n13423), .A2(n12901), .ZN(n17784) );
  NOR2_X2 U11309 ( .A1(n17787), .A2(n17786), .ZN(n17788) );
  NOR2_X2 U11310 ( .A1(n13426), .A2(n12473), .ZN(n17786) );
  NOR2_X2 U11311 ( .A1(n13431), .A2(n12472), .ZN(n17787) );
  AOI21_X2 U11312 ( .B1(n13196), .B2(REG_FILE_reg_out_22__22_), .A(n17809), 
        .ZN(n17810) );
  NOR2_X2 U11313 ( .A1(n17808), .A2(n13452), .ZN(n17809) );
  NOR2_X2 U11314 ( .A1(n11021), .A2(n13174), .ZN(n14811) );
  NOR2_X2 U11315 ( .A1(n11031), .A2(n13169), .ZN(n14457) );
  NAND2_X2 U11316 ( .A1(n17683), .A2(n18641), .ZN(n17685) );
  NOR2_X2 U11317 ( .A1(n17957), .A2(n13452), .ZN(n17958) );
  NOR2_X2 U11318 ( .A1(n17934), .A2(n17933), .ZN(n17939) );
  NOR2_X2 U11319 ( .A1(n13421), .A2(n12474), .ZN(n17934) );
  NOR2_X2 U11320 ( .A1(n13424), .A2(n12903), .ZN(n17933) );
  NOR2_X2 U11321 ( .A1(n17936), .A2(n17935), .ZN(n17937) );
  NOR2_X2 U11322 ( .A1(n13426), .A2(n12476), .ZN(n17935) );
  NOR2_X2 U11323 ( .A1(n13431), .A2(n12475), .ZN(n17936) );
  NOR2_X2 U11324 ( .A1(n14074), .A2(n14077), .ZN(n14065) );
  NOR2_X2 U11325 ( .A1(n12109), .A2(n13174), .ZN(n14941) );
  NOR2_X2 U11326 ( .A1(n12120), .A2(n13169), .ZN(n14600) );
  NOR2_X2 U11327 ( .A1(n18047), .A2(n13452), .ZN(n18048) );
  NOR2_X2 U11328 ( .A1(n18024), .A2(n18023), .ZN(n18029) );
  NOR2_X2 U11329 ( .A1(n13421), .A2(n12477), .ZN(n18024) );
  NOR2_X2 U11330 ( .A1(n13423), .A2(n12905), .ZN(n18023) );
  NOR2_X2 U11331 ( .A1(n18026), .A2(n18025), .ZN(n18027) );
  NOR2_X2 U11332 ( .A1(n13426), .A2(n12479), .ZN(n18025) );
  NOR2_X2 U11333 ( .A1(n13431), .A2(n12478), .ZN(n18026) );
  NOR2_X2 U11334 ( .A1(n18090), .A2(n13452), .ZN(n18091) );
  NOR2_X2 U11335 ( .A1(n18067), .A2(n18066), .ZN(n18072) );
  NOR2_X2 U11336 ( .A1(n13421), .A2(n12480), .ZN(n18067) );
  NOR2_X2 U11337 ( .A1(n13424), .A2(n12907), .ZN(n18066) );
  NOR2_X2 U11338 ( .A1(n18069), .A2(n18068), .ZN(n18070) );
  NOR2_X2 U11339 ( .A1(n13426), .A2(n12482), .ZN(n18068) );
  NOR2_X2 U11340 ( .A1(n13431), .A2(n12481), .ZN(n18069) );
  NOR2_X2 U11341 ( .A1(n18135), .A2(n13452), .ZN(n18136) );
  NOR2_X2 U11342 ( .A1(n18112), .A2(n18111), .ZN(n18117) );
  NOR2_X2 U11343 ( .A1(n13421), .A2(n12483), .ZN(n18112) );
  NOR2_X2 U11344 ( .A1(n13423), .A2(n12909), .ZN(n18111) );
  NOR2_X2 U11345 ( .A1(n18114), .A2(n18113), .ZN(n18115) );
  NOR2_X2 U11346 ( .A1(n13426), .A2(n12485), .ZN(n18113) );
  NOR2_X2 U11347 ( .A1(n13431), .A2(n12484), .ZN(n18114) );
  NOR2_X2 U11348 ( .A1(n18176), .A2(n13452), .ZN(n18177) );
  NOR2_X2 U11349 ( .A1(n18153), .A2(n18152), .ZN(n18158) );
  NOR2_X2 U11350 ( .A1(n13421), .A2(n12486), .ZN(n18153) );
  NOR2_X2 U11351 ( .A1(n13424), .A2(n12911), .ZN(n18152) );
  NOR2_X2 U11352 ( .A1(n18155), .A2(n18154), .ZN(n18156) );
  NOR2_X2 U11353 ( .A1(n13426), .A2(n12488), .ZN(n18154) );
  NOR2_X2 U11354 ( .A1(n13431), .A2(n12487), .ZN(n18155) );
  NOR2_X2 U11355 ( .A1(n18221), .A2(n13452), .ZN(n18222) );
  NOR2_X2 U11356 ( .A1(n18198), .A2(n18197), .ZN(n18203) );
  NOR2_X2 U11357 ( .A1(n13421), .A2(n12489), .ZN(n18198) );
  NOR2_X2 U11358 ( .A1(n13424), .A2(n12913), .ZN(n18197) );
  NOR2_X2 U11359 ( .A1(n18200), .A2(n18199), .ZN(n18201) );
  NOR2_X2 U11360 ( .A1(n13426), .A2(n12491), .ZN(n18199) );
  NOR2_X2 U11361 ( .A1(n13431), .A2(n12490), .ZN(n18200) );
  NOR2_X2 U11362 ( .A1(n12107), .A2(n13174), .ZN(n14921) );
  NOR2_X2 U11363 ( .A1(n12118), .A2(n13169), .ZN(n14578) );
  NOR2_X2 U11364 ( .A1(n12108), .A2(n13174), .ZN(n14931) );
  NOR2_X2 U11365 ( .A1(n12119), .A2(n13169), .ZN(n14589) );
  NAND2_X1 U11366 ( .A1(n10160), .A2(n15603), .ZN(n14972) );
  NOR2_X2 U11367 ( .A1(n12106), .A2(n13174), .ZN(n14911) );
  NOR2_X2 U11368 ( .A1(n12117), .A2(n13169), .ZN(n14567) );
  INV_X4 U11369 ( .A(n11905), .ZN(n13509) );
  NAND2_X1 U11370 ( .A1(n10160), .A2(n15603), .ZN(n13172) );
  NOR2_X2 U11371 ( .A1(n12110), .A2(n13174), .ZN(n14951) );
  NOR2_X2 U11372 ( .A1(n12121), .A2(n13169), .ZN(n14611) );
  NOR2_X2 U11373 ( .A1(n18429), .A2(n13452), .ZN(n18430) );
  NOR2_X2 U11374 ( .A1(n18406), .A2(n18405), .ZN(n18411) );
  NOR2_X2 U11375 ( .A1(n13421), .A2(n12492), .ZN(n18406) );
  NOR2_X2 U11376 ( .A1(n13423), .A2(n12915), .ZN(n18405) );
  NOR2_X2 U11377 ( .A1(n18408), .A2(n18407), .ZN(n18409) );
  NOR2_X2 U11378 ( .A1(n13426), .A2(n12494), .ZN(n18407) );
  NOR2_X2 U11379 ( .A1(n13431), .A2(n12493), .ZN(n18408) );
  INV_X4 U11380 ( .A(n13504), .ZN(n13503) );
  INV_X4 U11381 ( .A(n10835), .ZN(n13260) );
  INV_X4 U11382 ( .A(n10836), .ZN(n13258) );
  NOR2_X2 U11383 ( .A1(n11025), .A2(n13174), .ZN(n14961) );
  INV_X4 U11384 ( .A(n11832), .ZN(n13262) );
  NOR2_X2 U11385 ( .A1(n11035), .A2(n13169), .ZN(n14622) );
  INV_X4 U11386 ( .A(n13193), .ZN(n18493) );
  NOR2_X2 U11387 ( .A1(n18510), .A2(n13452), .ZN(n18511) );
  NAND2_X1 U11388 ( .A1(n15610), .A2(n15609), .ZN(n18727) );
  NAND2_X2 U11389 ( .A1(n15608), .A2(n15613), .ZN(n18726) );
  NOR2_X2 U11390 ( .A1(n18486), .A2(n18485), .ZN(n18487) );
  NOR2_X2 U11391 ( .A1(n13431), .A2(n12496), .ZN(n18486) );
  NOR2_X2 U11392 ( .A1(n18484), .A2(n18483), .ZN(n18489) );
  NOR2_X2 U11393 ( .A1(n13421), .A2(n12495), .ZN(n18484) );
  NOR2_X2 U11394 ( .A1(n13424), .A2(n12917), .ZN(n18483) );
  NAND3_X2 U11395 ( .A1(n18249), .A2(n18248), .A3(n18247), .ZN(n18539) );
  INV_X8 U11396 ( .A(n18928), .ZN(n13090) );
  INV_X4 U11397 ( .A(n13504), .ZN(n13502) );
  INV_X4 U11398 ( .A(n13257), .ZN(n13256) );
  INV_X4 U11399 ( .A(n10835), .ZN(n13261) );
  INV_X4 U11400 ( .A(n10836), .ZN(n13259) );
  INV_X4 U11401 ( .A(n11905), .ZN(n13510) );
  NAND2_X1 U11402 ( .A1(n10160), .A2(n15603), .ZN(n13173) );
  NOR2_X2 U11403 ( .A1(n11024), .A2(n13174), .ZN(n14841) );
  INV_X4 U11404 ( .A(n11832), .ZN(n13263) );
  NOR2_X2 U11405 ( .A1(n11034), .A2(n13169), .ZN(n14490) );
  AOI21_X2 U11406 ( .B1(n18606), .B2(n18605), .A(n18616), .ZN(n18607) );
  OAI21_X2 U11407 ( .B1(n19318), .B2(n15508), .A(net230387), .ZN(n15505) );
  INV_X4 U11408 ( .A(n13454), .ZN(n13452) );
  INV_X4 U11409 ( .A(n13457), .ZN(n13455) );
  INV_X4 U11410 ( .A(n13200), .ZN(n13201) );
  INV_X4 U11411 ( .A(n13198), .ZN(n13199) );
  INV_X4 U11412 ( .A(n10834), .ZN(n13474) );
  INV_X4 U11413 ( .A(n10833), .ZN(n13470) );
  INV_X4 U11414 ( .A(n13469), .ZN(n13468) );
  NOR2_X2 U11415 ( .A1(n13021), .A2(net222531), .ZN(net222353) );
  NAND2_X1 U11416 ( .A1(n14288), .A2(n14998), .ZN(n14633) );
  NOR2_X2 U11417 ( .A1(n11036), .A2(n13169), .ZN(n14635) );
  NAND3_X2 U11418 ( .A1(n16773), .A2(n16795), .A3(n16772), .ZN(n17697) );
  NAND3_X2 U11419 ( .A1(n17514), .A2(n17993), .A3(n17513), .ZN(n18338) );
  NOR2_X2 U11420 ( .A1(n19089), .A2(net232817), .ZN(n17989) );
  INV_X4 U11422 ( .A(n13940), .ZN(n13939) );
  NAND2_X2 U11423 ( .A1(n5909), .A2(n10817), .ZN(n5812) );
  INV_X4 U11424 ( .A(n13954), .ZN(n13933) );
  NAND3_X2 U11425 ( .A1(MEM_WB_OUT[109]), .A2(MEM_WB_OUT[110]), .A3(n5851), 
        .ZN(n5770) );
  NAND3_X2 U11426 ( .A1(n10802), .A2(n10353), .A3(n5890), .ZN(n5764) );
  NAND3_X2 U11427 ( .A1(n10802), .A2(n10353), .A3(n5851), .ZN(n5676) );
  NAND3_X2 U11428 ( .A1(MEM_WB_OUT[110]), .A2(n10802), .A3(n5890), .ZN(n5724)
         );
  NAND3_X2 U11429 ( .A1(MEM_WB_OUT[109]), .A2(n10353), .A3(n5890), .ZN(n5718)
         );
  NAND3_X2 U11430 ( .A1(MEM_WB_OUT[109]), .A2(MEM_WB_OUT[110]), .A3(n5890), 
        .ZN(n5680) );
  INV_X4 U11431 ( .A(n13953), .ZN(n13934) );
  NAND3_X2 U11432 ( .A1(MEM_WB_OUT[110]), .A2(n10802), .A3(n5851), .ZN(n5669)
         );
  NAND3_X2 U11433 ( .A1(MEM_WB_OUT[109]), .A2(n10353), .A3(n5851), .ZN(n5663)
         );
  INV_X4 U11434 ( .A(n13954), .ZN(n13935) );
  NOR2_X1 U11435 ( .A1(n19317), .A2(n19320), .ZN(n164) );
  NOR3_X2 U11436 ( .A1(n14971), .A2(n14970), .A3(n14969), .ZN(n2598) );
  NOR2_X2 U11437 ( .A1(n13259), .A2(n11673), .ZN(n14970) );
  NOR2_X2 U11438 ( .A1(n13261), .A2(n11496), .ZN(n14969) );
  NOR2_X2 U11439 ( .A1(n13256), .A2(n11641), .ZN(n14971) );
  NOR3_X2 U11440 ( .A1(n14900), .A2(n14899), .A3(n14898), .ZN(n2854) );
  NOR2_X2 U11441 ( .A1(n13258), .A2(n11665), .ZN(n14898) );
  NOR2_X2 U11442 ( .A1(n13260), .A2(n12073), .ZN(n14899) );
  NOR2_X2 U11443 ( .A1(n13256), .A2(n11633), .ZN(n14900) );
  NOR3_X2 U11444 ( .A1(n14890), .A2(n14889), .A3(n14888), .ZN(n2889) );
  NOR2_X2 U11445 ( .A1(n13259), .A2(n11664), .ZN(n14888) );
  NOR2_X2 U11446 ( .A1(n13261), .A2(n12381), .ZN(n14889) );
  NOR2_X2 U11447 ( .A1(n13256), .A2(n11632), .ZN(n14890) );
  NOR3_X2 U11448 ( .A1(n14850), .A2(n14849), .A3(n14848), .ZN(n3025) );
  NOR2_X2 U11449 ( .A1(n13259), .A2(n11659), .ZN(n14848) );
  NOR2_X2 U11450 ( .A1(n13261), .A2(n12373), .ZN(n14849) );
  NOR2_X2 U11451 ( .A1(n13256), .A2(n11627), .ZN(n14850) );
  NOR3_X2 U11452 ( .A1(n14880), .A2(n14879), .A3(n14878), .ZN(n2923) );
  NOR2_X2 U11453 ( .A1(n13259), .A2(n11663), .ZN(n14878) );
  NOR2_X2 U11454 ( .A1(n13261), .A2(n12379), .ZN(n14879) );
  NOR2_X2 U11455 ( .A1(n13256), .A2(n11631), .ZN(n14880) );
  NOR3_X2 U11456 ( .A1(n14870), .A2(n14869), .A3(n14868), .ZN(n2957) );
  NOR2_X2 U11457 ( .A1(n13259), .A2(n11662), .ZN(n14868) );
  NOR2_X2 U11458 ( .A1(n13261), .A2(n12377), .ZN(n14869) );
  NOR2_X2 U11459 ( .A1(n13256), .A2(n11630), .ZN(n14870) );
  NOR2_X2 U11460 ( .A1(n14523), .A2(n14522), .ZN(n14524) );
  NOR2_X2 U11461 ( .A1(n12377), .A2(n13171), .ZN(n14522) );
  NOR3_X2 U11462 ( .A1(n14860), .A2(n14859), .A3(n14858), .ZN(n2991) );
  NOR2_X2 U11463 ( .A1(n13259), .A2(n11661), .ZN(n14858) );
  NOR2_X2 U11464 ( .A1(n13261), .A2(n12375), .ZN(n14859) );
  NOR2_X2 U11465 ( .A1(n13256), .A2(n11629), .ZN(n14860) );
  NOR2_X2 U11466 ( .A1(n14512), .A2(n14511), .ZN(n14513) );
  NOR2_X2 U11467 ( .A1(n12375), .A2(n13170), .ZN(n14511) );
  NOR3_X2 U11468 ( .A1(n14699), .A2(n14698), .A3(n14697), .ZN(n3536) );
  NOR2_X2 U11469 ( .A1(n14968), .A2(n11643), .ZN(n14699) );
  NOR2_X2 U11470 ( .A1(n13258), .A2(n11675), .ZN(n14697) );
  NOR2_X2 U11471 ( .A1(n13260), .A2(n11686), .ZN(n14698) );
  NOR3_X2 U11472 ( .A1(n15600), .A2(n15599), .A3(n15598), .ZN(n15607) );
  NOR2_X1 U11473 ( .A1(n18662), .A2(n13453), .ZN(n15599) );
  NOR2_X2 U11474 ( .A1(n10861), .A2(n13197), .ZN(n15598) );
  NOR2_X2 U11475 ( .A1(n10959), .A2(n13195), .ZN(n15600) );
  NOR2_X2 U11476 ( .A1(n15602), .A2(n15601), .ZN(n15605) );
  NOR2_X2 U11477 ( .A1(n13458), .A2(n12413), .ZN(n15602) );
  NOR2_X2 U11478 ( .A1(n13461), .A2(n12828), .ZN(n15601) );
  NOR3_X2 U11479 ( .A1(n15590), .A2(n15589), .A3(n15588), .ZN(n15594) );
  NOR3_X2 U11480 ( .A1(n15587), .A2(n15586), .A3(n15585), .ZN(n15596) );
  NOR2_X2 U11481 ( .A1(n15592), .A2(n15591), .ZN(n15593) );
  NOR2_X2 U11482 ( .A1(n10958), .A2(n13447), .ZN(n15592) );
  NOR2_X2 U11483 ( .A1(n12767), .A2(n13450), .ZN(n15591) );
  NOR2_X2 U11484 ( .A1(n15615), .A2(n15614), .ZN(n15626) );
  NOR2_X2 U11485 ( .A1(n10245), .A2(n13202), .ZN(n15615) );
  NOR2_X2 U11486 ( .A1(n10949), .A2(n13204), .ZN(n15614) );
  NOR2_X2 U11487 ( .A1(n15612), .A2(n15611), .ZN(n15627) );
  NOR2_X2 U11488 ( .A1(n11881), .A2(n13199), .ZN(n15612) );
  NOR2_X2 U11489 ( .A1(n10371), .A2(n13201), .ZN(n15611) );
  NOR2_X2 U11490 ( .A1(n15623), .A2(n15622), .ZN(n15624) );
  NOR2_X2 U11491 ( .A1(n10871), .A2(n13474), .ZN(n15622) );
  NOR2_X2 U11492 ( .A1(n10870), .A2(n13473), .ZN(n15623) );
  NOR2_X2 U11493 ( .A1(n15619), .A2(n15618), .ZN(n15625) );
  NOR2_X2 U11494 ( .A1(n10869), .A2(n13468), .ZN(n15619) );
  NOR2_X2 U11495 ( .A1(n12937), .A2(n13470), .ZN(n15618) );
  NOR2_X2 U11496 ( .A1(nextPC_ex_out[5]), .A2(nextPC_ex_out[4]), .ZN(net226995) );
  NOR2_X2 U11497 ( .A1(nextPC_ex_out[3]), .A2(nextPC_ex_out[2]), .ZN(n15570)
         );
  OAI21_X1 U11498 ( .B1(n19076), .B2(n13491), .A(n15748), .ZN(n15750) );
  NOR2_X2 U11499 ( .A1(n19114), .A2(n11939), .ZN(n15749) );
  NOR2_X2 U11500 ( .A1(n18678), .A2(n13213), .ZN(n15727) );
  NOR3_X2 U11501 ( .A1(n14830), .A2(n14829), .A3(n14828), .ZN(n3093) );
  NOR2_X2 U11502 ( .A1(n13259), .A2(n11657), .ZN(n14828) );
  NOR2_X2 U11503 ( .A1(n13261), .A2(n12369), .ZN(n14829) );
  NOR2_X2 U11504 ( .A1(n13256), .A2(n11625), .ZN(n14830) );
  NOR3_X2 U11505 ( .A1(n14749), .A2(n14748), .A3(n14747), .ZN(n3366) );
  NOR2_X2 U11506 ( .A1(n13258), .A2(n11680), .ZN(n14747) );
  NOR2_X2 U11507 ( .A1(n13260), .A2(n11691), .ZN(n14748) );
  NOR2_X2 U11508 ( .A1(n13256), .A2(n11648), .ZN(n14749) );
  NOR3_X2 U11509 ( .A1(n14780), .A2(n14779), .A3(n14778), .ZN(n3264) );
  NOR2_X2 U11510 ( .A1(n13259), .A2(n11652), .ZN(n14778) );
  NOR2_X2 U11511 ( .A1(n13261), .A2(n12359), .ZN(n14779) );
  NOR2_X2 U11512 ( .A1(n13256), .A2(n11620), .ZN(n14780) );
  NOR3_X2 U11513 ( .A1(n14719), .A2(n14718), .A3(n14717), .ZN(n3468) );
  NOR2_X2 U11514 ( .A1(n13258), .A2(n11677), .ZN(n14717) );
  NOR2_X2 U11515 ( .A1(n13260), .A2(n11688), .ZN(n14718) );
  NOR2_X2 U11516 ( .A1(n13256), .A2(n11645), .ZN(n14719) );
  NOR3_X2 U11517 ( .A1(n14709), .A2(n14708), .A3(n14707), .ZN(n3502) );
  NOR2_X2 U11518 ( .A1(n13258), .A2(n11676), .ZN(n14707) );
  NOR2_X2 U11519 ( .A1(n13260), .A2(n11687), .ZN(n14708) );
  NOR2_X2 U11520 ( .A1(n13256), .A2(n11644), .ZN(n14709) );
  NOR3_X2 U11521 ( .A1(n15981), .A2(n15980), .A3(n15979), .ZN(n15987) );
  NOR2_X2 U11522 ( .A1(n15978), .A2(n13453), .ZN(n15980) );
  NOR2_X2 U11523 ( .A1(n10862), .A2(n13197), .ZN(n15979) );
  NOR2_X2 U11524 ( .A1(n10983), .A2(n13195), .ZN(n15981) );
  NOR2_X2 U11525 ( .A1(n15983), .A2(n15982), .ZN(n15985) );
  NOR2_X2 U11526 ( .A1(n13460), .A2(n12832), .ZN(n15982) );
  NOR2_X2 U11527 ( .A1(n13458), .A2(n12414), .ZN(n15983) );
  NOR2_X2 U11528 ( .A1(n15991), .A2(n15990), .ZN(n15998) );
  NOR2_X2 U11529 ( .A1(n10250), .A2(n13202), .ZN(n15991) );
  NOR2_X2 U11530 ( .A1(n10968), .A2(n13204), .ZN(n15990) );
  NOR2_X2 U11531 ( .A1(n15989), .A2(n15988), .ZN(n15999) );
  NOR2_X2 U11532 ( .A1(n11884), .A2(n13199), .ZN(n15989) );
  NOR2_X2 U11533 ( .A1(n10385), .A2(n13201), .ZN(n15988) );
  NOR2_X2 U11534 ( .A1(n15995), .A2(n15994), .ZN(n15996) );
  NOR2_X2 U11535 ( .A1(n10882), .A2(n13474), .ZN(n15994) );
  NOR2_X2 U11536 ( .A1(n10881), .A2(n13473), .ZN(n15995) );
  NOR2_X2 U11537 ( .A1(n15993), .A2(n15992), .ZN(n15997) );
  NOR2_X2 U11538 ( .A1(n10880), .A2(n13468), .ZN(n15993) );
  NOR2_X2 U11539 ( .A1(n12940), .A2(n13470), .ZN(n15992) );
  NOR3_X2 U11540 ( .A1(n15971), .A2(n15970), .A3(n15969), .ZN(n15975) );
  NOR3_X2 U11541 ( .A1(n15968), .A2(n15967), .A3(n15966), .ZN(n15977) );
  NOR2_X2 U11542 ( .A1(n15973), .A2(n15972), .ZN(n15974) );
  NOR2_X2 U11543 ( .A1(n10982), .A2(n13447), .ZN(n15973) );
  NOR2_X2 U11544 ( .A1(n12770), .A2(n13450), .ZN(n15972) );
  NOR3_X2 U11545 ( .A1(n16104), .A2(n16103), .A3(n16102), .ZN(n16110) );
  NOR2_X2 U11546 ( .A1(n16130), .A2(n13453), .ZN(n16103) );
  NOR2_X2 U11547 ( .A1(n10857), .A2(n13197), .ZN(n16102) );
  NOR2_X2 U11548 ( .A1(n10985), .A2(n13195), .ZN(n16104) );
  NOR2_X2 U11549 ( .A1(n16106), .A2(n16105), .ZN(n16108) );
  NOR2_X2 U11550 ( .A1(n13458), .A2(n12415), .ZN(n16106) );
  NOR2_X2 U11551 ( .A1(n13461), .A2(n12836), .ZN(n16105) );
  NOR2_X2 U11552 ( .A1(n16114), .A2(n16113), .ZN(n16121) );
  NOR2_X2 U11553 ( .A1(n10372), .A2(n13202), .ZN(n16114) );
  NOR2_X2 U11554 ( .A1(n10969), .A2(n13204), .ZN(n16113) );
  NOR2_X2 U11555 ( .A1(n16112), .A2(n16111), .ZN(n16122) );
  NOR2_X2 U11556 ( .A1(n12418), .A2(n13199), .ZN(n16112) );
  NOR2_X2 U11557 ( .A1(n10848), .A2(n13201), .ZN(n16111) );
  NOR2_X2 U11558 ( .A1(n16118), .A2(n16117), .ZN(n16119) );
  NOR2_X2 U11559 ( .A1(n10885), .A2(n13474), .ZN(n16117) );
  NOR2_X2 U11560 ( .A1(n10884), .A2(n13473), .ZN(n16118) );
  NOR2_X2 U11561 ( .A1(n16116), .A2(n16115), .ZN(n16120) );
  NOR2_X2 U11562 ( .A1(n10883), .A2(n13468), .ZN(n16116) );
  NOR2_X2 U11563 ( .A1(n12945), .A2(n13470), .ZN(n16115) );
  NOR3_X2 U11564 ( .A1(n16095), .A2(n16094), .A3(n16093), .ZN(n16099) );
  NOR3_X2 U11565 ( .A1(n16092), .A2(n16091), .A3(n16090), .ZN(n16101) );
  NOR2_X2 U11566 ( .A1(n16097), .A2(n16096), .ZN(n16098) );
  NOR2_X2 U11567 ( .A1(n10984), .A2(n13447), .ZN(n16097) );
  NOR2_X2 U11568 ( .A1(n12746), .A2(n13450), .ZN(n16096) );
  AOI21_X2 U11569 ( .B1(n13378), .B2(REG_FILE_reg_out_9__6_), .A(n16131), .ZN(
        n16132) );
  NOR2_X2 U11570 ( .A1(n16130), .A2(n13362), .ZN(n16131) );
  NOR2_X2 U11571 ( .A1(n13281), .A2(n11588), .ZN(n15067) );
  NOR2_X2 U11572 ( .A1(n12629), .A2(n13279), .ZN(n15066) );
  NOR3_X2 U11573 ( .A1(n14739), .A2(n14738), .A3(n14737), .ZN(n3400) );
  NOR2_X2 U11574 ( .A1(n13258), .A2(n11679), .ZN(n14737) );
  NOR2_X2 U11575 ( .A1(n13260), .A2(n11690), .ZN(n14738) );
  NOR2_X2 U11576 ( .A1(n13256), .A2(n11647), .ZN(n14739) );
  NOR3_X2 U11577 ( .A1(n16179), .A2(n16178), .A3(n16177), .ZN(n16185) );
  NOR2_X2 U11578 ( .A1(n16176), .A2(n13453), .ZN(n16178) );
  NOR2_X2 U11579 ( .A1(n10863), .A2(n13197), .ZN(n16177) );
  NOR2_X2 U11580 ( .A1(n10987), .A2(n13195), .ZN(n16179) );
  NOR2_X2 U11581 ( .A1(n16181), .A2(n16180), .ZN(n16183) );
  NOR2_X2 U11582 ( .A1(n13458), .A2(n12419), .ZN(n16181) );
  NOR2_X2 U11583 ( .A1(n13461), .A2(n12840), .ZN(n16180) );
  NOR2_X2 U11584 ( .A1(n16189), .A2(n16188), .ZN(n16196) );
  NOR2_X2 U11585 ( .A1(n10374), .A2(n13202), .ZN(n16189) );
  NOR2_X2 U11586 ( .A1(n10970), .A2(n13204), .ZN(n16188) );
  NOR2_X2 U11587 ( .A1(n16187), .A2(n16186), .ZN(n16197) );
  NOR2_X2 U11588 ( .A1(n11886), .A2(n13199), .ZN(n16187) );
  NOR2_X2 U11589 ( .A1(n10850), .A2(n13201), .ZN(n16186) );
  NOR2_X2 U11590 ( .A1(n16193), .A2(n16192), .ZN(n16194) );
  NOR2_X2 U11591 ( .A1(n10891), .A2(n13474), .ZN(n16192) );
  NOR2_X2 U11592 ( .A1(n10890), .A2(n13473), .ZN(n16193) );
  NOR2_X2 U11593 ( .A1(n16191), .A2(n16190), .ZN(n16195) );
  NOR2_X2 U11594 ( .A1(n10889), .A2(n13468), .ZN(n16191) );
  NOR2_X2 U11595 ( .A1(n12942), .A2(n13470), .ZN(n16190) );
  NOR3_X2 U11596 ( .A1(n16169), .A2(n16168), .A3(n16167), .ZN(n16173) );
  NOR3_X2 U11597 ( .A1(n16166), .A2(n16165), .A3(n16164), .ZN(n16175) );
  NOR2_X2 U11598 ( .A1(n16171), .A2(n16170), .ZN(n16172) );
  NOR2_X2 U11599 ( .A1(n10986), .A2(n13447), .ZN(n16171) );
  NOR2_X2 U11600 ( .A1(n12772), .A2(n13450), .ZN(n16170) );
  NOR3_X2 U11601 ( .A1(n14759), .A2(n14758), .A3(n14757), .ZN(n3332) );
  NOR2_X2 U11602 ( .A1(n13258), .A2(n11650), .ZN(n14757) );
  NOR2_X2 U11603 ( .A1(n13260), .A2(n11682), .ZN(n14758) );
  NOR2_X2 U11604 ( .A1(n13256), .A2(n11618), .ZN(n14759) );
  NOR3_X2 U11605 ( .A1(n16253), .A2(n16252), .A3(n16251), .ZN(n16259) );
  NOR2_X2 U11606 ( .A1(n16279), .A2(n13453), .ZN(n16252) );
  NOR2_X2 U11607 ( .A1(n10858), .A2(n13197), .ZN(n16251) );
  NOR2_X2 U11608 ( .A1(n10989), .A2(n13195), .ZN(n16253) );
  NOR2_X2 U11609 ( .A1(n16255), .A2(n16254), .ZN(n16257) );
  NOR2_X2 U11610 ( .A1(n13458), .A2(n12420), .ZN(n16255) );
  NOR2_X2 U11611 ( .A1(n13461), .A2(n12844), .ZN(n16254) );
  NOR2_X2 U11612 ( .A1(n16263), .A2(n16262), .ZN(n16270) );
  NOR2_X2 U11613 ( .A1(n10376), .A2(n13202), .ZN(n16263) );
  NOR2_X2 U11614 ( .A1(n10971), .A2(n13204), .ZN(n16262) );
  NOR2_X2 U11615 ( .A1(n16261), .A2(n16260), .ZN(n16271) );
  NOR2_X2 U11616 ( .A1(n12423), .A2(n13199), .ZN(n16261) );
  NOR2_X2 U11617 ( .A1(n10852), .A2(n13201), .ZN(n16260) );
  NOR2_X2 U11618 ( .A1(n16267), .A2(n16266), .ZN(n16268) );
  NOR2_X2 U11619 ( .A1(n10895), .A2(n13474), .ZN(n16266) );
  NOR2_X2 U11620 ( .A1(n10894), .A2(n13473), .ZN(n16267) );
  NOR2_X2 U11621 ( .A1(n16265), .A2(n16264), .ZN(n16269) );
  NOR2_X2 U11622 ( .A1(n10391), .A2(n13468), .ZN(n16265) );
  NOR2_X2 U11623 ( .A1(n12946), .A2(n13470), .ZN(n16264) );
  NOR3_X2 U11624 ( .A1(n16244), .A2(n16243), .A3(n16242), .ZN(n16248) );
  NOR3_X2 U11625 ( .A1(n16241), .A2(n16240), .A3(n16239), .ZN(n16250) );
  NOR2_X2 U11626 ( .A1(n16246), .A2(n16245), .ZN(n16247) );
  NOR2_X2 U11627 ( .A1(n10988), .A2(n13447), .ZN(n16246) );
  NOR2_X2 U11628 ( .A1(n12747), .A2(n13450), .ZN(n16245) );
  AOI21_X2 U11629 ( .B1(n13378), .B2(REG_FILE_reg_out_9__10_), .A(n16280), 
        .ZN(n16281) );
  NOR2_X2 U11630 ( .A1(n16279), .A2(n13362), .ZN(n16280) );
  NOR2_X2 U11631 ( .A1(n13281), .A2(n11590), .ZN(n15109) );
  NOR2_X2 U11632 ( .A1(n12631), .A2(n13279), .ZN(n15108) );
  NOR3_X2 U11633 ( .A1(n14770), .A2(n14769), .A3(n14768), .ZN(n3298) );
  NOR2_X2 U11634 ( .A1(n13258), .A2(n11651), .ZN(n14768) );
  NOR2_X2 U11635 ( .A1(n13260), .A2(n12357), .ZN(n14769) );
  NOR2_X2 U11636 ( .A1(n13256), .A2(n11619), .ZN(n14770) );
  NOR3_X2 U11637 ( .A1(n16353), .A2(n16352), .A3(n16351), .ZN(n16359) );
  NOR2_X2 U11638 ( .A1(n16413), .A2(n13453), .ZN(n16352) );
  NOR2_X2 U11639 ( .A1(n10859), .A2(n13197), .ZN(n16351) );
  NOR2_X2 U11640 ( .A1(n10991), .A2(n13195), .ZN(n16353) );
  NOR2_X2 U11641 ( .A1(n16355), .A2(n16354), .ZN(n16357) );
  NOR2_X2 U11642 ( .A1(n13458), .A2(n12424), .ZN(n16355) );
  NOR2_X2 U11643 ( .A1(n13461), .A2(n12848), .ZN(n16354) );
  NOR2_X2 U11644 ( .A1(n16363), .A2(n16362), .ZN(n16370) );
  NOR2_X2 U11645 ( .A1(n10377), .A2(n13202), .ZN(n16363) );
  NOR2_X2 U11646 ( .A1(n10972), .A2(n13204), .ZN(n16362) );
  NOR2_X2 U11647 ( .A1(n16361), .A2(n16360), .ZN(n16371) );
  NOR2_X2 U11648 ( .A1(n12427), .A2(n13199), .ZN(n16361) );
  NOR2_X2 U11649 ( .A1(n10853), .A2(n13201), .ZN(n16360) );
  NOR2_X2 U11650 ( .A1(n16367), .A2(n16366), .ZN(n16368) );
  NOR2_X2 U11651 ( .A1(n10897), .A2(n13474), .ZN(n16366) );
  NOR2_X2 U11652 ( .A1(n10896), .A2(n13473), .ZN(n16367) );
  NOR2_X2 U11653 ( .A1(n16365), .A2(n16364), .ZN(n16369) );
  NOR2_X2 U11654 ( .A1(n10392), .A2(n13468), .ZN(n16365) );
  NOR2_X2 U11655 ( .A1(n12947), .A2(n13470), .ZN(n16364) );
  NOR3_X2 U11656 ( .A1(n16343), .A2(n16342), .A3(n16341), .ZN(n16347) );
  NOR3_X2 U11657 ( .A1(n16340), .A2(n16339), .A3(n16338), .ZN(n16349) );
  NOR2_X2 U11658 ( .A1(n16345), .A2(n16344), .ZN(n16346) );
  NOR2_X2 U11659 ( .A1(n10990), .A2(n13447), .ZN(n16345) );
  NOR2_X2 U11660 ( .A1(n12748), .A2(n13450), .ZN(n16344) );
  AOI21_X2 U11661 ( .B1(n13378), .B2(REG_FILE_reg_out_9__11_), .A(n16379), 
        .ZN(n16380) );
  NOR2_X2 U11662 ( .A1(n16413), .A2(n13361), .ZN(n16379) );
  NOR2_X2 U11663 ( .A1(n13281), .A2(n11591), .ZN(n15114) );
  NOR2_X2 U11664 ( .A1(n12632), .A2(n13279), .ZN(n15113) );
  NOR3_X2 U11665 ( .A1(n14729), .A2(n14728), .A3(n14727), .ZN(n3434) );
  NOR2_X2 U11666 ( .A1(n13258), .A2(n11678), .ZN(n14727) );
  NOR2_X2 U11667 ( .A1(n13260), .A2(n11689), .ZN(n14728) );
  NOR2_X2 U11668 ( .A1(n13256), .A2(n11646), .ZN(n14729) );
  NOR3_X2 U11669 ( .A1(n16444), .A2(n16443), .A3(n16442), .ZN(n16450) );
  NOR2_X2 U11670 ( .A1(n16441), .A2(n13453), .ZN(n16443) );
  NOR2_X2 U11671 ( .A1(n10864), .A2(n13197), .ZN(n16442) );
  NOR2_X2 U11672 ( .A1(n10993), .A2(n13195), .ZN(n16444) );
  NOR2_X2 U11673 ( .A1(n16446), .A2(n16445), .ZN(n16448) );
  NOR2_X2 U11674 ( .A1(n13460), .A2(n12852), .ZN(n16445) );
  NOR2_X2 U11675 ( .A1(n13458), .A2(n12428), .ZN(n16446) );
  NOR2_X2 U11676 ( .A1(n16454), .A2(n16453), .ZN(n16461) );
  NOR2_X2 U11677 ( .A1(n10373), .A2(n13202), .ZN(n16454) );
  NOR2_X2 U11678 ( .A1(n10973), .A2(n13204), .ZN(n16453) );
  NOR2_X2 U11679 ( .A1(n16452), .A2(n16451), .ZN(n16462) );
  NOR2_X2 U11680 ( .A1(n11885), .A2(n13199), .ZN(n16452) );
  NOR2_X2 U11681 ( .A1(n10849), .A2(n13201), .ZN(n16451) );
  NOR2_X2 U11682 ( .A1(n16458), .A2(n16457), .ZN(n16459) );
  NOR2_X2 U11683 ( .A1(n10888), .A2(n13474), .ZN(n16457) );
  NOR2_X2 U11684 ( .A1(n10887), .A2(n13473), .ZN(n16458) );
  NOR2_X2 U11685 ( .A1(n16456), .A2(n16455), .ZN(n16460) );
  NOR2_X2 U11686 ( .A1(n10886), .A2(n13468), .ZN(n16456) );
  NOR2_X2 U11687 ( .A1(n12941), .A2(n13470), .ZN(n16455) );
  NOR3_X2 U11688 ( .A1(n16434), .A2(n16433), .A3(n16432), .ZN(n16438) );
  NOR3_X2 U11689 ( .A1(n16431), .A2(n16430), .A3(n16429), .ZN(n16440) );
  NOR2_X2 U11690 ( .A1(n16436), .A2(n16435), .ZN(n16437) );
  NOR2_X2 U11691 ( .A1(n10992), .A2(n13447), .ZN(n16436) );
  NOR2_X2 U11692 ( .A1(n12771), .A2(n13450), .ZN(n16435) );
  OAI21_X1 U11693 ( .B1(EXEC_STAGE_imm26_32[10]), .B2(net227290), .A(net232877), .ZN(net225906) );
  NOR3_X2 U11694 ( .A1(n16497), .A2(n16496), .A3(n16495), .ZN(n16503) );
  NOR2_X2 U11695 ( .A1(n16494), .A2(n13453), .ZN(n16496) );
  NOR2_X2 U11696 ( .A1(n10865), .A2(n13197), .ZN(n16495) );
  NOR2_X2 U11697 ( .A1(n10995), .A2(n13195), .ZN(n16497) );
  NOR2_X2 U11698 ( .A1(n16499), .A2(n16498), .ZN(n16501) );
  NOR2_X2 U11699 ( .A1(n13458), .A2(n12429), .ZN(n16499) );
  NOR2_X2 U11700 ( .A1(n13461), .A2(n12856), .ZN(n16498) );
  NOR2_X2 U11701 ( .A1(n16507), .A2(n16506), .ZN(n16514) );
  NOR2_X2 U11702 ( .A1(n10378), .A2(n13202), .ZN(n16507) );
  NOR2_X2 U11703 ( .A1(n10974), .A2(n13204), .ZN(n16506) );
  NOR2_X2 U11704 ( .A1(n16505), .A2(n16504), .ZN(n16515) );
  NOR2_X2 U11705 ( .A1(n12773), .A2(n13199), .ZN(n16505) );
  NOR2_X2 U11706 ( .A1(n10854), .A2(n13201), .ZN(n16504) );
  NOR2_X2 U11707 ( .A1(n16511), .A2(n16510), .ZN(n16512) );
  NOR2_X2 U11708 ( .A1(n10899), .A2(n13474), .ZN(n16510) );
  NOR2_X2 U11709 ( .A1(n10898), .A2(n13473), .ZN(n16511) );
  NOR2_X2 U11710 ( .A1(n16509), .A2(n16508), .ZN(n16513) );
  NOR2_X2 U11711 ( .A1(n10393), .A2(n13468), .ZN(n16509) );
  NOR2_X2 U11712 ( .A1(n12943), .A2(n13470), .ZN(n16508) );
  NOR3_X2 U11713 ( .A1(n16487), .A2(n16486), .A3(n16485), .ZN(n16491) );
  NOR3_X2 U11714 ( .A1(n16484), .A2(n16483), .A3(n16482), .ZN(n16493) );
  NOR2_X2 U11715 ( .A1(n16489), .A2(n16488), .ZN(n16490) );
  NOR2_X2 U11716 ( .A1(n10994), .A2(n13447), .ZN(n16489) );
  NOR2_X2 U11717 ( .A1(n12774), .A2(n13450), .ZN(n16488) );
  OAI21_X1 U11718 ( .B1(EXEC_STAGE_imm26_32[12]), .B2(net227290), .A(net232877), .ZN(net227071) );
  NOR3_X2 U11719 ( .A1(n14820), .A2(n14819), .A3(n14818), .ZN(n3127) );
  NOR2_X2 U11720 ( .A1(n13259), .A2(n11656), .ZN(n14818) );
  NOR2_X2 U11721 ( .A1(n13261), .A2(n12367), .ZN(n14819) );
  NOR2_X2 U11722 ( .A1(n13256), .A2(n11624), .ZN(n14820) );
  OAI21_X1 U11723 ( .B1(EXEC_STAGE_imm26_32[13]), .B2(net227290), .A(net232877), .ZN(net225778) );
  NOR3_X2 U11724 ( .A1(n16581), .A2(n16580), .A3(n16579), .ZN(n16587) );
  NOR2_X2 U11725 ( .A1(n17608), .A2(n13453), .ZN(n16580) );
  NOR2_X2 U11726 ( .A1(n10252), .A2(n13197), .ZN(n16579) );
  NOR2_X2 U11727 ( .A1(n10997), .A2(n13195), .ZN(n16581) );
  NOR2_X2 U11728 ( .A1(n16583), .A2(n16582), .ZN(n16585) );
  NOR2_X2 U11729 ( .A1(n13458), .A2(n12430), .ZN(n16583) );
  NOR2_X2 U11730 ( .A1(n13461), .A2(n12860), .ZN(n16582) );
  NOR2_X2 U11731 ( .A1(n16591), .A2(n16590), .ZN(n16598) );
  NOR2_X2 U11732 ( .A1(n10379), .A2(n13202), .ZN(n16591) );
  NOR2_X2 U11733 ( .A1(n10975), .A2(n13204), .ZN(n16590) );
  NOR2_X2 U11734 ( .A1(n16589), .A2(n16588), .ZN(n16599) );
  NOR2_X2 U11735 ( .A1(n12433), .A2(n13199), .ZN(n16589) );
  NOR2_X2 U11736 ( .A1(n10855), .A2(n13201), .ZN(n16588) );
  NOR2_X2 U11737 ( .A1(n16595), .A2(n16594), .ZN(n16596) );
  NOR2_X2 U11738 ( .A1(n10901), .A2(n13474), .ZN(n16594) );
  NOR2_X2 U11739 ( .A1(n10900), .A2(n13473), .ZN(n16595) );
  NOR2_X2 U11740 ( .A1(n16593), .A2(n16592), .ZN(n16597) );
  NOR2_X2 U11741 ( .A1(n10394), .A2(n13468), .ZN(n16593) );
  NOR2_X2 U11742 ( .A1(n12948), .A2(n13470), .ZN(n16592) );
  NOR3_X2 U11743 ( .A1(n16571), .A2(n16570), .A3(n16569), .ZN(n16575) );
  NOR3_X2 U11744 ( .A1(n16568), .A2(n16567), .A3(n16566), .ZN(n16577) );
  NOR2_X2 U11745 ( .A1(n16573), .A2(n16572), .ZN(n16574) );
  NOR2_X2 U11746 ( .A1(n10996), .A2(n13447), .ZN(n16573) );
  NOR2_X2 U11747 ( .A1(n12749), .A2(n13450), .ZN(n16572) );
  AOI21_X2 U11748 ( .B1(n13378), .B2(REG_FILE_reg_out_9__13_), .A(n16607), 
        .ZN(n16608) );
  NOR2_X2 U11749 ( .A1(n17608), .A2(n13361), .ZN(n16607) );
  NOR2_X2 U11750 ( .A1(n13282), .A2(n11594), .ZN(n15135) );
  NOR2_X2 U11751 ( .A1(n12635), .A2(n13278), .ZN(n15134) );
  NOR3_X2 U11752 ( .A1(n16642), .A2(n16641), .A3(n16640), .ZN(n16648) );
  NOR2_X2 U11753 ( .A1(n16639), .A2(n13453), .ZN(n16641) );
  NOR2_X2 U11754 ( .A1(n10866), .A2(n13197), .ZN(n16640) );
  NOR2_X2 U11755 ( .A1(n10999), .A2(n13195), .ZN(n16642) );
  NOR2_X2 U11756 ( .A1(n16644), .A2(n16643), .ZN(n16646) );
  NOR2_X2 U11757 ( .A1(n13458), .A2(n12434), .ZN(n16644) );
  NOR2_X2 U11758 ( .A1(n13461), .A2(n12864), .ZN(n16643) );
  NOR2_X2 U11759 ( .A1(n16652), .A2(n16651), .ZN(n16659) );
  NOR2_X2 U11760 ( .A1(n10380), .A2(n13202), .ZN(n16652) );
  NOR2_X2 U11761 ( .A1(n10976), .A2(n13204), .ZN(n16651) );
  NOR2_X2 U11762 ( .A1(n16650), .A2(n16649), .ZN(n16660) );
  NOR2_X2 U11763 ( .A1(n11887), .A2(n13199), .ZN(n16650) );
  NOR2_X2 U11764 ( .A1(n10856), .A2(n13201), .ZN(n16649) );
  NOR2_X2 U11765 ( .A1(n16656), .A2(n16655), .ZN(n16657) );
  NOR2_X2 U11766 ( .A1(n10903), .A2(n13474), .ZN(n16655) );
  NOR2_X2 U11767 ( .A1(n10902), .A2(n13473), .ZN(n16656) );
  NOR2_X2 U11768 ( .A1(n16654), .A2(n16653), .ZN(n16658) );
  NOR2_X2 U11769 ( .A1(n10395), .A2(n13468), .ZN(n16654) );
  NOR2_X2 U11770 ( .A1(n12944), .A2(n13470), .ZN(n16653) );
  NOR3_X2 U11771 ( .A1(n16632), .A2(n16631), .A3(n16630), .ZN(n16636) );
  NOR3_X2 U11772 ( .A1(n16629), .A2(n16628), .A3(n16627), .ZN(n16638) );
  NOR2_X2 U11773 ( .A1(n16634), .A2(n16633), .ZN(n16635) );
  NOR2_X2 U11774 ( .A1(n10998), .A2(n13447), .ZN(n16634) );
  NOR2_X2 U11775 ( .A1(n12775), .A2(n13450), .ZN(n16633) );
  NOR3_X2 U11776 ( .A1(n16685), .A2(n16684), .A3(n16683), .ZN(n16691) );
  NOR2_X2 U11777 ( .A1(n10253), .A2(n13197), .ZN(n16683) );
  NOR2_X2 U11778 ( .A1(n11000), .A2(n13195), .ZN(n16685) );
  NOR2_X2 U11779 ( .A1(n16687), .A2(n16686), .ZN(n16689) );
  NOR2_X2 U11780 ( .A1(n13458), .A2(n12435), .ZN(n16687) );
  NOR2_X2 U11781 ( .A1(n13461), .A2(n12868), .ZN(n16686) );
  NOR2_X2 U11782 ( .A1(n16695), .A2(n16694), .ZN(n16702) );
  NOR2_X2 U11783 ( .A1(n10846), .A2(n13202), .ZN(n16695) );
  NOR2_X2 U11784 ( .A1(n12080), .A2(n13204), .ZN(n16694) );
  NOR2_X2 U11785 ( .A1(n16693), .A2(n16692), .ZN(n16703) );
  NOR2_X2 U11786 ( .A1(n12438), .A2(n13199), .ZN(n16693) );
  NOR2_X2 U11787 ( .A1(n12024), .A2(n13201), .ZN(n16692) );
  NOR2_X2 U11788 ( .A1(n16699), .A2(n16698), .ZN(n16700) );
  NOR2_X2 U11789 ( .A1(n10905), .A2(n13474), .ZN(n16698) );
  NOR2_X2 U11790 ( .A1(n10904), .A2(n13473), .ZN(n16699) );
  NOR2_X2 U11791 ( .A1(n16697), .A2(n16696), .ZN(n16701) );
  NOR2_X2 U11792 ( .A1(n10396), .A2(n13468), .ZN(n16697) );
  NOR2_X2 U11793 ( .A1(n12952), .A2(n13470), .ZN(n16696) );
  NOR3_X2 U11794 ( .A1(n16676), .A2(n16675), .A3(n16674), .ZN(n16680) );
  NOR3_X2 U11795 ( .A1(n16673), .A2(n16672), .A3(n16671), .ZN(n16682) );
  NOR2_X2 U11796 ( .A1(n16678), .A2(n16677), .ZN(n16679) );
  NOR2_X2 U11797 ( .A1(n12082), .A2(n13447), .ZN(n16678) );
  NOR2_X2 U11798 ( .A1(n12750), .A2(n13450), .ZN(n16677) );
  AOI21_X2 U11799 ( .B1(n13378), .B2(REG_FILE_reg_out_9__15_), .A(n16712), 
        .ZN(n16713) );
  NOR2_X2 U11800 ( .A1(n13282), .A2(n11596), .ZN(n15156) );
  NOR2_X2 U11801 ( .A1(n12637), .A2(n13278), .ZN(n15155) );
  NOR3_X2 U11802 ( .A1(n16738), .A2(n16737), .A3(n16736), .ZN(n16764) );
  NAND3_X2 U11803 ( .A1(n16735), .A2(n16734), .A3(n16733), .ZN(n16738) );
  NOR3_X2 U11804 ( .A1(n14679), .A2(n14678), .A3(n14677), .ZN(n3605) );
  NOR2_X2 U11805 ( .A1(n14968), .A2(n11639), .ZN(n14679) );
  NOR2_X2 U11806 ( .A1(n13258), .A2(n11671), .ZN(n14677) );
  NOR2_X2 U11807 ( .A1(n13260), .A2(n11684), .ZN(n14678) );
  NOR3_X2 U11808 ( .A1(n16847), .A2(n16846), .A3(n16845), .ZN(n16853) );
  NOR2_X2 U11809 ( .A1(n16844), .A2(n13453), .ZN(n16846) );
  NOR2_X2 U11810 ( .A1(n10867), .A2(n13197), .ZN(n16845) );
  NOR2_X2 U11811 ( .A1(n12083), .A2(n13195), .ZN(n16847) );
  NOR2_X2 U11812 ( .A1(n16849), .A2(n16848), .ZN(n16851) );
  NOR2_X2 U11813 ( .A1(n13459), .A2(n12442), .ZN(n16849) );
  NOR2_X2 U11814 ( .A1(n13460), .A2(n12874), .ZN(n16848) );
  NOR3_X2 U11815 ( .A1(n16837), .A2(n16836), .A3(n16835), .ZN(n16841) );
  NOR3_X2 U11816 ( .A1(n16834), .A2(n16833), .A3(n16832), .ZN(n16843) );
  NOR2_X2 U11817 ( .A1(n16839), .A2(n16838), .ZN(n16840) );
  NOR2_X2 U11818 ( .A1(n11001), .A2(n13448), .ZN(n16839) );
  NOR2_X2 U11819 ( .A1(n12769), .A2(n13451), .ZN(n16838) );
  NOR2_X2 U11820 ( .A1(n16857), .A2(n16856), .ZN(n16864) );
  NOR2_X2 U11821 ( .A1(n10247), .A2(n13202), .ZN(n16857) );
  NOR2_X2 U11822 ( .A1(n10977), .A2(n13204), .ZN(n16856) );
  NOR2_X2 U11823 ( .A1(n16855), .A2(n16854), .ZN(n16865) );
  NOR2_X2 U11824 ( .A1(n11883), .A2(n13199), .ZN(n16855) );
  NOR2_X2 U11825 ( .A1(n10382), .A2(n13201), .ZN(n16854) );
  NOR2_X2 U11826 ( .A1(n16859), .A2(n16858), .ZN(n16863) );
  NOR2_X2 U11827 ( .A1(n10387), .A2(n13467), .ZN(n16859) );
  NOR2_X2 U11828 ( .A1(n12939), .A2(n13471), .ZN(n16858) );
  NOR2_X2 U11829 ( .A1(n16861), .A2(n16860), .ZN(n16862) );
  NOR2_X2 U11830 ( .A1(n10874), .A2(n13472), .ZN(n16861) );
  NOR2_X2 U11831 ( .A1(n10875), .A2(n13475), .ZN(n16860) );
  NOR3_X2 U11832 ( .A1(n16921), .A2(n16920), .A3(n16919), .ZN(n16927) );
  NOR2_X2 U11833 ( .A1(n17570), .A2(n13453), .ZN(n16920) );
  NOR2_X2 U11834 ( .A1(n10254), .A2(n13197), .ZN(n16919) );
  NOR2_X2 U11835 ( .A1(n12084), .A2(n13195), .ZN(n16921) );
  NOR2_X2 U11836 ( .A1(n16923), .A2(n16922), .ZN(n16925) );
  NOR2_X2 U11837 ( .A1(n13459), .A2(n12443), .ZN(n16923) );
  NOR2_X2 U11838 ( .A1(n13460), .A2(n12878), .ZN(n16922) );
  NOR3_X2 U11839 ( .A1(n16911), .A2(n16910), .A3(n16909), .ZN(n16915) );
  NOR3_X2 U11840 ( .A1(n16908), .A2(n16907), .A3(n16906), .ZN(n16917) );
  NOR2_X2 U11841 ( .A1(n16913), .A2(n16912), .ZN(n16914) );
  NOR2_X2 U11842 ( .A1(n11002), .A2(n13448), .ZN(n16913) );
  NOR2_X2 U11843 ( .A1(n12752), .A2(n13451), .ZN(n16912) );
  NOR2_X2 U11844 ( .A1(n16931), .A2(n16930), .ZN(n16938) );
  NOR2_X2 U11845 ( .A1(n10248), .A2(n13202), .ZN(n16931) );
  NOR2_X2 U11846 ( .A1(n10978), .A2(n13204), .ZN(n16930) );
  NOR2_X2 U11847 ( .A1(n16929), .A2(n16928), .ZN(n16939) );
  NOR2_X2 U11848 ( .A1(n12446), .A2(n13199), .ZN(n16929) );
  NOR2_X2 U11849 ( .A1(n10383), .A2(n13201), .ZN(n16928) );
  NOR2_X2 U11850 ( .A1(n16933), .A2(n16932), .ZN(n16937) );
  NOR2_X2 U11851 ( .A1(n10388), .A2(n13467), .ZN(n16933) );
  NOR2_X2 U11852 ( .A1(n12949), .A2(n13471), .ZN(n16932) );
  NOR2_X2 U11853 ( .A1(n16935), .A2(n16934), .ZN(n16936) );
  NOR2_X2 U11854 ( .A1(n10876), .A2(n13472), .ZN(n16935) );
  NOR2_X2 U11855 ( .A1(n10877), .A2(n13475), .ZN(n16934) );
  AOI21_X2 U11856 ( .B1(n13376), .B2(REG_FILE_reg_out_9__3_), .A(n16947), .ZN(
        n16948) );
  NOR2_X2 U11857 ( .A1(n17570), .A2(n13361), .ZN(n16947) );
  NOR2_X2 U11858 ( .A1(n13281), .A2(n12390), .ZN(n15041) );
  NOR2_X2 U11859 ( .A1(n12639), .A2(n13279), .ZN(n15040) );
  NOR3_X2 U11860 ( .A1(n16994), .A2(n16993), .A3(n16992), .ZN(n17000) );
  NOR2_X2 U11861 ( .A1(n17020), .A2(n13453), .ZN(n16993) );
  NOR2_X2 U11862 ( .A1(n10255), .A2(n13197), .ZN(n16992) );
  NOR2_X2 U11863 ( .A1(n12085), .A2(n13195), .ZN(n16994) );
  NOR2_X2 U11864 ( .A1(n16996), .A2(n16995), .ZN(n16998) );
  NOR2_X2 U11865 ( .A1(n13459), .A2(n12447), .ZN(n16996) );
  NOR2_X2 U11866 ( .A1(n13460), .A2(n12882), .ZN(n16995) );
  NOR3_X2 U11867 ( .A1(n16985), .A2(n16984), .A3(n16983), .ZN(n16989) );
  NOR3_X2 U11868 ( .A1(n16982), .A2(n16981), .A3(n16980), .ZN(n16991) );
  NOR2_X2 U11869 ( .A1(n16987), .A2(n16986), .ZN(n16988) );
  NOR2_X2 U11870 ( .A1(n11003), .A2(n13448), .ZN(n16987) );
  NOR2_X2 U11871 ( .A1(n12753), .A2(n13451), .ZN(n16986) );
  NOR2_X2 U11872 ( .A1(n17004), .A2(n17003), .ZN(n17011) );
  NOR2_X2 U11873 ( .A1(n10375), .A2(n13202), .ZN(n17004) );
  NOR2_X2 U11874 ( .A1(n10979), .A2(n13204), .ZN(n17003) );
  NOR2_X2 U11875 ( .A1(n17002), .A2(n17001), .ZN(n17012) );
  NOR2_X2 U11876 ( .A1(n12450), .A2(n13199), .ZN(n17002) );
  NOR2_X2 U11877 ( .A1(n10851), .A2(n13201), .ZN(n17001) );
  NOR2_X2 U11878 ( .A1(n17006), .A2(n17005), .ZN(n17010) );
  NOR2_X2 U11879 ( .A1(n10390), .A2(n13467), .ZN(n17006) );
  NOR2_X2 U11880 ( .A1(n12950), .A2(n13471), .ZN(n17005) );
  NOR2_X2 U11881 ( .A1(n17008), .A2(n17007), .ZN(n17009) );
  NOR2_X2 U11882 ( .A1(n10892), .A2(n13472), .ZN(n17008) );
  NOR2_X2 U11883 ( .A1(n10893), .A2(n13475), .ZN(n17007) );
  AOI21_X2 U11884 ( .B1(n13376), .B2(REG_FILE_reg_out_9__9_), .A(n17021), .ZN(
        n17022) );
  NOR2_X2 U11885 ( .A1(n17020), .A2(n13361), .ZN(n17021) );
  NOR2_X2 U11886 ( .A1(n13281), .A2(n12398), .ZN(n15104) );
  NOR2_X2 U11887 ( .A1(n12640), .A2(n13279), .ZN(n15103) );
  NOR2_X2 U11888 ( .A1(nextPC_ex_out[10]), .A2(net227065), .ZN(net227064) );
  NOR3_X2 U11889 ( .A1(n17079), .A2(n17078), .A3(n17077), .ZN(n17105) );
  NAND3_X2 U11890 ( .A1(n17076), .A2(n17075), .A3(n17074), .ZN(n17079) );
  NAND3_X2 U11891 ( .A1(net227105), .A2(net227106), .A3(n13010), .ZN(net224954) );
  NAND2_X1 U11892 ( .A1(n13358), .A2(n13151), .ZN(n16815) );
  NOR3_X2 U11893 ( .A1(n14669), .A2(n14668), .A3(n14667), .ZN(n3639) );
  NOR2_X2 U11894 ( .A1(n14968), .A2(n11628), .ZN(n14669) );
  NOR2_X2 U11895 ( .A1(n13258), .A2(n11660), .ZN(n14667) );
  NOR2_X2 U11896 ( .A1(n13260), .A2(n11683), .ZN(n14668) );
  NOR3_X2 U11897 ( .A1(n17171), .A2(n17170), .A3(n17169), .ZN(n17177) );
  NOR2_X2 U11898 ( .A1(n17168), .A2(n13453), .ZN(n17170) );
  NOR2_X2 U11899 ( .A1(n10868), .A2(n13197), .ZN(n17169) );
  NOR2_X2 U11900 ( .A1(n12086), .A2(n13195), .ZN(n17171) );
  NOR2_X2 U11901 ( .A1(n17173), .A2(n17172), .ZN(n17175) );
  NOR2_X2 U11902 ( .A1(n13459), .A2(n12454), .ZN(n17173) );
  NOR2_X2 U11903 ( .A1(n13460), .A2(n12888), .ZN(n17172) );
  NOR3_X2 U11904 ( .A1(n17161), .A2(n17160), .A3(n17159), .ZN(n17165) );
  NOR3_X2 U11905 ( .A1(n17158), .A2(n17157), .A3(n17156), .ZN(n17167) );
  NOR2_X2 U11906 ( .A1(n17163), .A2(n17162), .ZN(n17164) );
  NOR2_X2 U11907 ( .A1(n11004), .A2(n13448), .ZN(n17163) );
  NOR2_X2 U11908 ( .A1(n12768), .A2(n13451), .ZN(n17162) );
  NOR2_X2 U11909 ( .A1(n17181), .A2(n17180), .ZN(n17188) );
  NOR2_X2 U11910 ( .A1(n10246), .A2(n13202), .ZN(n17181) );
  NOR2_X2 U11911 ( .A1(n10980), .A2(n13204), .ZN(n17180) );
  NOR2_X2 U11912 ( .A1(n17179), .A2(n17178), .ZN(n17189) );
  NOR2_X2 U11913 ( .A1(n11882), .A2(n13199), .ZN(n17179) );
  NOR2_X2 U11914 ( .A1(n10381), .A2(n13201), .ZN(n17178) );
  NOR2_X2 U11915 ( .A1(n17183), .A2(n17182), .ZN(n17187) );
  NOR2_X2 U11916 ( .A1(n10386), .A2(n13467), .ZN(n17183) );
  NOR2_X2 U11917 ( .A1(n12938), .A2(n13471), .ZN(n17182) );
  NOR2_X2 U11918 ( .A1(n17185), .A2(n17184), .ZN(n17186) );
  NOR2_X2 U11919 ( .A1(n10872), .A2(n13472), .ZN(n17185) );
  NOR2_X2 U11920 ( .A1(n10873), .A2(n13475), .ZN(n17184) );
  INV_X4 U11921 ( .A(n13180), .ZN(n19157) );
  NOR3_X2 U11922 ( .A1(n17245), .A2(n17244), .A3(n17243), .ZN(n17251) );
  NOR2_X2 U11923 ( .A1(n17313), .A2(n13453), .ZN(n17244) );
  NOR2_X2 U11924 ( .A1(n10256), .A2(n13197), .ZN(n17243) );
  NOR2_X2 U11925 ( .A1(n12087), .A2(n13195), .ZN(n17245) );
  NOR2_X2 U11926 ( .A1(n17247), .A2(n17246), .ZN(n17249) );
  NOR2_X2 U11927 ( .A1(n13459), .A2(n12455), .ZN(n17247) );
  NOR2_X2 U11928 ( .A1(n13460), .A2(n12892), .ZN(n17246) );
  NOR3_X2 U11929 ( .A1(n17232), .A2(n17231), .A3(n17230), .ZN(n17241) );
  NOR2_X2 U11930 ( .A1(n17237), .A2(n17236), .ZN(n17238) );
  NOR2_X2 U11931 ( .A1(n11005), .A2(n13448), .ZN(n17237) );
  NOR2_X2 U11932 ( .A1(n12755), .A2(n13451), .ZN(n17236) );
  NOR2_X2 U11933 ( .A1(n17255), .A2(n17254), .ZN(n17262) );
  NOR2_X2 U11934 ( .A1(n10249), .A2(n13202), .ZN(n17255) );
  NOR2_X2 U11935 ( .A1(n17253), .A2(n17252), .ZN(n17263) );
  NOR2_X2 U11936 ( .A1(n12458), .A2(n13199), .ZN(n17253) );
  NOR2_X2 U11937 ( .A1(n10384), .A2(n13201), .ZN(n17252) );
  NOR2_X2 U11938 ( .A1(n17257), .A2(n17256), .ZN(n17261) );
  NOR2_X2 U11939 ( .A1(n10389), .A2(n13467), .ZN(n17257) );
  NOR2_X2 U11940 ( .A1(n12951), .A2(n13471), .ZN(n17256) );
  NOR2_X2 U11941 ( .A1(n17259), .A2(n17258), .ZN(n17260) );
  NOR2_X2 U11942 ( .A1(n10878), .A2(n13472), .ZN(n17259) );
  NOR2_X2 U11943 ( .A1(n10879), .A2(n13475), .ZN(n17258) );
  AOI21_X2 U11944 ( .B1(n13378), .B2(REG_FILE_reg_out_9__4_), .A(n17274), .ZN(
        n17275) );
  NOR2_X2 U11945 ( .A1(n17313), .A2(n13361), .ZN(n17274) );
  INV_X4 U11946 ( .A(n13178), .ZN(n19159) );
  NOR2_X2 U11947 ( .A1(n13281), .A2(n12391), .ZN(n15046) );
  NOR2_X2 U11948 ( .A1(n12642), .A2(n13279), .ZN(n15045) );
  NAND3_X2 U11949 ( .A1(n16311), .A2(n18252), .A3(n16019), .ZN(n17300) );
  NOR3_X2 U11950 ( .A1(n17349), .A2(n17348), .A3(n17347), .ZN(n17374) );
  NAND3_X2 U11951 ( .A1(n17346), .A2(n17345), .A3(n17344), .ZN(n17349) );
  NOR3_X2 U11952 ( .A1(n17400), .A2(n17399), .A3(n17398), .ZN(n17425) );
  NAND3_X2 U11953 ( .A1(n17397), .A2(n17396), .A3(n17395), .ZN(n17400) );
  NAND3_X2 U11954 ( .A1(n17474), .A2(n17473), .A3(n17472), .ZN(n17477) );
  NOR3_X2 U11955 ( .A1(n17455), .A2(n17454), .A3(n17453), .ZN(n17481) );
  NAND3_X2 U11956 ( .A1(n17452), .A2(n17451), .A3(n17450), .ZN(n17455) );
  NOR2_X1 U11957 ( .A1(n13209), .A2(n17544), .ZN(n17545) );
  NOR3_X2 U11958 ( .A1(n14689), .A2(n14688), .A3(n14687), .ZN(n3571) );
  NOR2_X2 U11959 ( .A1(n14968), .A2(n11642), .ZN(n14689) );
  NOR2_X2 U11960 ( .A1(n13258), .A2(n11674), .ZN(n14687) );
  NOR2_X2 U11961 ( .A1(n13260), .A2(n11685), .ZN(n14688) );
  NOR3_X2 U11962 ( .A1(n14790), .A2(n14789), .A3(n14788), .ZN(n3230) );
  NOR2_X2 U11963 ( .A1(n13259), .A2(n11653), .ZN(n14788) );
  NOR2_X2 U11964 ( .A1(n13261), .A2(n12361), .ZN(n14789) );
  NOR2_X2 U11965 ( .A1(n13256), .A2(n11621), .ZN(n14790) );
  NOR3_X2 U11966 ( .A1(n14800), .A2(n14799), .A3(n14798), .ZN(n3195) );
  NOR2_X2 U11967 ( .A1(n13259), .A2(n11654), .ZN(n14798) );
  NOR2_X2 U11968 ( .A1(n13261), .A2(n12363), .ZN(n14799) );
  NOR2_X2 U11969 ( .A1(n13256), .A2(n11622), .ZN(n14800) );
  INV_X4 U11970 ( .A(n13384), .ZN(n13383) );
  INV_X4 U11971 ( .A(n13375), .ZN(n13374) );
  INV_X4 U11972 ( .A(n13372), .ZN(n13370) );
  NAND3_X2 U11973 ( .A1(n17993), .A2(n17696), .A3(n17695), .ZN(n18329) );
  NOR2_X2 U11974 ( .A1(n17694), .A2(net224151), .ZN(n17695) );
  NOR2_X2 U11975 ( .A1(n13021), .A2(net232817), .ZN(net224151) );
  NAND3_X2 U11976 ( .A1(n17530), .A2(n17993), .A3(n17529), .ZN(n18328) );
  NOR3_X2 U11977 ( .A1(n14810), .A2(n14809), .A3(n14808), .ZN(n3161) );
  NOR2_X2 U11978 ( .A1(n13259), .A2(n11655), .ZN(n14808) );
  NOR2_X2 U11979 ( .A1(n13261), .A2(n12365), .ZN(n14809) );
  NOR2_X2 U11980 ( .A1(n13256), .A2(n11623), .ZN(n14810) );
  NOR3_X2 U11981 ( .A1(n14940), .A2(n14939), .A3(n14938), .ZN(n2718) );
  NOR2_X2 U11982 ( .A1(n13258), .A2(n11669), .ZN(n14938) );
  NOR2_X2 U11983 ( .A1(n13260), .A2(n12077), .ZN(n14939) );
  NOR2_X2 U11984 ( .A1(n13256), .A2(n11637), .ZN(n14940) );
  NOR3_X2 U11985 ( .A1(n14920), .A2(n14919), .A3(n14918), .ZN(n2786) );
  NOR2_X2 U11986 ( .A1(n13258), .A2(n11667), .ZN(n14918) );
  NOR2_X2 U11987 ( .A1(n13260), .A2(n12075), .ZN(n14919) );
  NOR2_X2 U11988 ( .A1(n13256), .A2(n11635), .ZN(n14920) );
  NOR3_X2 U11989 ( .A1(n14930), .A2(n14929), .A3(n14928), .ZN(n2752) );
  NOR2_X2 U11990 ( .A1(n13259), .A2(n11668), .ZN(n14928) );
  NOR2_X2 U11991 ( .A1(n13261), .A2(n12076), .ZN(n14929) );
  NOR2_X2 U11992 ( .A1(n13256), .A2(n11636), .ZN(n14930) );
  NOR3_X2 U11993 ( .A1(n14910), .A2(n14909), .A3(n14908), .ZN(n2820) );
  NOR2_X2 U11994 ( .A1(n13259), .A2(n11666), .ZN(n14908) );
  NOR2_X2 U11995 ( .A1(n13261), .A2(n12074), .ZN(n14909) );
  NOR2_X2 U11996 ( .A1(n13256), .A2(n11634), .ZN(n14910) );
  NAND3_X2 U11997 ( .A1(n15785), .A2(n13044), .A3(n14098), .ZN(n14044) );
  NOR3_X2 U11998 ( .A1(n14950), .A2(n14949), .A3(n14948), .ZN(n2684) );
  NOR2_X2 U11999 ( .A1(n13259), .A2(n11670), .ZN(n14948) );
  NOR2_X2 U12000 ( .A1(n13261), .A2(n12078), .ZN(n14949) );
  NOR2_X2 U12001 ( .A1(n13256), .A2(n11638), .ZN(n14950) );
  INV_X4 U12002 ( .A(n13479), .ZN(n13478) );
  INV_X4 U12003 ( .A(n18845), .ZN(n13479) );
  NOR3_X2 U12004 ( .A1(n14960), .A2(n14959), .A3(n14958), .ZN(n2650) );
  NOR2_X2 U12005 ( .A1(n13258), .A2(n11672), .ZN(n14958) );
  NOR2_X2 U12006 ( .A1(n13260), .A2(n11494), .ZN(n14959) );
  NOR2_X2 U12007 ( .A1(n13256), .A2(n11640), .ZN(n14960) );
  NOR2_X1 U12008 ( .A1(n18534), .A2(net222304), .ZN(n18538) );
  NAND3_X2 U12009 ( .A1(n13993), .A2(n13992), .A3(n13991), .ZN(n15700) );
  NAND3_X1 U12010 ( .A1(MEM_WB_OUT[67]), .A2(n14078), .A3(n13880), .ZN(n13992)
         );
  INV_X8 U12011 ( .A(n15836), .ZN(n18927) );
  NOR3_X2 U12012 ( .A1(n14840), .A2(n14839), .A3(n14838), .ZN(n3059) );
  NOR2_X2 U12013 ( .A1(n13259), .A2(n11658), .ZN(n14838) );
  NOR2_X2 U12014 ( .A1(n13261), .A2(n12371), .ZN(n14839) );
  NOR2_X2 U12015 ( .A1(n13256), .A2(n11626), .ZN(n14840) );
  NAND3_X2 U12016 ( .A1(n17993), .A2(n17125), .A3(n17124), .ZN(n17994) );
  NOR2_X2 U12017 ( .A1(n17123), .A2(n17122), .ZN(n17124) );
  INV_X4 U12018 ( .A(n13394), .ZN(n13393) );
  NOR2_X2 U12019 ( .A1(n16791), .A2(net232817), .ZN(n16792) );
  NAND3_X2 U12020 ( .A1(n17519), .A2(n17993), .A3(n17518), .ZN(n18296) );
  NOR2_X2 U12021 ( .A1(n17517), .A2(n17516), .ZN(n17518) );
  NOR2_X2 U12022 ( .A1(n18658), .A2(n18657), .ZN(n18659) );
  AOI21_X2 U12023 ( .B1(n18656), .B2(n18655), .A(n18668), .ZN(n18657) );
  OAI21_X1 U12024 ( .B1(n18662), .B2(n18661), .A(n18660), .ZN(n18663) );
  OAI21_X1 U12025 ( .B1(n13218), .B2(n11913), .A(n6741), .ZN(n6625) );
  NAND3_X1 U12026 ( .A1(n13218), .A2(n11913), .A3(ID_EXEC_OUT[156]), .ZN(n6741) );
  NOR3_X2 U12027 ( .A1(n15695), .A2(n17517), .A3(n15694), .ZN(n15696) );
  OAI21_X1 U12028 ( .B1(n18635), .B2(n19101), .A(n18634), .ZN(n18640) );
  NOR2_X1 U12029 ( .A1(n18630), .A2(net232817), .ZN(n18631) );
  NOR2_X1 U12030 ( .A1(n18638), .A2(n18637), .ZN(n18639) );
  OAI21_X2 U12031 ( .B1(n15735), .B2(n15734), .A(n15733), .ZN(n15746) );
  NOR2_X2 U12032 ( .A1(n15744), .A2(n15743), .ZN(n15745) );
  NAND2_X2 U12033 ( .A1(n14293), .A2(n14982), .ZN(n14632) );
  INV_X4 U12034 ( .A(n13170), .ZN(n14400) );
  INV_X4 U12035 ( .A(n13384), .ZN(n13382) );
  INV_X8 U12036 ( .A(n13378), .ZN(n13377) );
  INV_X4 U12037 ( .A(n17270), .ZN(n13187) );
  NAND2_X1 U12038 ( .A1(n14991), .A2(n2506), .ZN(n17270) );
  NOR3_X2 U12039 ( .A1(n18717), .A2(n18716), .A3(n18715), .ZN(n18725) );
  NOR2_X1 U12040 ( .A1(n18930), .A2(n13452), .ZN(n18716) );
  NOR2_X2 U12041 ( .A1(n10367), .A2(n13197), .ZN(n18715) );
  NOR2_X2 U12042 ( .A1(n10257), .A2(n13195), .ZN(n18717) );
  NOR2_X2 U12043 ( .A1(n18720), .A2(n18719), .ZN(n18723) );
  NOR2_X2 U12044 ( .A1(n13458), .A2(n12498), .ZN(n18720) );
  NOR2_X2 U12045 ( .A1(n13461), .A2(n12920), .ZN(n18719) );
  NOR3_X2 U12046 ( .A1(n18704), .A2(n18703), .A3(n18702), .ZN(n18709) );
  NOR3_X2 U12047 ( .A1(n18696), .A2(n18695), .A3(n18694), .ZN(n18711) );
  NAND3_X2 U12048 ( .A1(n18693), .A2(n18692), .A3(n18691), .ZN(n18694) );
  NOR2_X2 U12049 ( .A1(n18707), .A2(n18706), .ZN(n18708) );
  NOR2_X2 U12050 ( .A1(n12025), .A2(n13447), .ZN(n18707) );
  NOR2_X2 U12051 ( .A1(n12785), .A2(n13450), .ZN(n18706) );
  NOR2_X2 U12052 ( .A1(n18732), .A2(n18731), .ZN(n18740) );
  NOR2_X2 U12053 ( .A1(n12412), .A2(n13202), .ZN(n18732) );
  NOR2_X2 U12054 ( .A1(n12088), .A2(n13204), .ZN(n18731) );
  NOR2_X2 U12055 ( .A1(n18729), .A2(n18728), .ZN(n18741) );
  NOR2_X2 U12056 ( .A1(n12063), .A2(n13199), .ZN(n18729) );
  NOR2_X2 U12057 ( .A1(n12411), .A2(n13201), .ZN(n18728) );
  NOR2_X2 U12058 ( .A1(n18737), .A2(n18736), .ZN(n18738) );
  NOR2_X2 U12059 ( .A1(n12081), .A2(n13474), .ZN(n18736) );
  NOR2_X2 U12060 ( .A1(n10847), .A2(n13473), .ZN(n18737) );
  NOR2_X2 U12061 ( .A1(n18735), .A2(n18734), .ZN(n18739) );
  NOR2_X2 U12062 ( .A1(n10251), .A2(n13468), .ZN(n18735) );
  NOR2_X2 U12063 ( .A1(n12062), .A2(n13470), .ZN(n18734) );
  INV_X4 U12064 ( .A(net231353), .ZN(net231333) );
  NOR3_X2 U12065 ( .A1(n18849), .A2(n18848), .A3(n18847), .ZN(n19059) );
  AOI21_X2 U12066 ( .B1(n13492), .B2(n19113), .A(n19112), .ZN(n19120) );
  NOR2_X2 U12067 ( .A1(n18314), .A2(n13207), .ZN(n18315) );
  INV_X4 U12068 ( .A(n13127), .ZN(n13148) );
  INV_X4 U12069 ( .A(n13124), .ZN(n13154) );
  INV_X16 U12070 ( .A(n13351), .ZN(n13349) );
  INV_X16 U12071 ( .A(n13346), .ZN(n13344) );
  INV_X4 U12072 ( .A(reset), .ZN(n13956) );
  INV_X4 U12073 ( .A(reset), .ZN(n13955) );
  NOR2_X2 U12074 ( .A1(EXEC_STAGE_mul_ex_CurrentState_0_), .A2(
        EXEC_STAGE_mul_ex_CurrentState_2_), .ZN(n7289) );
  NOR2_X2 U12075 ( .A1(n13245), .A2(n12342), .ZN(n14528) );
  NOR2_X2 U12076 ( .A1(net231243), .A2(n11956), .ZN(n14526) );
  NOR2_X2 U12077 ( .A1(n13245), .A2(n12341), .ZN(n14517) );
  NOR2_X2 U12078 ( .A1(net231239), .A2(n10812), .ZN(n14515) );
  NOR2_X2 U12079 ( .A1(n14988), .A2(n14987), .ZN(n2502) );
  NOR2_X2 U12080 ( .A1(n12826), .A2(n13272), .ZN(n14988) );
  NOR2_X2 U12081 ( .A1(n12827), .A2(n13269), .ZN(n14987) );
  NOR3_X2 U12082 ( .A1(n14994), .A2(n14993), .A3(n14992), .ZN(n15004) );
  NOR2_X2 U12083 ( .A1(n2522), .A2(n14989), .ZN(n15006) );
  NOR3_X2 U12084 ( .A1(n14985), .A2(n14984), .A3(n14983), .ZN(n2509) );
  NOR2_X2 U12085 ( .A1(n13281), .A2(n11586), .ZN(n14985) );
  NOR2_X2 U12086 ( .A1(n12627), .A2(n13279), .ZN(n14984) );
  AOI21_X1 U12087 ( .B1(net231615), .B2(n18870), .A(n15649), .ZN(n15650) );
  NOR2_X2 U12088 ( .A1(net231249), .A2(n12122), .ZN(n15649) );
  NOR2_X2 U12089 ( .A1(n13244), .A2(n12326), .ZN(n14351) );
  NOR2_X2 U12090 ( .A1(net231217), .A2(n11931), .ZN(n14349) );
  NOR2_X2 U12091 ( .A1(n4510), .A2(n4511), .ZN(n4495) );
  NOR2_X2 U12092 ( .A1(n15053), .A2(n15052), .ZN(n2402) );
  NOR2_X2 U12093 ( .A1(n12830), .A2(n13272), .ZN(n15053) );
  NOR2_X2 U12094 ( .A1(n12831), .A2(n13269), .ZN(n15052) );
  NOR3_X2 U12095 ( .A1(n15057), .A2(n15056), .A3(n15055), .ZN(n15062) );
  NOR2_X2 U12096 ( .A1(n2412), .A2(n15054), .ZN(n15064) );
  NOR3_X2 U12097 ( .A1(n15051), .A2(n15050), .A3(n15049), .ZN(n2403) );
  NOR2_X2 U12098 ( .A1(n13281), .A2(n11587), .ZN(n15051) );
  NOR2_X2 U12099 ( .A1(n12628), .A2(n13279), .ZN(n15050) );
  NOR2_X1 U12100 ( .A1(n19031), .A2(n13491), .ZN(n16084) );
  NAND3_X2 U12101 ( .A1(n16058), .A2(n16057), .A3(n16056), .ZN(n16076) );
  AOI21_X2 U12102 ( .B1(n16073), .B2(n16072), .A(n16071), .ZN(n16074) );
  NOR2_X2 U12103 ( .A1(n15090), .A2(n15089), .ZN(n2341) );
  NOR2_X2 U12104 ( .A1(n12838), .A2(n13272), .ZN(n15090) );
  NOR2_X2 U12105 ( .A1(n12839), .A2(n13269), .ZN(n15089) );
  NOR3_X2 U12106 ( .A1(n15094), .A2(n15093), .A3(n15092), .ZN(n15099) );
  NOR2_X2 U12107 ( .A1(n2351), .A2(n15091), .ZN(n15101) );
  NOR3_X2 U12108 ( .A1(n15088), .A2(n15087), .A3(n15086), .ZN(n2342) );
  NOR2_X2 U12109 ( .A1(n13281), .A2(n11589), .ZN(n15088) );
  NOR2_X2 U12110 ( .A1(n12630), .A2(n13279), .ZN(n15087) );
  NOR2_X2 U12111 ( .A1(n13211), .A2(n16316), .ZN(n16317) );
  NAND3_X2 U12112 ( .A1(n16309), .A2(n16308), .A3(n16307), .ZN(n16318) );
  OAI21_X1 U12113 ( .B1(n16298), .B2(n16297), .A(n19016), .ZN(n16308) );
  NOR2_X1 U12114 ( .A1(n19011), .A2(n13491), .ZN(n16326) );
  NOR2_X2 U12115 ( .A1(n15074), .A2(n15073), .ZN(n2362) );
  NOR2_X2 U12116 ( .A1(n12850), .A2(n13272), .ZN(n15074) );
  NOR2_X2 U12117 ( .A1(n12851), .A2(n13269), .ZN(n15073) );
  NOR3_X2 U12118 ( .A1(n15078), .A2(n15077), .A3(n15076), .ZN(n15083) );
  NOR2_X2 U12119 ( .A1(n2372), .A2(n15075), .ZN(n15085) );
  NOR3_X2 U12120 ( .A1(n15072), .A2(n15071), .A3(n15070), .ZN(n2363) );
  NOR2_X2 U12121 ( .A1(n13281), .A2(n11592), .ZN(n15072) );
  NOR2_X2 U12122 ( .A1(n12633), .A2(n13279), .ZN(n15071) );
  OAI21_X1 U12123 ( .B1(n15413), .B2(IMEM_BUS_OUT[11]), .A(n15412), .ZN(n16474) );
  OAI21_X2 U12124 ( .B1(EXEC_STAGE_imm26_32[11]), .B2(net227290), .A(net232877), .ZN(net225894) );
  NOR2_X2 U12125 ( .A1(n15121), .A2(n15120), .ZN(n2261) );
  NOR2_X2 U12126 ( .A1(n12854), .A2(n13273), .ZN(n15121) );
  NOR2_X2 U12127 ( .A1(n12855), .A2(n13270), .ZN(n15120) );
  NOR3_X2 U12128 ( .A1(n15125), .A2(n15124), .A3(n15123), .ZN(n15130) );
  NOR2_X2 U12129 ( .A1(n2271), .A2(n15122), .ZN(n15132) );
  NOR3_X2 U12130 ( .A1(n15119), .A2(n15118), .A3(n15117), .ZN(n2262) );
  NOR2_X2 U12131 ( .A1(n13282), .A2(n11593), .ZN(n15119) );
  NOR2_X2 U12132 ( .A1(n12634), .A2(n13278), .ZN(n15118) );
  NAND3_X2 U12133 ( .A1(n16542), .A2(n16541), .A3(n16540), .ZN(n16551) );
  NAND3_X2 U12134 ( .A1(n16528), .A2(n16527), .A3(n16526), .ZN(n17617) );
  AOI21_X2 U12135 ( .B1(n15420), .B2(IMEM_BUS_OUT[14]), .A(IMEM_BUS_OUT[13]), 
        .ZN(n15416) );
  NOR2_X2 U12136 ( .A1(n15142), .A2(n15141), .ZN(n2221) );
  NOR2_X2 U12137 ( .A1(n12862), .A2(n13273), .ZN(n15142) );
  NOR2_X2 U12138 ( .A1(n12863), .A2(n13270), .ZN(n15141) );
  NOR3_X2 U12139 ( .A1(n15146), .A2(n15145), .A3(n15144), .ZN(n15151) );
  NOR2_X2 U12140 ( .A1(n2231), .A2(n15143), .ZN(n15153) );
  NOR3_X2 U12141 ( .A1(n15140), .A2(n15139), .A3(n15138), .ZN(n2222) );
  NOR2_X2 U12142 ( .A1(n13282), .A2(n11595), .ZN(n15140) );
  NOR2_X2 U12143 ( .A1(n12636), .A2(n13278), .ZN(n15139) );
  AOI222_X1 U12144 ( .A1(n19153), .A2(REG_FILE_reg_out_14__16_), .B1(n13499), 
        .B2(REG_FILE_reg_out_4__16_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__16_), .ZN(n2172) );
  NOR3_X2 U12145 ( .A1(n15170), .A2(n15169), .A3(n15168), .ZN(n15171) );
  NOR2_X2 U12146 ( .A1(n12751), .A2(n13382), .ZN(n15169) );
  OAI21_X2 U12147 ( .B1(n13364), .B2(n12870), .A(n12922), .ZN(n15170) );
  NOR2_X1 U12148 ( .A1(n12797), .A2(n13377), .ZN(n15168) );
  NOR3_X2 U12149 ( .A1(n15167), .A2(n15166), .A3(n15165), .ZN(n15172) );
  NOR2_X2 U12150 ( .A1(n10942), .A2(n13371), .ZN(n15166) );
  NOR2_X2 U12151 ( .A1(n11854), .A2(n13373), .ZN(n15165) );
  NOR3_X2 U12152 ( .A1(n15161), .A2(n15160), .A3(n15159), .ZN(n2179) );
  NOR2_X2 U12153 ( .A1(n15027), .A2(n15026), .ZN(n2462) );
  NOR2_X2 U12154 ( .A1(n12872), .A2(n13272), .ZN(n15027) );
  NOR2_X2 U12155 ( .A1(n12873), .A2(n13269), .ZN(n15026) );
  NOR3_X2 U12156 ( .A1(n15031), .A2(n15030), .A3(n15029), .ZN(n15036) );
  NOR2_X2 U12157 ( .A1(n2472), .A2(n15028), .ZN(n15038) );
  NOR3_X2 U12158 ( .A1(n15025), .A2(n15024), .A3(n15023), .ZN(n2463) );
  NOR2_X2 U12159 ( .A1(n13281), .A2(n12387), .ZN(n15025) );
  NOR2_X2 U12160 ( .A1(n12638), .A2(n13279), .ZN(n15024) );
  AOI211_X2 U12161 ( .C1(n18644), .C2(n17561), .A(n16894), .B(n16893), .ZN(
        n16895) );
  AOI21_X1 U12162 ( .B1(n18360), .B2(n16876), .A(n16875), .ZN(n16897) );
  OAI21_X1 U12163 ( .B1(n13021), .B2(net223104), .A(n13022), .ZN(net225203) );
  INV_X4 U12164 ( .A(n16970), .ZN(n13080) );
  INV_X4 U12165 ( .A(net231273), .ZN(net231253) );
  AOI21_X1 U12166 ( .B1(n15435), .B2(IMEM_BUS_OUT[10]), .A(IMEM_BUS_OUT[9]), 
        .ZN(n15436) );
  NOR2_X1 U12167 ( .A1(n12802), .A2(n13377), .ZN(n17110) );
  OAI21_X2 U12168 ( .B1(n13364), .B2(n12884), .A(n12929), .ZN(n17108) );
  NOR3_X2 U12169 ( .A1(n15175), .A2(n15174), .A3(n15173), .ZN(n2159) );
  NOR2_X2 U12170 ( .A1(n15011), .A2(n15010), .ZN(n2482) );
  NOR2_X2 U12171 ( .A1(n12886), .A2(n13272), .ZN(n15011) );
  NOR2_X2 U12172 ( .A1(n12887), .A2(n13269), .ZN(n15010) );
  NOR3_X2 U12173 ( .A1(n15015), .A2(n15014), .A3(n15013), .ZN(n15020) );
  NOR2_X2 U12174 ( .A1(n2492), .A2(n15012), .ZN(n15022) );
  NOR3_X2 U12175 ( .A1(n15009), .A2(n15008), .A3(n15007), .ZN(n2483) );
  NOR2_X2 U12176 ( .A1(n13281), .A2(n12384), .ZN(n15009) );
  NOR2_X2 U12177 ( .A1(n12641), .A2(n13278), .ZN(n15008) );
  AOI21_X1 U12178 ( .B1(net231615), .B2(n18872), .A(n17220), .ZN(n17221) );
  NOR2_X2 U12179 ( .A1(net231227), .A2(n12125), .ZN(n17220) );
  NOR2_X2 U12180 ( .A1(nextPC_ex_out[3]), .A2(net224713), .ZN(n17217) );
  INV_X4 U12181 ( .A(n15634), .ZN(n17267) );
  AOI21_X2 U12182 ( .B1(n15633), .B2(n18754), .A(n16766), .ZN(n15634) );
  NOR2_X2 U12183 ( .A1(n13221), .A2(n12020), .ZN(n15633) );
  AOI21_X1 U12184 ( .B1(net231615), .B2(n18867), .A(n17286), .ZN(n17288) );
  NAND3_X2 U12185 ( .A1(net224704), .A2(nextPC_ex_out[4]), .A3(
        nextPC_ex_out[5]), .ZN(n17287) );
  NOR2_X2 U12186 ( .A1(net231231), .A2(n12126), .ZN(n17286) );
  NOR3_X2 U12187 ( .A1(nextPC_ex_out[5]), .A2(n11914), .A3(net231915), .ZN(
        n17290) );
  OAI21_X2 U12188 ( .B1(nextPC_ex_out[4]), .B2(net224709), .A(net224710), .ZN(
        net224707) );
  NOR3_X2 U12189 ( .A1(nextPC_ex_out[4]), .A2(n10355), .A3(net224713), .ZN(
        n17285) );
  NOR2_X1 U12190 ( .A1(n12806), .A2(n13377), .ZN(n17334) );
  OAI21_X2 U12191 ( .B1(n13364), .B2(n12894), .A(n12930), .ZN(n17332) );
  AOI222_X2 U12192 ( .A1(n19153), .A2(REG_FILE_reg_out_14__18_), .B1(n13499), 
        .B2(REG_FILE_reg_out_4__18_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__18_), .ZN(n2131) );
  NOR2_X1 U12193 ( .A1(n12808), .A2(n13377), .ZN(n17385) );
  OAI21_X2 U12194 ( .B1(n13364), .B2(n12896), .A(n12931), .ZN(n17383) );
  AOI222_X2 U12195 ( .A1(n19153), .A2(REG_FILE_reg_out_14__19_), .B1(n13499), 
        .B2(REG_FILE_reg_out_4__19_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__19_), .ZN(n2111) );
  INV_X4 U12196 ( .A(net231273), .ZN(net231255) );
  NOR2_X1 U12197 ( .A1(n12810), .A2(n13377), .ZN(n17440) );
  OAI21_X2 U12198 ( .B1(n13364), .B2(n12898), .A(n12932), .ZN(n17438) );
  AOI222_X2 U12199 ( .A1(n19153), .A2(REG_FILE_reg_out_14__20_), .B1(n13498), 
        .B2(REG_FILE_reg_out_4__20_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__20_), .ZN(n2091) );
  NAND3_X2 U12200 ( .A1(n17590), .A2(n17589), .A3(n17588), .ZN(n17742) );
  NOR2_X1 U12201 ( .A1(n12812), .A2(n13377), .ZN(n17625) );
  OAI21_X2 U12202 ( .B1(n13364), .B2(n12900), .A(n12933), .ZN(n17623) );
  AOI222_X2 U12203 ( .A1(n19153), .A2(REG_FILE_reg_out_14__21_), .B1(n13498), 
        .B2(REG_FILE_reg_out_4__21_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__21_), .ZN(n2071) );
  NOR3_X2 U12204 ( .A1(n17647), .A2(n17646), .A3(n17645), .ZN(n17664) );
  NOR3_X2 U12205 ( .A1(n17661), .A2(n17660), .A3(n17659), .ZN(n17662) );
  AOI21_X1 U12206 ( .B1(n15467), .B2(IMEM_BUS_OUT[22]), .A(IMEM_BUS_OUT[21]), 
        .ZN(n15463) );
  NAND3_X1 U12207 ( .A1(n17828), .A2(n10810), .A3(n17827), .ZN(net224173) );
  NOR2_X1 U12208 ( .A1(n12814), .A2(n13377), .ZN(n17778) );
  OAI21_X2 U12209 ( .B1(n12902), .B2(n13365), .A(n12934), .ZN(n17770) );
  AOI222_X2 U12210 ( .A1(n19153), .A2(REG_FILE_reg_out_14__22_), .B1(n13498), 
        .B2(REG_FILE_reg_out_4__22_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__22_), .ZN(n2051) );
  NOR3_X2 U12211 ( .A1(n17807), .A2(n17806), .A3(n17805), .ZN(n17817) );
  NOR3_X2 U12212 ( .A1(n17800), .A2(n17799), .A3(n17798), .ZN(n17818) );
  AOI222_X2 U12213 ( .A1(n19153), .A2(REG_FILE_reg_out_14__23_), .B1(n13498), 
        .B2(REG_FILE_reg_out_4__23_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__23_), .ZN(n2031) );
  NOR3_X2 U12214 ( .A1(n15223), .A2(n15222), .A3(n15221), .ZN(n15224) );
  OAI21_X2 U12215 ( .B1(n12904), .B2(n13365), .A(n12718), .ZN(n15223) );
  NOR2_X2 U12216 ( .A1(n12758), .A2(n13382), .ZN(n15222) );
  NOR2_X1 U12217 ( .A1(n12816), .A2(n13377), .ZN(n15221) );
  NOR3_X2 U12218 ( .A1(n15220), .A2(n15219), .A3(n15218), .ZN(n15225) );
  NOR2_X2 U12219 ( .A1(n10533), .A2(n13371), .ZN(n15219) );
  NOR2_X2 U12220 ( .A1(n11873), .A2(n13373), .ZN(n15218) );
  NOR3_X2 U12221 ( .A1(n15214), .A2(n15213), .A3(n15212), .ZN(n2038) );
  NOR3_X2 U12222 ( .A1(n17956), .A2(n17955), .A3(n17954), .ZN(n17966) );
  NOR3_X2 U12223 ( .A1(n17964), .A2(n17963), .A3(n17962), .ZN(n17965) );
  NOR3_X2 U12224 ( .A1(n17949), .A2(n17948), .A3(n17947), .ZN(n17967) );
  OAI21_X1 U12225 ( .B1(n15470), .B2(IMEM_BUS_OUT[23]), .A(n15469), .ZN(n17973) );
  AOI222_X2 U12226 ( .A1(n19153), .A2(REG_FILE_reg_out_14__24_), .B1(n13498), 
        .B2(REG_FILE_reg_out_4__24_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__24_), .ZN(n2011) );
  NOR3_X2 U12227 ( .A1(n15237), .A2(n15236), .A3(n15235), .ZN(n15238) );
  OAI21_X2 U12228 ( .B1(n12906), .B2(n13365), .A(n12923), .ZN(n15237) );
  NOR2_X2 U12229 ( .A1(n12759), .A2(n13382), .ZN(n15236) );
  NOR2_X1 U12230 ( .A1(n12817), .A2(n13377), .ZN(n15235) );
  NOR3_X2 U12231 ( .A1(n15234), .A2(n15233), .A3(n15232), .ZN(n15239) );
  NOR2_X2 U12232 ( .A1(n10534), .A2(n13371), .ZN(n15233) );
  NOR2_X2 U12233 ( .A1(n11874), .A2(n13373), .ZN(n15232) );
  NOR3_X2 U12234 ( .A1(n15228), .A2(n15227), .A3(n15226), .ZN(n2018) );
  NOR3_X2 U12235 ( .A1(n18046), .A2(n18045), .A3(n18044), .ZN(n18056) );
  NOR3_X2 U12236 ( .A1(n18039), .A2(n18038), .A3(n18037), .ZN(n18057) );
  NOR3_X2 U12237 ( .A1(n18054), .A2(n18053), .A3(n18052), .ZN(n18055) );
  NOR3_X2 U12238 ( .A1(n15248), .A2(n15247), .A3(n15246), .ZN(n15253) );
  NOR2_X2 U12239 ( .A1(n10535), .A2(n13371), .ZN(n15247) );
  NOR2_X2 U12240 ( .A1(n11875), .A2(n13373), .ZN(n15246) );
  NOR3_X2 U12241 ( .A1(n15251), .A2(n15250), .A3(n15249), .ZN(n15252) );
  OAI21_X2 U12242 ( .B1(n12908), .B2(n13365), .A(n12720), .ZN(n15251) );
  NOR2_X2 U12243 ( .A1(n12760), .A2(n13382), .ZN(n15250) );
  NOR2_X1 U12244 ( .A1(n12818), .A2(n13377), .ZN(n15249) );
  AOI222_X2 U12245 ( .A1(n19153), .A2(REG_FILE_reg_out_14__25_), .B1(n13498), 
        .B2(REG_FILE_reg_out_4__25_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__25_), .ZN(n1991) );
  NOR3_X2 U12246 ( .A1(n15245), .A2(n15244), .A3(n15243), .ZN(n1999) );
  NOR3_X2 U12247 ( .A1(n18089), .A2(n18088), .A3(n18087), .ZN(n18099) );
  NOR3_X2 U12248 ( .A1(n18097), .A2(n18096), .A3(n18095), .ZN(n18098) );
  NOR3_X2 U12249 ( .A1(n18082), .A2(n18081), .A3(n18080), .ZN(n18100) );
  INV_X4 U12250 ( .A(net231271), .ZN(net231257) );
  NOR3_X2 U12251 ( .A1(n15263), .A2(n15262), .A3(n15261), .ZN(n15268) );
  NOR2_X2 U12252 ( .A1(n10536), .A2(n13371), .ZN(n15262) );
  NOR2_X2 U12253 ( .A1(n11876), .A2(n13373), .ZN(n15261) );
  NOR3_X2 U12254 ( .A1(n15266), .A2(n15265), .A3(n15264), .ZN(n15267) );
  NOR2_X2 U12255 ( .A1(n12761), .A2(n13382), .ZN(n15265) );
  OAI21_X2 U12256 ( .B1(n12910), .B2(n13364), .A(n12924), .ZN(n15266) );
  NOR2_X1 U12257 ( .A1(n12819), .A2(n13377), .ZN(n15264) );
  AOI222_X2 U12258 ( .A1(n19153), .A2(REG_FILE_reg_out_14__26_), .B1(n13498), 
        .B2(REG_FILE_reg_out_4__26_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__26_), .ZN(n1971) );
  NOR3_X2 U12259 ( .A1(n15260), .A2(n15259), .A3(n15258), .ZN(n1979) );
  NOR3_X2 U12260 ( .A1(n18134), .A2(n18133), .A3(n18132), .ZN(n18144) );
  NOR3_X2 U12261 ( .A1(n18127), .A2(n18126), .A3(n18125), .ZN(n18145) );
  NOR3_X2 U12262 ( .A1(n18142), .A2(n18141), .A3(n18140), .ZN(n18143) );
  NOR3_X2 U12263 ( .A1(n15277), .A2(n15276), .A3(n15275), .ZN(n15282) );
  NOR2_X2 U12264 ( .A1(n10537), .A2(n13371), .ZN(n15276) );
  NOR2_X2 U12265 ( .A1(n11877), .A2(n13373), .ZN(n15275) );
  NOR3_X2 U12266 ( .A1(n15280), .A2(n15279), .A3(n15278), .ZN(n15281) );
  NOR2_X2 U12267 ( .A1(n12762), .A2(n13382), .ZN(n15279) );
  OAI21_X2 U12268 ( .B1(n12912), .B2(n13364), .A(n12925), .ZN(n15280) );
  NOR2_X1 U12269 ( .A1(n12820), .A2(n13377), .ZN(n15278) );
  AOI222_X2 U12270 ( .A1(n19153), .A2(REG_FILE_reg_out_14__27_), .B1(n13498), 
        .B2(REG_FILE_reg_out_4__27_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__27_), .ZN(n1951) );
  NOR3_X2 U12271 ( .A1(n15271), .A2(n15270), .A3(n15269), .ZN(n1958) );
  NOR3_X2 U12272 ( .A1(n18175), .A2(n18174), .A3(n18173), .ZN(n18185) );
  NOR3_X2 U12273 ( .A1(n18168), .A2(n18167), .A3(n18166), .ZN(n18186) );
  NOR3_X2 U12274 ( .A1(n18183), .A2(n18182), .A3(n18181), .ZN(n18184) );
  NOR3_X2 U12275 ( .A1(n15293), .A2(n15292), .A3(n15291), .ZN(n15298) );
  NOR2_X2 U12276 ( .A1(n10538), .A2(n13371), .ZN(n15292) );
  NOR2_X2 U12277 ( .A1(n11878), .A2(n13373), .ZN(n15291) );
  NOR3_X2 U12278 ( .A1(n15296), .A2(n15295), .A3(n15294), .ZN(n15297) );
  NOR2_X2 U12279 ( .A1(n12763), .A2(n13382), .ZN(n15295) );
  OAI21_X2 U12280 ( .B1(n12914), .B2(n13364), .A(n12926), .ZN(n15296) );
  NOR2_X1 U12281 ( .A1(n12821), .A2(n13377), .ZN(n15294) );
  AOI222_X2 U12282 ( .A1(n19153), .A2(REG_FILE_reg_out_14__28_), .B1(n13498), 
        .B2(REG_FILE_reg_out_4__28_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__28_), .ZN(n1930) );
  NOR3_X2 U12283 ( .A1(n15285), .A2(n15284), .A3(n15283), .ZN(n1937) );
  NOR3_X2 U12284 ( .A1(n18220), .A2(n18219), .A3(n18218), .ZN(n18230) );
  NOR3_X2 U12285 ( .A1(n18228), .A2(n18227), .A3(n18226), .ZN(n18229) );
  NOR3_X2 U12286 ( .A1(n18213), .A2(n18212), .A3(n18211), .ZN(n18231) );
  NOR3_X2 U12287 ( .A1(n15307), .A2(n15306), .A3(n15305), .ZN(n15312) );
  NOR2_X2 U12288 ( .A1(n10539), .A2(n13371), .ZN(n15306) );
  NOR2_X2 U12289 ( .A1(n11879), .A2(n13373), .ZN(n15305) );
  NOR3_X2 U12290 ( .A1(n15310), .A2(n15309), .A3(n15308), .ZN(n15311) );
  NOR2_X2 U12291 ( .A1(n12764), .A2(n13382), .ZN(n15309) );
  OAI21_X2 U12292 ( .B1(n12916), .B2(n13364), .A(n12719), .ZN(n15310) );
  NOR2_X1 U12293 ( .A1(n12822), .A2(n13377), .ZN(n15308) );
  AOI222_X2 U12294 ( .A1(n19153), .A2(REG_FILE_reg_out_14__29_), .B1(n13498), 
        .B2(REG_FILE_reg_out_4__29_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__29_), .ZN(n1910) );
  NOR3_X2 U12295 ( .A1(n15301), .A2(n15300), .A3(n15299), .ZN(n1917) );
  NOR3_X2 U12296 ( .A1(n18428), .A2(n18427), .A3(n18426), .ZN(n18438) );
  NOR3_X2 U12297 ( .A1(n18436), .A2(n18435), .A3(n18434), .ZN(n18437) );
  NOR3_X2 U12298 ( .A1(n18421), .A2(n18420), .A3(n18419), .ZN(n18439) );
  INV_X4 U12299 ( .A(net231329), .ZN(net231323) );
  NOR3_X2 U12300 ( .A1(n15321), .A2(n15320), .A3(n15319), .ZN(n15326) );
  NOR2_X2 U12301 ( .A1(n10540), .A2(n13371), .ZN(n15320) );
  NOR2_X2 U12302 ( .A1(n11880), .A2(n13373), .ZN(n15319) );
  NOR3_X2 U12303 ( .A1(n15324), .A2(n15323), .A3(n15322), .ZN(n15325) );
  NOR2_X2 U12304 ( .A1(n12765), .A2(n13382), .ZN(n15323) );
  OAI21_X2 U12305 ( .B1(n12918), .B2(n13364), .A(n12927), .ZN(n15324) );
  NOR2_X1 U12306 ( .A1(n12823), .A2(n13377), .ZN(n15322) );
  AOI222_X2 U12307 ( .A1(n19153), .A2(REG_FILE_reg_out_14__30_), .B1(n13498), 
        .B2(REG_FILE_reg_out_4__30_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__30_), .ZN(n1890) );
  NOR3_X2 U12308 ( .A1(n15315), .A2(n15314), .A3(n15313), .ZN(n1897) );
  NOR3_X2 U12309 ( .A1(n18509), .A2(n18508), .A3(n18507), .ZN(n18519) );
  NOR3_X2 U12310 ( .A1(n18517), .A2(n18516), .A3(n18515), .ZN(n18518) );
  NOR3_X2 U12311 ( .A1(n18501), .A2(n18500), .A3(n18499), .ZN(n18520) );
  INV_X4 U12312 ( .A(net231335), .ZN(net231309) );
  INV_X4 U12313 ( .A(net231337), .ZN(net231303) );
  INV_X4 U12314 ( .A(net231335), .ZN(net231305) );
  INV_X4 U12315 ( .A(net231337), .ZN(net231301) );
  NOR3_X2 U12316 ( .A1(n15342), .A2(n15341), .A3(n15340), .ZN(n15347) );
  NOR2_X2 U12317 ( .A1(n10367), .A2(n13371), .ZN(n15341) );
  NOR2_X2 U12318 ( .A1(n12079), .A2(n13373), .ZN(n15340) );
  NOR3_X2 U12319 ( .A1(n15345), .A2(n15344), .A3(n15343), .ZN(n15346) );
  NOR2_X2 U12320 ( .A1(n12498), .A2(n13382), .ZN(n15344) );
  OAI21_X2 U12321 ( .B1(n12920), .B2(n13364), .A(n12928), .ZN(n15345) );
  NOR2_X1 U12322 ( .A1(n12824), .A2(n13377), .ZN(n15343) );
  AOI222_X2 U12323 ( .A1(n19153), .A2(REG_FILE_reg_out_14__31_), .B1(n13498), 
        .B2(REG_FILE_reg_out_4__31_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__31_), .ZN(n1842) );
  NOR3_X2 U12324 ( .A1(n15333), .A2(n15332), .A3(n15331), .ZN(n1860) );
  NOR3_X1 U12325 ( .A1(n5546), .A2(n18766), .A3(n18781), .ZN(n18767) );
  INV_X4 U12326 ( .A(net231341), .ZN(net231291) );
  INV_X4 U12327 ( .A(net231271), .ZN(net231259) );
  NAND3_X2 U12328 ( .A1(n18774), .A2(net230387), .A3(n18788), .ZN(n18787) );
  INV_X4 U12329 ( .A(reset), .ZN(n13947) );
  INV_X4 U12330 ( .A(reset), .ZN(n13951) );
  INV_X4 U12331 ( .A(net231271), .ZN(net231261) );
  INV_X4 U12332 ( .A(reset), .ZN(n13941) );
  INV_X4 U12333 ( .A(reset), .ZN(n13953) );
  INV_X4 U12334 ( .A(reset), .ZN(n13940) );
  AOI21_X1 U12335 ( .B1(ID_EXEC_OUT[156]), .B2(n13493), .A(n11913), .ZN(n19145) );
  OAI21_X1 U12336 ( .B1(n13480), .B2(n18831), .A(n18830), .ZN(n7971) );
  OAI21_X1 U12337 ( .B1(n13480), .B2(n18815), .A(n18814), .ZN(n7956) );
  OAI21_X1 U12338 ( .B1(n13480), .B2(n18812), .A(n18811), .ZN(n7955) );
  OAI21_X1 U12339 ( .B1(n12033), .B2(net231235), .A(n1266), .ZN(n8002) );
  OAI21_X1 U12340 ( .B1(n12067), .B2(net231211), .A(n1250), .ZN(n8010) );
  OAI21_X1 U12341 ( .B1(n12066), .B2(net231211), .A(n1252), .ZN(n8009) );
  OAI21_X2 U12342 ( .B1(n12031), .B2(net231235), .A(n1256), .ZN(n8007) );
  OAI21_X2 U12343 ( .B1(n12032), .B2(net231233), .A(n1254), .ZN(n8008) );
  OAI21_X1 U12344 ( .B1(n12071), .B2(net231211), .A(n1238), .ZN(n7865) );
  OAI21_X1 U12345 ( .B1(n12068), .B2(net231211), .A(n1244), .ZN(n7868) );
  OAI21_X1 U12346 ( .B1(n12070), .B2(net231211), .A(n1240), .ZN(n7866) );
  OAI21_X1 U12347 ( .B1(n12069), .B2(net231211), .A(n1242), .ZN(n7867) );
  NOR2_X2 U12348 ( .A1(n5520), .A2(n14266), .ZN(n14267) );
  AOI211_X2 U12349 ( .C1(n18644), .C2(n17149), .A(n16825), .B(n16824), .ZN(
        n16826) );
  NOR2_X2 U12350 ( .A1(n18287), .A2(n18286), .ZN(n18288) );
  AOI21_X1 U12351 ( .B1(n17924), .B2(n18367), .A(n18366), .ZN(n18380) );
  OAI21_X1 U12352 ( .B1(n19295), .B2(net231211), .A(n1258), .ZN(n8006) );
  OAI21_X1 U12353 ( .B1(n19298), .B2(net231235), .A(n1264), .ZN(n8003) );
  OAI21_X2 U12354 ( .B1(n19296), .B2(net231233), .A(n1260), .ZN(n8005) );
  AOI21_X2 U12355 ( .B1(n18465), .B2(n18360), .A(n18464), .ZN(n18479) );
  NOR2_X2 U12356 ( .A1(n18391), .A2(n18390), .ZN(n18403) );
  OAI21_X1 U12357 ( .B1(n13480), .B2(n18827), .A(n18826), .ZN(n7965) );
  NOR2_X2 U12358 ( .A1(n16418), .A2(n16417), .ZN(n16424) );
  AOI211_X2 U12359 ( .C1(n19118), .C2(n16422), .A(n16421), .B(n16420), .ZN(
        n16423) );
  OAI21_X1 U12360 ( .B1(n13480), .B2(n18823), .A(n18822), .ZN(n7962) );
  OAI21_X1 U12361 ( .B1(n13480), .B2(n18819), .A(n18818), .ZN(n7959) );
  OAI21_X1 U12362 ( .B1(n13480), .B2(n18807), .A(n18806), .ZN(n7951) );
  AOI211_X2 U12363 ( .C1(n17924), .C2(n18368), .A(n18353), .B(n18352), .ZN(
        n18354) );
  OAI21_X2 U12364 ( .B1(net137549), .B2(net231211), .A(n18832), .ZN(n7973) );
  OAI21_X2 U12365 ( .B1(n19299), .B2(net231235), .A(n1270), .ZN(n8001) );
  OAI21_X2 U12366 ( .B1(net230379), .B2(n18763), .A(n18762), .ZN(n7840) );
  OAI21_X1 U12367 ( .B1(n13480), .B2(n18803), .A(n18802), .ZN(n7948) );
  OAI21_X1 U12368 ( .B1(n13480), .B2(n18809), .A(n18808), .ZN(n7954) );
  NOR2_X2 U12369 ( .A1(n13956), .A2(n7286), .ZN(EXEC_STAGE_mul_ex_N16) );
  AOI21_X2 U12370 ( .B1(n7284), .B2(n7288), .A(n13956), .ZN(
        EXEC_STAGE_mul_ex_N15) );
  NOR2_X2 U12371 ( .A1(n7291), .A2(n13955), .ZN(EXEC_STAGE_mul_ex_N14) );
  AOI21_X2 U12372 ( .B1(n7289), .B2(EXEC_MEM_IN_250), .A(n13541), .ZN(n7291)
         );
  NOR2_X2 U12373 ( .A1(n2602), .A2(n2603), .ZN(n2567) );
  NOR2_X2 U12374 ( .A1(n3685), .A2(n3686), .ZN(n3656) );
  NOR2_X2 U12375 ( .A1(n2855), .A2(n2856), .ZN(n2837) );
  NOR3_X2 U12376 ( .A1(n14561), .A2(n14560), .A3(n14559), .ZN(n3940) );
  NOR2_X2 U12377 ( .A1(n3957), .A2(n3958), .ZN(n3942) );
  NOR2_X2 U12378 ( .A1(n2890), .A2(n2891), .ZN(n2872) );
  NOR3_X2 U12379 ( .A1(n14550), .A2(n14549), .A3(n14548), .ZN(n3969) );
  NOR2_X2 U12380 ( .A1(n3986), .A2(n3987), .ZN(n3971) );
  NOR2_X2 U12381 ( .A1(n3026), .A2(n3027), .ZN(n3008) );
  NOR3_X2 U12382 ( .A1(n14506), .A2(n14505), .A3(n14504), .ZN(n4085) );
  NOR2_X2 U12383 ( .A1(n4102), .A2(n4103), .ZN(n4087) );
  NOR2_X2 U12384 ( .A1(n2924), .A2(n2925), .ZN(n2906) );
  NOR3_X2 U12385 ( .A1(n14539), .A2(n14538), .A3(n14537), .ZN(n3998) );
  NOR2_X2 U12386 ( .A1(n4015), .A2(n4016), .ZN(n4000) );
  NOR2_X2 U12387 ( .A1(n2958), .A2(n2959), .ZN(n2940) );
  NOR2_X2 U12388 ( .A1(n2992), .A2(n2993), .ZN(n2974) );
  NOR2_X2 U12389 ( .A1(n3537), .A2(n3538), .ZN(n3519) );
  NOR3_X2 U12390 ( .A1(n14340), .A2(n14339), .A3(n14338), .ZN(n4522) );
  OAI21_X2 U12391 ( .B1(n15565), .B2(n15564), .A(n15563), .ZN(n15580) );
  NOR2_X2 U12392 ( .A1(n13492), .A2(n15932), .ZN(n15933) );
  NOR2_X2 U12393 ( .A1(n3094), .A2(n3095), .ZN(n3076) );
  NOR3_X2 U12394 ( .A1(n14484), .A2(n14483), .A3(n14482), .ZN(n4143) );
  NOR2_X2 U12395 ( .A1(n4160), .A2(n4161), .ZN(n4145) );
  NOR2_X2 U12396 ( .A1(n3367), .A2(n3368), .ZN(n3349) );
  NOR3_X2 U12397 ( .A1(n14395), .A2(n14394), .A3(n14393), .ZN(n4376) );
  NOR2_X2 U12398 ( .A1(n3265), .A2(n3266), .ZN(n3247) );
  NOR3_X2 U12399 ( .A1(n14429), .A2(n14428), .A3(n14427), .ZN(n4289) );
  NOR2_X2 U12400 ( .A1(n4306), .A2(n4307), .ZN(n4291) );
  NOR2_X2 U12401 ( .A1(n3469), .A2(n3470), .ZN(n3451) );
  NOR3_X2 U12402 ( .A1(n14362), .A2(n14361), .A3(n14360), .ZN(n4463) );
  NOR2_X2 U12403 ( .A1(n3503), .A2(n3504), .ZN(n3485) );
  AOI21_X2 U12404 ( .B1(ID_EXEC_OUT[209]), .B2(n13216), .A(n16006), .ZN(n16041) );
  NOR3_X2 U12405 ( .A1(n16039), .A2(n16038), .A3(n16037), .ZN(n16040) );
  AOI21_X2 U12406 ( .B1(n13492), .B2(n16005), .A(n16004), .ZN(n16042) );
  NOR2_X2 U12407 ( .A1(n2393), .A2(n2392), .ZN(n16138) );
  AOI211_X1 U12408 ( .C1(n17924), .C2(n16157), .A(n16156), .B(n16155), .ZN(
        n16158) );
  NOR2_X2 U12409 ( .A1(n3401), .A2(n3402), .ZN(n3383) );
  NOR3_X2 U12410 ( .A1(n14384), .A2(n14383), .A3(n14382), .ZN(n4405) );
  NOR3_X2 U12411 ( .A1(n16218), .A2(n16217), .A3(n16216), .ZN(n16231) );
  NOR2_X2 U12412 ( .A1(n3333), .A2(n3334), .ZN(n3315) );
  NOR3_X2 U12413 ( .A1(n14407), .A2(n14406), .A3(n14405), .ZN(n4347) );
  NOR2_X2 U12414 ( .A1(n2312), .A2(n2311), .ZN(n16287) );
  NOR2_X2 U12415 ( .A1(n3299), .A2(n3300), .ZN(n3281) );
  NOR3_X2 U12416 ( .A1(n14418), .A2(n14417), .A3(n14416), .ZN(n4318) );
  NOR2_X2 U12417 ( .A1(n4335), .A2(n4336), .ZN(n4320) );
  NOR2_X2 U12418 ( .A1(n2292), .A2(n2291), .ZN(n16386) );
  NOR2_X2 U12419 ( .A1(n3435), .A2(n3436), .ZN(n3417) );
  NOR3_X2 U12420 ( .A1(n14373), .A2(n14372), .A3(n14371), .ZN(n4434) );
  NOR2_X2 U12421 ( .A1(n3128), .A2(n3129), .ZN(n3110) );
  NOR3_X2 U12422 ( .A1(n14473), .A2(n14472), .A3(n14471), .ZN(n4172) );
  NOR2_X2 U12423 ( .A1(n4189), .A2(n4190), .ZN(n4174) );
  NOR2_X2 U12424 ( .A1(n2252), .A2(n2251), .ZN(n16614) );
  NOR2_X2 U12425 ( .A1(n2212), .A2(n2211), .ZN(n16719) );
  NOR2_X2 U12426 ( .A1(n3606), .A2(n3607), .ZN(n3588) );
  NOR3_X2 U12427 ( .A1(n14318), .A2(n14317), .A3(n14316), .ZN(n4580) );
  NOR2_X2 U12428 ( .A1(n2453), .A2(n2452), .ZN(n16954) );
  AOI21_X1 U12429 ( .B1(net231615), .B2(n19038), .A(n16964), .ZN(n16965) );
  NOR2_X2 U12430 ( .A1(n2332), .A2(n2331), .ZN(n17028) );
  OAI221_X2 U12431 ( .B1(net231227), .B2(n10946), .C1(n17035), .C2(net231915), 
        .A(n17034), .ZN(n7517) );
  OAI21_X1 U12432 ( .B1(n17048), .B2(n17047), .A(n19012), .ZN(n17064) );
  AOI211_X2 U12433 ( .C1(n18360), .C2(n17149), .A(n17148), .B(n17147), .ZN(
        n17150) );
  AOI21_X2 U12434 ( .B1(n19118), .B2(n17145), .A(n17144), .ZN(n17151) );
  NOR2_X2 U12435 ( .A1(n3640), .A2(n3641), .ZN(n3622) );
  NOR3_X2 U12436 ( .A1(n14307), .A2(n14306), .A3(n14305), .ZN(n4609) );
  AOI21_X1 U12437 ( .B1(net231615), .B2(n18873), .A(n17195), .ZN(n17210) );
  NOR2_X2 U12438 ( .A1(n2433), .A2(n2432), .ZN(n17281) );
  INV_X4 U12439 ( .A(n13943), .ZN(n13888) );
  AOI211_X2 U12440 ( .C1(n18644), .C2(n17322), .A(n17321), .B(n17320), .ZN(
        n17323) );
  AOI21_X2 U12441 ( .B1(ID_EXEC_OUT[224]), .B2(n13216), .A(n17508), .ZN(n17554) );
  NOR2_X2 U12442 ( .A1(n3572), .A2(n3573), .ZN(n3554) );
  NOR3_X2 U12443 ( .A1(n14329), .A2(n14328), .A3(n14327), .ZN(n4551) );
  OAI21_X2 U12444 ( .B1(n17573), .B2(n13213), .A(n17572), .ZN(n17579) );
  NOR2_X2 U12445 ( .A1(n3231), .A2(n3232), .ZN(n3213) );
  NOR3_X2 U12446 ( .A1(n14440), .A2(n14439), .A3(n14438), .ZN(n4260) );
  NOR2_X2 U12447 ( .A1(n4277), .A2(n4278), .ZN(n4262) );
  INV_X4 U12448 ( .A(n13951), .ZN(n13921) );
  AOI211_X2 U12449 ( .C1(n17692), .C2(n18985), .A(n17691), .B(n17690), .ZN(
        n17718) );
  NOR2_X2 U12450 ( .A1(n3196), .A2(n3197), .ZN(n3178) );
  NOR3_X2 U12451 ( .A1(n14451), .A2(n14450), .A3(n14449), .ZN(n4231) );
  NOR2_X2 U12452 ( .A1(n4248), .A2(n4249), .ZN(n4233) );
  AOI211_X2 U12453 ( .C1(n13490), .C2(n18852), .A(n17763), .B(n17762), .ZN(
        n17764) );
  NOR3_X2 U12454 ( .A1(n17862), .A2(n17861), .A3(n17860), .ZN(n17863) );
  NOR2_X2 U12455 ( .A1(n3162), .A2(n3163), .ZN(n3144) );
  NOR3_X2 U12456 ( .A1(n14462), .A2(n14461), .A3(n14460), .ZN(n4202) );
  NOR2_X2 U12457 ( .A1(n4219), .A2(n4220), .ZN(n4204) );
  AOI21_X2 U12458 ( .B1(n17900), .B2(n17899), .A(n17898), .ZN(n17902) );
  AOI211_X2 U12459 ( .C1(n13490), .C2(n18014), .A(n18013), .B(n18012), .ZN(
        n18015) );
  NOR2_X2 U12460 ( .A1(n2719), .A2(n2720), .ZN(n2701) );
  NOR3_X2 U12461 ( .A1(n14605), .A2(n14604), .A3(n14603), .ZN(n3823) );
  NOR2_X2 U12462 ( .A1(n3840), .A2(n3841), .ZN(n3825) );
  NOR2_X2 U12463 ( .A1(n2787), .A2(n2788), .ZN(n2769) );
  NOR3_X2 U12464 ( .A1(n14583), .A2(n14582), .A3(n14581), .ZN(n3881) );
  NOR2_X2 U12465 ( .A1(n3898), .A2(n3899), .ZN(n3883) );
  NOR2_X2 U12466 ( .A1(n2753), .A2(n2754), .ZN(n2735) );
  NOR3_X2 U12467 ( .A1(n14594), .A2(n14593), .A3(n14592), .ZN(n3852) );
  NOR2_X2 U12468 ( .A1(n3869), .A2(n3870), .ZN(n3854) );
  NOR2_X2 U12469 ( .A1(n2821), .A2(n2822), .ZN(n2803) );
  NOR3_X2 U12470 ( .A1(n14572), .A2(n14571), .A3(n14570), .ZN(n3911) );
  NOR2_X2 U12471 ( .A1(n3928), .A2(n3929), .ZN(n3913) );
  NOR2_X2 U12472 ( .A1(n2685), .A2(n2686), .ZN(n2667) );
  NOR3_X2 U12473 ( .A1(n14616), .A2(n14615), .A3(n14614), .ZN(n3794) );
  NOR2_X2 U12474 ( .A1(n3811), .A2(n3812), .ZN(n3796) );
  NOR2_X2 U12475 ( .A1(n2651), .A2(n2652), .ZN(n2633) );
  NOR3_X2 U12476 ( .A1(n14627), .A2(n14626), .A3(n14625), .ZN(n3765) );
  NOR2_X2 U12477 ( .A1(n3782), .A2(n3783), .ZN(n3767) );
  AOI21_X1 U12478 ( .B1(n19107), .B2(n18531), .A(n18530), .ZN(n18555) );
  AOI211_X1 U12479 ( .C1(n17924), .C2(n19117), .A(n18553), .B(n18552), .ZN(
        n18554) );
  NOR2_X2 U12480 ( .A1(n3060), .A2(n3061), .ZN(n3042) );
  NOR3_X2 U12481 ( .A1(n14495), .A2(n14494), .A3(n14493), .ZN(n4114) );
  NOR2_X2 U12482 ( .A1(n4131), .A2(n4132), .ZN(n4116) );
  INV_X4 U12483 ( .A(n13947), .ZN(n13900) );
  AOI21_X1 U12484 ( .B1(n17924), .B2(n18575), .A(n18574), .ZN(n18583) );
  NOR2_X2 U12485 ( .A1(n18682), .A2(n18681), .ZN(n18683) );
  INV_X4 U12486 ( .A(n13944), .ZN(n13894) );
  NOR3_X2 U12487 ( .A1(n14296), .A2(n14295), .A3(n14294), .ZN(n4638) );
  INV_X4 U12488 ( .A(n13946), .ZN(n13899) );
  INV_X4 U12489 ( .A(n13941), .ZN(n13883) );
  INV_X4 U12490 ( .A(n13947), .ZN(n13901) );
  INV_X4 U12491 ( .A(n13949), .ZN(n13915) );
  INV_X4 U12492 ( .A(n13944), .ZN(n13926) );
  INV_X4 U12493 ( .A(n13943), .ZN(n13893) );
  INV_X4 U12494 ( .A(n13946), .ZN(n13898) );
  NAND3_X2 U12495 ( .A1(n18750), .A2(n18749), .A3(n18748), .ZN(n7834) );
  NOR3_X2 U12496 ( .A1(n12569), .A2(n14253), .A3(n14252), .ZN(n5499) );
  NOR3_X2 U12497 ( .A1(n5516), .A2(n5478), .A3(n5484), .ZN(n5518) );
  INV_X4 U12498 ( .A(n13945), .ZN(n13896) );
  OAI21_X2 U12499 ( .B1(net231245), .B2(n12052), .A(n5535), .ZN(n7846) );
  NAND3_X2 U12500 ( .A1(n10359), .A2(n12129), .A3(n12133), .ZN(n18765) );
  OAI21_X2 U12501 ( .B1(n12050), .B2(net231233), .A(n1236), .ZN(n7864) );
  OAI21_X2 U12502 ( .B1(n10906), .B2(net231211), .A(n12219), .ZN(n7869) );
  OAI21_X2 U12503 ( .B1(net231245), .B2(n12051), .A(n5555), .ZN(n7872) );
  NOR2_X2 U12504 ( .A1(n14214), .A2(n14213), .ZN(n14215) );
  OAI21_X2 U12505 ( .B1(net231245), .B2(n19318), .A(n5549), .ZN(n7877) );
  AOI21_X2 U12506 ( .B1(n10359), .B2(n18784), .A(n18783), .ZN(n18785) );
  NOR2_X2 U12507 ( .A1(n12064), .A2(net231241), .ZN(n18783) );
  OAI21_X2 U12508 ( .B1(n10933), .B2(net231211), .A(n18789), .ZN(n7905) );
  NAND3_X2 U12509 ( .A1(n18788), .A2(n12129), .A3(n10359), .ZN(n18789) );
  INV_X4 U12510 ( .A(n13948), .ZN(n13924) );
  OAI21_X2 U12511 ( .B1(net231245), .B2(n10939), .A(n2555), .ZN(n7918) );
  INV_X4 U12512 ( .A(n13941), .ZN(n13884) );
  OAI21_X2 U12513 ( .B1(net231245), .B2(n10938), .A(n2557), .ZN(n7924) );
  OAI21_X2 U12514 ( .B1(net231245), .B2(n10937), .A(n2559), .ZN(n7930) );
  OAI21_X2 U12515 ( .B1(net231245), .B2(n12551), .A(n2559), .ZN(n7931) );
  OAI21_X2 U12516 ( .B1(net231233), .B2(n12072), .A(n2559), .ZN(n7932) );
  INV_X4 U12517 ( .A(n13952), .ZN(n13925) );
  INV_X4 U12518 ( .A(n13947), .ZN(n13902) );
  INV_X4 U12519 ( .A(n13951), .ZN(n13920) );
  OAI21_X2 U12520 ( .B1(net231245), .B2(n10936), .A(n2562), .ZN(n7936) );
  INV_X4 U12521 ( .A(n13951), .ZN(n13919) );
  OAI21_X2 U12522 ( .B1(net231245), .B2(n12058), .A(n2564), .ZN(n7940) );
  INV_X4 U12523 ( .A(n13942), .ZN(n13892) );
  OAI21_X2 U12524 ( .B1(net231245), .B2(n10935), .A(n2564), .ZN(n7944) );
  OAI21_X2 U12525 ( .B1(n12065), .B2(net231211), .A(n18801), .ZN(n7946) );
  INV_X4 U12526 ( .A(n13942), .ZN(n13916) );
  OAI21_X2 U12527 ( .B1(n12054), .B2(net231211), .A(n18805), .ZN(n7949) );
  OAI21_X2 U12528 ( .B1(n12055), .B2(net231211), .A(n18817), .ZN(n7957) );
  INV_X4 U12529 ( .A(n13941), .ZN(n13885) );
  OAI21_X2 U12530 ( .B1(n12056), .B2(net231235), .A(n18821), .ZN(n7960) );
  OAI21_X2 U12531 ( .B1(n12057), .B2(net231211), .A(n18825), .ZN(n7963) );
  INV_X4 U12532 ( .A(n13948), .ZN(n13922) );
  INV_X4 U12533 ( .A(n13945), .ZN(n13897) );
  INV_X4 U12534 ( .A(n13952), .ZN(n13931) );
  OAI21_X2 U12535 ( .B1(n19297), .B2(net231237), .A(n1262), .ZN(n8004) );
  OAI21_X2 U12536 ( .B1(n19294), .B2(net231235), .A(n1248), .ZN(n8011) );
  INV_X4 U12537 ( .A(n13940), .ZN(n13881) );
  INV_X4 U12538 ( .A(n13953), .ZN(n13932) );
  INV_X4 U12539 ( .A(n13949), .ZN(n13891) );
  NOR2_X2 U12540 ( .A1(n6892), .A2(n6893), .ZN(n6891) );
  INV_X4 U12541 ( .A(n13940), .ZN(n13882) );
  INV_X4 U12542 ( .A(n13950), .ZN(n13914) );
  NOR3_X2 U12543 ( .A1(n14640), .A2(n14639), .A3(n14638), .ZN(n3704) );
  NOR2_X2 U12544 ( .A1(n3738), .A2(n3739), .ZN(n3706) );
  INV_X4 U12545 ( .A(net239630), .ZN(net239631) );
  INV_X1 U12546 ( .A(net227219), .ZN(net239815) );
  OAI22_X1 U12547 ( .A1(net231245), .A2(net239744), .B1(n12300), .B2(net230379), .ZN(n7991) );
  NAND3_X4 U12548 ( .A1(net223442), .A2(net227259), .A3(net227248), .ZN(
        net227245) );
  INV_X4 U12549 ( .A(net224699), .ZN(net239673) );
  NAND2_X4 U12550 ( .A1(net223666), .A2(net239761), .ZN(net227189) );
  XNOR2_X2 U12551 ( .A(n10149), .B(net239083), .ZN(n15531) );
  INV_X8 U12552 ( .A(net227200), .ZN(net233180) );
  NAND2_X2 U12553 ( .A1(nextPC_ex_out[26]), .A2(n10148), .ZN(net239533) );
  OAI21_X2 U12554 ( .B1(net227156), .B2(net227157), .A(net227158), .ZN(
        net227137) );
  NAND3_X4 U12555 ( .A1(n13006), .A2(net227220), .A3(net227219), .ZN(net227200) );
  INV_X4 U12556 ( .A(net231313), .ZN(net231337) );
  INV_X4 U12557 ( .A(net231333), .ZN(net231311) );
  INV_X4 U12558 ( .A(net231333), .ZN(net231315) );
  INV_X4 U12559 ( .A(net230403), .ZN(net230399) );
  INV_X8 U12560 ( .A(net230399), .ZN(net230393) );
  INV_X4 U12561 ( .A(net231353), .ZN(net231341) );
  INV_X4 U12562 ( .A(net231277), .ZN(net231241) );
  INV_X4 U12563 ( .A(net231279), .ZN(net231233) );
  INV_X4 U12564 ( .A(net231279), .ZN(net231237) );
  INV_X4 U12565 ( .A(reset), .ZN(n13945) );
  INV_X4 U12566 ( .A(n13942), .ZN(n13887) );
  INV_X4 U12567 ( .A(n13942), .ZN(n13913) );
  INV_X4 U12568 ( .A(reset), .ZN(n13946) );
  INV_X4 U12569 ( .A(n13942), .ZN(n13886) );
  INV_X4 U12570 ( .A(n13942), .ZN(n13912) );
  INV_X4 U12571 ( .A(net231275), .ZN(net231249) );
  INV_X4 U12572 ( .A(net231277), .ZN(net231239) );
  INV_X4 U12573 ( .A(net231341), .ZN(net231289) );
  INV_X4 U12574 ( .A(net231283), .ZN(net231221) );
  INV_X4 U12575 ( .A(net231275), .ZN(net231245) );
  INV_X4 U12576 ( .A(reset), .ZN(n13942) );
  INV_X4 U12577 ( .A(n13949), .ZN(n13918) );
  INV_X4 U12578 ( .A(n13949), .ZN(n13917) );
  INV_X4 U12579 ( .A(net231345), .ZN(net231275) );
  INV_X4 U12580 ( .A(net231345), .ZN(net231279) );
  INV_X4 U12581 ( .A(n13950), .ZN(n13889) );
  INV_X4 U12582 ( .A(n13950), .ZN(n13907) );
  INV_X8 U12583 ( .A(n13215), .ZN(n18360) );
  INV_X4 U12584 ( .A(net231283), .ZN(net231227) );
  INV_X4 U12585 ( .A(n13949), .ZN(n13906) );
  INV_X4 U12586 ( .A(n13949), .ZN(n13905) );
  INV_X4 U12587 ( .A(n13943), .ZN(n13890) );
  INV_X2 U12588 ( .A(net230399), .ZN(net230387) );
  INV_X4 U12589 ( .A(net231283), .ZN(net231223) );
  INV_X4 U12590 ( .A(net231275), .ZN(net231247) );
  INV_X4 U12591 ( .A(net231279), .ZN(net231211) );
  OAI21_X2 U12592 ( .B1(n5662), .B2(n5676), .A(n13934), .ZN(n5729) );
  OAI21_X2 U12593 ( .B1(n5662), .B2(n5724), .A(n13934), .ZN(n5727) );
  OAI21_X2 U12594 ( .B1(n5668), .B2(n5724), .A(n13934), .ZN(n5723) );
  OAI21_X2 U12595 ( .B1(n5662), .B2(n5669), .A(n13935), .ZN(n5673) );
  OAI21_X2 U12596 ( .B1(n5668), .B2(n5669), .A(n13935), .ZN(n5667) );
  OAI21_X2 U12597 ( .B1(n5718), .B2(n5816), .A(n13933), .ZN(n5891) );
  AND2_X4 U12598 ( .A1(n14644), .A2(n18813), .ZN(n10160) );
  INV_X4 U12599 ( .A(net230387), .ZN(net230383) );
  INV_X4 U12600 ( .A(net230387), .ZN(net230381) );
  AND2_X4 U12601 ( .A1(n14647), .A2(n10824), .ZN(n10161) );
  NAND2_X2 U12602 ( .A1(ID_EXEC_OUT[275]), .A2(net230393), .ZN(n19114) );
  INV_X4 U12603 ( .A(net231275), .ZN(net231217) );
  INV_X4 U12604 ( .A(net231275), .ZN(net231231) );
  INV_X4 U12605 ( .A(net231283), .ZN(net231225) );
  INV_X4 U12606 ( .A(reset), .ZN(n13949) );
  INV_X4 U12607 ( .A(n13952), .ZN(n13929) );
  INV_X4 U12608 ( .A(n13944), .ZN(n13895) );
  INV_X4 U12609 ( .A(n13949), .ZN(n13923) );
  NAND2_X4 U12610 ( .A1(n164), .A2(n10262), .ZN(n10162) );
  NAND2_X4 U12611 ( .A1(n10258), .A2(n94), .ZN(n10163) );
  NAND2_X4 U12612 ( .A1(n10322), .A2(n129), .ZN(n10164) );
  NAND2_X4 U12613 ( .A1(n10323), .A2(n164), .ZN(n10165) );
  NAND2_X4 U12614 ( .A1(n200), .A2(n10259), .ZN(n10166) );
  NAND2_X4 U12615 ( .A1(n164), .A2(n10259), .ZN(n10167) );
  OAI21_X2 U12616 ( .B1(n5770), .B2(n5812), .A(n13932), .ZN(n5905) );
  OAI21_X2 U12617 ( .B1(n5680), .B2(n5812), .A(n13933), .ZN(n5888) );
  OAI21_X2 U12618 ( .B1(n5676), .B2(n5812), .A(n13932), .ZN(n5910) );
  OAI21_X2 U12619 ( .B1(n5663), .B2(n5816), .A(n13932), .ZN(n5907) );
  OAI21_X2 U12620 ( .B1(n5764), .B2(n5812), .A(n13933), .ZN(n5901) );
  OAI21_X2 U12621 ( .B1(n5764), .B2(n5816), .A(n13933), .ZN(n5899) );
  OAI21_X2 U12622 ( .B1(n5724), .B2(n5812), .A(n13933), .ZN(n5897) );
  OAI21_X2 U12623 ( .B1(n5724), .B2(n5816), .A(n13933), .ZN(n5895) );
  OAI21_X2 U12624 ( .B1(n5718), .B2(n5812), .A(n13933), .ZN(n5893) );
  OAI21_X2 U12625 ( .B1(n5676), .B2(n5816), .A(n13933), .ZN(n5886) );
  OAI21_X2 U12626 ( .B1(n5669), .B2(n5812), .A(n13933), .ZN(n5818) );
  OAI21_X2 U12627 ( .B1(n5669), .B2(n5816), .A(n13933), .ZN(n5813) );
  OAI21_X2 U12628 ( .B1(n5663), .B2(n5812), .A(n13934), .ZN(n5777) );
  INV_X8 U12629 ( .A(n13466), .ZN(n13465) );
  INV_X4 U12630 ( .A(n11952), .ZN(n13287) );
  INV_X4 U12631 ( .A(n11952), .ZN(n13286) );
  INV_X4 U12632 ( .A(n11997), .ZN(n13285) );
  INV_X4 U12633 ( .A(n11997), .ZN(n13284) );
  INV_X4 U12634 ( .A(n12004), .ZN(n13329) );
  INV_X4 U12635 ( .A(n12004), .ZN(n13328) );
  INV_X4 U12636 ( .A(n12010), .ZN(n13353) );
  INV_X4 U12637 ( .A(n12010), .ZN(n13352) );
  AND3_X4 U12638 ( .A1(offset_26_id[8]), .A2(n12953), .A3(n12984), .ZN(n10197)
         );
  OR3_X1 U12639 ( .A1(EXEC_MEM_OUT_141), .A2(ID_EXEC_OUT[276]), .A3(net231289), 
        .ZN(n10198) );
  INV_X8 U12640 ( .A(n18677), .ZN(n13210) );
  INV_X4 U12641 ( .A(n14103), .ZN(n14019) );
  AND2_X2 U12642 ( .A1(n15728), .A2(n11913), .ZN(n10199) );
  INV_X1 U12643 ( .A(net231361), .ZN(net231357) );
  INV_X4 U12644 ( .A(net139963), .ZN(net231361) );
  INV_X4 U12645 ( .A(net231345), .ZN(net231283) );
  AND2_X2 U12646 ( .A1(n10199), .A2(n18651), .ZN(n10235) );
  INV_X4 U12647 ( .A(reset), .ZN(n13943) );
  INV_X4 U12648 ( .A(n13948), .ZN(n13911) );
  INV_X4 U12649 ( .A(n13948), .ZN(n13904) );
  INV_X4 U12650 ( .A(n13948), .ZN(n13903) );
  INV_X4 U12651 ( .A(n13439), .ZN(n13438) );
  AND3_X4 U12652 ( .A1(offset_26_id[9]), .A2(offset_26_id[8]), .A3(n13220), 
        .ZN(n10241) );
  INV_X4 U12653 ( .A(n11946), .ZN(n13289) );
  INV_X4 U12654 ( .A(n11946), .ZN(n13288) );
  INV_X4 U12655 ( .A(n11951), .ZN(n13291) );
  INV_X4 U12656 ( .A(n11951), .ZN(n13290) );
  INV_X4 U12657 ( .A(n11953), .ZN(n13297) );
  INV_X4 U12658 ( .A(n11953), .ZN(n13296) );
  INV_X4 U12659 ( .A(n11954), .ZN(n13299) );
  INV_X4 U12660 ( .A(n11954), .ZN(n13298) );
  INV_X4 U12661 ( .A(n11978), .ZN(n13295) );
  INV_X4 U12662 ( .A(n11978), .ZN(n13294) );
  INV_X4 U12663 ( .A(n11979), .ZN(n13301) );
  INV_X4 U12664 ( .A(n11979), .ZN(n13300) );
  INV_X4 U12665 ( .A(n11948), .ZN(n13293) );
  INV_X4 U12666 ( .A(n11948), .ZN(n13292) );
  INV_X4 U12667 ( .A(n11988), .ZN(n13303) );
  INV_X4 U12668 ( .A(n11988), .ZN(n13302) );
  INV_X4 U12669 ( .A(n11999), .ZN(n13315) );
  INV_X4 U12670 ( .A(n11999), .ZN(n13314) );
  INV_X4 U12671 ( .A(n12000), .ZN(n13321) );
  INV_X4 U12672 ( .A(n12000), .ZN(n13320) );
  INV_X4 U12673 ( .A(n12001), .ZN(n13323) );
  INV_X4 U12674 ( .A(n12001), .ZN(n13322) );
  INV_X4 U12675 ( .A(n12003), .ZN(n13327) );
  INV_X4 U12676 ( .A(n12003), .ZN(n13326) );
  INV_X4 U12677 ( .A(n12002), .ZN(n13325) );
  INV_X4 U12678 ( .A(n12002), .ZN(n13324) );
  INV_X4 U12679 ( .A(n12005), .ZN(n13333) );
  INV_X4 U12680 ( .A(n12005), .ZN(n13332) );
  INV_X4 U12681 ( .A(n11925), .ZN(n13335) );
  INV_X4 U12682 ( .A(n11925), .ZN(n13334) );
  INV_X4 U12683 ( .A(n12006), .ZN(n13337) );
  INV_X4 U12684 ( .A(n12006), .ZN(n13336) );
  INV_X4 U12685 ( .A(n11926), .ZN(n13343) );
  INV_X4 U12686 ( .A(n11926), .ZN(n13342) );
  INV_X4 U12687 ( .A(n12009), .ZN(n13348) );
  INV_X4 U12688 ( .A(n12009), .ZN(n13347) );
  INV_X4 U12689 ( .A(n12008), .ZN(n13341) );
  INV_X4 U12690 ( .A(n12008), .ZN(n13340) );
  INV_X4 U12691 ( .A(n11924), .ZN(n13330) );
  INV_X4 U12692 ( .A(n11924), .ZN(n13331) );
  INV_X4 U12693 ( .A(n12007), .ZN(n13339) );
  INV_X4 U12694 ( .A(n12007), .ZN(n13338) );
  AND3_X4 U12695 ( .A1(n13220), .A2(n12982), .A3(n12984), .ZN(n10244) );
  INV_X16 U12697 ( .A(n13355), .ZN(n13354) );
  INV_X4 U12698 ( .A(n15490), .ZN(n13355) );
  INV_X4 U12699 ( .A(n11974), .ZN(n13787) );
  INV_X4 U12700 ( .A(n11974), .ZN(n13786) );
  INV_X4 U12701 ( .A(n11984), .ZN(n13442) );
  INV_X4 U12702 ( .A(n11984), .ZN(n13443) );
  INV_X4 U12703 ( .A(n11923), .ZN(n13306) );
  INV_X4 U12704 ( .A(n11923), .ZN(n13307) );
  AND2_X4 U12705 ( .A1(n15354), .A2(n15349), .ZN(n10258) );
  AND2_X4 U12706 ( .A1(n12274), .A2(n15354), .ZN(n10259) );
  AND2_X4 U12707 ( .A1(n15349), .A2(n10837), .ZN(n10262) );
  AND2_X4 U12708 ( .A1(n15351), .A2(n10837), .ZN(n10322) );
  AND2_X4 U12709 ( .A1(n15353), .A2(n15354), .ZN(n10323) );
  INV_X16 U12710 ( .A(n13483), .ZN(n13480) );
  INV_X4 U12711 ( .A(n18532), .ZN(n16207) );
  OAI22_X2 U12712 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[156]), .B1(
        MEM_WB_OUT[124]), .B2(n12978), .ZN(n5808) );
  OAI22_X2 U12713 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[157]), .B1(
        MEM_WB_OUT[125]), .B2(n12978), .ZN(n5807) );
  OAI22_X2 U12714 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[158]), .B1(
        MEM_WB_OUT[126]), .B2(n12978), .ZN(n5806) );
  OAI22_X2 U12715 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[159]), .B1(
        MEM_WB_OUT[127]), .B2(n12978), .ZN(n5805) );
  OAI22_X2 U12716 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[160]), .B1(
        MEM_WB_OUT[128]), .B2(n12978), .ZN(n5804) );
  OAI22_X2 U12717 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[162]), .B1(
        MEM_WB_OUT[130]), .B2(n12978), .ZN(n5802) );
  OAI22_X2 U12718 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[163]), .B1(
        MEM_WB_OUT[131]), .B2(n12978), .ZN(n5801) );
  OAI22_X2 U12719 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[146]), .B1(
        MEM_WB_OUT[114]), .B2(n12978), .ZN(n5799) );
  OAI22_X2 U12720 ( .A1(n13876), .A2(MEM_WB_OUT[145]), .B1(MEM_WB_OUT[113]), 
        .B2(n13875), .ZN(n5810) );
  OAI22_X2 U12721 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[155]), .B1(
        MEM_WB_OUT[123]), .B2(n13874), .ZN(n5809) );
  OAI22_X2 U12722 ( .A1(n13876), .A2(MEM_WB_OUT[161]), .B1(MEM_WB_OUT[129]), 
        .B2(n13874), .ZN(n5803) );
  OAI22_X2 U12723 ( .A1(n13876), .A2(MEM_WB_OUT[166]), .B1(MEM_WB_OUT[134]), 
        .B2(n13874), .ZN(n5797) );
  OAI22_X2 U12724 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[167]), .B1(
        MEM_WB_OUT[135]), .B2(n13874), .ZN(n5796) );
  OAI22_X2 U12725 ( .A1(n13876), .A2(MEM_WB_OUT[168]), .B1(MEM_WB_OUT[136]), 
        .B2(n13874), .ZN(n5795) );
  OAI22_X2 U12726 ( .A1(n13876), .A2(MEM_WB_OUT[169]), .B1(MEM_WB_OUT[137]), 
        .B2(n13874), .ZN(n5794) );
  OAI22_X2 U12727 ( .A1(n13876), .A2(MEM_WB_OUT[170]), .B1(MEM_WB_OUT[138]), 
        .B2(n13874), .ZN(n5793) );
  OAI22_X2 U12728 ( .A1(n13876), .A2(MEM_WB_OUT[171]), .B1(MEM_WB_OUT[139]), 
        .B2(n13874), .ZN(n5792) );
  OAI22_X2 U12729 ( .A1(n13876), .A2(MEM_WB_OUT[172]), .B1(MEM_WB_OUT[140]), 
        .B2(n13874), .ZN(n5791) );
  OAI22_X2 U12730 ( .A1(n13876), .A2(MEM_WB_OUT[173]), .B1(MEM_WB_OUT[141]), 
        .B2(n13874), .ZN(n5790) );
  OAI22_X2 U12731 ( .A1(n13876), .A2(MEM_WB_OUT[174]), .B1(MEM_WB_OUT[142]), 
        .B2(n13874), .ZN(n5789) );
  OAI22_X2 U12732 ( .A1(n13876), .A2(MEM_WB_OUT[147]), .B1(MEM_WB_OUT[115]), 
        .B2(n13875), .ZN(n5788) );
  OAI22_X2 U12733 ( .A1(n13876), .A2(MEM_WB_OUT[175]), .B1(MEM_WB_OUT[143]), 
        .B2(n13875), .ZN(n5787) );
  OAI22_X2 U12734 ( .A1(n13876), .A2(MEM_WB_OUT[176]), .B1(MEM_WB_OUT[144]), 
        .B2(n13875), .ZN(n5786) );
  OAI22_X2 U12735 ( .A1(n13876), .A2(MEM_WB_OUT[148]), .B1(MEM_WB_OUT[116]), 
        .B2(n13875), .ZN(n5785) );
  OAI22_X2 U12736 ( .A1(n13876), .A2(MEM_WB_OUT[149]), .B1(MEM_WB_OUT[117]), 
        .B2(n13875), .ZN(n5784) );
  OAI22_X2 U12737 ( .A1(n13876), .A2(MEM_WB_OUT[150]), .B1(MEM_WB_OUT[118]), 
        .B2(n13875), .ZN(n5783) );
  OAI22_X2 U12738 ( .A1(n13876), .A2(MEM_WB_OUT[151]), .B1(MEM_WB_OUT[119]), 
        .B2(n13875), .ZN(n5782) );
  OAI22_X2 U12739 ( .A1(n13876), .A2(MEM_WB_OUT[152]), .B1(MEM_WB_OUT[120]), 
        .B2(n13875), .ZN(n5781) );
  OAI22_X2 U12740 ( .A1(n13876), .A2(MEM_WB_OUT[153]), .B1(MEM_WB_OUT[121]), 
        .B2(n13875), .ZN(n5780) );
  OAI22_X2 U12741 ( .A1(n13876), .A2(MEM_WB_OUT[154]), .B1(MEM_WB_OUT[122]), 
        .B2(n13875), .ZN(n5779) );
  INV_X16 U12742 ( .A(n13428), .ZN(n13427) );
  INV_X2 U12743 ( .A(net231357), .ZN(net231353) );
  INV_X4 U12744 ( .A(net231331), .ZN(net231321) );
  INV_X4 U12745 ( .A(net231333), .ZN(net231313) );
  INV_X4 U12746 ( .A(n10235), .ZN(n13215) );
  INV_X4 U12747 ( .A(n17775), .ZN(n13381) );
  INV_X4 U12748 ( .A(n13381), .ZN(n13380) );
  AND2_X4 U12749 ( .A1(n14986), .A2(n2506), .ZN(n10349) );
  INV_X4 U12750 ( .A(n13547), .ZN(n13546) );
  INV_X4 U12751 ( .A(reset), .ZN(n13950) );
  AND2_X4 U12752 ( .A1(n15620), .A2(n10197), .ZN(n10350) );
  OAI21_X2 U12753 ( .B1(n5663), .B2(n5668), .A(n13934), .ZN(n5776) );
  OAI21_X2 U12754 ( .B1(n5662), .B2(n5764), .A(n13934), .ZN(n5767) );
  OAI21_X2 U12755 ( .B1(n5668), .B2(n5764), .A(n13934), .ZN(n5732) );
  OAI21_X2 U12756 ( .B1(n5662), .B2(n5718), .A(n13934), .ZN(n5721) );
  OAI21_X2 U12757 ( .B1(n5668), .B2(n5718), .A(n13934), .ZN(n5717) );
  OAI21_X2 U12758 ( .B1(n5668), .B2(n5676), .A(n13935), .ZN(n5675) );
  OAI21_X2 U12759 ( .B1(n5662), .B2(n5663), .A(n13935), .ZN(n5630) );
  AND2_X4 U12760 ( .A1(n19162), .A2(n10197), .ZN(n10352) );
  AND2_X4 U12761 ( .A1(n2511), .A2(n14999), .ZN(n10354) );
  INV_X4 U12762 ( .A(n11912), .ZN(n13305) );
  INV_X4 U12763 ( .A(n11912), .ZN(n13304) );
  AND2_X2 U12764 ( .A1(IF_ID_OUT[32]), .A2(net230387), .ZN(n10359) );
  AND2_X2 U12765 ( .A1(net230393), .A2(n10948), .ZN(n10361) );
  AND2_X4 U12766 ( .A1(n16061), .A2(n13386), .ZN(n10363) );
  INV_X4 U12767 ( .A(n14658), .ZN(n13506) );
  INV_X4 U12768 ( .A(n14658), .ZN(n13505) );
  INV_X4 U12769 ( .A(n11996), .ZN(n13419) );
  INV_X4 U12770 ( .A(n11996), .ZN(n13420) );
  INV_X4 U12771 ( .A(n11972), .ZN(n13826) );
  INV_X4 U12772 ( .A(n11972), .ZN(n13825) );
  INV_X4 U12773 ( .A(n11976), .ZN(n13830) );
  INV_X4 U12774 ( .A(n11976), .ZN(n13829) );
  AND2_X2 U12775 ( .A1(n15613), .A2(n15603), .ZN(n11989) );
  INV_X4 U12776 ( .A(n11989), .ZN(n13417) );
  INV_X4 U12777 ( .A(n11989), .ZN(n13418) );
  INV_X8 U12778 ( .A(n13191), .ZN(n13192) );
  INV_X4 U12779 ( .A(n18701), .ZN(n13191) );
  AND2_X4 U12782 ( .A1(n12274), .A2(n10837), .ZN(n10397) );
  AND3_X4 U12783 ( .A1(ID_EXEC_OUT[156]), .A2(ID_EXEC_OUT[157]), .A3(
        ID_EXEC_OUT[158]), .ZN(n10398) );
  INV_X4 U12784 ( .A(n14657), .ZN(n13507) );
  INV_X4 U12785 ( .A(n14657), .ZN(n13508) );
  AND2_X4 U12786 ( .A1(n15353), .A2(n10837), .ZN(n10531) );
  AND2_X4 U12787 ( .A1(n13936), .A2(n787), .ZN(n10532) );
  NAND2_X1 U12788 ( .A1(n10160), .A2(n15616), .ZN(n14646) );
  NAND2_X1 U12789 ( .A1(n10160), .A2(n10244), .ZN(n14648) );
  AND2_X4 U12790 ( .A1(n13936), .A2(n272), .ZN(n10541) );
  INV_X4 U12791 ( .A(n13463), .ZN(n13464) );
  AND2_X4 U12792 ( .A1(n13937), .A2(n27), .ZN(n10542) );
  INV_X4 U12793 ( .A(net230393), .ZN(net230373) );
  INV_X4 U12794 ( .A(net230387), .ZN(net230377) );
  INV_X4 U12795 ( .A(net230387), .ZN(net230379) );
  AND2_X4 U12796 ( .A1(n13935), .A2(n1135), .ZN(n10544) );
  AND2_X4 U12797 ( .A1(n13935), .A2(n1028), .ZN(n10545) );
  AND2_X4 U12798 ( .A1(n13936), .A2(n719), .ZN(n10546) );
  AND2_X4 U12799 ( .A1(n13936), .A2(n581), .ZN(n10547) );
  AND2_X4 U12800 ( .A1(n13936), .A2(n235), .ZN(n10548) );
  AND2_X4 U12801 ( .A1(n13935), .A2(n959), .ZN(n10549) );
  AND2_X4 U12802 ( .A1(n13936), .A2(n651), .ZN(n10550) );
  AND2_X4 U12803 ( .A1(n13936), .A2(n376), .ZN(n10551) );
  AND2_X4 U12804 ( .A1(n13936), .A2(n342), .ZN(n10552) );
  AND2_X4 U12805 ( .A1(n13936), .A2(n685), .ZN(n10553) );
  AND2_X4 U12806 ( .A1(n13937), .A2(n201), .ZN(n10554) );
  AND2_X4 U12807 ( .A1(n13937), .A2(n95), .ZN(n10555) );
  AND2_X4 U12808 ( .A1(n13935), .A2(n924), .ZN(n10556) );
  AND2_X4 U12809 ( .A1(n13936), .A2(n616), .ZN(n10557) );
  OR2_X4 U12810 ( .A1(n15507), .A2(n15505), .ZN(n10558) );
  AND2_X4 U12811 ( .A1(n19124), .A2(n18651), .ZN(n10559) );
  OAI22_X2 U12812 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[164]), .B1(
        MEM_WB_OUT[132]), .B2(n12978), .ZN(n5800) );
  OAI22_X2 U12813 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[165]), .B1(
        MEM_WB_OUT[133]), .B2(n13874), .ZN(n5798) );
  INV_X4 U12814 ( .A(n16207), .ZN(n13394) );
  AND4_X4 U12815 ( .A1(n17968), .A2(n17967), .A3(n17966), .A4(n17965), .ZN(
        n10773) );
  AND4_X4 U12816 ( .A1(n18058), .A2(n18057), .A3(n18056), .A4(n18055), .ZN(
        n10774) );
  AND4_X4 U12817 ( .A1(n18101), .A2(n18100), .A3(n18099), .A4(n18098), .ZN(
        n10775) );
  AND4_X4 U12818 ( .A1(n18146), .A2(n18145), .A3(n18144), .A4(n18143), .ZN(
        n10776) );
  AND4_X4 U12819 ( .A1(n18232), .A2(n18231), .A3(n18230), .A4(n18229), .ZN(
        n10777) );
  AND4_X4 U12820 ( .A1(n18440), .A2(n18439), .A3(n18438), .A4(n18437), .ZN(
        n10778) );
  AND4_X4 U12821 ( .A1(n18521), .A2(n18520), .A3(n18519), .A4(n18518), .ZN(
        n10779) );
  AND4_X4 U12822 ( .A1(n18187), .A2(n18186), .A3(n18185), .A4(n18184), .ZN(
        n10780) );
  AND2_X4 U12823 ( .A1(n2508), .A2(n14999), .ZN(n10782) );
  INV_X4 U12824 ( .A(n10198), .ZN(n13550) );
  AND2_X4 U12825 ( .A1(n14995), .A2(n2506), .ZN(n10801) );
  INV_X2 U12826 ( .A(n10235), .ZN(n13214) );
  INV_X1 U12827 ( .A(net231357), .ZN(net231349) );
  INV_X4 U12828 ( .A(net231349), .ZN(net231345) );
  INV_X4 U12829 ( .A(net231321), .ZN(net231339) );
  INV_X4 U12830 ( .A(n12714), .ZN(n13430) );
  INV_X4 U12831 ( .A(n13430), .ZN(n13433) );
  INV_X4 U12832 ( .A(reset), .ZN(n13948) );
  INV_X4 U12833 ( .A(n13950), .ZN(n13910) );
  INV_X4 U12834 ( .A(n13950), .ZN(n13909) );
  INV_X4 U12835 ( .A(n13950), .ZN(n13908) );
  AND2_X4 U12836 ( .A1(n15608), .A2(n15620), .ZN(n10803) );
  AND2_X4 U12837 ( .A1(n10244), .A2(n15620), .ZN(n10804) );
  AND2_X4 U12838 ( .A1(n10241), .A2(n15617), .ZN(n10805) );
  INV_X4 U12839 ( .A(n18637), .ZN(n16300) );
  AND2_X4 U12840 ( .A1(n2527), .A2(net231359), .ZN(n10808) );
  AND2_X4 U12841 ( .A1(n14644), .A2(n10824), .ZN(n10809) );
  INV_X4 U12842 ( .A(n14283), .ZN(n13238) );
  INV_X4 U12843 ( .A(n14283), .ZN(n13239) );
  NAND2_X1 U12844 ( .A1(n10808), .A2(n14998), .ZN(n14282) );
  INV_X4 U12845 ( .A(n14282), .ZN(n13236) );
  INV_X4 U12846 ( .A(n14282), .ZN(n13237) );
  INV_X1 U12847 ( .A(n16295), .ZN(n16279) );
  INV_X16 U12848 ( .A(n13187), .ZN(n13188) );
  AND2_X4 U12849 ( .A1(n15613), .A2(n10197), .ZN(n10827) );
  AND2_X4 U12850 ( .A1(n12540), .A2(n10398), .ZN(n10829) );
  AND2_X2 U12852 ( .A1(n2511), .A2(n14991), .ZN(n10831) );
  AND2_X2 U12853 ( .A1(n2506), .A2(n14990), .ZN(n10832) );
  AND2_X4 U12854 ( .A1(n10244), .A2(n15617), .ZN(n10833) );
  AND2_X4 U12855 ( .A1(n15621), .A2(n15620), .ZN(n10834) );
  AND2_X2 U12856 ( .A1(n19162), .A2(n15603), .ZN(n10835) );
  AND2_X4 U12857 ( .A1(n10809), .A2(n10197), .ZN(n10836) );
  INV_X4 U12858 ( .A(n11929), .ZN(n13753) );
  INV_X4 U12859 ( .A(n11929), .ZN(n13752) );
  INV_X4 U12860 ( .A(n11970), .ZN(n13779) );
  INV_X4 U12861 ( .A(n11970), .ZN(n13778) );
  INV_X4 U12862 ( .A(n11971), .ZN(n13818) );
  INV_X4 U12863 ( .A(n11971), .ZN(n13817) );
  INV_X4 U12864 ( .A(n11973), .ZN(n13775) );
  INV_X4 U12865 ( .A(n11973), .ZN(n13774) );
  INV_X4 U12866 ( .A(n11975), .ZN(n13814) );
  INV_X4 U12867 ( .A(n11975), .ZN(n13813) );
  AND2_X2 U12868 ( .A1(RegWrite_wb_out), .A2(n19315), .ZN(n10837) );
  INV_X4 U12869 ( .A(n12015), .ZN(n13822) );
  INV_X4 U12870 ( .A(n12015), .ZN(n13821) );
  INV_X4 U12871 ( .A(n12011), .ZN(n13770) );
  INV_X4 U12872 ( .A(n12011), .ZN(n13771) );
  INV_X4 U12873 ( .A(n12012), .ZN(n13840) );
  INV_X4 U12874 ( .A(n12012), .ZN(n13839) );
  INV_X4 U12875 ( .A(n12013), .ZN(n13634) );
  INV_X4 U12876 ( .A(n12013), .ZN(n13635) );
  INV_X4 U12877 ( .A(n12014), .ZN(n13658) );
  INV_X4 U12878 ( .A(n12014), .ZN(n13659) );
  INV_X4 U12879 ( .A(n11998), .ZN(n13678) );
  INV_X4 U12880 ( .A(n11998), .ZN(n13679) );
  INV_X1 U12881 ( .A(n17774), .ZN(n13376) );
  AND2_X2 U12882 ( .A1(n16872), .A2(n13938), .ZN(n10839) );
  INV_X4 U12883 ( .A(n18727), .ZN(n13200) );
  INV_X8 U12884 ( .A(n13194), .ZN(n13195) );
  INV_X4 U12885 ( .A(n18712), .ZN(n13194) );
  INV_X4 U12886 ( .A(n18726), .ZN(n13198) );
  INV_X8 U12887 ( .A(n13203), .ZN(n13204) );
  INV_X4 U12888 ( .A(n18730), .ZN(n13203) );
  INV_X8 U12889 ( .A(n13189), .ZN(n13190) );
  INV_X4 U12890 ( .A(n18700), .ZN(n13189) );
  AND2_X2 U12891 ( .A1(n15617), .A2(n15603), .ZN(n10841) );
  AND2_X2 U12892 ( .A1(n2508), .A2(n14997), .ZN(n10842) );
  AND2_X4 U12893 ( .A1(n18309), .A2(n18641), .ZN(n10843) );
  AND2_X2 U12894 ( .A1(n16918), .A2(n13938), .ZN(n10907) );
  AND2_X2 U12895 ( .A1(n17242), .A2(n13938), .ZN(n10908) );
  AND2_X2 U12896 ( .A1(n17045), .A2(n13938), .ZN(n10909) );
  AND2_X2 U12897 ( .A1(n15718), .A2(n13938), .ZN(n10934) );
  OR4_X4 U12898 ( .A1(n15508), .A2(net230373), .A3(n19318), .A4(n15507), .ZN(
        n10943) );
  AND2_X2 U12899 ( .A1(n15610), .A2(n15603), .ZN(n10944) );
  AND2_X4 U12900 ( .A1(n5811), .A2(n19306), .ZN(n10950) );
  AND2_X4 U12901 ( .A1(n5811), .A2(n19308), .ZN(n10951) );
  AND2_X4 U12902 ( .A1(n5811), .A2(n19302), .ZN(n10952) );
  AND2_X4 U12903 ( .A1(n5811), .A2(n19303), .ZN(n10953) );
  AND2_X4 U12904 ( .A1(n5811), .A2(n19304), .ZN(n10954) );
  AND2_X4 U12905 ( .A1(n5811), .A2(n19305), .ZN(n10955) );
  AND2_X4 U12906 ( .A1(n5811), .A2(n19309), .ZN(n10956) );
  AND2_X4 U12907 ( .A1(n5811), .A2(n19307), .ZN(n10957) );
  AND2_X4 U12908 ( .A1(n5815), .A2(n19307), .ZN(n10960) );
  AND2_X4 U12909 ( .A1(n5815), .A2(n19308), .ZN(n10961) );
  AND2_X4 U12910 ( .A1(n5815), .A2(n19302), .ZN(n10962) );
  AND2_X4 U12911 ( .A1(n5815), .A2(n19303), .ZN(n10963) );
  AND2_X4 U12912 ( .A1(n5815), .A2(n19304), .ZN(n10964) );
  AND2_X4 U12913 ( .A1(n5815), .A2(n19306), .ZN(n10965) );
  AND2_X4 U12914 ( .A1(n5815), .A2(n19305), .ZN(n10966) );
  AND2_X4 U12915 ( .A1(n5815), .A2(n19309), .ZN(n10967) );
  AND2_X4 U12916 ( .A1(net225077), .A2(n10357), .ZN(n11016) );
  AND2_X4 U12917 ( .A1(n5670), .A2(n19307), .ZN(n11037) );
  AND2_X4 U12918 ( .A1(n5670), .A2(n19309), .ZN(n11038) );
  AND2_X4 U12919 ( .A1(n10160), .A2(n15608), .ZN(n11039) );
  AND2_X4 U12920 ( .A1(n10160), .A2(n10241), .ZN(n11040) );
  AND2_X2 U12921 ( .A1(n2503), .A2(n14991), .ZN(n11042) );
  AND2_X4 U12922 ( .A1(n15608), .A2(n19162), .ZN(n11043) );
  AND2_X4 U12923 ( .A1(n15608), .A2(n10809), .ZN(n11044) );
  AND2_X4 U12924 ( .A1(n15616), .A2(n19162), .ZN(n11046) );
  AND2_X4 U12925 ( .A1(n15616), .A2(n10809), .ZN(n11047) );
  AND2_X2 U12926 ( .A1(n14293), .A2(n14998), .ZN(n11048) );
  AND2_X4 U12927 ( .A1(n15609), .A2(n10161), .ZN(n11049) );
  AND2_X4 U12928 ( .A1(n15609), .A2(n19162), .ZN(n11050) );
  AND2_X4 U12929 ( .A1(n19162), .A2(n10241), .ZN(n11051) );
  AND2_X4 U12930 ( .A1(n14999), .A2(n10808), .ZN(n11052) );
  AND2_X4 U12931 ( .A1(n14986), .A2(n10808), .ZN(n11053) );
  AND2_X4 U12932 ( .A1(n10244), .A2(n10809), .ZN(n11054) );
  AND2_X4 U12933 ( .A1(n10244), .A2(n19162), .ZN(n11055) );
  AND2_X4 U12934 ( .A1(n10197), .A2(n10160), .ZN(n11056) );
  AND2_X4 U12935 ( .A1(n10808), .A2(n14997), .ZN(n11057) );
  AND2_X4 U12936 ( .A1(n10808), .A2(n14982), .ZN(n11058) );
  AND2_X4 U12937 ( .A1(n10161), .A2(n15608), .ZN(n11059) );
  AND2_X4 U12938 ( .A1(n10161), .A2(n10241), .ZN(n11060) );
  AND2_X2 U12939 ( .A1(n10809), .A2(n15603), .ZN(n11061) );
  AND2_X4 U12940 ( .A1(n10809), .A2(n10241), .ZN(n11062) );
  AND2_X4 U12941 ( .A1(n14991), .A2(n10808), .ZN(n11063) );
  AND2_X4 U12942 ( .A1(n19308), .A2(n5670), .ZN(n11064) );
  AND2_X4 U12943 ( .A1(n19303), .A2(n5670), .ZN(n11065) );
  AND2_X4 U12944 ( .A1(n19304), .A2(n5670), .ZN(n11066) );
  AND2_X4 U12945 ( .A1(n19305), .A2(n5670), .ZN(n11067) );
  AND2_X4 U12946 ( .A1(n19306), .A2(n5670), .ZN(n11068) );
  AND2_X4 U12947 ( .A1(n19308), .A2(n5664), .ZN(n11069) );
  AND2_X4 U12948 ( .A1(n19302), .A2(n5664), .ZN(n11070) );
  AND2_X4 U12949 ( .A1(n19306), .A2(n5664), .ZN(n11071) );
  AND2_X4 U12950 ( .A1(n19303), .A2(n5664), .ZN(n11072) );
  AND2_X4 U12951 ( .A1(n19304), .A2(n5664), .ZN(n11073) );
  AND2_X4 U12952 ( .A1(n19309), .A2(n5664), .ZN(n11074) );
  INV_X4 U12953 ( .A(n13168), .ZN(n13169) );
  INV_X4 U12954 ( .A(n14632), .ZN(n13168) );
  NOR2_X2 U12955 ( .A1(n14281), .A2(n14277), .ZN(n11075) );
  NOR2_X2 U12956 ( .A1(n14281), .A2(n14271), .ZN(n11076) );
  NOR2_X2 U12957 ( .A1(n14281), .A2(n14274), .ZN(n11077) );
  NOR2_X2 U12958 ( .A1(n14281), .A2(n14276), .ZN(n11078) );
  NOR2_X2 U12959 ( .A1(n14281), .A2(n14280), .ZN(n11079) );
  NOR2_X2 U12960 ( .A1(n14279), .A2(n14275), .ZN(n11080) );
  NOR2_X2 U12961 ( .A1(n14279), .A2(n14278), .ZN(n11081) );
  AND2_X2 U12962 ( .A1(n13167), .A2(net230387), .ZN(n11083) );
  AND2_X4 U12963 ( .A1(n13936), .A2(n13787), .ZN(n11084) );
  AND2_X4 U12964 ( .A1(n13936), .A2(n13814), .ZN(n11085) );
  AND2_X4 U12965 ( .A1(n13936), .A2(n13818), .ZN(n11086) );
  AND2_X4 U12966 ( .A1(n13936), .A2(n13822), .ZN(n11087) );
  AND2_X4 U12967 ( .A1(n13936), .A2(n13826), .ZN(n11088) );
  AND2_X4 U12968 ( .A1(n13936), .A2(n13830), .ZN(n11089) );
  AND2_X4 U12969 ( .A1(n13935), .A2(n13753), .ZN(n11090) );
  AND2_X4 U12970 ( .A1(n13935), .A2(n10162), .ZN(n11091) );
  AND2_X4 U12971 ( .A1(n13935), .A2(n10163), .ZN(n11092) );
  AND2_X4 U12972 ( .A1(n13935), .A2(n13775), .ZN(n11093) );
  AND2_X4 U12973 ( .A1(n13935), .A2(n13779), .ZN(n11094) );
  AND2_X4 U12974 ( .A1(n13937), .A2(n10166), .ZN(n11095) );
  AND2_X4 U12975 ( .A1(n13937), .A2(n10167), .ZN(n11096) );
  INV_X4 U12976 ( .A(n12978), .ZN(n13876) );
  INV_X4 U12977 ( .A(MEM_WB_OUT[178]), .ZN(n13875) );
  INV_X4 U12978 ( .A(MEM_WB_OUT[178]), .ZN(n13874) );
  NAND2_X1 U12979 ( .A1(ID_EXEC_OUT[276]), .A2(net230387), .ZN(n18586) );
  OR2_X4 U12980 ( .A1(n13365), .A2(n12836), .ZN(n11461) );
  OR2_X4 U12981 ( .A1(n13365), .A2(n12844), .ZN(n11462) );
  OR2_X4 U12982 ( .A1(n13365), .A2(n12848), .ZN(n11463) );
  OR2_X4 U12983 ( .A1(n13365), .A2(n12860), .ZN(n11464) );
  OR2_X4 U12984 ( .A1(n13365), .A2(n12868), .ZN(n11465) );
  OR2_X4 U12985 ( .A1(n13365), .A2(n12878), .ZN(n11466) );
  OR2_X4 U12986 ( .A1(n13365), .A2(n12882), .ZN(n11467) );
  OR2_X4 U12987 ( .A1(n13365), .A2(n12892), .ZN(n11468) );
  INV_X4 U12988 ( .A(n1746), .ZN(net230403) );
  AND2_X4 U12989 ( .A1(n15608), .A2(n15610), .ZN(n11572) );
  INV_X4 U12990 ( .A(n17771), .ZN(n13369) );
  INV_X4 U12991 ( .A(n719), .ZN(n13791) );
  INV_X4 U12992 ( .A(n13791), .ZN(n13790) );
  INV_X4 U12993 ( .A(n651), .ZN(n13801) );
  INV_X4 U12994 ( .A(n13801), .ZN(n13800) );
  INV_X4 U12995 ( .A(n13801), .ZN(n13799) );
  INV_X4 U12996 ( .A(n685), .ZN(n13796) );
  INV_X4 U12997 ( .A(n13796), .ZN(n13795) );
  INV_X4 U12998 ( .A(n13796), .ZN(n13794) );
  INV_X4 U12999 ( .A(n616), .ZN(n13806) );
  INV_X4 U13000 ( .A(n13806), .ZN(n13805) );
  INV_X4 U13001 ( .A(n13806), .ZN(n13804) );
  XNOR2_X2 U13002 ( .A(n19313), .B(offset_26_id[6]), .ZN(n11583) );
  NAND2_X1 U13003 ( .A1(net230393), .A2(EXEC_MEM_IN[102]), .ZN(net223104) );
  NAND2_X2 U13004 ( .A1(n5774), .A2(n10817), .ZN(n5662) );
  NAND2_X2 U13005 ( .A1(MEM_WB_OUT[111]), .A2(n5774), .ZN(n5668) );
  NAND2_X2 U13006 ( .A1(MEM_WB_OUT[111]), .A2(n5909), .ZN(n5816) );
  NAND2_X2 U13007 ( .A1(n10160), .A2(n15609), .ZN(n11832) );
  INV_X4 U13008 ( .A(n12061), .ZN(n13457) );
  INV_X4 U13009 ( .A(n13457), .ZN(n13456) );
  NAND2_X2 U13010 ( .A1(n14288), .A2(n14997), .ZN(n11833) );
  NAND2_X2 U13011 ( .A1(n14288), .A2(n14995), .ZN(n11834) );
  NAND2_X2 U13012 ( .A1(n14288), .A2(n14986), .ZN(n11835) );
  NAND2_X2 U13013 ( .A1(n14288), .A2(n14982), .ZN(n11836) );
  NAND2_X2 U13014 ( .A1(n14288), .A2(n14990), .ZN(n11837) );
  NAND2_X2 U13015 ( .A1(n14293), .A2(n14991), .ZN(n11896) );
  NAND2_X2 U13016 ( .A1(n14293), .A2(n14999), .ZN(n11897) );
  NAND2_X2 U13017 ( .A1(n14293), .A2(n14990), .ZN(n11898) );
  NAND2_X2 U13018 ( .A1(n14293), .A2(n14995), .ZN(n11899) );
  NAND2_X2 U13019 ( .A1(n14293), .A2(n14997), .ZN(n11900) );
  NAND2_X2 U13020 ( .A1(n10808), .A2(n14995), .ZN(n11901) );
  NAND2_X2 U13021 ( .A1(n10808), .A2(n14990), .ZN(n11902) );
  NAND2_X2 U13022 ( .A1(n10161), .A2(n15616), .ZN(n11903) );
  NAND2_X2 U13023 ( .A1(n10161), .A2(n10244), .ZN(n11904) );
  NAND2_X2 U13024 ( .A1(n10161), .A2(n10197), .ZN(n11905) );
  NAND2_X2 U13025 ( .A1(n10809), .A2(n15621), .ZN(n11906) );
  NAND2_X2 U13026 ( .A1(n10809), .A2(n15609), .ZN(n11907) );
  INV_X4 U13027 ( .A(n10558), .ZN(n13411) );
  INV_X4 U13028 ( .A(n10558), .ZN(n13412) );
  NAND2_X2 U13029 ( .A1(n14273), .A2(n14999), .ZN(n11908) );
  INV_X4 U13030 ( .A(n2182), .ZN(n13731) );
  NAND2_X2 U13031 ( .A1(n14273), .A2(n14991), .ZN(n11909) );
  NAND2_X1 U13032 ( .A1(n14273), .A2(n14998), .ZN(n11910) );
  NAND2_X1 U13033 ( .A1(n15507), .A2(net230387), .ZN(n11911) );
  INV_X4 U13034 ( .A(n18705), .ZN(n13449) );
  INV_X2 U13035 ( .A(n18532), .ZN(n16059) );
  INV_X4 U13036 ( .A(net231355), .ZN(net231329) );
  INV_X2 U13037 ( .A(net231345), .ZN(net231271) );
  INV_X4 U13038 ( .A(net231331), .ZN(net231317) );
  INV_X4 U13039 ( .A(net231345), .ZN(net231277) );
  NAND3_X2 U13040 ( .A1(EXEC_STAGE_mul_ex_CurrentState_1_), .A2(n10159), .A3(
        EXEC_STAGE_mul_ex_CurrentState_2_), .ZN(n7286) );
  NAND3_X2 U13041 ( .A1(n10159), .A2(n10543), .A3(
        EXEC_STAGE_mul_ex_CurrentState_2_), .ZN(n7288) );
  INV_X4 U13042 ( .A(reset), .ZN(n13952) );
  AND2_X2 U13043 ( .A1(n17868), .A2(n13938), .ZN(n11912) );
  AND2_X4 U13044 ( .A1(n13125), .A2(n13938), .ZN(n11923) );
  AND2_X2 U13045 ( .A1(n17981), .A2(n13937), .ZN(n11924) );
  AND2_X2 U13046 ( .A1(n13101), .A2(n13937), .ZN(n11925) );
  AND2_X2 U13047 ( .A1(n15686), .A2(n13937), .ZN(n11926) );
  INV_X1 U13048 ( .A(n17045), .ZN(n17020) );
  AND2_X4 U13049 ( .A1(n200), .A2(n10262), .ZN(n11929) );
  AND2_X2 U13050 ( .A1(n16147), .A2(n13939), .ZN(n11946) );
  AND2_X2 U13051 ( .A1(n16295), .A2(n13938), .ZN(n11948) );
  AND2_X2 U13052 ( .A1(n16222), .A2(n13938), .ZN(n11951) );
  AND2_X2 U13053 ( .A1(n16031), .A2(n13939), .ZN(n11952) );
  AND2_X2 U13054 ( .A1(n16070), .A2(n13938), .ZN(n11953) );
  AND2_X2 U13055 ( .A1(n16539), .A2(n13938), .ZN(n11954) );
  AND2_X4 U13056 ( .A1(n10322), .A2(n200), .ZN(n11970) );
  AND2_X4 U13057 ( .A1(n10531), .A2(n200), .ZN(n11971) );
  AND2_X4 U13058 ( .A1(n10323), .A2(n129), .ZN(n11972) );
  AND2_X4 U13059 ( .A1(n10322), .A2(n94), .ZN(n11973) );
  AND2_X4 U13060 ( .A1(n10397), .A2(n94), .ZN(n11974) );
  AND2_X4 U13061 ( .A1(n10531), .A2(n94), .ZN(n11975) );
  AND2_X4 U13062 ( .A1(n10323), .A2(n94), .ZN(n11976) );
  AND2_X2 U13063 ( .A1(n16350), .A2(n13938), .ZN(n11978) );
  AND2_X2 U13064 ( .A1(n16578), .A2(n13938), .ZN(n11979) );
  NAND2_X2 U13065 ( .A1(IMEM_BUS_OUT[5]), .A2(n15402), .ZN(n15451) );
  AND2_X4 U13066 ( .A1(n15610), .A2(n10197), .ZN(n11984) );
  AND2_X2 U13067 ( .A1(n17737), .A2(n13938), .ZN(n11988) );
  AND4_X1 U13068 ( .A1(ID_STAGE_imm16_aluA[26]), .A2(ID_STAGE_imm16_aluA[27]), 
        .A3(ID_STAGE_imm16_aluA[29]), .A4(n10840), .ZN(n11991) );
  AND2_X2 U13069 ( .A1(n15621), .A2(n15613), .ZN(n11992) );
  AND2_X4 U13070 ( .A1(net225187), .A2(nextPC_ex_out[8]), .ZN(n11994) );
  AND2_X4 U13071 ( .A1(n15609), .A2(n15613), .ZN(n11996) );
  AND2_X2 U13072 ( .A1(n18623), .A2(n13939), .ZN(n11997) );
  AND2_X4 U13073 ( .A1(n5664), .A2(n19307), .ZN(n11998) );
  AND2_X2 U13074 ( .A1(n17094), .A2(n13938), .ZN(n11999) );
  AND2_X2 U13075 ( .A1(n17331), .A2(n13938), .ZN(n12000) );
  AND2_X2 U13076 ( .A1(n17382), .A2(n13938), .ZN(n12001) );
  AND2_X2 U13077 ( .A1(n17546), .A2(n13937), .ZN(n12002) );
  AND2_X2 U13078 ( .A1(n17622), .A2(n13937), .ZN(n12003) );
  AND2_X2 U13079 ( .A1(n17840), .A2(n13937), .ZN(n12004) );
  AND2_X2 U13080 ( .A1(n15770), .A2(n13937), .ZN(n12005) );
  AND2_X2 U13081 ( .A1(n15837), .A2(n13937), .ZN(n12006) );
  AND2_X2 U13082 ( .A1(n15682), .A2(n13937), .ZN(n12007) );
  AND2_X2 U13083 ( .A1(n15678), .A2(n13937), .ZN(n12008) );
  AND2_X2 U13084 ( .A1(n15700), .A2(n13937), .ZN(n12009) );
  AND2_X2 U13085 ( .A1(n10118), .A2(n13937), .ZN(n12010) );
  AND2_X4 U13086 ( .A1(n13935), .A2(n10164), .ZN(n12011) );
  AND2_X4 U13087 ( .A1(n13936), .A2(n10165), .ZN(n12012) );
  AND2_X4 U13088 ( .A1(n19302), .A2(n5670), .ZN(n12013) );
  AND2_X4 U13089 ( .A1(n19305), .A2(n5664), .ZN(n12014) );
  AND2_X4 U13090 ( .A1(n10531), .A2(n164), .ZN(n12015) );
  AND2_X4 U13091 ( .A1(nextPC_ex_out[10]), .A2(nextPC_ex_out[9]), .ZN(n12019)
         );
  AND2_X4 U13092 ( .A1(n15351), .A2(n15354), .ZN(n12022) );
  AND2_X2 U13093 ( .A1(ID_EXEC_OUT[156]), .A2(n11913), .ZN(n12030) );
  OR2_X1 U13094 ( .A1(ID_EXEC_OUT[275]), .A2(EXEC_MEM_OUT_141), .ZN(n12035) );
  XNOR2_X1 U13095 ( .A(n10828), .B(n10351), .ZN(n12053) );
  INV_X2 U13097 ( .A(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[20]), .ZN(n19296)
         );
  AND2_X2 U13098 ( .A1(n10244), .A2(n15613), .ZN(n12061) );
  INV_X4 U13099 ( .A(n17768), .ZN(n13363) );
  INV_X4 U13100 ( .A(n13363), .ZN(n13362) );
  INV_X4 U13101 ( .A(n18733), .ZN(n13469) );
  INV_X8 U13102 ( .A(n10804), .ZN(n13473) );
  INV_X4 U13103 ( .A(n15334), .ZN(n13277) );
  INV_X8 U13104 ( .A(n13277), .ZN(n13276) );
  INV_X8 U13105 ( .A(n13277), .ZN(n13275) );
  INV_X4 U13106 ( .A(n15335), .ZN(n13280) );
  INV_X8 U13107 ( .A(n13280), .ZN(n13279) );
  INV_X8 U13108 ( .A(n13280), .ZN(n13278) );
  AND2_X4 U13109 ( .A1(nextPC_ex_out[14]), .A2(nextPC_ex_out[15]), .ZN(n12127)
         );
  NAND2_X2 U13110 ( .A1(net223742), .A2(n11950), .ZN(net227186) );
  INV_X4 U13111 ( .A(net227186), .ZN(net227216) );
  OR2_X2 U13112 ( .A1(ID_STAGE_imm16_aluA[22]), .A2(ID_STAGE_imm16_aluA[23]), 
        .ZN(n12128) );
  INV_X4 U13113 ( .A(n18718), .ZN(n13462) );
  INV_X4 U13114 ( .A(n13462), .ZN(n13461) );
  INV_X4 U13115 ( .A(n13462), .ZN(n13460) );
  INV_X4 U13116 ( .A(n10841), .ZN(n13424) );
  INV_X8 U13117 ( .A(n10841), .ZN(n13423) );
  INV_X4 U13118 ( .A(n19097), .ZN(n13489) );
  INV_X4 U13119 ( .A(n13489), .ZN(n13488) );
  AND2_X4 U13120 ( .A1(n19076), .A2(n19075), .ZN(n12132) );
  AND2_X2 U13121 ( .A1(n5506), .A2(n12555), .ZN(n12133) );
  OR2_X4 U13122 ( .A1(net227048), .A2(net227012), .ZN(n12205) );
  OR2_X4 U13123 ( .A1(net230377), .A2(n18769), .ZN(n12219) );
  NAND2_X2 U13124 ( .A1(n19300), .A2(n10157), .ZN(n1866) );
  AND2_X4 U13125 ( .A1(n19025), .A2(n19026), .ZN(n12253) );
  AND2_X2 U13126 ( .A1(n19313), .A2(n19311), .ZN(n12274) );
  INV_X4 U13127 ( .A(n10943), .ZN(n13415) );
  INV_X4 U13128 ( .A(n10943), .ZN(n13416) );
  AND2_X2 U13129 ( .A1(net225529), .A2(nextPC_ex_out[14]), .ZN(n12309) );
  NAND2_X1 U13130 ( .A1(n15498), .A2(n19359), .ZN(n15506) );
  INV_X4 U13131 ( .A(n15330), .ZN(n13274) );
  AND2_X2 U13132 ( .A1(MEM_WB_OUT[31]), .A2(n13878), .ZN(n12501) );
  OR2_X4 U13133 ( .A1(n13184), .A2(n12418), .ZN(n12526) );
  OR2_X4 U13134 ( .A1(n13184), .A2(n12423), .ZN(n12527) );
  OR2_X4 U13135 ( .A1(n13184), .A2(n12427), .ZN(n12528) );
  OR2_X4 U13136 ( .A1(n13184), .A2(n12433), .ZN(n12529) );
  OR2_X4 U13137 ( .A1(n13184), .A2(n12438), .ZN(n12530) );
  OR2_X4 U13138 ( .A1(n13184), .A2(n12446), .ZN(n12531) );
  OR2_X4 U13139 ( .A1(n13184), .A2(n12450), .ZN(n12532) );
  OR2_X4 U13140 ( .A1(n13184), .A2(n12458), .ZN(n12533) );
  XNOR2_X1 U13141 ( .A(n19317), .B(offset_26_id[3]), .ZN(n12539) );
  AND3_X4 U13142 ( .A1(n18654), .A2(n10157), .A3(n12017), .ZN(n12540) );
  INV_X4 U13143 ( .A(n10842), .ZN(n13743) );
  INV_X4 U13144 ( .A(n11048), .ZN(n13244) );
  INV_X4 U13145 ( .A(n11048), .ZN(n13245) );
  INV_X4 U13146 ( .A(n14968), .ZN(n13257) );
  INV_X4 U13147 ( .A(n11059), .ZN(n13251) );
  INV_X4 U13148 ( .A(n11059), .ZN(n13250) );
  INV_X4 U13149 ( .A(n11039), .ZN(n13253) );
  INV_X4 U13150 ( .A(n11039), .ZN(n13252) );
  INV_X16 U13151 ( .A(n13357), .ZN(n13356) );
  INV_X4 U13152 ( .A(n11051), .ZN(n13709) );
  INV_X4 U13153 ( .A(n11051), .ZN(n13708) );
  INV_X4 U13154 ( .A(n11053), .ZN(n13689) );
  INV_X4 U13155 ( .A(n11053), .ZN(n13688) );
  INV_X4 U13156 ( .A(n1871), .ZN(n13737) );
  INV_X4 U13157 ( .A(n11042), .ZN(n13745) );
  INV_X4 U13158 ( .A(n11042), .ZN(n13744) );
  INV_X4 U13159 ( .A(n11040), .ZN(n13713) );
  INV_X4 U13160 ( .A(n11040), .ZN(n13712) );
  INV_X4 U13161 ( .A(n11050), .ZN(n13717) );
  INV_X4 U13162 ( .A(n11050), .ZN(n13716) );
  INV_X4 U13163 ( .A(n11056), .ZN(n13721) );
  INV_X4 U13164 ( .A(n11056), .ZN(n13720) );
  INV_X4 U13165 ( .A(n11047), .ZN(n13725) );
  INV_X4 U13166 ( .A(n11047), .ZN(n13724) );
  INV_X4 U13167 ( .A(n18713), .ZN(n13454) );
  INV_X4 U13168 ( .A(n13454), .ZN(n13453) );
  INV_X4 U13169 ( .A(n11075), .ZN(n13685) );
  INV_X4 U13170 ( .A(n11075), .ZN(n13684) );
  INV_X4 U13171 ( .A(n11078), .ZN(n13693) );
  INV_X4 U13172 ( .A(n11078), .ZN(n13692) );
  INV_X4 U13173 ( .A(n11079), .ZN(n13697) );
  INV_X4 U13174 ( .A(n11079), .ZN(n13696) );
  INV_X4 U13175 ( .A(n10361), .ZN(net231915) );
  INV_X4 U13176 ( .A(n959), .ZN(n13765) );
  INV_X4 U13177 ( .A(n13765), .ZN(n13764) );
  INV_X4 U13178 ( .A(n376), .ZN(n13834) );
  INV_X4 U13179 ( .A(n13834), .ZN(n13833) );
  INV_X4 U13180 ( .A(n342), .ZN(n13838) );
  INV_X4 U13181 ( .A(n13838), .ZN(n13837) );
  INV_X4 U13182 ( .A(n1028), .ZN(n13759) );
  INV_X4 U13183 ( .A(n13759), .ZN(n13758) );
  INV_X4 U13184 ( .A(n581), .ZN(n13810) );
  INV_X4 U13185 ( .A(n13810), .ZN(n13809) );
  INV_X4 U13186 ( .A(n1135), .ZN(n13747) );
  INV_X4 U13187 ( .A(n13747), .ZN(n13746) );
  INV_X4 U13188 ( .A(n235), .ZN(n13848) );
  INV_X4 U13189 ( .A(n13848), .ZN(n13847) );
  INV_X4 U13190 ( .A(n201), .ZN(n13852) );
  INV_X4 U13191 ( .A(n13852), .ZN(n13851) );
  OR2_X4 U13192 ( .A1(net227186), .A2(net227187), .ZN(n12558) );
  INV_X4 U13193 ( .A(n95), .ZN(n13860) );
  INV_X4 U13194 ( .A(n13860), .ZN(n13859) );
  INV_X4 U13195 ( .A(n27), .ZN(n13864) );
  INV_X4 U13196 ( .A(n13864), .ZN(n13863) );
  INV_X4 U13197 ( .A(n787), .ZN(n13783) );
  INV_X4 U13198 ( .A(n13783), .ZN(n13782) );
  INV_X4 U13199 ( .A(n924), .ZN(n13769) );
  INV_X4 U13200 ( .A(n13769), .ZN(n13768) );
  INV_X4 U13201 ( .A(n272), .ZN(n13844) );
  INV_X4 U13202 ( .A(n13844), .ZN(n13843) );
  INV_X4 U13203 ( .A(n11043), .ZN(n13703) );
  INV_X4 U13204 ( .A(n11043), .ZN(n13702) );
  INV_X4 U13205 ( .A(n11046), .ZN(n13707) );
  INV_X4 U13206 ( .A(n11046), .ZN(n13706) );
  INV_X4 U13207 ( .A(n11086), .ZN(n13816) );
  INV_X4 U13208 ( .A(n11086), .ZN(n13815) );
  INV_X4 U13209 ( .A(n11057), .ZN(n13247) );
  INV_X4 U13210 ( .A(n11057), .ZN(n13246) );
  INV_X4 U13211 ( .A(n11063), .ZN(n13681) );
  INV_X4 U13212 ( .A(n11063), .ZN(n13680) );
  INV_X4 U13213 ( .A(n11061), .ZN(n13254) );
  INV_X4 U13214 ( .A(n11061), .ZN(n13255) );
  NAND3_X2 U13215 ( .A1(n18350), .A2(n18349), .A3(n18348), .ZN(n18397) );
  INV_X4 U13216 ( .A(n10839), .ZN(n13309) );
  INV_X4 U13217 ( .A(n10839), .ZN(n13308) );
  INV_X4 U13218 ( .A(n10907), .ZN(n13311) );
  INV_X4 U13219 ( .A(n10907), .ZN(n13310) );
  INV_X4 U13220 ( .A(n10909), .ZN(n13313) );
  INV_X4 U13221 ( .A(n10909), .ZN(n13312) );
  INV_X4 U13222 ( .A(n10934), .ZN(n13317) );
  INV_X4 U13223 ( .A(n10934), .ZN(n13316) );
  INV_X4 U13224 ( .A(n10908), .ZN(n13319) );
  INV_X4 U13225 ( .A(n10908), .ZN(n13318) );
  INV_X4 U13226 ( .A(n11083), .ZN(n13476) );
  INV_X4 U13227 ( .A(n11083), .ZN(n13477) );
  OR2_X4 U13228 ( .A1(n18759), .A2(n14257), .ZN(n12569) );
  INV_X4 U13229 ( .A(n11060), .ZN(n13710) );
  INV_X4 U13230 ( .A(n11060), .ZN(n13711) );
  INV_X4 U13231 ( .A(n11049), .ZN(n13714) );
  INV_X4 U13232 ( .A(n11049), .ZN(n13715) );
  INV_X4 U13233 ( .A(n11054), .ZN(n13718) );
  INV_X4 U13234 ( .A(n11054), .ZN(n13719) );
  INV_X4 U13235 ( .A(n11055), .ZN(n13722) );
  INV_X4 U13236 ( .A(n11055), .ZN(n13723) );
  OR2_X4 U13237 ( .A1(n18980), .A2(n18888), .ZN(n12600) );
  AND3_X4 U13238 ( .A1(ID_EXEC_OUT[63]), .A2(n13049), .A3(n13055), .ZN(n12602)
         );
  INV_X4 U13239 ( .A(n11076), .ZN(n13686) );
  INV_X4 U13240 ( .A(n11076), .ZN(n13687) );
  INV_X4 U13241 ( .A(n11080), .ZN(n13694) );
  INV_X4 U13242 ( .A(n11080), .ZN(n13695) );
  INV_X4 U13243 ( .A(n11077), .ZN(n13690) );
  INV_X4 U13244 ( .A(n11077), .ZN(n13691) );
  INV_X4 U13245 ( .A(n11081), .ZN(n13698) );
  INV_X4 U13246 ( .A(n11081), .ZN(n13699) );
  INV_X4 U13247 ( .A(n10556), .ZN(n13766) );
  INV_X4 U13248 ( .A(n10556), .ZN(n13767) );
  INV_X4 U13249 ( .A(n10950), .ZN(n13552) );
  INV_X4 U13250 ( .A(n10950), .ZN(n13553) );
  INV_X4 U13251 ( .A(n10960), .ZN(n13556) );
  INV_X4 U13252 ( .A(n10960), .ZN(n13557) );
  INV_X4 U13253 ( .A(n10951), .ZN(n13560) );
  INV_X4 U13254 ( .A(n10951), .ZN(n13561) );
  INV_X4 U13255 ( .A(n10961), .ZN(n13564) );
  INV_X4 U13256 ( .A(n10961), .ZN(n13565) );
  INV_X4 U13257 ( .A(n10952), .ZN(n13568) );
  INV_X4 U13258 ( .A(n10952), .ZN(n13569) );
  INV_X4 U13259 ( .A(n10962), .ZN(n13572) );
  INV_X4 U13260 ( .A(n10962), .ZN(n13573) );
  INV_X4 U13261 ( .A(n10953), .ZN(n13576) );
  INV_X4 U13262 ( .A(n10953), .ZN(n13577) );
  INV_X4 U13263 ( .A(n10963), .ZN(n13580) );
  INV_X4 U13264 ( .A(n10963), .ZN(n13581) );
  INV_X4 U13265 ( .A(n10954), .ZN(n13584) );
  INV_X4 U13266 ( .A(n10954), .ZN(n13585) );
  INV_X4 U13267 ( .A(n10964), .ZN(n13588) );
  INV_X4 U13268 ( .A(n10964), .ZN(n13589) );
  INV_X4 U13269 ( .A(n10955), .ZN(n13592) );
  INV_X4 U13270 ( .A(n10955), .ZN(n13593) );
  INV_X4 U13271 ( .A(n10965), .ZN(n13596) );
  INV_X4 U13272 ( .A(n10965), .ZN(n13597) );
  INV_X4 U13273 ( .A(n10966), .ZN(n13600) );
  INV_X4 U13274 ( .A(n10966), .ZN(n13601) );
  INV_X4 U13275 ( .A(n10956), .ZN(n13604) );
  INV_X4 U13276 ( .A(n10956), .ZN(n13605) );
  INV_X4 U13277 ( .A(n10967), .ZN(n13608) );
  INV_X4 U13278 ( .A(n10967), .ZN(n13609) );
  INV_X4 U13279 ( .A(n10544), .ZN(n13748) );
  INV_X4 U13280 ( .A(n10544), .ZN(n13749) );
  INV_X4 U13281 ( .A(n11091), .ZN(n13754) );
  INV_X4 U13282 ( .A(n11091), .ZN(n13755) );
  INV_X4 U13283 ( .A(n11092), .ZN(n13760) );
  INV_X4 U13284 ( .A(n11092), .ZN(n13761) );
  INV_X4 U13285 ( .A(n10549), .ZN(n13762) );
  INV_X4 U13286 ( .A(n10549), .ZN(n13763) );
  INV_X4 U13287 ( .A(n11084), .ZN(n13784) );
  INV_X4 U13288 ( .A(n11084), .ZN(n13785) );
  INV_X4 U13289 ( .A(n10546), .ZN(n13788) );
  INV_X4 U13290 ( .A(n10546), .ZN(n13789) );
  INV_X4 U13291 ( .A(n10553), .ZN(n13792) );
  INV_X4 U13292 ( .A(n10553), .ZN(n13793) );
  INV_X4 U13293 ( .A(n11087), .ZN(n13819) );
  INV_X4 U13294 ( .A(n11087), .ZN(n13820) );
  INV_X4 U13295 ( .A(n11088), .ZN(n13823) );
  INV_X4 U13296 ( .A(n11088), .ZN(n13824) );
  INV_X4 U13297 ( .A(n11089), .ZN(n13827) );
  INV_X4 U13298 ( .A(n11089), .ZN(n13828) );
  INV_X4 U13299 ( .A(n10551), .ZN(n13831) );
  INV_X4 U13300 ( .A(n10551), .ZN(n13832) );
  INV_X4 U13301 ( .A(n10552), .ZN(n13835) );
  INV_X4 U13302 ( .A(n10552), .ZN(n13836) );
  INV_X4 U13303 ( .A(n10541), .ZN(n13841) );
  INV_X4 U13304 ( .A(n10541), .ZN(n13842) );
  INV_X4 U13305 ( .A(n10548), .ZN(n13845) );
  INV_X4 U13306 ( .A(n10548), .ZN(n13846) );
  INV_X4 U13307 ( .A(n10554), .ZN(n13849) );
  INV_X4 U13308 ( .A(n10554), .ZN(n13850) );
  INV_X4 U13309 ( .A(n11095), .ZN(n13853) );
  INV_X4 U13310 ( .A(n11095), .ZN(n13854) );
  INV_X4 U13311 ( .A(n11096), .ZN(n13855) );
  INV_X4 U13312 ( .A(n11096), .ZN(n13856) );
  INV_X4 U13313 ( .A(n18698), .ZN(n13446) );
  INV_X4 U13314 ( .A(n13446), .ZN(n13444) );
  INV_X4 U13315 ( .A(n13446), .ZN(n13445) );
  INV_X4 U13316 ( .A(n15328), .ZN(n13268) );
  INV_X8 U13317 ( .A(n13268), .ZN(n13266) );
  INV_X8 U13318 ( .A(n13268), .ZN(n13267) );
  INV_X4 U13319 ( .A(n11058), .ZN(n13248) );
  INV_X4 U13320 ( .A(n11058), .ZN(n13249) );
  INV_X4 U13321 ( .A(n11037), .ZN(n13618) );
  INV_X4 U13322 ( .A(n11037), .ZN(n13619) );
  INV_X4 U13323 ( .A(n11038), .ZN(n13674) );
  INV_X4 U13324 ( .A(n11038), .ZN(n13675) );
  INV_X4 U13325 ( .A(n11069), .ZN(n13622) );
  INV_X4 U13326 ( .A(n11069), .ZN(n13623) );
  INV_X4 U13327 ( .A(n11064), .ZN(n13626) );
  INV_X4 U13328 ( .A(n11064), .ZN(n13627) );
  INV_X4 U13329 ( .A(n11070), .ZN(n13630) );
  INV_X4 U13330 ( .A(n11070), .ZN(n13631) );
  INV_X4 U13331 ( .A(n11071), .ZN(n13638) );
  INV_X4 U13332 ( .A(n11071), .ZN(n13639) );
  INV_X4 U13333 ( .A(n11072), .ZN(n13642) );
  INV_X4 U13334 ( .A(n11072), .ZN(n13643) );
  INV_X4 U13335 ( .A(n11065), .ZN(n13646) );
  INV_X4 U13336 ( .A(n11065), .ZN(n13647) );
  INV_X4 U13337 ( .A(n11073), .ZN(n13650) );
  INV_X4 U13338 ( .A(n11073), .ZN(n13651) );
  INV_X4 U13339 ( .A(n11066), .ZN(n13654) );
  INV_X4 U13340 ( .A(n11066), .ZN(n13655) );
  INV_X4 U13341 ( .A(n11067), .ZN(n13662) );
  INV_X4 U13342 ( .A(n11067), .ZN(n13663) );
  INV_X4 U13343 ( .A(n11068), .ZN(n13666) );
  INV_X4 U13344 ( .A(n11068), .ZN(n13667) );
  INV_X4 U13345 ( .A(n11074), .ZN(n13670) );
  INV_X4 U13346 ( .A(n11074), .ZN(n13671) );
  INV_X4 U13347 ( .A(n11052), .ZN(n13682) );
  INV_X4 U13348 ( .A(n11052), .ZN(n13683) );
  INV_X4 U13349 ( .A(n11085), .ZN(n13812) );
  INV_X4 U13350 ( .A(n11085), .ZN(n13811) );
  INV_X4 U13351 ( .A(n10550), .ZN(n13798) );
  INV_X4 U13352 ( .A(n10550), .ZN(n13797) );
  INV_X4 U13353 ( .A(n10557), .ZN(n13803) );
  INV_X4 U13354 ( .A(n10557), .ZN(n13802) );
  INV_X4 U13355 ( .A(n10555), .ZN(n13858) );
  INV_X4 U13356 ( .A(n10555), .ZN(n13857) );
  INV_X4 U13357 ( .A(n10542), .ZN(n13862) );
  INV_X4 U13358 ( .A(n10542), .ZN(n13861) );
  INV_X4 U13359 ( .A(n11090), .ZN(n13751) );
  INV_X4 U13360 ( .A(n11090), .ZN(n13750) );
  INV_X4 U13361 ( .A(n10545), .ZN(n13757) );
  INV_X4 U13362 ( .A(n10545), .ZN(n13756) );
  INV_X4 U13363 ( .A(n11093), .ZN(n13773) );
  INV_X4 U13364 ( .A(n11093), .ZN(n13772) );
  INV_X4 U13365 ( .A(n11094), .ZN(n13777) );
  INV_X4 U13366 ( .A(n11094), .ZN(n13776) );
  INV_X4 U13367 ( .A(n10532), .ZN(n13781) );
  INV_X4 U13368 ( .A(n10532), .ZN(n13780) );
  INV_X4 U13369 ( .A(n10547), .ZN(n13807) );
  INV_X4 U13370 ( .A(n10547), .ZN(n13808) );
  INV_X4 U13371 ( .A(n10957), .ZN(n13612) );
  INV_X4 U13372 ( .A(n10957), .ZN(n13613) );
  INV_X4 U13373 ( .A(n11062), .ZN(n13700) );
  INV_X4 U13374 ( .A(n11062), .ZN(n13701) );
  INV_X4 U13375 ( .A(n11044), .ZN(n13704) );
  INV_X4 U13376 ( .A(n11044), .ZN(n13705) );
  OR2_X1 U13377 ( .A1(n5513), .A2(n14239), .ZN(n12690) );
  AND2_X2 U13378 ( .A1(n15620), .A2(n15603), .ZN(n12713) );
  AND2_X4 U13379 ( .A1(n15617), .A2(n10197), .ZN(n12714) );
  INV_X4 U13380 ( .A(n11903), .ZN(n13518) );
  INV_X4 U13381 ( .A(n11903), .ZN(n13517) );
  INV_X4 U13382 ( .A(n11904), .ZN(n13514) );
  INV_X4 U13383 ( .A(n11904), .ZN(n13513) );
  INV_X4 U13384 ( .A(n11899), .ZN(n13536) );
  INV_X4 U13385 ( .A(n11899), .ZN(n13535) );
  OR2_X1 U13386 ( .A1(n17957), .A2(n13362), .ZN(n12718) );
  OR2_X1 U13387 ( .A1(n18429), .A2(n13362), .ZN(n12719) );
  OR2_X1 U13388 ( .A1(n18090), .A2(n13362), .ZN(n12720) );
  INV_X4 U13389 ( .A(n5776), .ZN(n13617) );
  INV_X4 U13390 ( .A(n13617), .ZN(n13616) );
  INV_X4 U13391 ( .A(n5727), .ZN(n13641) );
  INV_X4 U13392 ( .A(n13641), .ZN(n13640) );
  INV_X4 U13393 ( .A(n5723), .ZN(n13645) );
  INV_X4 U13394 ( .A(n13645), .ZN(n13644) );
  INV_X4 U13395 ( .A(n5673), .ZN(n13669) );
  INV_X4 U13396 ( .A(n13669), .ZN(n13668) );
  INV_X4 U13397 ( .A(n5667), .ZN(n13673) );
  INV_X4 U13398 ( .A(n13673), .ZN(n13672) );
  INV_X4 U13399 ( .A(n5773), .ZN(n13621) );
  INV_X4 U13400 ( .A(n13621), .ZN(n13620) );
  OAI21_X2 U13401 ( .B1(n5662), .B2(n5770), .A(n13934), .ZN(n5773) );
  INV_X4 U13402 ( .A(n5769), .ZN(n13625) );
  INV_X4 U13403 ( .A(n13625), .ZN(n13624) );
  OAI21_X2 U13404 ( .B1(n5668), .B2(n5770), .A(n13934), .ZN(n5769) );
  INV_X4 U13405 ( .A(n5721), .ZN(n13649) );
  INV_X4 U13406 ( .A(n13649), .ZN(n13648) );
  INV_X4 U13407 ( .A(n5717), .ZN(n13653) );
  INV_X4 U13408 ( .A(n13653), .ZN(n13652) );
  INV_X4 U13409 ( .A(n5684), .ZN(n13657) );
  INV_X4 U13410 ( .A(n13657), .ZN(n13656) );
  OAI21_X2 U13411 ( .B1(n5662), .B2(n5680), .A(n13934), .ZN(n5684) );
  INV_X4 U13412 ( .A(n5679), .ZN(n13661) );
  INV_X4 U13413 ( .A(n13661), .ZN(n13660) );
  OAI21_X2 U13414 ( .B1(n5668), .B2(n5680), .A(n13935), .ZN(n5679) );
  INV_X4 U13415 ( .A(n5630), .ZN(n13677) );
  INV_X4 U13416 ( .A(n13677), .ZN(n13676) );
  INV_X4 U13417 ( .A(n5897), .ZN(n13579) );
  INV_X4 U13418 ( .A(n13579), .ZN(n13578) );
  INV_X4 U13419 ( .A(n5895), .ZN(n13583) );
  INV_X4 U13420 ( .A(n13583), .ZN(n13582) );
  INV_X4 U13421 ( .A(n5818), .ZN(n13607) );
  INV_X4 U13422 ( .A(n13607), .ZN(n13606) );
  INV_X4 U13423 ( .A(n5813), .ZN(n13611) );
  INV_X4 U13424 ( .A(n13611), .ZN(n13610) );
  INV_X4 U13425 ( .A(n5907), .ZN(n13559) );
  INV_X4 U13426 ( .A(n13559), .ZN(n13558) );
  INV_X4 U13427 ( .A(n5905), .ZN(n13563) );
  INV_X4 U13428 ( .A(n13563), .ZN(n13562) );
  INV_X4 U13429 ( .A(n5903), .ZN(n13567) );
  INV_X4 U13430 ( .A(n13567), .ZN(n13566) );
  OAI21_X2 U13431 ( .B1(n5770), .B2(n5816), .A(n13933), .ZN(n5903) );
  INV_X4 U13432 ( .A(n5893), .ZN(n13587) );
  INV_X4 U13433 ( .A(n13587), .ZN(n13586) );
  INV_X4 U13434 ( .A(n5891), .ZN(n13591) );
  INV_X4 U13435 ( .A(n13591), .ZN(n13590) );
  INV_X4 U13436 ( .A(n5888), .ZN(n13595) );
  INV_X4 U13437 ( .A(n13595), .ZN(n13594) );
  INV_X4 U13438 ( .A(n5853), .ZN(n13603) );
  INV_X4 U13439 ( .A(n13603), .ZN(n13602) );
  OAI21_X2 U13440 ( .B1(n5680), .B2(n5816), .A(n13933), .ZN(n5853) );
  INV_X4 U13441 ( .A(n5777), .ZN(n13615) );
  INV_X4 U13442 ( .A(n13615), .ZN(n13614) );
  INV_X4 U13443 ( .A(n5767), .ZN(n13629) );
  INV_X4 U13444 ( .A(n13629), .ZN(n13628) );
  INV_X4 U13445 ( .A(n5732), .ZN(n13633) );
  INV_X4 U13446 ( .A(n13633), .ZN(n13632) );
  INV_X4 U13447 ( .A(n5729), .ZN(n13637) );
  INV_X4 U13448 ( .A(n13637), .ZN(n13636) );
  INV_X4 U13449 ( .A(n5675), .ZN(n13665) );
  INV_X4 U13450 ( .A(n13665), .ZN(n13664) );
  INV_X4 U13451 ( .A(n5910), .ZN(n13555) );
  INV_X4 U13452 ( .A(n13555), .ZN(n13554) );
  INV_X4 U13453 ( .A(n5901), .ZN(n13571) );
  INV_X4 U13454 ( .A(n13571), .ZN(n13570) );
  INV_X4 U13455 ( .A(n5899), .ZN(n13575) );
  INV_X4 U13456 ( .A(n13575), .ZN(n13574) );
  INV_X4 U13457 ( .A(n5886), .ZN(n13599) );
  INV_X4 U13458 ( .A(n13599), .ZN(n13598) );
  AND2_X4 U13459 ( .A1(net224704), .A2(nextPC_ex_out[3]), .ZN(n12745) );
  INV_X4 U13460 ( .A(n14646), .ZN(n13519) );
  INV_X4 U13461 ( .A(n14646), .ZN(n13520) );
  INV_X4 U13462 ( .A(n14648), .ZN(n13515) );
  INV_X4 U13463 ( .A(n14648), .ZN(n13516) );
  OR2_X4 U13464 ( .A1(IMEM_BUS_IN[1]), .A2(IMEM_BUS_IN[2]), .ZN(n12921) );
  INV_X4 U13465 ( .A(n11909), .ZN(n13532) );
  INV_X4 U13466 ( .A(n11909), .ZN(n13531) );
  INV_X4 U13467 ( .A(n11900), .ZN(n13528) );
  INV_X4 U13468 ( .A(n11900), .ZN(n13527) );
  INV_X4 U13469 ( .A(n11837), .ZN(n13524) );
  INV_X4 U13470 ( .A(n11837), .ZN(n13523) );
  INV_X4 U13471 ( .A(n11833), .ZN(n13227) );
  INV_X4 U13472 ( .A(n11833), .ZN(n13226) );
  INV_X4 U13473 ( .A(n11896), .ZN(n13231) );
  INV_X4 U13474 ( .A(n11896), .ZN(n13230) );
  INV_X4 U13475 ( .A(n11902), .ZN(n13533) );
  INV_X4 U13476 ( .A(n11902), .ZN(n13534) );
  INV_X4 U13477 ( .A(n1882), .ZN(n13734) );
  INV_X16 U13478 ( .A(n13734), .ZN(n13733) );
  INV_X16 U13479 ( .A(n13734), .ZN(n13732) );
  INV_X4 U13480 ( .A(net223104), .ZN(net231615) );
  INV_X8 U13481 ( .A(n10944), .ZN(n13463) );
  INV_X4 U13482 ( .A(n11908), .ZN(n13529) );
  INV_X4 U13483 ( .A(n11908), .ZN(n13530) );
  INV_X4 U13484 ( .A(n11835), .ZN(n13525) );
  INV_X4 U13485 ( .A(n11835), .ZN(n13526) );
  INV_X4 U13486 ( .A(n11836), .ZN(n13521) );
  INV_X4 U13487 ( .A(n11836), .ZN(n13522) );
  INV_X4 U13488 ( .A(n11910), .ZN(n13228) );
  INV_X4 U13489 ( .A(n11910), .ZN(n13229) );
  INV_X4 U13490 ( .A(n11897), .ZN(n13232) );
  INV_X4 U13491 ( .A(n11897), .ZN(n13233) );
  INV_X4 U13492 ( .A(n11907), .ZN(n13511) );
  INV_X4 U13493 ( .A(n11907), .ZN(n13512) );
  INV_X8 U13494 ( .A(n10369), .ZN(net232877) );
  OR2_X4 U13495 ( .A1(n16753), .A2(n13362), .ZN(n12922) );
  OR2_X1 U13496 ( .A1(n18047), .A2(n13362), .ZN(n12923) );
  OR2_X1 U13497 ( .A1(n18135), .A2(n13362), .ZN(n12924) );
  OR2_X1 U13498 ( .A1(n18176), .A2(n13362), .ZN(n12925) );
  OR2_X1 U13499 ( .A1(n18221), .A2(n13362), .ZN(n12926) );
  OR2_X1 U13500 ( .A1(n18510), .A2(n13362), .ZN(n12927) );
  OR2_X4 U13501 ( .A1(n18930), .A2(n13362), .ZN(n12928) );
  INV_X8 U13502 ( .A(n10350), .ZN(n13440) );
  INV_X4 U13503 ( .A(n13440), .ZN(n13441) );
  OR2_X1 U13504 ( .A1(n17141), .A2(n13361), .ZN(n12929) );
  OR2_X1 U13505 ( .A1(n18570), .A2(n13361), .ZN(n12930) );
  OR2_X1 U13506 ( .A1(n17905), .A2(n13361), .ZN(n12931) );
  OR2_X1 U13507 ( .A1(n17470), .A2(n13361), .ZN(n12932) );
  OR2_X1 U13508 ( .A1(n17681), .A2(n13361), .ZN(n12933) );
  OR2_X1 U13509 ( .A1(n17808), .A2(n13361), .ZN(n12934) );
  INV_X8 U13510 ( .A(n18271), .ZN(n13387) );
  INV_X8 U13511 ( .A(n13387), .ZN(n13385) );
  AND2_X2 U13512 ( .A1(n13493), .A2(n12030), .ZN(n12935) );
  INV_X4 U13513 ( .A(n11911), .ZN(n13414) );
  INV_X4 U13514 ( .A(n11911), .ZN(n13413) );
  AND2_X4 U13515 ( .A1(n15644), .A2(n15643), .ZN(n12936) );
  INV_X4 U13516 ( .A(n11834), .ZN(n13234) );
  INV_X4 U13517 ( .A(n11834), .ZN(n13235) );
  INV_X4 U13518 ( .A(n11901), .ZN(n13242) );
  INV_X4 U13519 ( .A(n11901), .ZN(n13243) );
  INV_X4 U13520 ( .A(n11898), .ZN(n13240) );
  INV_X4 U13521 ( .A(n11898), .ZN(n13241) );
  INV_X4 U13522 ( .A(n11906), .ZN(n13264) );
  INV_X4 U13523 ( .A(n11906), .ZN(n13265) );
  NAND3_X1 U13524 ( .A1(n18774), .A2(n13221), .A3(n12016), .ZN(n14242) );
  AND2_X2 U13525 ( .A1(n19130), .A2(n19128), .ZN(n12954) );
  INV_X8 U13526 ( .A(n10833), .ZN(n13471) );
  INV_X8 U13527 ( .A(n10827), .ZN(n13422) );
  AND2_X4 U13528 ( .A1(n14265), .A2(n14264), .ZN(n12955) );
  INV_X4 U13529 ( .A(n18586), .ZN(n13410) );
  INV_X4 U13530 ( .A(n18586), .ZN(n13409) );
  INV_X4 U13531 ( .A(n15329), .ZN(n13271) );
  INV_X8 U13532 ( .A(n13271), .ZN(n13270) );
  OR2_X4 U13533 ( .A1(n1866), .A2(n12023), .ZN(n12956) );
  OR2_X4 U13534 ( .A1(n1866), .A2(n12027), .ZN(n12957) );
  INV_X4 U13535 ( .A(n2184), .ZN(n13728) );
  OR2_X1 U13536 ( .A1(n1866), .A2(n12300), .ZN(n12958) );
  INV_X4 U13537 ( .A(n17776), .ZN(n13384) );
  OR2_X4 U13538 ( .A1(n1866), .A2(n10816), .ZN(n12959) );
  INV_X1 U13540 ( .A(n13159), .ZN(n18462) );
  OR2_X4 U13541 ( .A1(n1866), .A2(n12021), .ZN(n12960) );
  OR2_X4 U13542 ( .A1(n1866), .A2(n11983), .ZN(n12961) );
  AND2_X4 U13543 ( .A1(n10840), .A2(n12039), .ZN(n12962) );
  OR2_X4 U13544 ( .A1(n1866), .A2(n18790), .ZN(n12963) );
  OR2_X4 U13545 ( .A1(n18662), .A2(n13362), .ZN(n12964) );
  OR2_X4 U13546 ( .A1(n18616), .A2(n18615), .ZN(n12965) );
  OR2_X4 U13547 ( .A1(n1866), .A2(n12039), .ZN(n12966) );
  OR2_X4 U13548 ( .A1(n1866), .A2(n18794), .ZN(n12967) );
  INV_X8 U13549 ( .A(n16816), .ZN(n13360) );
  INV_X16 U13550 ( .A(n13360), .ZN(n13358) );
  OR2_X4 U13551 ( .A1(n1866), .A2(n12028), .ZN(n12968) );
  OR2_X4 U13552 ( .A1(n1866), .A2(n10838), .ZN(n12969) );
  OR2_X4 U13553 ( .A1(n16844), .A2(n13362), .ZN(n12970) );
  OR2_X4 U13554 ( .A1(n15978), .A2(n13362), .ZN(n12971) );
  OR2_X4 U13555 ( .A1(n16441), .A2(n13362), .ZN(n12972) );
  OR2_X4 U13556 ( .A1(n16176), .A2(n13362), .ZN(n12973) );
  OR2_X4 U13557 ( .A1(n16494), .A2(n13362), .ZN(n12974) );
  INV_X1 U13558 ( .A(n13216), .ZN(n13217) );
  OR2_X4 U13559 ( .A1(n17168), .A2(n13362), .ZN(n12975) );
  OR2_X4 U13560 ( .A1(n16639), .A2(n13362), .ZN(n12976) );
  INV_X4 U13561 ( .A(n13205), .ZN(n13206) );
  INV_X4 U13562 ( .A(n18745), .ZN(n13205) );
  INV_X1 U13563 ( .A(n13207), .ZN(n17908) );
  INV_X8 U13564 ( .A(n13164), .ZN(n13165) );
  NAND2_X1 U13565 ( .A1(net239344), .A2(net224404), .ZN(n12977) );
  INV_X1 U13566 ( .A(n13213), .ZN(n18302) );
  INV_X4 U13567 ( .A(n18697), .ZN(n13439) );
  INV_X4 U13568 ( .A(n18721), .ZN(n13466) );
  INV_X4 U13569 ( .A(n10198), .ZN(n13551) );
  INV_X4 U13570 ( .A(n10198), .ZN(n13548) );
  INV_X4 U13571 ( .A(n10198), .ZN(n13549) );
  INV_X1 U13572 ( .A(net231361), .ZN(net231359) );
  INV_X2 U13573 ( .A(net231283), .ZN(net231263) );
  INV_X4 U13574 ( .A(reset), .ZN(n13944) );
  INV_X4 U13575 ( .A(n13953), .ZN(n13930) );
  INV_X4 U13576 ( .A(n13952), .ZN(n13928) );
  INV_X4 U13577 ( .A(n13944), .ZN(n13927) );
  INV_X4 U13578 ( .A(EXEC_STAGE_mul_ex_N378), .ZN(n13867) );
  INV_X4 U13579 ( .A(n13867), .ZN(n13866) );
  INV_X4 U13580 ( .A(n13867), .ZN(n13865) );
  INV_X4 U13581 ( .A(EXEC_STAGE_mul_ex_N444), .ZN(n13873) );
  INV_X4 U13582 ( .A(n13873), .ZN(n13871) );
  INV_X4 U13583 ( .A(n13873), .ZN(n13872) );
  INV_X4 U13584 ( .A(EXEC_STAGE_mul_ex_N411), .ZN(n13870) );
  INV_X4 U13585 ( .A(n13870), .ZN(n13868) );
  INV_X4 U13586 ( .A(n13870), .ZN(n13869) );
  INV_X4 U13587 ( .A(n7283), .ZN(n13542) );
  INV_X4 U13588 ( .A(n7283), .ZN(n13543) );
  INV_X4 U13589 ( .A(n10106), .ZN(n13547) );
  NOR3_X2 U13590 ( .A1(EXEC_STAGE_mul_ex_CurrentState_1_), .A2(
        EXEC_STAGE_mul_ex_CurrentState_2_), .A3(n10159), .ZN(n10106) );
  INV_X4 U13591 ( .A(n13547), .ZN(n13544) );
  INV_X4 U13592 ( .A(n13547), .ZN(n13545) );
  INV_X4 U13593 ( .A(n7284), .ZN(n13541) );
  INV_X4 U13594 ( .A(n7286), .ZN(n13537) );
  INV_X4 U13595 ( .A(n7286), .ZN(n13538) );
  INV_X4 U13596 ( .A(n7288), .ZN(n13539) );
  INV_X4 U13597 ( .A(n7288), .ZN(n13540) );
  NAND3_X2 U13598 ( .A1(n14203), .A2(n14204), .A3(n14202), .ZN(n14210) );
  INV_X8 U13599 ( .A(n18777), .ZN(n15379) );
  OAI22_X1 U13600 ( .A1(n12306), .A2(net231261), .B1(net230377), .B2(n18777), 
        .ZN(n7890) );
  INV_X8 U13601 ( .A(n15489), .ZN(n15491) );
  NOR2_X1 U13602 ( .A1(n13186), .A2(n12937), .ZN(n14993) );
  NOR2_X1 U13603 ( .A1(n13186), .A2(n12938), .ZN(n15014) );
  NOR2_X1 U13604 ( .A1(n13186), .A2(n12939), .ZN(n15030) );
  NOR2_X1 U13605 ( .A1(n13186), .A2(n12940), .ZN(n15056) );
  NOR2_X1 U13606 ( .A1(n13186), .A2(n12941), .ZN(n15077) );
  NOR2_X1 U13607 ( .A1(n13186), .A2(n12942), .ZN(n15093) );
  NOR2_X1 U13608 ( .A1(n13186), .A2(n12943), .ZN(n15124) );
  NOR2_X1 U13609 ( .A1(n13186), .A2(n12944), .ZN(n15145) );
  NOR2_X1 U13610 ( .A1(n13186), .A2(n12945), .ZN(n16128) );
  NOR2_X1 U13611 ( .A1(n13186), .A2(n12946), .ZN(n16277) );
  NOR2_X1 U13612 ( .A1(n13186), .A2(n12947), .ZN(n16377) );
  NOR2_X1 U13613 ( .A1(n13186), .A2(n12948), .ZN(n16605) );
  NOR2_X1 U13614 ( .A1(n13186), .A2(n12949), .ZN(n16945) );
  NOR2_X1 U13615 ( .A1(n13186), .A2(n12950), .ZN(n17018) );
  NOR2_X1 U13616 ( .A1(n13186), .A2(n12951), .ZN(n17272) );
  NOR2_X1 U13617 ( .A1(n13186), .A2(n12952), .ZN(n16709) );
  INV_X8 U13618 ( .A(n17269), .ZN(n13185) );
  AND2_X4 U13619 ( .A1(n2532), .A2(n1790), .ZN(n2528) );
  AND2_X2 U13620 ( .A1(IMEM_BUS_OUT[19]), .A2(IMEM_BUS_OUT[20]), .ZN(n12980)
         );
  INV_X8 U13621 ( .A(n15464), .ZN(n12979) );
  AND2_X2 U13622 ( .A1(n12979), .A2(IMEM_BUS_OUT[20]), .ZN(n15459) );
  NAND2_X4 U13623 ( .A1(n13359), .A2(n17712), .ZN(net223079) );
  OAI211_X1 U13624 ( .C1(n17541), .C2(n17540), .A(n17539), .B(n17538), .ZN(
        n17542) );
  INV_X8 U13625 ( .A(n17685), .ZN(n18310) );
  OAI21_X1 U13626 ( .B1(n15432), .B2(IMEM_BUS_OUT[7]), .A(n15431), .ZN(n16467)
         );
  INV_X1 U13627 ( .A(n15431), .ZN(n15429) );
  INV_X1 U13628 ( .A(n14210), .ZN(n14211) );
  NAND2_X1 U13629 ( .A1(n15438), .A2(n15437), .ZN(n17031) );
  NOR2_X1 U13631 ( .A1(n12318), .A2(n15437), .ZN(n15432) );
  XNOR2_X1 U13632 ( .A(n15437), .B(n12318), .ZN(n16974) );
  INV_X8 U13633 ( .A(destReg_wb_out[4]), .ZN(n19320) );
  INV_X32 U13634 ( .A(n13186), .ZN(n19152) );
  OAI211_X2 U13635 ( .C1(n19099), .C2(n18641), .A(n18474), .B(n18473), .ZN(
        n18529) );
  NAND2_X1 U13636 ( .A1(n15632), .A2(n1790), .ZN(n18745) );
  INV_X1 U13637 ( .A(n1790), .ZN(n19300) );
  NAND3_X1 U13638 ( .A1(n14996), .A2(n10157), .A3(n1790), .ZN(n17768) );
  NAND2_X4 U13639 ( .A1(n5506), .A2(n14235), .ZN(n1790) );
  AOI222_X2 U13640 ( .A1(n19153), .A2(REG_FILE_reg_out_14__17_), .B1(n13499), 
        .B2(REG_FILE_reg_out_4__17_), .C1(n19152), .C2(
        REG_FILE_reg_out_20__17_), .ZN(n2152) );
  OAI21_X2 U13641 ( .B1(IMEM_BUS_OUT[4]), .B2(n15403), .A(n15452), .ZN(n17284)
         );
  INV_X8 U13642 ( .A(n18775), .ZN(n15375) );
  OAI22_X1 U13643 ( .A1(n12307), .A2(net231261), .B1(net230377), .B2(n18775), 
        .ZN(n7884) );
  INV_X8 U13644 ( .A(n15631), .ZN(n13166) );
  INV_X1 U13645 ( .A(n13167), .ZN(n15356) );
  INV_X1 U13646 ( .A(n13167), .ZN(n15358) );
  INV_X1 U13647 ( .A(n13167), .ZN(n15365) );
  OAI21_X1 U13648 ( .B1(IMEM_BUS_OUT[5]), .B2(n15402), .A(n15451), .ZN(n16958)
         );
  AOI21_X2 U13649 ( .B1(n13492), .B2(n18399), .A(n18398), .ZN(n18400) );
  NAND3_X2 U13650 ( .A1(n15603), .A2(n14998), .A3(n12016), .ZN(n14194) );
  OAI21_X1 U13651 ( .B1(IMEM_BUS_OUT[6]), .B2(n15429), .A(n15428), .ZN(n16968)
         );
  NOR3_X2 U13652 ( .A1(ID_STAGE_imm16_aluA[28]), .A2(offset_26_id[1]), .A3(
        offset_26_id[5]), .ZN(n14196) );
  NOR3_X1 U13653 ( .A1(offset_26_id[0]), .A2(offset_26_id[1]), .A3(
        EXEC_MEM_OUT_141), .ZN(n2527) );
  NOR3_X1 U13654 ( .A1(EXEC_MEM_OUT_141), .A2(offset_26_id[1]), .A3(n10360), 
        .ZN(n2530) );
  AND2_X4 U13655 ( .A1(n2527), .A2(n2528), .ZN(n2511) );
  OAI21_X2 U13656 ( .B1(n13220), .B2(n15370), .A(n15369), .ZN(n18776) );
  NAND2_X4 U13657 ( .A1(n13166), .A2(n5558), .ZN(n15370) );
  NAND3_X1 U13658 ( .A1(IMEM_BUS_OUT[15]), .A2(IMEM_BUS_OUT[16]), .A3(n12992), 
        .ZN(n12983) );
  AOI22_X1 U13659 ( .A1(net231311), .A2(EXEC_STAGE_imm16_32[31]), .B1(
        ID_STAGE_imm16_aluA[31]), .B2(net230393), .ZN(n5586) );
  NAND2_X1 U13660 ( .A1(n14265), .A2(ID_STAGE_imm16_aluA[31]), .ZN(n14251) );
  NAND2_X1 U13661 ( .A1(ID_STAGE_imm16_aluA[31]), .A2(n12027), .ZN(n14233) );
  NAND3_X2 U13662 ( .A1(n14255), .A2(n18768), .A3(n18771), .ZN(n14191) );
  NAND3_X1 U13663 ( .A1(net230387), .A2(IF_ID_OUT[37]), .A3(n14217), .ZN(n5535) );
  OAI22_X1 U13664 ( .A1(n12212), .A2(net231261), .B1(IF_ID_OUT[37]), .B2(
        n18787), .ZN(n7878) );
  NAND3_X1 U13665 ( .A1(n18780), .A2(IF_ID_OUT[37]), .A3(n12016), .ZN(n18782)
         );
  NAND4_X1 U13666 ( .A1(n19163), .A2(IF_ID_OUT[37]), .A3(n18768), .A4(n18767), 
        .ZN(n18846) );
  NAND3_X1 U13667 ( .A1(n14255), .A2(n13221), .A3(n14254), .ZN(n14260) );
  AOI21_X1 U13668 ( .B1(n14243), .B2(n14255), .A(n19300), .ZN(n14230) );
  NAND3_X1 U13669 ( .A1(IF_ID_OUT[37]), .A2(n12029), .A3(n13221), .ZN(n5513)
         );
  INV_X2 U13670 ( .A(n14255), .ZN(n14225) );
  NAND2_X1 U13671 ( .A1(IF_ID_OUT[37]), .A2(n12016), .ZN(n15392) );
  AND2_X4 U13672 ( .A1(n2530), .A2(n2528), .ZN(n2503) );
  OAI21_X1 U13673 ( .B1(n17873), .B2(n18003), .A(n17759), .ZN(n17760) );
  INV_X1 U13674 ( .A(n15398), .ZN(n12985) );
  XNOR2_X2 U13675 ( .A(n16536), .B(n16537), .ZN(n16538) );
  NOR2_X2 U13676 ( .A1(n13154), .A2(n13877), .ZN(n13963) );
  NAND3_X1 U13677 ( .A1(n5529), .A2(ID_STAGE_imm16_aluA[29]), .A3(n13167), 
        .ZN(n14246) );
  NOR2_X2 U13678 ( .A1(ID_STAGE_imm16_aluA[29]), .A2(n10840), .ZN(n14219) );
  NOR2_X2 U13679 ( .A1(offset_26_id[0]), .A2(ID_STAGE_imm16_aluA[29]), .ZN(
        n14189) );
  NAND2_X1 U13680 ( .A1(net230387), .A2(ID_STAGE_imm16_aluA[29]), .ZN(n14187)
         );
  XNOR2_X1 U13681 ( .A(n18562), .B(n18561), .ZN(n18563) );
  OAI21_X2 U13682 ( .B1(n17131), .B2(n17130), .A(n16786), .ZN(n16788) );
  AOI21_X2 U13683 ( .B1(n18316), .B2(n13492), .A(n18315), .ZN(n18317) );
  INV_X1 U13684 ( .A(n12983), .ZN(n15420) );
  INV_X1 U13685 ( .A(n19351), .ZN(n15417) );
  OAI21_X4 U13686 ( .B1(n15796), .B2(n15795), .A(n17895), .ZN(n15801) );
  OAI22_X2 U13687 ( .A1(n17875), .A2(n17874), .B1(n17873), .B2(n18008), .ZN(
        n17876) );
  AND2_X4 U13688 ( .A1(n2533), .A2(n2528), .ZN(n2506) );
  NAND2_X1 U13689 ( .A1(offset_26_id[2]), .A2(net231271), .ZN(n18826) );
  NAND2_X1 U13690 ( .A1(offset_26_id[2]), .A2(net230387), .ZN(n18825) );
  NAND3_X1 U13691 ( .A1(offset_26_id[2]), .A2(n10844), .A3(n10368), .ZN(n14271) );
  NAND2_X1 U13692 ( .A1(n15418), .A2(n15417), .ZN(n16617) );
  NOR2_X1 U13693 ( .A1(n12317), .A2(n15417), .ZN(n15413) );
  XNOR2_X1 U13694 ( .A(n15417), .B(n12317), .ZN(n16520) );
  NAND3_X2 U13695 ( .A1(n17891), .A2(n17890), .A3(n17889), .ZN(n7632) );
  NAND2_X1 U13696 ( .A1(offset_26_id[9]), .A2(net231325), .ZN(n18802) );
  NAND2_X1 U13697 ( .A1(offset_26_id[9]), .A2(net230387), .ZN(n18801) );
  NAND3_X1 U13698 ( .A1(offset_26_id[9]), .A2(n12953), .A3(n12982), .ZN(n14649) );
  NAND3_X1 U13699 ( .A1(offset_26_id[9]), .A2(n13220), .A3(n12982), .ZN(n14645) );
  XOR2_X1 U13700 ( .A(n19320), .B(offset_26_id[9]), .Z(n5464) );
  OAI21_X1 U13701 ( .B1(n15423), .B2(IMEM_BUS_OUT[15]), .A(n12983), .ZN(n16722) );
  AOI22_X1 U13702 ( .A1(net231301), .A2(EXEC_STAGE_imm26_32[27]), .B1(
        ID_STAGE_imm16_aluA[27]), .B2(net230393), .ZN(n5608) );
  AOI22_X1 U13703 ( .A1(net231311), .A2(EXEC_STAGE_imm16_32[27]), .B1(
        ID_STAGE_imm16_aluA[27]), .B2(net230393), .ZN(n5590) );
  NOR3_X1 U13704 ( .A1(ID_STAGE_imm16_aluA[26]), .A2(ID_STAGE_imm16_aluA[28]), 
        .A3(ID_STAGE_imm16_aluA[27]), .ZN(n5529) );
  NOR2_X1 U13705 ( .A1(ID_STAGE_imm16_aluA[27]), .A2(n19300), .ZN(n18189) );
  NOR3_X2 U13706 ( .A1(ID_STAGE_imm16_aluA[24]), .A2(ID_STAGE_imm16_aluA[26]), 
        .A3(ID_STAGE_imm16_aluA[27]), .ZN(n14195) );
  OAI22_X4 U13707 ( .A1(n15391), .A2(n15390), .B1(n15389), .B2(n15388), .ZN(
        n15397) );
  AND2_X2 U13708 ( .A1(n16395), .A2(n16396), .ZN(n12990) );
  NAND2_X1 U13709 ( .A1(n15874), .A2(net222497), .ZN(n16396) );
  OAI21_X4 U13710 ( .B1(n18662), .B2(n14123), .A(n18665), .ZN(n18653) );
  NAND3_X2 U13711 ( .A1(IMEM_BUS_OUT[15]), .A2(IMEM_BUS_OUT[16]), .A3(n12992), 
        .ZN(n15422) );
  INV_X1 U13712 ( .A(n12992), .ZN(n15440) );
  NAND2_X1 U13713 ( .A1(n18771), .A2(n11991), .ZN(n18772) );
  NAND2_X1 U13714 ( .A1(ID_STAGE_imm16_aluA[30]), .A2(net230387), .ZN(n18832)
         );
  NAND3_X1 U13715 ( .A1(n18756), .A2(ID_STAGE_imm16_aluA[30]), .A3(n12962), 
        .ZN(n18757) );
  NAND3_X1 U13716 ( .A1(n14256), .A2(n18771), .A3(ID_STAGE_imm16_aluA[28]), 
        .ZN(n14259) );
  NAND2_X1 U13717 ( .A1(n14231), .A2(n18771), .ZN(n14229) );
  AOI21_X1 U13718 ( .B1(n14223), .B2(n18771), .A(n14226), .ZN(n14227) );
  NAND2_X1 U13719 ( .A1(ID_STAGE_imm16_aluA[31]), .A2(ID_STAGE_imm16_aluA[30]), 
        .ZN(n14245) );
  NAND2_X1 U13720 ( .A1(ID_STAGE_imm16_aluA[30]), .A2(n12023), .ZN(n18766) );
  INV_X1 U13721 ( .A(n18665), .ZN(n18667) );
  NAND2_X4 U13722 ( .A1(n13356), .A2(ID_EXEC_OUT[32]), .ZN(n18665) );
  NAND2_X1 U13723 ( .A1(net223324), .A2(n19068), .ZN(n18244) );
  NAND2_X1 U13724 ( .A1(n19107), .A2(n19068), .ZN(n18634) );
  INV_X8 U13725 ( .A(n18587), .ZN(n19068) );
  NAND3_X2 U13726 ( .A1(n18768), .A2(IF_ID_OUT[36]), .A3(n12016), .ZN(n14208)
         );
  NAND2_X1 U13727 ( .A1(IF_ID_OUT[36]), .A2(n12020), .ZN(n5520) );
  AOI22_X1 U13728 ( .A1(n14247), .A2(n14255), .B1(n14265), .B2(n18771), .ZN(
        n14263) );
  NOR2_X1 U13729 ( .A1(IF_ID_OUT[36]), .A2(n12020), .ZN(n14236) );
  NAND3_X2 U13730 ( .A1(n17927), .A2(n17926), .A3(n17925), .ZN(n17930) );
  NOR2_X4 U13731 ( .A1(n12993), .A2(n15455), .ZN(n12992) );
  NAND2_X1 U13732 ( .A1(offset_26_id[3]), .A2(net231271), .ZN(n18822) );
  NAND2_X1 U13733 ( .A1(offset_26_id[3]), .A2(net230387), .ZN(n18821) );
  NAND3_X1 U13734 ( .A1(offset_26_id[3]), .A2(n12026), .A3(n10368), .ZN(n14280) );
  NAND2_X1 U13735 ( .A1(offset_26_id[3]), .A2(offset_26_id[2]), .ZN(n14269) );
  NAND2_X1 U13736 ( .A1(n15475), .A2(n12985), .ZN(n18106) );
  NOR2_X1 U13737 ( .A1(n12319), .A2(n12985), .ZN(n15470) );
  XNOR2_X1 U13738 ( .A(n12985), .B(n12319), .ZN(n18063) );
  NAND2_X4 U13740 ( .A1(n16325), .A2(n16324), .ZN(n17040) );
  AOI21_X2 U13741 ( .B1(n16327), .B2(n13492), .A(n16326), .ZN(n16328) );
  NAND3_X2 U13742 ( .A1(n15480), .A2(IMEM_BUS_OUT[25]), .A3(IMEM_BUS_OUT[26]), 
        .ZN(n15474) );
  INV_X1 U13743 ( .A(n15459), .ZN(n15460) );
  NAND2_X4 U13744 ( .A1(IMEM_BUS_OUT[6]), .A2(n15401), .ZN(n15428) );
  INV_X8 U13745 ( .A(n15431), .ZN(n15401) );
  OAI21_X1 U13746 ( .B1(IMEM_BUS_OUT[18]), .B2(n15399), .A(n15455), .ZN(n17381) );
  INV_X1 U13747 ( .A(n15455), .ZN(n15441) );
  NAND2_X4 U13748 ( .A1(IMEM_BUS_OUT[18]), .A2(n15399), .ZN(n15455) );
  NAND3_X2 U13749 ( .A1(n16042), .A2(n16041), .A3(n16040), .ZN(n7367) );
  INV_X2 U13750 ( .A(n18547), .ZN(n18549) );
  NAND2_X1 U13751 ( .A1(n13484), .A2(n18653), .ZN(n18656) );
  OAI21_X2 U13752 ( .B1(n15725), .B2(n19101), .A(n18679), .ZN(n15726) );
  NOR2_X1 U13753 ( .A1(n18679), .A2(n18652), .ZN(n18658) );
  NAND2_X4 U13754 ( .A1(n19068), .A2(ID_EXEC_OUT[157]), .ZN(n18679) );
  OAI21_X1 U13755 ( .B1(n13218), .B2(n19105), .A(n13151), .ZN(n15829) );
  INV_X2 U13756 ( .A(n18322), .ZN(n18323) );
  XNOR2_X2 U13757 ( .A(n17979), .B(n13100), .ZN(n17980) );
  NAND2_X4 U13758 ( .A1(IMEM_BUS_OUT[4]), .A2(n15403), .ZN(n15452) );
  NAND2_X4 U13759 ( .A1(net239508), .A2(net233102), .ZN(n16557) );
  INV_X2 U13760 ( .A(n15447), .ZN(n15444) );
  NAND2_X4 U13761 ( .A1(IMEM_BUS_OUT[3]), .A2(n15448), .ZN(n15447) );
  NAND2_X4 U13762 ( .A1(n18322), .A2(n18324), .ZN(n17896) );
  OAI21_X2 U13763 ( .B1(n17582), .B2(n18550), .A(n17581), .ZN(n7592) );
  NAND2_X4 U13764 ( .A1(net223324), .A2(n16879), .ZN(n17993) );
  INV_X8 U13765 ( .A(n18679), .ZN(n16879) );
  AOI21_X2 U13766 ( .B1(n14105), .B2(
        WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[20]), .A(n14104), .ZN(n14001)
         );
  AOI21_X2 U13767 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[21]), .B2(
        n14105), .A(n14104), .ZN(n14006) );
  AOI21_X2 U13769 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[18]), .B2(
        n14105), .A(n14104), .ZN(n14026) );
  AOI21_X2 U13770 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[19]), .B2(
        n14019), .A(n14104), .ZN(n14031) );
  OAI22_X1 U13772 ( .A1(n12310), .A2(net231259), .B1(IMEM_BUS_OUT[29]), .B2(
        n13480), .ZN(n7728) );
  XNOR2_X1 U13773 ( .A(IMEM_BUS_OUT[28]), .B(IMEM_BUS_OUT[29]), .ZN(n18237) );
  NAND2_X4 U13774 ( .A1(IMEM_BUS_OUT[28]), .A2(IMEM_BUS_OUT[29]), .ZN(n15479)
         );
  OAI21_X1 U13775 ( .B1(IMEM_BUS_OUT[19]), .B2(n15459), .A(n15457), .ZN(n17432) );
  NAND2_X4 U13776 ( .A1(n12979), .A2(n12980), .ZN(n15457) );
  OAI21_X4 U13777 ( .B1(n13000), .B2(n15801), .A(n15800), .ZN(n17892) );
  INV_X8 U13778 ( .A(n15897), .ZN(n15907) );
  NAND3_X1 U13779 ( .A1(n16780), .A2(n17721), .A3(n17722), .ZN(n16782) );
  NAND3_X1 U13780 ( .A1(n17721), .A2(n17720), .A3(n17722), .ZN(n17726) );
  INV_X4 U13781 ( .A(n17721), .ZN(n15869) );
  INV_X2 U13782 ( .A(n18303), .ZN(n18307) );
  NAND2_X4 U13783 ( .A1(n17706), .A2(n17705), .ZN(n18303) );
  OAI21_X2 U13784 ( .B1(n17836), .B2(n13100), .A(n17835), .ZN(n17838) );
  NAND2_X4 U13785 ( .A1(n17722), .A2(n15850), .ZN(n15868) );
  AOI21_X2 U13786 ( .B1(n17714), .B2(n13492), .A(n17713), .ZN(n17715) );
  NOR2_X4 U13787 ( .A1(n14066), .A2(n14065), .ZN(n14067) );
  NAND2_X1 U13788 ( .A1(offset_26_id[4]), .A2(net231325), .ZN(n18818) );
  XOR2_X1 U13789 ( .A(n19320), .B(offset_26_id[4]), .Z(n2536) );
  NAND2_X1 U13790 ( .A1(offset_26_id[4]), .A2(net230387), .ZN(n18817) );
  NAND2_X1 U13791 ( .A1(n14272), .A2(offset_26_id[4]), .ZN(n14274) );
  NAND3_X1 U13792 ( .A1(offset_26_id[4]), .A2(offset_26_id[3]), .A3(n12026), 
        .ZN(n14277) );
  NAND3_X1 U13793 ( .A1(offset_26_id[4]), .A2(n12026), .A3(n10844), .ZN(n14276) );
  NAND3_X1 U13794 ( .A1(offset_26_id[4]), .A2(offset_26_id[2]), .A3(n10844), 
        .ZN(n14275) );
  INV_X16 U13795 ( .A(n15488), .ZN(n13351) );
  NAND2_X4 U13796 ( .A1(n15407), .A2(n13939), .ZN(n15488) );
  NOR2_X4 U13797 ( .A1(n12999), .A2(n18306), .ZN(n15780) );
  NAND2_X4 U13798 ( .A1(n18303), .A2(n17707), .ZN(n18304) );
  INV_X1 U13799 ( .A(n12994), .ZN(n16325) );
  AOI21_X1 U13800 ( .B1(n15480), .B2(IMEM_BUS_OUT[26]), .A(IMEM_BUS_OUT[25]), 
        .ZN(n15473) );
  XNOR2_X1 U13801 ( .A(IMEM_BUS_OUT[26]), .B(n15480), .ZN(n18151) );
  INV_X1 U13802 ( .A(n15480), .ZN(n15481) );
  AOI21_X4 U13803 ( .B1(n16395), .B2(n12996), .A(n12995), .ZN(n12994) );
  AND2_X2 U13804 ( .A1(n16396), .A2(n16397), .ZN(n12996) );
  NAND3_X4 U13805 ( .A1(n16077), .A2(n16080), .A3(n16078), .ZN(n15897) );
  XOR2_X1 U13806 ( .A(n18466), .B(n18467), .Z(n18477) );
  NAND2_X4 U13807 ( .A1(n18627), .A2(n19070), .ZN(n13097) );
  AND3_X4 U13808 ( .A1(n15671), .A2(n14098), .A3(n13055), .ZN(n12997) );
  XNOR2_X2 U13809 ( .A(n18621), .B(n13218), .ZN(n12998) );
  INV_X2 U13810 ( .A(n15791), .ZN(n15796) );
  AOI21_X4 U13811 ( .B1(n18622), .B2(n13492), .A(n13490), .ZN(n18627) );
  INV_X8 U13812 ( .A(n17558), .ZN(n16899) );
  NAND2_X4 U13813 ( .A1(n15913), .A2(n15914), .ZN(n17558) );
  AOI21_X4 U13814 ( .B1(n16903), .B2(n16904), .A(n16902), .ZN(n19149) );
  INV_X1 U13815 ( .A(n18306), .ZN(n17707) );
  NOR2_X2 U13816 ( .A1(n13000), .A2(n17500), .ZN(n17501) );
  INV_X4 U13817 ( .A(n13000), .ZN(n17893) );
  NAND2_X4 U13818 ( .A1(n14084), .A2(n14083), .ZN(n15671) );
  NAND2_X4 U13819 ( .A1(net239598), .A2(net239667), .ZN(n16469) );
  AOI21_X2 U13820 ( .B1(n18307), .B2(n18306), .A(n18305), .ZN(n18316) );
  OAI21_X4 U13821 ( .B1(net239454), .B2(n16963), .A(net225183), .ZN(n16966) );
  OAI21_X4 U13822 ( .B1(n16967), .B2(n16966), .A(n16965), .ZN(n7499) );
  NAND2_X2 U13824 ( .A1(n17285), .A2(net224699), .ZN(n17293) );
  INV_X2 U13825 ( .A(net224708), .ZN(net224699) );
  INV_X2 U13826 ( .A(n19108), .ZN(n19109) );
  OAI21_X1 U13827 ( .B1(IMEM_BUS_OUT[17]), .B2(n15441), .A(n15440), .ZN(n17116) );
  NOR2_X1 U13828 ( .A1(n12542), .A2(n15440), .ZN(n15423) );
  XNOR2_X1 U13829 ( .A(n15440), .B(n12542), .ZN(n16768) );
  OAI21_X1 U13830 ( .B1(IMEM_BUS_OUT[2]), .B2(n15444), .A(n15443), .ZN(n17211)
         );
  NAND2_X4 U13831 ( .A1(IMEM_BUS_OUT[2]), .A2(n15404), .ZN(n15443) );
  NOR3_X2 U13832 ( .A1(net225172), .A2(net225192), .A3(n16960), .ZN(n16967) );
  NAND2_X2 U13833 ( .A1(net239673), .A2(net224707), .ZN(n17292) );
  INV_X2 U13834 ( .A(n15769), .ZN(n12999) );
  NOR2_X4 U13835 ( .A1(n17502), .A2(n13001), .ZN(n13000) );
  AND3_X4 U13836 ( .A1(n17705), .A2(n15790), .A3(n15789), .ZN(n13001) );
  INV_X8 U13837 ( .A(net225172), .ZN(net239454) );
  NAND2_X4 U13838 ( .A1(n17213), .A2(n17214), .ZN(n17228) );
  OAI22_X1 U13839 ( .A1(n19313), .A2(net231263), .B1(net231313), .B2(n19312), 
        .ZN(n7888) );
  NOR3_X1 U13840 ( .A1(n10122), .A2(n19318), .A3(n10860), .ZN(n15498) );
  NAND2_X1 U13841 ( .A1(offset_26_id[8]), .A2(net231325), .ZN(n18806) );
  XOR2_X1 U13842 ( .A(n19317), .B(offset_26_id[8]), .Z(n5463) );
  NAND2_X1 U13843 ( .A1(offset_26_id[8]), .A2(net230387), .ZN(n18805) );
  NAND3_X1 U13844 ( .A1(offset_26_id[9]), .A2(offset_26_id[8]), .A3(n12953), 
        .ZN(n14656) );
  NAND3_X1 U13845 ( .A1(offset_26_id[8]), .A2(n13220), .A3(n12984), .ZN(n14641) );
  INV_X16 U13846 ( .A(n15485), .ZN(n13346) );
  NAND2_X4 U13847 ( .A1(n13482), .A2(n13939), .ZN(n15485) );
  NAND2_X4 U13848 ( .A1(net227255), .A2(net233181), .ZN(net239616) );
  NAND3_X2 U13849 ( .A1(net239616), .A2(net227207), .A3(net227192), .ZN(
        net227205) );
  INV_X16 U13850 ( .A(net233180), .ZN(net233181) );
  NAND3_X4 U13851 ( .A1(n10148), .A2(net239553), .A3(n13002), .ZN(net227221)
         );
  INV_X4 U13852 ( .A(n13007), .ZN(n13002) );
  NAND3_X1 U13853 ( .A1(n13002), .A2(net239553), .A3(n10148), .ZN(net239475)
         );
  XNOR2_X1 U13854 ( .A(nextPC_ex_out[27]), .B(n13002), .ZN(net223440) );
  MUX2_X2 U13855 ( .A(n11082), .B(n12258), .S(net239627), .Z(n13007) );
  MUX2_X2 U13856 ( .A(n11082), .B(n12258), .S(net239767), .Z(net227243) );
  INV_X8 U13857 ( .A(net233141), .ZN(net233142) );
  XNOR2_X2 U13858 ( .A(net227254), .B(net239756), .ZN(net223663) );
  NAND2_X2 U13859 ( .A1(net233181), .A2(net227255), .ZN(net239722) );
  NAND4_X4 U13860 ( .A1(n13018), .A2(n10124), .A3(n13005), .A4(net223447), 
        .ZN(net227220) );
  NAND3_X4 U13861 ( .A1(net227220), .A2(net227219), .A3(net227265), .ZN(
        net239254) );
  NAND4_X2 U13862 ( .A1(net227219), .A2(net227220), .A3(net227239), .A4(
        net227240), .ZN(net227213) );
  INV_X2 U13863 ( .A(nextPC_ex_out[27]), .ZN(net223447) );
  OAI22_X2 U13864 ( .A1(n11107), .A2(net231259), .B1(net230381), .B2(net223447), .ZN(n7682) );
  NAND4_X4 U13865 ( .A1(net227261), .A2(net239477), .A3(net222980), .A4(
        net223447), .ZN(net227219) );
  INV_X8 U13866 ( .A(n13003), .ZN(n13004) );
  NAND2_X4 U13867 ( .A1(net223366), .A2(net239220), .ZN(n13003) );
  NAND3_X4 U13868 ( .A1(net227089), .A2(net227088), .A3(net227087), .ZN(
        net227069) );
  OAI21_X4 U13869 ( .B1(net227075), .B2(n11934), .A(net227069), .ZN(net239017)
         );
  INV_X4 U13870 ( .A(net225778), .ZN(net227087) );
  NAND3_X4 U13871 ( .A1(net227079), .A2(net225684), .A3(net227090), .ZN(
        net227089) );
  NAND3_X4 U13872 ( .A1(net227094), .A2(net227095), .A3(n13009), .ZN(net227088) );
  NOR2_X4 U13873 ( .A1(nextPC_ex_out[13]), .A2(n13008), .ZN(n13009) );
  INV_X4 U13874 ( .A(net227077), .ZN(n13008) );
  XNOR2_X2 U13875 ( .A(n13008), .B(n11993), .ZN(net225681) );
  XNOR2_X2 U13876 ( .A(net225778), .B(n11934), .ZN(net225777) );
  OAI221_X4 U13877 ( .B1(net239767), .B2(net239371), .C1(n10111), .C2(
        net239628), .A(nextPC_ex_out[31]), .ZN(net222698) );
  NAND2_X1 U13878 ( .A1(n10140), .A2(net231325), .ZN(net222642) );
  INV_X16 U13879 ( .A(net233241), .ZN(net233242) );
  INV_X4 U13880 ( .A(net233216), .ZN(net233241) );
  INV_X8 U13881 ( .A(net233242), .ZN(net239782) );
  NAND3_X4 U13882 ( .A1(net227079), .A2(net225684), .A3(n11993), .ZN(net227081) );
  NAND3_X4 U13883 ( .A1(net227094), .A2(net227095), .A3(net227077), .ZN(
        net225780) );
  NAND3_X4 U13884 ( .A1(net227103), .A2(net227102), .A3(net227101), .ZN(
        net227093) );
  NAND2_X1 U13885 ( .A1(net239674), .A2(net224954), .ZN(net224953) );
  INV_X4 U13886 ( .A(net227117), .ZN(n13010) );
  NAND3_X4 U13887 ( .A1(net227105), .A2(n15552), .A3(n13010), .ZN(net227128)
         );
  XNOR2_X2 U13888 ( .A(nextPC_ex_out[18]), .B(n13010), .ZN(net224658) );
  NAND3_X2 U13889 ( .A1(net239404), .A2(net224491), .A3(net227119), .ZN(
        net227105) );
  NAND3_X2 U13890 ( .A1(net224660), .A2(net224661), .A3(nextPC_ex_out[18]), 
        .ZN(net224955) );
  NAND2_X2 U13891 ( .A1(n13011), .A2(net227121), .ZN(net224660) );
  INV_X8 U13892 ( .A(n13012), .ZN(n13011) );
  NAND2_X4 U13893 ( .A1(n13011), .A2(net227121), .ZN(net239473) );
  NAND2_X4 U13894 ( .A1(n13011), .A2(net227121), .ZN(net227122) );
  OAI21_X4 U13895 ( .B1(net227139), .B2(net227135), .A(net224493), .ZN(n13012)
         );
  NAND3_X4 U13896 ( .A1(net224491), .A2(net227143), .A3(n10242), .ZN(net239459) );
  NAND3_X2 U13897 ( .A1(net227143), .A2(net224491), .A3(net227119), .ZN(
        net227115) );
  NAND2_X1 U13898 ( .A1(nextPC_ex_out[19]), .A2(nextPC_ex_out[20]), .ZN(
        net239030) );
  NAND2_X2 U13899 ( .A1(net224404), .A2(nextPC_ex_out[19]), .ZN(net227135) );
  NAND3_X2 U13900 ( .A1(net227093), .A2(net227098), .A3(n11955), .ZN(net227084) );
  NAND2_X4 U13901 ( .A1(net227093), .A2(net227098), .ZN(net225528) );
  NAND3_X2 U13902 ( .A1(net227093), .A2(net227098), .A3(n11955), .ZN(net227086) );
  INV_X4 U13903 ( .A(net225450), .ZN(net227101) );
  NAND3_X4 U13904 ( .A1(net227107), .A2(net227108), .A3(n13014), .ZN(net227102) );
  NOR2_X4 U13905 ( .A1(nextPC_ex_out[16]), .A2(n13013), .ZN(n13014) );
  INV_X4 U13906 ( .A(net227110), .ZN(n13013) );
  XNOR2_X2 U13907 ( .A(n13013), .B(n11995), .ZN(net224952) );
  OAI21_X4 U13908 ( .B1(EXEC_STAGE_imm26_32[16]), .B2(net227290), .A(net232877), .ZN(net225450) );
  XNOR2_X2 U13909 ( .A(net225450), .B(n11928), .ZN(net225449) );
  NAND3_X4 U13910 ( .A1(net239459), .A2(net227122), .A3(n13015), .ZN(net227107) );
  NAND3_X4 U13911 ( .A1(net227108), .A2(net227107), .A3(net227110), .ZN(
        net225452) );
  NAND2_X4 U13912 ( .A1(net227205), .A2(net227204), .ZN(net224181) );
  INV_X8 U13913 ( .A(net224181), .ZN(net227201) );
  INV_X4 U13914 ( .A(net227208), .ZN(net227204) );
  NAND2_X2 U13915 ( .A1(net227216), .A2(n11985), .ZN(net227208) );
  NAND2_X2 U13916 ( .A1(nextPC_ex_out[22]), .A2(net227208), .ZN(net227231) );
  NAND2_X2 U13917 ( .A1(net223743), .A2(n11985), .ZN(net227236) );
  OAI22_X2 U13918 ( .A1(n11106), .A2(net231257), .B1(net230377), .B2(n11985), 
        .ZN(n7640) );
  NAND2_X1 U13919 ( .A1(net227216), .A2(net233131), .ZN(net223796) );
  NAND3_X4 U13920 ( .A1(n13017), .A2(net223442), .A3(net227259), .ZN(net227199) );
  INV_X2 U13921 ( .A(net227199), .ZN(net239630) );
  NAND2_X4 U13922 ( .A1(net227199), .A2(net239572), .ZN(net227214) );
  NOR2_X4 U13923 ( .A1(net227262), .A2(n13016), .ZN(n13017) );
  NAND2_X2 U13924 ( .A1(nextPC_ex_out[27]), .A2(net223444), .ZN(n13016) );
  BUF_X32 U13925 ( .A(net227262), .Z(net239669) );
  NAND3_X4 U13926 ( .A1(net233133), .A2(net227261), .A3(net239477), .ZN(
        net227259) );
  NAND3_X4 U13927 ( .A1(net227259), .A2(net223442), .A3(net227269), .ZN(
        net223666) );
  NAND3_X4 U13928 ( .A1(net227261), .A2(net239477), .A3(net239390), .ZN(
        net223442) );
  NAND2_X4 U13929 ( .A1(net227275), .A2(net223368), .ZN(net227274) );
  NAND2_X4 U13930 ( .A1(net223365), .A2(nextPC_ex_out[28]), .ZN(net227275) );
  NAND3_X2 U13931 ( .A1(net239329), .A2(net227277), .A3(net227276), .ZN(
        net223366) );
  INV_X8 U13932 ( .A(net222698), .ZN(net227282) );
  INV_X1 U13933 ( .A(n10135), .ZN(net239823) );
  NOR2_X4 U13934 ( .A1(net233106), .A2(net224709), .ZN(n13019) );
  NOR3_X4 U13935 ( .A1(net225204), .A2(n13019), .A3(net225203), .ZN(net225202)
         );
  NAND2_X2 U13936 ( .A1(net224704), .A2(n10355), .ZN(net224709) );
  OAI21_X4 U13937 ( .B1(net233078), .B2(net225207), .A(net225209), .ZN(
        net224708) );
  NOR2_X2 U13938 ( .A1(net225206), .A2(net224708), .ZN(net225204) );
  INV_X8 U13939 ( .A(net225210), .ZN(net225207) );
  AOI22_X2 U13940 ( .A1(net225184), .A2(net225185), .B1(net225186), .B2(
        net224713), .ZN(net225183) );
  NAND2_X4 U13941 ( .A1(net225214), .A2(net225209), .ZN(net239507) );
  NAND3_X2 U13942 ( .A1(nextPC_ex_out[4]), .A2(nextPC_ex_out[5]), .A3(
        net225209), .ZN(net227048) );
  NAND2_X4 U13943 ( .A1(net227086), .A2(net225529), .ZN(net227079) );
  NAND2_X4 U13944 ( .A1(net225528), .A2(nextPC_ex_out[15]), .ZN(net225684) );
  XNOR2_X2 U13945 ( .A(net225529), .B(nextPC_ex_out[15]), .ZN(net225526) );
  NAND2_X4 U13946 ( .A1(net225528), .A2(n12127), .ZN(net227095) );
  OAI21_X4 U13947 ( .B1(net239767), .B2(net239806), .A(n13020), .ZN(net227254)
         );
  NAND2_X4 U13948 ( .A1(net227270), .A2(net227271), .ZN(net223444) );
  NAND3_X1 U13949 ( .A1(n10137), .A2(net239828), .A3(net223444), .ZN(net223439) );
  INV_X4 U13950 ( .A(nextPC_ex_out[28]), .ZN(net227271) );
  INV_X4 U13951 ( .A(net223365), .ZN(net227270) );
  NAND3_X4 U13952 ( .A1(net227270), .A2(net239554), .A3(net239555), .ZN(
        net239553) );
  INV_X1 U13953 ( .A(net227270), .ZN(net239528) );
  NAND2_X1 U13954 ( .A1(nextPC_ex_out[25]), .A2(net227254), .ZN(net223742) );
  INV_X4 U13955 ( .A(nextPC_ex_out[28]), .ZN(net137317) );
  NAND2_X2 U13957 ( .A1(EXEC_MEM_OUT_114), .A2(net231323), .ZN(n13022) );
  NAND2_X2 U13958 ( .A1(EXEC_MEM_IN_250), .A2(n13023), .ZN(net139963) );
  INV_X4 U13959 ( .A(EXEC_STAGE_mul_done), .ZN(n13023) );
  INV_X4 U13960 ( .A(net225212), .ZN(n13021) );
  OAI221_X2 U13961 ( .B1(n13021), .B2(net222304), .C1(net232817), .C2(
        net223078), .A(net223079), .ZN(net223077) );
  NAND2_X2 U13962 ( .A1(net224704), .A2(nextPC_ex_out[5]), .ZN(net225206) );
  NAND2_X4 U13963 ( .A1(net227010), .A2(net227009), .ZN(net233078) );
  INV_X4 U13964 ( .A(net224847), .ZN(net227009) );
  AOI211_X4 U13965 ( .C1(net227009), .C2(n10357), .A(net225191), .B(net227048), 
        .ZN(net227040) );
  NAND3_X2 U13966 ( .A1(net224841), .A2(net224842), .A3(net224843), .ZN(
        net227010) );
  INV_X4 U13967 ( .A(net227012), .ZN(net224843) );
  NAND3_X2 U13968 ( .A1(net224843), .A2(net224841), .A3(net224842), .ZN(
        net224840) );
  NAND2_X2 U13969 ( .A1(n13025), .A2(net225188), .ZN(net224847) );
  NAND2_X2 U13970 ( .A1(net227033), .A2(nextPC_ex_out[6]), .ZN(n13025) );
  INV_X4 U13971 ( .A(net224816), .ZN(net227033) );
  AOI21_X2 U13972 ( .B1(net239379), .B2(net224853), .A(net227033), .ZN(
        net227035) );
  NAND2_X2 U13973 ( .A1(net227033), .A2(n10361), .ZN(net225185) );
  NAND3_X2 U13974 ( .A1(net224844), .A2(net224845), .A3(net224846), .ZN(
        net224841) );
  NAND3_X2 U13975 ( .A1(net227024), .A2(net225908), .A3(n12019), .ZN(n13026)
         );
  NAND3_X2 U13976 ( .A1(net227024), .A2(net225908), .A3(n12019), .ZN(net227015) );
  INV_X4 U13977 ( .A(net225076), .ZN(net227013) );
  NAND2_X2 U13978 ( .A1(net227053), .A2(net227047), .ZN(net239380) );
  NAND2_X2 U13979 ( .A1(n13024), .A2(net225187), .ZN(net227012) );
  INV_X4 U13980 ( .A(net225195), .ZN(n13024) );
  XNOR2_X2 U13981 ( .A(n13024), .B(n10357), .ZN(net225160) );
  NAND3_X4 U13982 ( .A1(net227128), .A2(n13027), .A3(n11995), .ZN(net225453)
         );
  NAND3_X4 U13984 ( .A1(net239459), .A2(net239473), .A3(nextPC_ex_out[18]), 
        .ZN(n13027) );
  NAND3_X4 U13985 ( .A1(net225893), .A2(net227063), .A3(n12018), .ZN(net225908) );
  OAI22_X2 U13986 ( .A1(n11538), .A2(net231251), .B1(net230381), .B2(n12018), 
        .ZN(n7421) );
  NAND2_X4 U13987 ( .A1(net239017), .A2(nextPC_ex_out[12]), .ZN(net227063) );
  NAND2_X4 U13988 ( .A1(net227068), .A2(net225824), .ZN(net225893) );
  NAND3_X4 U13989 ( .A1(net227073), .A2(net225893), .A3(n13028), .ZN(net227047) );
  INV_X4 U13990 ( .A(net227071), .ZN(net225824) );
  XNOR2_X2 U13991 ( .A(net225824), .B(nextPC_ex_out[12]), .ZN(net225821) );
  XNOR2_X2 U13992 ( .A(net225894), .B(nextPC_ex_out[11]), .ZN(net225889) );
  NAND2_X4 U13993 ( .A1(net239017), .A2(net227072), .ZN(net227044) );
  OAI21_X4 U13994 ( .B1(n11934), .B2(net227075), .A(net239414), .ZN(net225823)
         );
  OAI22_X2 U13995 ( .A1(n11539), .A2(net231253), .B1(net230379), .B2(n11934), 
        .ZN(n7446) );
  NAND2_X2 U13996 ( .A1(net227192), .A2(n10139), .ZN(net227217) );
  OAI221_X4 U13997 ( .B1(net227189), .B2(net227188), .C1(net239737), .C2(
        net227191), .A(net227192), .ZN(net223741) );
  NAND2_X2 U13998 ( .A1(n10361), .A2(net224816), .ZN(net224713) );
  NAND3_X2 U13999 ( .A1(net224844), .A2(net224845), .A3(net227042), .ZN(
        net227041) );
  NAND2_X4 U14000 ( .A1(net227047), .A2(net227053), .ZN(net227014) );
  NAND3_X4 U14001 ( .A1(net225076), .A2(net227047), .A3(net227046), .ZN(
        net227026) );
  NAND2_X4 U14002 ( .A1(net227047), .A2(net227046), .ZN(net227045) );
  OAI21_X4 U14003 ( .B1(net225194), .B2(net225195), .A(net225196), .ZN(
        net225172) );
  NAND2_X4 U14004 ( .A1(net223589), .A2(n11962), .ZN(net227192) );
  NAND4_X2 U14005 ( .A1(nextPC_ex_out[22]), .A2(net239722), .A3(net227207), 
        .A4(net227192), .ZN(net227230) );
  AOI21_X1 U14006 ( .B1(net223664), .B2(net239761), .A(net223665), .ZN(
        net223662) );
  XNOR2_X1 U14007 ( .A(net137303), .B(net239761), .ZN(net223586) );
  NAND3_X4 U14008 ( .A1(net227044), .A2(net227043), .A3(net225894), .ZN(
        net227024) );
  NAND3_X4 U14009 ( .A1(net227044), .A2(net227043), .A3(net227064), .ZN(
        net225076) );
  INV_X4 U14010 ( .A(net225894), .ZN(net227065) );
  OAI21_X4 U14011 ( .B1(net227145), .B2(net227144), .A(net239356), .ZN(
        net224403) );
  NAND2_X4 U14012 ( .A1(net224403), .A2(net239031), .ZN(net227121) );
  BUF_X32 U14013 ( .A(net224403), .Z(net233124) );
  NAND2_X4 U14014 ( .A1(net224403), .A2(nextPC_ex_out[20]), .ZN(net227143) );
  INV_X8 U14015 ( .A(net224174), .ZN(net227144) );
  AOI21_X4 U14016 ( .B1(n13031), .B2(n13032), .A(net227148), .ZN(net227145) );
  NAND3_X2 U14017 ( .A1(net227150), .A2(net233131), .A3(net227216), .ZN(n13031) );
  NAND2_X2 U14018 ( .A1(net227216), .A2(net227167), .ZN(net227166) );
  CLKBUF_X3 U14019 ( .A(n10108), .Z(net233131) );
  NAND2_X1 U14020 ( .A1(net233131), .A2(n10107), .ZN(net223740) );
  NAND2_X4 U14021 ( .A1(net227136), .A2(net227137), .ZN(net227142) );
  NAND2_X1 U14022 ( .A1(net224173), .A2(net224174), .ZN(net224170) );
  OAI22_X4 U14023 ( .A1(net239496), .A2(net227180), .B1(n13033), .B2(net227148), .ZN(net227136) );
  AOI21_X4 U14024 ( .B1(net227182), .B2(net227149), .A(net227183), .ZN(n13033)
         );
  NAND2_X2 U14025 ( .A1(net227150), .A2(n11927), .ZN(net227187) );
  INV_X8 U14026 ( .A(net223741), .ZN(net227165) );
  NAND2_X4 U14027 ( .A1(net227081), .A2(net225780), .ZN(net227075) );
  NAND3_X4 U14028 ( .A1(net227081), .A2(net225780), .A3(nextPC_ex_out[13]), 
        .ZN(net227070) );
  OAI21_X4 U14029 ( .B1(net227156), .B2(net227157), .A(net227158), .ZN(
        net239356) );
  INV_X4 U14030 ( .A(n10154), .ZN(net227156) );
  INV_X4 U14031 ( .A(n10154), .ZN(net239496) );
  AOI21_X4 U14032 ( .B1(net227230), .B2(net227231), .A(net224182), .ZN(
        net227229) );
  OAI21_X4 U14033 ( .B1(net227174), .B2(net227175), .A(net227176), .ZN(
        net227157) );
  NAND2_X2 U14034 ( .A1(net224816), .A2(n10356), .ZN(net225209) );
  NAND3_X4 U14035 ( .A1(net225163), .A2(net224850), .A3(n11994), .ZN(net225210) );
  NAND2_X2 U14036 ( .A1(net224850), .A2(n11994), .ZN(net224838) );
  AOI21_X2 U14038 ( .B1(net225198), .B2(net224850), .A(nextPC_ex_out[8]), .ZN(
        net225194) );
  NAND3_X4 U14039 ( .A1(net239032), .A2(n11920), .A3(net227026), .ZN(net224850) );
  NAND2_X4 U14040 ( .A1(net227142), .A2(net224404), .ZN(net224491) );
  INV_X4 U14041 ( .A(net227153), .ZN(net224404) );
  XNOR2_X2 U14042 ( .A(net224404), .B(n11927), .ZN(net224402) );
  MUX2_X2 U14043 ( .A(n11564), .B(n12561), .S(net239782), .Z(net227153) );
  NAND2_X2 U14044 ( .A1(EXEC_STAGE_imm16_32[20]), .A2(net231325), .ZN(
        net222629) );
  NAND2_X2 U14045 ( .A1(EXEC_STAGE_imm26_32[20]), .A2(net231325), .ZN(
        net222628) );
  OAI22_X4 U14046 ( .A1(net227159), .A2(net227160), .B1(net227201), .B2(n13036), .ZN(net227158) );
  INV_X4 U14047 ( .A(n13039), .ZN(n13034) );
  NAND3_X4 U14048 ( .A1(net227163), .A2(net227164), .A3(n13034), .ZN(net224182) );
  XNOR2_X2 U14049 ( .A(nextPC_ex_out[23]), .B(n13034), .ZN(net223794) );
  MUX2_X2 U14050 ( .A(n11558), .B(n12556), .S(net239782), .Z(n13039) );
  INV_X4 U14051 ( .A(n13037), .ZN(n13035) );
  NAND2_X2 U14052 ( .A1(nextPC_ex_out[23]), .A2(n13035), .ZN(net227170) );
  OAI21_X4 U14053 ( .B1(nextPC_ex_out[21]), .B2(nextPC_ex_out[22]), .A(n13035), 
        .ZN(net227167) );
  XNOR2_X2 U14054 ( .A(nextPC_ex_out[21]), .B(n13035), .ZN(net224171) );
  MUX2_X2 U14055 ( .A(n11559), .B(n12557), .S(net239782), .Z(n13037) );
  BUF_X32 U14056 ( .A(net227201), .Z(net239424) );
  NOR3_X4 U14057 ( .A1(net227201), .A2(net227202), .A3(n13038), .ZN(net227148)
         );
  INV_X1 U14059 ( .A(net227174), .ZN(net239846) );
  XNOR2_X2 U14060 ( .A(n18884), .B(n18885), .ZN(n13040) );
  INV_X8 U14062 ( .A(n18962), .ZN(n13041) );
  NAND2_X4 U14063 ( .A1(ID_EXEC_OUT[92]), .A2(n13403), .ZN(n15681) );
  XNOR2_X2 U14064 ( .A(n18858), .B(n18967), .ZN(n13043) );
  NAND3_X2 U14065 ( .A1(n13973), .A2(n13972), .A3(n19355), .ZN(n13044) );
  INV_X16 U14066 ( .A(n14099), .ZN(n18654) );
  INV_X2 U14067 ( .A(net239815), .ZN(net239816) );
  XNOR2_X1 U14068 ( .A(n18921), .B(n13493), .ZN(n13046) );
  AOI21_X1 U14069 ( .B1(n6890), .B2(n10140), .A(ID_EXEC_OUT[145]), .ZN(n6889)
         );
  NAND3_X2 U14070 ( .A1(net227277), .A2(net239329), .A3(net227276), .ZN(
        net239805) );
  NAND2_X2 U14071 ( .A1(DMEM_BUS_OUT[22]), .A2(n13484), .ZN(n15767) );
  NAND2_X1 U14072 ( .A1(DMEM_BUS_OUT[24]), .A2(n18927), .ZN(n15772) );
  NAND2_X1 U14073 ( .A1(DMEM_BUS_OUT[26]), .A2(n18927), .ZN(n15839) );
  NAND3_X2 U14074 ( .A1(n15773), .A2(n15772), .A3(n15771), .ZN(n18924) );
  BUF_X4 U14076 ( .A(n14178), .Z(n13047) );
  BUF_X8 U14077 ( .A(n14178), .Z(n13048) );
  NAND2_X2 U14078 ( .A1(n14125), .A2(n13963), .ZN(n14178) );
  NAND2_X4 U14079 ( .A1(n13980), .A2(n13981), .ZN(n13049) );
  NOR3_X2 U14081 ( .A1(n18865), .A2(n18864), .A3(n18863), .ZN(n19057) );
  XNOR2_X1 U14082 ( .A(n18921), .B(n18922), .ZN(n18978) );
  NAND2_X1 U14083 ( .A1(n17987), .A2(n18921), .ZN(n18017) );
  INV_X1 U14084 ( .A(n18921), .ZN(n18923) );
  OAI21_X2 U14085 ( .B1(n18978), .B2(n18977), .A(n18976), .ZN(n18983) );
  INV_X1 U14086 ( .A(net239035), .ZN(net239776) );
  BUF_X32 U14087 ( .A(net233133), .Z(net239774) );
  BUF_X32 U14088 ( .A(n18951), .Z(n13052) );
  XNOR2_X2 U14089 ( .A(n13053), .B(n13132), .ZN(n15494) );
  OR2_X4 U14090 ( .A1(net233242), .A2(n13062), .ZN(n15529) );
  NAND2_X4 U14091 ( .A1(n13401), .A2(n15686), .ZN(n15687) );
  INV_X1 U14092 ( .A(n15686), .ZN(n18429) );
  NAND2_X2 U14093 ( .A1(n18968), .A2(n13043), .ZN(n18956) );
  OAI21_X4 U14094 ( .B1(n18964), .B2(n18965), .A(n18963), .ZN(n18971) );
  NAND3_X2 U14096 ( .A1(n13973), .A2(n13972), .A3(n13971), .ZN(n13055) );
  NAND3_X2 U14097 ( .A1(n13972), .A2(n13973), .A3(n19355), .ZN(n13056) );
  INV_X2 U14098 ( .A(n13137), .ZN(n13057) );
  AOI21_X2 U14099 ( .B1(net224699), .B2(n17290), .A(n17289), .ZN(n17291) );
  NAND2_X1 U14100 ( .A1(ID_EXEC_OUT[201]), .A2(net231325), .ZN(n18804) );
  INV_X2 U14101 ( .A(net233181), .ZN(net227190) );
  INV_X8 U14104 ( .A(n18385), .ZN(n18967) );
  INV_X8 U14105 ( .A(n18966), .ZN(n18858) );
  OR2_X2 U14106 ( .A1(n13134), .A2(n13044), .ZN(n13983) );
  INV_X8 U14107 ( .A(n13402), .ZN(n13401) );
  NAND2_X1 U14108 ( .A1(n18861), .A2(n10130), .ZN(n13067) );
  OAI22_X1 U14109 ( .A1(n13221), .A2(n4685), .B1(net231263), .B2(n13045), .ZN(
        n7899) );
  NAND3_X4 U14110 ( .A1(n13148), .A2(n13073), .A3(n14124), .ZN(n14103) );
  NOR3_X2 U14111 ( .A1(n11116), .A2(n13878), .A3(n13073), .ZN(n13962) );
  NAND3_X2 U14112 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[31]), .A2(
        n13880), .A3(n13073), .ZN(n14073) );
  INV_X4 U14113 ( .A(n13133), .ZN(n13058) );
  BUF_X32 U14114 ( .A(n18293), .Z(n13060) );
  CLKBUF_X3 U14115 ( .A(n15785), .Z(n13101) );
  NAND2_X1 U14117 ( .A1(n15645), .A2(net224816), .ZN(n15644) );
  NAND2_X4 U14118 ( .A1(n17216), .A2(n17222), .ZN(n17213) );
  NAND2_X4 U14119 ( .A1(RegWrite_wb_out), .A2(n13045), .ZN(n13976) );
  NAND2_X4 U14120 ( .A1(n13400), .A2(n13101), .ZN(n15786) );
  NAND3_X2 U14121 ( .A1(n18918), .A2(n18916), .A3(n18917), .ZN(n13061) );
  NAND3_X2 U14122 ( .A1(n18918), .A2(n18916), .A3(n18917), .ZN(n18995) );
  NOR4_X2 U14123 ( .A1(n14116), .A2(n10126), .A3(n13877), .A4(n11472), .ZN(
        n14066) );
  NOR3_X2 U14124 ( .A1(n11557), .A2(n10126), .A3(n13877), .ZN(n13959) );
  NOR3_X2 U14125 ( .A1(n10126), .A2(n13877), .A3(n11555), .ZN(n14080) );
  NOR3_X1 U14126 ( .A1(n13878), .A2(n13153), .A3(n12071), .ZN(n13986) );
  NOR3_X2 U14127 ( .A1(n10126), .A2(n13877), .A3(n11556), .ZN(n13990) );
  NAND3_X1 U14128 ( .A1(n13486), .A2(n15671), .A3(n18929), .ZN(n15672) );
  NAND3_X2 U14129 ( .A1(n18601), .A2(n18588), .A3(n18610), .ZN(n15913) );
  AOI21_X2 U14130 ( .B1(n14064), .B2(n13219), .A(n14063), .ZN(n14069) );
  NAND3_X2 U14131 ( .A1(n13219), .A2(n13880), .A3(MEM_WB_OUT[59]), .ZN(n14015)
         );
  BUF_X16 U14132 ( .A(net227024), .Z(net239667) );
  INV_X8 U14133 ( .A(net227214), .ZN(net227232) );
  NAND2_X4 U14134 ( .A1(n18281), .A2(n17495), .ZN(n18362) );
  NAND2_X4 U14135 ( .A1(n18280), .A2(n17494), .ZN(n18281) );
  NAND2_X4 U14136 ( .A1(n17493), .A2(n17492), .ZN(n18280) );
  NAND2_X4 U14137 ( .A1(n18466), .A2(n18467), .ZN(n17493) );
  NOR2_X4 U14138 ( .A1(n17673), .A2(n15542), .ZN(n15543) );
  NAND2_X1 U14139 ( .A1(MEM_WB_OUT[64]), .A2(n13223), .ZN(n14048) );
  NOR2_X2 U14140 ( .A1(n14103), .A2(n12068), .ZN(n14045) );
  NAND2_X1 U14141 ( .A1(n15844), .A2(n13041), .ZN(n17496) );
  INV_X8 U14142 ( .A(n18861), .ZN(n18962) );
  INV_X8 U14143 ( .A(n13090), .ZN(n13092) );
  INV_X16 U14144 ( .A(n18624), .ZN(n13402) );
  NAND2_X4 U14145 ( .A1(DMEM_BUS_OUT[27]), .A2(n13485), .ZN(n15684) );
  INV_X2 U14146 ( .A(n18960), .ZN(n13066) );
  NAND2_X2 U14147 ( .A1(n12935), .A2(n19140), .ZN(n19129) );
  NAND2_X1 U14148 ( .A1(ID_EXEC_OUT[196]), .A2(net231277), .ZN(n18820) );
  INV_X1 U14149 ( .A(n17892), .ZN(n17900) );
  NAND4_X2 U14150 ( .A1(net227256), .A2(net227192), .A3(net239816), .A4(
        net239825), .ZN(n15536) );
  INV_X8 U14151 ( .A(n13063), .ZN(n13149) );
  INV_X1 U14152 ( .A(net239669), .ZN(net239621) );
  NOR2_X4 U14153 ( .A1(n18293), .A2(n13064), .ZN(n13063) );
  AND2_X2 U14154 ( .A1(DMEM_BUS_OUT[24]), .A2(n13157), .ZN(n13064) );
  OAI211_X2 U14155 ( .C1(n18902), .C2(n18901), .A(n13094), .B(n18900), .ZN(
        n18904) );
  NOR3_X4 U14156 ( .A1(n15541), .A2(net227197), .A3(net227198), .ZN(n13065) );
  NAND2_X1 U14157 ( .A1(n15776), .A2(n18980), .ZN(n15789) );
  NAND2_X2 U14158 ( .A1(n18962), .A2(n13066), .ZN(n13068) );
  NAND2_X4 U14159 ( .A1(n18610), .A2(n18588), .ZN(n17294) );
  NAND2_X4 U14160 ( .A1(net227040), .A2(net227041), .ZN(n15554) );
  NAND2_X2 U14161 ( .A1(n12998), .A2(n13492), .ZN(n18628) );
  NAND3_X2 U14162 ( .A1(ID_EXEC_OUT[86]), .A2(n13092), .A3(n13098), .ZN(n15768) );
  NAND2_X4 U14163 ( .A1(net227084), .A2(n12309), .ZN(net227094) );
  INV_X1 U14164 ( .A(n19364), .ZN(n13069) );
  INV_X4 U14165 ( .A(n13069), .ZN(n13070) );
  NAND2_X4 U14166 ( .A1(n18445), .A2(nextPC_ex_out[29]), .ZN(net223368) );
  NAND2_X2 U14167 ( .A1(n13073), .A2(n13961), .ZN(n14036) );
  NAND2_X4 U14168 ( .A1(net239767), .A2(n13078), .ZN(net227277) );
  NAND3_X4 U14169 ( .A1(n13045), .A2(n13099), .A3(MEM_WB_REG_MEM_WB_REG_N77), 
        .ZN(n15665) );
  AND2_X4 U14170 ( .A1(n15533), .A2(n10107), .ZN(net239572) );
  INV_X1 U14171 ( .A(n13148), .ZN(n13961) );
  INV_X8 U14172 ( .A(net239553), .ZN(net227242) );
  INV_X8 U14173 ( .A(n13118), .ZN(n13880) );
  OAI21_X4 U14175 ( .B1(n11980), .B2(n13879), .A(n13047), .ZN(n13072) );
  INV_X8 U14176 ( .A(n13999), .ZN(n14102) );
  NAND2_X4 U14177 ( .A1(n19063), .A2(n19062), .ZN(n13074) );
  INV_X1 U14178 ( .A(n13073), .ZN(n14078) );
  NAND2_X4 U14179 ( .A1(n13407), .A2(n17737), .ZN(n14174) );
  INV_X2 U14180 ( .A(n13408), .ZN(n13407) );
  OAI211_X2 U14181 ( .C1(n12071), .C2(n13165), .A(n13048), .B(n14172), .ZN(
        n17737) );
  AOI22_X1 U14182 ( .A1(MEM_WB_OUT[51]), .A2(n13222), .B1(MEM_WB_OUT[14]), 
        .B2(n13877), .ZN(n14172) );
  INV_X2 U14183 ( .A(n13075), .ZN(n13076) );
  XNOR2_X1 U14184 ( .A(n15792), .B(n18966), .ZN(n18395) );
  NAND2_X1 U14185 ( .A1(n18967), .A2(n18966), .ZN(n18970) );
  OAI211_X1 U14186 ( .C1(n12070), .C2(n13165), .A(n13048), .B(n14153), .ZN(
        n16578) );
  OAI211_X1 U14187 ( .C1(n12068), .C2(n13165), .A(n13048), .B(n14145), .ZN(
        n16350) );
  OAI211_X1 U14188 ( .C1(n12069), .C2(n13165), .A(n13048), .B(n14156), .ZN(
        n16539) );
  INV_X2 U14189 ( .A(n13077), .ZN(n13078) );
  NAND2_X4 U14190 ( .A1(n13073), .A2(n13880), .ZN(n13998) );
  INV_X1 U14191 ( .A(n13140), .ZN(n13079) );
  NAND3_X4 U14192 ( .A1(n15849), .A2(n17893), .A3(n15848), .ZN(n17722) );
  NAND2_X2 U14193 ( .A1(n15780), .A2(n15779), .ZN(n15781) );
  NAND2_X4 U14194 ( .A1(n15548), .A2(n15547), .ZN(n15549) );
  OAI21_X4 U14195 ( .B1(n19036), .B2(n19037), .A(n19035), .ZN(n19043) );
  AOI22_X1 U14196 ( .A1(n13490), .A2(n13060), .B1(n10829), .B2(
        DMEM_BUS_OUT[24]), .ZN(n18294) );
  INV_X2 U14197 ( .A(n18968), .ZN(n18969) );
  INV_X4 U14198 ( .A(net223797), .ZN(net227174) );
  NAND2_X2 U14199 ( .A1(n16970), .A2(net225172), .ZN(n13081) );
  NAND2_X4 U14200 ( .A1(n13082), .A2(n13081), .ZN(n16973) );
  NAND2_X4 U14201 ( .A1(n19027), .A2(n12253), .ZN(n19034) );
  NOR2_X4 U14203 ( .A1(n15502), .A2(n19361), .ZN(n15663) );
  NAND2_X1 U14205 ( .A1(n13131), .A2(n13059), .ZN(n13087) );
  INV_X4 U14206 ( .A(n13131), .ZN(n13085) );
  INV_X2 U14207 ( .A(n13059), .ZN(n13086) );
  NAND2_X1 U14208 ( .A1(n19024), .A2(n19023), .ZN(n19026) );
  NAND2_X4 U14210 ( .A1(n10113), .A2(n15566), .ZN(net225198) );
  NAND2_X4 U14211 ( .A1(n13049), .A2(n14099), .ZN(n13997) );
  NAND3_X2 U14212 ( .A1(ID_EXEC_OUT[57]), .A2(n13049), .A3(n13044), .ZN(n14043) );
  NAND3_X4 U14213 ( .A1(n15500), .A2(n15499), .A3(RegWrite_wb_out), .ZN(n15501) );
  NOR2_X2 U14214 ( .A1(n13116), .A2(n17204), .ZN(n17225) );
  INV_X8 U14216 ( .A(n15677), .ZN(n18625) );
  INV_X4 U14217 ( .A(n17219), .ZN(n17218) );
  XNOR2_X2 U14218 ( .A(n13086), .B(n13138), .ZN(n13979) );
  NOR3_X2 U14219 ( .A1(n19060), .A2(ID_EXEC_OUT[156]), .A3(ID_EXEC_OUT[158]), 
        .ZN(n19133) );
  OAI221_X4 U14220 ( .B1(n13098), .B2(n11938), .C1(n16753), .C2(n15811), .A(
        n15810), .ZN(n16823) );
  NAND3_X2 U14221 ( .A1(n13092), .A2(n13098), .A3(ID_EXEC_OUT[80]), .ZN(n15810) );
  INV_X1 U14222 ( .A(net239424), .ZN(net239415) );
  INV_X2 U14223 ( .A(n19092), .ZN(n13089) );
  INV_X16 U14224 ( .A(n13090), .ZN(n13091) );
  AOI21_X4 U14225 ( .B1(n18988), .B2(n18989), .A(n18987), .ZN(n18998) );
  INV_X1 U14226 ( .A(nextPC_ex_out[25]), .ZN(net223591) );
  NAND3_X4 U14227 ( .A1(n15788), .A2(n15787), .A3(n15786), .ZN(n18385) );
  INV_X8 U14228 ( .A(n15538), .ZN(n13111) );
  NAND2_X1 U14229 ( .A1(ID_EXEC_OUT[89]), .A2(n18625), .ZN(n15788) );
  NOR3_X4 U14230 ( .A1(n19148), .A2(n19147), .A3(n19146), .ZN(n19151) );
  OAI21_X2 U14231 ( .B1(n17222), .B2(n17223), .A(n17221), .ZN(n17224) );
  INV_X1 U14232 ( .A(n10143), .ZN(n18446) );
  INV_X1 U14233 ( .A(net227188), .ZN(net239374) );
  INV_X4 U14234 ( .A(n13145), .ZN(n13131) );
  INV_X2 U14235 ( .A(net239370), .ZN(net239371) );
  NAND3_X2 U14236 ( .A1(net239082), .A2(net239356), .A3(net224493), .ZN(n15548) );
  NAND3_X2 U14237 ( .A1(n18893), .A2(n18891), .A3(n18892), .ZN(n13094) );
  NAND3_X4 U14238 ( .A1(n14148), .A2(n14149), .A3(n14150), .ZN(n17868) );
  NAND2_X2 U14239 ( .A1(n13222), .A2(MEM_WB_OUT[52]), .ZN(n14149) );
  OAI21_X4 U14240 ( .B1(n18984), .B2(n18983), .A(n18982), .ZN(n18988) );
  INV_X16 U14241 ( .A(n13149), .ZN(n18925) );
  INV_X1 U14242 ( .A(n10142), .ZN(net239344) );
  OAI211_X1 U14243 ( .C1(n13165), .C2(n19298), .A(n13048), .B(n14132), .ZN(
        n16872) );
  OAI211_X1 U14244 ( .C1(n13165), .C2(n12067), .A(n13048), .B(n14139), .ZN(
        n17045) );
  OAI211_X1 U14245 ( .C1(n13165), .C2(n12220), .A(n13048), .B(n14136), .ZN(
        n16295) );
  NAND3_X2 U14246 ( .A1(n18887), .A2(n18891), .A3(n18893), .ZN(n18894) );
  INV_X1 U14248 ( .A(n10156), .ZN(net224180) );
  NOR2_X1 U14249 ( .A1(nextPC_ex_out[26]), .A2(n18107), .ZN(net223665) );
  NAND2_X1 U14250 ( .A1(nextPC_ex_out[26]), .A2(n18107), .ZN(net223664) );
  NAND3_X2 U14251 ( .A1(n15840), .A2(n15839), .A3(n15838), .ZN(n18958) );
  NAND3_X2 U14252 ( .A1(ID_EXEC_OUT[58]), .A2(n13049), .A3(n13055), .ZN(n13982) );
  INV_X1 U14253 ( .A(n19070), .ZN(n13095) );
  NAND2_X4 U14254 ( .A1(n15670), .A2(n15669), .ZN(n13098) );
  BUF_X32 U14255 ( .A(n17978), .Z(n13100) );
  INV_X16 U14256 ( .A(n18927), .ZN(n13486) );
  INV_X8 U14257 ( .A(n13486), .ZN(n13485) );
  NAND2_X2 U14258 ( .A1(n13046), .A2(n18922), .ZN(n17835) );
  INV_X2 U14259 ( .A(EXEC_STAGE_imm26_32[25]), .ZN(net137569) );
  NOR2_X2 U14260 ( .A1(n15654), .A2(n15653), .ZN(n15655) );
  AOI211_X1 U14261 ( .C1(n17858), .C2(n18979), .A(n17857), .B(n17856), .ZN(
        n17864) );
  INV_X1 U14262 ( .A(n18979), .ZN(n18981) );
  XNOR2_X1 U14263 ( .A(n18979), .B(n18980), .ZN(n18976) );
  INV_X4 U14264 ( .A(n18630), .ZN(n13102) );
  XNOR2_X2 U14265 ( .A(n13105), .B(n13123), .ZN(n13975) );
  NAND2_X1 U14267 ( .A1(net223796), .A2(net239846), .ZN(n17974) );
  XNOR2_X2 U14268 ( .A(n13160), .B(n18943), .ZN(n18949) );
  INV_X16 U14269 ( .A(n13160), .ZN(n13161) );
  INV_X16 U14271 ( .A(n18862), .ZN(n18943) );
  INV_X4 U14272 ( .A(n13128), .ZN(n13103) );
  XNOR2_X2 U14273 ( .A(n13158), .B(n18641), .ZN(n13104) );
  INV_X4 U14274 ( .A(n13104), .ZN(n18938) );
  XNOR2_X1 U14275 ( .A(net223662), .B(net239621), .ZN(n18065) );
  INV_X2 U14276 ( .A(n13121), .ZN(n13115) );
  NOR2_X1 U14277 ( .A1(net227242), .A2(net227243), .ZN(net227239) );
  INV_X16 U14278 ( .A(n14123), .ZN(n18664) );
  XOR2_X2 U14279 ( .A(n13079), .B(n13136), .Z(n13978) );
  NAND3_X2 U14280 ( .A1(n15770), .A2(n13056), .A3(n14098), .ZN(n14100) );
  INV_X16 U14281 ( .A(n13225), .ZN(n13223) );
  INV_X16 U14282 ( .A(n13225), .ZN(n13222) );
  INV_X4 U14283 ( .A(n13225), .ZN(n13224) );
  NAND2_X4 U14284 ( .A1(n13400), .A2(n17868), .ZN(n15816) );
  INV_X1 U14285 ( .A(ID_EXEC_OUT[193]), .ZN(n18829) );
  NOR2_X4 U14286 ( .A1(n14122), .A2(n13108), .ZN(n13106) );
  INV_X4 U14287 ( .A(n13106), .ZN(n14117) );
  INV_X1 U14288 ( .A(n19091), .ZN(n19092) );
  NAND2_X1 U14289 ( .A1(n18883), .A2(n19091), .ZN(n18900) );
  NOR3_X4 U14290 ( .A1(n13979), .A2(n13978), .A3(n13977), .ZN(n13980) );
  INV_X4 U14291 ( .A(net239776), .ZN(net239221) );
  NAND2_X4 U14292 ( .A1(n15543), .A2(n13093), .ZN(net227149) );
  NAND3_X2 U14293 ( .A1(n14067), .A2(n14068), .A3(n14069), .ZN(n17981) );
  NAND3_X1 U14294 ( .A1(n13208), .A2(n18641), .A3(n13159), .ZN(n18556) );
  INV_X1 U14295 ( .A(MEM_WB_REG_MEM_WB_REG_N147), .ZN(n19312) );
  AOI211_X1 U14296 ( .C1(n18642), .C2(n18641), .A(n18640), .B(n18639), .ZN(
        n18647) );
  OAI221_X1 U14297 ( .B1(n14011), .B2(n17685), .C1(n17537), .C2(n18641), .A(
        n17536), .ZN(n17907) );
  OAI211_X1 U14298 ( .C1(n15709), .C2(n18641), .A(n15708), .B(n15707), .ZN(
        n16876) );
  XNOR2_X1 U14299 ( .A(n15827), .B(n18641), .ZN(n18547) );
  XNOR2_X1 U14300 ( .A(n18641), .B(n13494), .ZN(n15830) );
  AOI21_X1 U14301 ( .B1(net231289), .B2(EXEC_STAGE_imm26_32[29]), .A(n19163), 
        .ZN(n5606) );
  AOI21_X1 U14302 ( .B1(net239805), .B2(n18447), .A(n10155), .ZN(n18239) );
  INV_X16 U14303 ( .A(n13402), .ZN(n13400) );
  INV_X16 U14304 ( .A(n13402), .ZN(n13399) );
  INV_X8 U14305 ( .A(n15550), .ZN(n15551) );
  NAND2_X4 U14306 ( .A1(n15549), .A2(n11917), .ZN(n15550) );
  NAND2_X2 U14307 ( .A1(n18885), .A2(n18884), .ZN(n18889) );
  AOI22_X1 U14308 ( .A1(net231301), .A2(EXEC_STAGE_imm26_32[31]), .B1(
        ID_STAGE_imm16_aluA[31]), .B2(net230393), .ZN(n5603) );
  NAND2_X4 U14309 ( .A1(n18664), .A2(n19347), .ZN(n14111) );
  NOR2_X4 U14310 ( .A1(n18961), .A2(n13110), .ZN(n18964) );
  INV_X8 U14312 ( .A(n14176), .ZN(n13225) );
  NAND3_X2 U14313 ( .A1(n14040), .A2(n14041), .A3(n14042), .ZN(n15785) );
  AND3_X4 U14314 ( .A1(n13142), .A2(n13143), .A3(n13144), .ZN(n13971) );
  NAND2_X4 U14315 ( .A1(n14037), .A2(n14124), .ZN(n14092) );
  INV_X4 U14316 ( .A(n14036), .ZN(n14037) );
  NOR2_X2 U14317 ( .A1(n16711), .A2(n13361), .ZN(n16712) );
  NOR2_X1 U14318 ( .A1(n16711), .A2(n13453), .ZN(n16684) );
  NOR2_X2 U14319 ( .A1(n14103), .A2(n12070), .ZN(n14054) );
  OAI22_X1 U14320 ( .A1(n12308), .A2(net231257), .B1(net230381), .B2(net223591), .ZN(n7665) );
  XOR2_X2 U14321 ( .A(n13112), .B(n13135), .Z(n13970) );
  NAND2_X4 U14322 ( .A1(ID_EXEC_OUT[148]), .A2(n15666), .ZN(n15667) );
  XNOR2_X2 U14324 ( .A(ID_EXEC_OUT[198]), .B(n13115), .ZN(n15495) );
  INV_X8 U14325 ( .A(n17216), .ZN(n17204) );
  INV_X4 U14326 ( .A(n13117), .ZN(n13118) );
  NOR2_X2 U14327 ( .A1(n14103), .A2(n12069), .ZN(n14085) );
  BUF_X32 U14328 ( .A(n18261), .Z(n13119) );
  NAND2_X2 U14329 ( .A1(n15651), .A2(n17216), .ZN(n17219) );
  OAI21_X2 U14330 ( .B1(n17222), .B2(n15652), .A(n15650), .ZN(n15653) );
  NAND2_X1 U14331 ( .A1(EXEC_STAGE_imm16_32[28]), .A2(net231311), .ZN(n18836)
         );
  XOR2_X1 U14332 ( .A(n13130), .B(n13120), .Z(n13974) );
  AOI21_X4 U14333 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[16]), .B2(
        n14105), .A(n14104), .ZN(n14106) );
  XOR2_X1 U14334 ( .A(net239528), .B(net137317), .Z(n18238) );
  INV_X1 U14335 ( .A(net239220), .ZN(net239150) );
  INV_X8 U14336 ( .A(n18944), .ZN(n13162) );
  NOR2_X2 U14337 ( .A1(n14036), .A2(n19298), .ZN(n13964) );
  INV_X2 U14338 ( .A(net227163), .ZN(net227202) );
  AOI22_X1 U14339 ( .A1(n10829), .A2(DMEM_BUS_OUT[25]), .B1(n13490), .B2(
        n13126), .ZN(n18386) );
  NAND2_X1 U14340 ( .A1(n15792), .A2(n18966), .ZN(n17705) );
  NAND2_X1 U14341 ( .A1(n16061), .A2(n17754), .ZN(n17755) );
  NAND2_X1 U14342 ( .A1(n13390), .A2(n17754), .ZN(n16819) );
  NAND2_X1 U14343 ( .A1(n13487), .A2(n17754), .ZN(n16548) );
  NAND2_X1 U14344 ( .A1(n13393), .A2(n17754), .ZN(n16293) );
  NAND2_X1 U14345 ( .A1(n13392), .A2(n16884), .ZN(n16889) );
  NAND2_X1 U14346 ( .A1(n13389), .A2(n16884), .ZN(n16203) );
  NAND2_X1 U14347 ( .A1(n13396), .A2(n16884), .ZN(n16047) );
  INV_X1 U14349 ( .A(n16753), .ZN(n13125) );
  BUF_X32 U14350 ( .A(n18384), .Z(n13126) );
  AOI21_X1 U14351 ( .B1(net231289), .B2(EXEC_STAGE_imm16_32[29]), .A(n19163), 
        .ZN(n5588) );
  XNOR2_X2 U14352 ( .A(n13128), .B(n13058), .ZN(n13977) );
  NAND2_X4 U14353 ( .A1(net227245), .A2(net227246), .ZN(n15532) );
  INV_X1 U14354 ( .A(n17981), .ZN(n17957) );
  INV_X1 U14355 ( .A(n17868), .ZN(n16711) );
  XOR2_X2 U14356 ( .A(n13132), .B(n13133), .Z(n13968) );
  NAND2_X1 U14357 ( .A1(n17982), .A2(n17868), .ZN(n17869) );
  XNOR2_X1 U14358 ( .A(n18862), .B(n13494), .ZN(n15834) );
  NAND2_X1 U14359 ( .A1(n18641), .A2(n18862), .ZN(n18532) );
  NAND3_X2 U14360 ( .A1(n13996), .A2(n13995), .A3(n13994), .ZN(n18939) );
  NAND2_X4 U14361 ( .A1(n13401), .A2(n15682), .ZN(n15683) );
  INV_X2 U14362 ( .A(n13135), .ZN(n13136) );
  AOI22_X1 U14363 ( .A1(n17983), .A2(ID_EXEC_OUT[48]), .B1(n17982), .B2(n13125), .ZN(n16812) );
  XOR2_X2 U14364 ( .A(n13137), .B(n13138), .Z(n13969) );
  NOR2_X1 U14365 ( .A1(n13050), .A2(n13491), .ZN(n17147) );
  NAND2_X1 U14366 ( .A1(net231615), .A2(n18966), .ZN(n18064) );
  NAND2_X1 U14367 ( .A1(n18310), .A2(n18966), .ZN(n17921) );
  NAND2_X1 U14368 ( .A1(n13385), .A2(n18966), .ZN(n18275) );
  NOR2_X1 U14369 ( .A1(n14092), .A2(n12060), .ZN(n14086) );
  NOR2_X1 U14370 ( .A1(n14092), .A2(n19297), .ZN(n14046) );
  NOR2_X2 U14371 ( .A1(n14092), .A2(n14122), .ZN(n14094) );
  NOR2_X2 U14372 ( .A1(n14092), .A2(n19295), .ZN(n14053) );
  NAND4_X1 U14373 ( .A1(n13880), .A2(n13073), .A3(
        WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[26]), .A4(n13985), .ZN(n13966)
         );
  NAND2_X4 U14374 ( .A1(n13106), .A2(n13147), .ZN(n14000) );
  INV_X1 U14375 ( .A(n17673), .ZN(n17674) );
  OAI21_X4 U14376 ( .B1(n16973), .B2(net231915), .A(n16972), .ZN(n7504) );
  NAND2_X1 U14377 ( .A1(n12977), .A2(n10136), .ZN(n17433) );
  AOI22_X1 U14378 ( .A1(MEM_WB_OUT[19]), .A2(n13878), .B1(MEM_WB_OUT[88]), 
        .B2(n14102), .ZN(n14033) );
  AOI22_X1 U14379 ( .A1(MEM_WB_OUT[20]), .A2(n13878), .B1(MEM_WB_OUT[89]), 
        .B2(n14102), .ZN(n14003) );
  AOI22_X1 U14380 ( .A1(MEM_WB_OUT[18]), .A2(n13877), .B1(MEM_WB_OUT[87]), 
        .B2(n14102), .ZN(n14028) );
  AOI22_X1 U14381 ( .A1(MEM_WB_OUT[21]), .A2(n13878), .B1(MEM_WB_OUT[90]), 
        .B2(n14102), .ZN(n14008) );
  INV_X2 U14383 ( .A(n13154), .ZN(n13960) );
  NAND2_X4 U14384 ( .A1(n13154), .A2(n13148), .ZN(n14116) );
  NAND2_X4 U14386 ( .A1(net227213), .A2(n15537), .ZN(n15538) );
  INV_X8 U14387 ( .A(n15532), .ZN(n15537) );
  NAND2_X4 U14389 ( .A1(net239631), .A2(net233181), .ZN(n15541) );
  NAND2_X4 U14390 ( .A1(n15790), .A2(n15789), .ZN(n15777) );
  AOI22_X4 U14391 ( .A1(MEM_WB_OUT[24]), .A2(n13877), .B1(MEM_WB_OUT[93]), 
        .B2(n14102), .ZN(n14097) );
  INV_X1 U14392 ( .A(n18883), .ZN(n13141) );
  INV_X1 U14393 ( .A(n10129), .ZN(n18883) );
  AOI22_X4 U14394 ( .A1(MEM_WB_OUT[25]), .A2(n13877), .B1(MEM_WB_OUT[94]), 
        .B2(n14102), .ZN(n14042) );
  NAND3_X4 U14395 ( .A1(n18929), .A2(n17840), .A3(n13098), .ZN(n15766) );
  NAND2_X1 U14396 ( .A1(n13409), .A2(n13041), .ZN(n18358) );
  NAND2_X1 U14397 ( .A1(n18346), .A2(n13041), .ZN(n18335) );
  OAI21_X1 U14398 ( .B1(n13491), .B2(n18372), .A(n18371), .ZN(n18374) );
  AOI22_X1 U14399 ( .A1(n10843), .A2(n18966), .B1(n18347), .B2(n13041), .ZN(
        n17854) );
  NAND2_X1 U14400 ( .A1(n13052), .A2(n18953), .ZN(n18864) );
  NOR4_X1 U14401 ( .A1(n18966), .A2(n13041), .A3(n13161), .A4(n18922), .ZN(
        n14113) );
  NAND2_X1 U14402 ( .A1(net232816), .A2(n13041), .ZN(n16013) );
  NAND2_X1 U14403 ( .A1(net223324), .A2(n13041), .ZN(n15737) );
  NAND2_X1 U14404 ( .A1(n13358), .A2(n13041), .ZN(n16543) );
  NAND2_X1 U14405 ( .A1(n13386), .A2(n13041), .ZN(n18270) );
  NAND2_X1 U14406 ( .A1(n13409), .A2(n13089), .ZN(n17867) );
  NAND2_X1 U14407 ( .A1(net231615), .A2(n13089), .ZN(n16723) );
  NOR4_X1 U14408 ( .A1(n13089), .A2(net222497), .A3(n19000), .A4(n19029), .ZN(
        n14184) );
  NAND2_X1 U14409 ( .A1(n13358), .A2(n13089), .ZN(n17992) );
  NAND2_X1 U14410 ( .A1(n13386), .A2(n13089), .ZN(n16772) );
  NAND2_X1 U14411 ( .A1(n15819), .A2(n19091), .ZN(n17732) );
  OAI211_X1 U14412 ( .C1(n19296), .C2(n13165), .A(n13048), .B(n14142), .ZN(
        n17242) );
  XNOR2_X1 U14413 ( .A(n15819), .B(n19091), .ZN(n17733) );
  OAI211_X1 U14414 ( .C1(n12031), .C2(n13165), .A(n13048), .B(n14126), .ZN(
        n16147) );
  OAI211_X1 U14415 ( .C1(n19295), .C2(n13165), .A(n13048), .B(n14168), .ZN(
        n16031) );
  OAI211_X1 U14416 ( .C1(n12032), .C2(n13165), .A(n13048), .B(n14164), .ZN(
        n16070) );
  OAI211_X1 U14417 ( .C1(n19297), .C2(n13165), .A(n13048), .B(n14129), .ZN(
        n16918) );
  OAI211_X1 U14418 ( .C1(n13165), .C2(n12066), .A(n13048), .B(n14160), .ZN(
        n16222) );
  NAND2_X1 U14419 ( .A1(n18930), .A2(n18929), .ZN(n18933) );
  NAND3_X2 U14420 ( .A1(n15770), .A2(n13098), .A3(n18929), .ZN(n15771) );
  NAND3_X1 U14421 ( .A1(n18929), .A2(n15837), .A3(n13098), .ZN(n15838) );
  INV_X8 U14422 ( .A(n15501), .ZN(n15662) );
  INV_X8 U14423 ( .A(n19046), .ZN(n19053) );
  NAND2_X4 U14425 ( .A1(n15775), .A2(n15774), .ZN(n15790) );
  INV_X8 U14426 ( .A(n15497), .ZN(n15669) );
  NOR3_X4 U14427 ( .A1(n18973), .A2(n18974), .A3(n18972), .ZN(n18984) );
  NAND3_X2 U14428 ( .A1(n15837), .A2(n13055), .A3(n14098), .ZN(n13984) );
  NOR2_X4 U14429 ( .A1(net227058), .A2(n12205), .ZN(n17196) );
  INV_X4 U14430 ( .A(net239030), .ZN(net239031) );
  NAND3_X2 U14431 ( .A1(net227024), .A2(net225908), .A3(nextPC_ex_out[10]), 
        .ZN(net239032) );
  NAND2_X4 U14432 ( .A1(n14098), .A2(n13056), .ZN(n14123) );
  NOR4_X4 U14433 ( .A1(n18957), .A2(n18956), .A3(n18955), .A4(n18954), .ZN(
        n18973) );
  NAND2_X2 U14434 ( .A1(n12954), .A2(n19129), .ZN(n19131) );
  NAND3_X1 U14435 ( .A1(n19088), .A2(n13493), .A3(n13151), .ZN(n19130) );
  NOR2_X1 U14436 ( .A1(n11915), .A2(n19134), .ZN(n19128) );
  NAND2_X4 U14437 ( .A1(n15779), .A2(n15769), .ZN(n17709) );
  OAI21_X1 U14438 ( .B1(n10128), .B2(n16797), .A(n17120), .ZN(n17754) );
  OAI211_X1 U14439 ( .C1(n10128), .C2(net232817), .A(n18274), .B(n16301), .ZN(
        n16884) );
  INV_X4 U14440 ( .A(MEM_WB_OUT[103]), .ZN(n13146) );
  INV_X8 U14441 ( .A(n13146), .ZN(n13147) );
  NAND2_X4 U14442 ( .A1(n18929), .A2(n15836), .ZN(n15811) );
  INV_X1 U14444 ( .A(n17591), .ZN(n17592) );
  NAND2_X4 U14445 ( .A1(n17591), .A2(n17593), .ZN(n16395) );
  INV_X1 U14446 ( .A(EXEC_STAGE_imm26_32[30]), .ZN(net137549) );
  INV_X16 U14447 ( .A(n14099), .ZN(n13157) );
  NAND2_X1 U14448 ( .A1(destReg_wb_out[0]), .A2(n19313), .ZN(n15350) );
  INV_X1 U14449 ( .A(destReg_wb_out[0]), .ZN(n19311) );
  XOR2_X1 U14450 ( .A(offset_26_id[5]), .B(destReg_wb_out[0]), .Z(n5467) );
  XOR2_X1 U14451 ( .A(offset_26_id[0]), .B(destReg_wb_out[0]), .Z(n2539) );
  NAND2_X4 U14452 ( .A1(n15493), .A2(n15492), .ZN(n15668) );
  XNOR2_X2 U14453 ( .A(ID_EXEC_OUT[200]), .B(n19348), .ZN(n15493) );
  XNOR2_X1 U14454 ( .A(n13051), .B(n13493), .ZN(n15858) );
  INV_X1 U14455 ( .A(EXEC_STAGE_imm16_32[30]), .ZN(net137550) );
  INV_X8 U14456 ( .A(n15811), .ZN(n18624) );
  INV_X1 U14458 ( .A(ID_EXEC_OUT[192]), .ZN(n15664) );
  NAND2_X1 U14459 ( .A1(n15663), .A2(n15662), .ZN(n15508) );
  NAND2_X4 U14460 ( .A1(DMEM_BUS_OUT[16]), .A2(n13157), .ZN(n14109) );
  AOI22_X1 U14461 ( .A1(net231311), .A2(ID_EXEC_OUT[200]), .B1(n13220), .B2(
        net230393), .ZN(n4674) );
  NAND2_X1 U14462 ( .A1(n18752), .A2(n18751), .ZN(n7837) );
  INV_X1 U14463 ( .A(MEM_WB_REG_MEM_WB_REG_N76), .ZN(n18779) );
  OAI221_X1 U14465 ( .B1(n10128), .B2(n18586), .C1(n12299), .C2(net231237), 
        .A(n6753), .ZN(n7714) );
  NOR2_X1 U14466 ( .A1(n10128), .A2(net222304), .ZN(n15735) );
  INV_X16 U14467 ( .A(n15712), .ZN(n13357) );
  INV_X1 U14468 ( .A(n18884), .ZN(n18630) );
  INV_X1 U14469 ( .A(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[16]), .ZN(n19299)
         );
  INV_X4 U14470 ( .A(n13103), .ZN(n19317) );
  NAND2_X4 U14471 ( .A1(ID_EXEC_OUT[47]), .A2(n15712), .ZN(n17871) );
  INV_X8 U14472 ( .A(n12602), .ZN(n13155) );
  INV_X1 U14473 ( .A(n13408), .ZN(n13405) );
  INV_X16 U14474 ( .A(n13408), .ZN(n13406) );
  NAND2_X4 U14475 ( .A1(ID_EXEC_OUT[48]), .A2(n15712), .ZN(n14110) );
  NOR2_X2 U14476 ( .A1(net227190), .A2(net227214), .ZN(n15539) );
  NAND2_X4 U14477 ( .A1(n19063), .A2(n19062), .ZN(n19074) );
  AOI211_X4 U14478 ( .C1(n13218), .C2(n19137), .A(n19144), .B(n19136), .ZN(
        n19147) );
  NAND2_X4 U14479 ( .A1(n13040), .A2(n18889), .ZN(n18893) );
  NAND2_X4 U14480 ( .A1(n17978), .A2(n17835), .ZN(n15779) );
  NAND4_X1 U14481 ( .A1(n13093), .A2(n17674), .A3(net223796), .A4(
        nextPC_ex_out[23]), .ZN(n17827) );
  NAND2_X1 U14482 ( .A1(n10151), .A2(net239374), .ZN(n18107) );
  OAI221_X4 U14483 ( .B1(n19083), .B2(n19082), .C1(n19081), .C2(n19080), .A(
        n19079), .ZN(n19084) );
  INV_X8 U14484 ( .A(n12997), .ZN(n13156) );
  NOR2_X1 U14485 ( .A1(n19317), .A2(destReg_wb_out[4]), .ZN(n200) );
  MUX2_X2 U14486 ( .A(n15531), .B(n15530), .S(net239627), .Z(net233133) );
  NOR2_X2 U14487 ( .A1(n13218), .A2(n19140), .ZN(n19060) );
  NAND2_X4 U14488 ( .A1(n13148), .A2(n13960), .ZN(n14074) );
  INV_X1 U14489 ( .A(MEM_WB_REG_MEM_WB_REG_N146), .ZN(n19314) );
  NAND2_X4 U14490 ( .A1(n17196), .A2(net224853), .ZN(n17197) );
  NOR2_X1 U14491 ( .A1(n10133), .A2(n13491), .ZN(n18337) );
  NAND3_X2 U14492 ( .A1(n15566), .A2(n13026), .A3(n11016), .ZN(net224853) );
  NAND2_X4 U14493 ( .A1(n14119), .A2(n14079), .ZN(n13999) );
  INV_X1 U14494 ( .A(n13101), .ZN(n18090) );
  NAND2_X4 U14495 ( .A1(n17892), .A2(n17897), .ZN(n17721) );
  NAND3_X2 U14496 ( .A1(net227024), .A2(net225908), .A3(nextPC_ex_out[10]), 
        .ZN(net224845) );
  NOR2_X1 U14497 ( .A1(n18938), .A2(n13491), .ZN(n18530) );
  NAND2_X1 U14498 ( .A1(n18938), .A2(n18949), .ZN(n18863) );
  INV_X1 U14499 ( .A(n10351), .ZN(n19313) );
  NAND3_X2 U14500 ( .A1(n15655), .A2(n15657), .A3(n15656), .ZN(n7333) );
  INV_X4 U14501 ( .A(n17199), .ZN(n17209) );
  NAND3_X2 U14502 ( .A1(n17291), .A2(n17292), .A3(n17293), .ZN(n7555) );
  INV_X1 U14503 ( .A(n13119), .ZN(n18262) );
  AOI22_X4 U14504 ( .A1(n18664), .A2(n15678), .B1(ID_EXEC_OUT[60]), .B2(n15712), .ZN(n18261) );
  NAND2_X1 U14505 ( .A1(ID_EXEC_OUT[195]), .A2(net231317), .ZN(n18824) );
  NAND2_X1 U14506 ( .A1(net231615), .A2(n13102), .ZN(n16770) );
  NAND2_X1 U14507 ( .A1(n13410), .A2(n13102), .ZN(n16556) );
  NOR4_X1 U14508 ( .A1(n13151), .A2(n13163), .A3(n13149), .A4(n13102), .ZN(
        n14112) );
  NAND2_X1 U14509 ( .A1(n13386), .A2(n13102), .ZN(n16790) );
  NAND2_X1 U14510 ( .A1(n16816), .A2(n13102), .ZN(n18245) );
  NAND2_X1 U14511 ( .A1(n15858), .A2(n18884), .ZN(n17728) );
  XNOR2_X1 U14512 ( .A(n15858), .B(n18884), .ZN(n16787) );
  AOI22_X4 U14513 ( .A1(n18664), .A2(n15682), .B1(ID_EXEC_OUT[59]), .B2(n15712), .ZN(n18372) );
  INV_X8 U14514 ( .A(n14116), .ZN(n14079) );
  OAI21_X1 U14515 ( .B1(n13154), .B2(n14117), .A(n14116), .ZN(n14118) );
  NAND3_X2 U14516 ( .A1(n17209), .A2(n17208), .A3(n17210), .ZN(n7542) );
  NOR2_X4 U14517 ( .A1(n17204), .A2(n17203), .ZN(n17205) );
  NOR2_X2 U14518 ( .A1(n15648), .A2(n15647), .ZN(n15654) );
  INV_X2 U14519 ( .A(n15648), .ZN(n15565) );
  NAND2_X4 U14520 ( .A1(n17218), .A2(n17217), .ZN(n17227) );
  NAND2_X1 U14521 ( .A1(net224180), .A2(net239415), .ZN(n17828) );
  NAND2_X4 U14522 ( .A1(net227015), .A2(net225077), .ZN(n15562) );
  INV_X1 U14523 ( .A(n13152), .ZN(n19315) );
  NAND3_X2 U14524 ( .A1(n18905), .A2(n18895), .A3(n18903), .ZN(n18906) );
  NAND3_X1 U14525 ( .A1(ID_EXEC_OUT[62]), .A2(n13049), .A3(n13056), .ZN(n13994) );
  NAND3_X1 U14526 ( .A1(ID_EXEC_OUT[56]), .A2(n13049), .A3(n13055), .ZN(n14101) );
  NAND2_X4 U14527 ( .A1(net225823), .A2(nextPC_ex_out[12]), .ZN(net227073) );
  NAND4_X1 U14528 ( .A1(n18963), .A2(n10133), .A3(n18968), .A4(n18978), .ZN(
        n18865) );
  OAI21_X2 U14529 ( .B1(net137550), .B2(net231247), .A(n18832), .ZN(n7974) );
  NAND2_X4 U14530 ( .A1(n14044), .A2(n14043), .ZN(n18384) );
  INV_X1 U14531 ( .A(n19140), .ZN(n19137) );
  NOR2_X1 U14532 ( .A1(n18886), .A2(n13491), .ZN(n16824) );
  AOI21_X2 U14533 ( .B1(n18916), .B2(n18910), .A(n18993), .ZN(n18920) );
  NAND3_X2 U14534 ( .A1(n18894), .A2(n18900), .A3(n18899), .ZN(n18905) );
  NAND3_X2 U14535 ( .A1(n15579), .A2(n15581), .A3(n15580), .ZN(n7325) );
  NAND2_X4 U14536 ( .A1(n16142), .A2(n15911), .ZN(n18588) );
  NAND2_X4 U14537 ( .A1(n15791), .A2(n15793), .ZN(n17502) );
  NAND2_X4 U14538 ( .A1(n17708), .A2(n15781), .ZN(n15791) );
  NAND2_X1 U14539 ( .A1(destReg_wb_out[0]), .A2(n10351), .ZN(n15352) );
  NAND2_X1 U14540 ( .A1(n19311), .A2(n10351), .ZN(n15348) );
  AOI21_X1 U14541 ( .B1(n13092), .B2(n12275), .A(n18927), .ZN(n18934) );
  NAND3_X1 U14542 ( .A1(ID_EXEC_OUT[95]), .A2(n13092), .A3(n13486), .ZN(n15673) );
  NAND3_X1 U14543 ( .A1(ID_EXEC_OUT[90]), .A2(n13092), .A3(n13098), .ZN(n15840) );
  NAND3_X1 U14544 ( .A1(ID_EXEC_OUT[88]), .A2(n13098), .A3(n13092), .ZN(n15773) );
  INV_X16 U14545 ( .A(n13091), .ZN(n18929) );
  NAND2_X4 U14546 ( .A1(net227068), .A2(net227067), .ZN(net227043) );
  NAND2_X4 U14547 ( .A1(n10113), .A2(n15566), .ZN(net225163) );
  NAND2_X4 U14548 ( .A1(net227002), .A2(n10112), .ZN(net225214) );
  OAI211_X1 U14549 ( .C1(nextPC_ex_out[31]), .C2(n18747), .A(net239823), .B(
        n10361), .ZN(n18749) );
  OAI211_X4 U14550 ( .C1(n19145), .C2(n19144), .A(n19143), .B(n19142), .ZN(
        n19146) );
  NOR2_X1 U14551 ( .A1(n13070), .A2(n13491), .ZN(n17880) );
  NAND3_X2 U14552 ( .A1(n19141), .A2(ID_EXEC_OUT[156]), .A3(n19140), .ZN(
        n19142) );
  NAND4_X1 U14553 ( .A1(n18895), .A2(n13050), .A3(n13070), .A4(n18886), .ZN(
        n18849) );
  NOR2_X1 U14554 ( .A1(n13103), .A2(destReg_wb_out[4]), .ZN(n129) );
  NOR2_X1 U14555 ( .A1(n19320), .A2(n13103), .ZN(n94) );
  NAND3_X2 U14556 ( .A1(n18912), .A2(n18913), .A3(n18906), .ZN(n18916) );
  OAI211_X2 U14557 ( .C1(n18915), .C2(n18914), .A(n18912), .B(n18913), .ZN(
        n18918) );
  NAND3_X2 U14558 ( .A1(n18893), .A2(n18892), .A3(n19364), .ZN(n18899) );
  NAND2_X4 U14559 ( .A1(n10123), .A2(n15540), .ZN(net227180) );
  XNOR2_X1 U14560 ( .A(net239774), .B(net239823), .ZN(n18528) );
  OAI21_X1 U14561 ( .B1(net239774), .B2(net239823), .A(net239150), .ZN(n18447)
         );
  NAND4_X1 U14562 ( .A1(n17896), .A2(n17895), .A3(n17894), .A4(n17893), .ZN(
        n17899) );
  XOR2_X1 U14564 ( .A(n13220), .B(n13152), .Z(n5466) );
  XOR2_X1 U14565 ( .A(offset_26_id[2]), .B(n13152), .Z(n2538) );
  NAND3_X1 U14566 ( .A1(n14098), .A2(n15686), .A3(n13055), .ZN(n14058) );
  NAND3_X1 U14567 ( .A1(n15700), .A2(n13055), .A3(n14098), .ZN(n13996) );
  NOR2_X1 U14568 ( .A1(n14098), .A2(n14051), .ZN(n14052) );
  NAND2_X1 U14569 ( .A1(n10116), .A2(net239459), .ZN(n17327) );
  NAND2_X4 U14570 ( .A1(n15642), .A2(n15641), .ZN(n17215) );
  NAND2_X4 U14571 ( .A1(net227052), .A2(net225076), .ZN(n15566) );
  NAND3_X2 U14572 ( .A1(n17216), .A2(n17222), .A3(n17201), .ZN(n17207) );
  OAI211_X4 U14573 ( .C1(net224837), .C2(net224838), .A(net224839), .B(
        net224840), .ZN(n17216) );
  OAI211_X4 U14574 ( .C1(n18998), .C2(n18997), .A(n18995), .B(n18996), .ZN(
        n19009) );
  NAND3_X2 U14575 ( .A1(n18905), .A2(n18904), .A3(n18903), .ZN(n18912) );
  NAND4_X4 U14576 ( .A1(n19056), .A2(n19058), .A3(n19057), .A4(n19059), .ZN(
        n19140) );
  NAND2_X4 U14577 ( .A1(n13981), .A2(n13980), .ZN(n14091) );
  INV_X8 U14578 ( .A(n18383), .ZN(n18966) );
  NAND2_X4 U14579 ( .A1(n18372), .A2(n14050), .ZN(n18861) );
  NAND2_X4 U14580 ( .A1(n14061), .A2(n14060), .ZN(n18942) );
  NAND2_X4 U14581 ( .A1(n18261), .A2(n14090), .ZN(n18944) );
  INV_X16 U14582 ( .A(n14192), .ZN(n15603) );
  INV_X32 U14583 ( .A(n13177), .ZN(n13178) );
  INV_X32 U14584 ( .A(n13179), .ZN(n13180) );
  INV_X32 U14585 ( .A(n13185), .ZN(n13186) );
  NAND2_X4 U14586 ( .A1(n14990), .A2(n2503), .ZN(n17269) );
  INV_X16 U14587 ( .A(n13182), .ZN(n19154) );
  NAND2_X4 U14588 ( .A1(n10244), .A2(n15610), .ZN(n18699) );
  NAND4_X4 U14589 ( .A1(n15662), .A2(n15664), .A3(ID_EXEC_OUT[148]), .A4(
        n15663), .ZN(n18928) );
  NAND2_X4 U14590 ( .A1(n15670), .A2(n15669), .ZN(n15836) );
  INV_X32 U14591 ( .A(net232816), .ZN(net232817) );
  INV_X8 U14592 ( .A(net222304), .ZN(net223324) );
  NAND2_X4 U14593 ( .A1(n15723), .A2(n18651), .ZN(n18677) );
  NAND2_X4 U14594 ( .A1(n16879), .A2(n16007), .ZN(n16064) );
  INV_X32 U14595 ( .A(n13212), .ZN(n13213) );
  NAND2_X4 U14596 ( .A1(n19088), .A2(n18651), .ZN(n18451) );
  INV_X4 U14597 ( .A(n19114), .ZN(n13216) );
  INV_X16 U14598 ( .A(n13213), .ZN(n19118) );
  INV_X16 U14599 ( .A(n18699), .ZN(n18494) );
  INV_X32 U14600 ( .A(n13346), .ZN(n13345) );
  INV_X32 U14601 ( .A(n13351), .ZN(n13350) );
  INV_X32 U14602 ( .A(n13360), .ZN(n13359) );
  INV_X32 U14603 ( .A(n13391), .ZN(n13388) );
  INV_X32 U14604 ( .A(n13391), .ZN(n13389) );
  INV_X32 U14605 ( .A(n13391), .ZN(n13390) );
  INV_X32 U14606 ( .A(n13395), .ZN(n13392) );
  INV_X32 U14607 ( .A(n13398), .ZN(n13396) );
  INV_X32 U14608 ( .A(n13482), .ZN(n13481) );
  INV_X16 U14609 ( .A(n13478), .ZN(n13482) );
  INV_X32 U14610 ( .A(n13486), .ZN(n13484) );
  INV_X32 U14611 ( .A(n13218), .ZN(n13493) );
  INV_X32 U14612 ( .A(n13218), .ZN(n13494) );
  NAND2_X2 U14613 ( .A1(net139963), .A2(n10157), .ZN(n1746) );
  NAND2_X2 U14614 ( .A1(MEM_WB_OUT[26]), .A2(n13878), .ZN(n13957) );
  INV_X4 U14615 ( .A(n13957), .ZN(n13958) );
  AOI21_X4 U14616 ( .B1(n13959), .B2(n14079), .A(n13958), .ZN(n13967) );
  INV_X4 U14617 ( .A(n14074), .ZN(n13985) );
  NAND3_X4 U14618 ( .A1(n13967), .A2(n13966), .A3(n13965), .ZN(n15837) );
  NOR2_X4 U14619 ( .A1(n13968), .A2(n15665), .ZN(n13973) );
  NOR2_X4 U14620 ( .A1(n13969), .A2(n13970), .ZN(n13972) );
  NAND3_X4 U14621 ( .A1(n13973), .A2(n13972), .A3(n13971), .ZN(n14099) );
  NAND3_X4 U14622 ( .A1(n13983), .A2(n13984), .A3(n13982), .ZN(n18345) );
  INV_X4 U14623 ( .A(n18345), .ZN(n14011) );
  NAND3_X4 U14624 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[22]), .A2(
        n13880), .A3(n13073), .ZN(n14012) );
  INV_X4 U14625 ( .A(n14012), .ZN(n13987) );
  NAND2_X2 U14627 ( .A1(MEM_WB_OUT[30]), .A2(n13878), .ZN(n13988) );
  INV_X4 U14628 ( .A(n13988), .ZN(n13989) );
  NAND2_X2 U14630 ( .A1(DMEM_BUS_OUT[30]), .A2(n13157), .ZN(n13995) );
  NAND2_X2 U14631 ( .A1(DMEM_BUS_OUT[20]), .A2(n18654), .ZN(n14005) );
  NAND2_X2 U14632 ( .A1(ID_EXEC_OUT[52]), .A2(n13356), .ZN(n17544) );
  INV_X4 U14633 ( .A(n13998), .ZN(n14119) );
  NAND2_X2 U14635 ( .A1(MEM_WB_OUT[57]), .A2(n13223), .ZN(n14002) );
  NOR2_X4 U14636 ( .A1(n13154), .A2(n12568), .ZN(n14124) );
  NAND3_X4 U14637 ( .A1(n14081), .A2(n13880), .A3(n14125), .ZN(n14068) );
  NAND2_X2 U14638 ( .A1(n13406), .A2(n17546), .ZN(n14004) );
  NAND3_X4 U14639 ( .A1(n14005), .A2(n17544), .A3(n14004), .ZN(n17505) );
  INV_X4 U14640 ( .A(n17505), .ZN(n18992) );
  NAND2_X2 U14641 ( .A1(DMEM_BUS_OUT[21]), .A2(n18654), .ZN(n14010) );
  NAND2_X2 U14642 ( .A1(ID_EXEC_OUT[53]), .A2(n13356), .ZN(n17680) );
  NAND2_X2 U14643 ( .A1(MEM_WB_OUT[58]), .A2(n13224), .ZN(n14007) );
  NAND2_X2 U14644 ( .A1(n13406), .A2(n17622), .ZN(n14009) );
  NAND3_X4 U14645 ( .A1(n14010), .A2(n17680), .A3(n14009), .ZN(n17712) );
  INV_X4 U14646 ( .A(n17712), .ZN(n18986) );
  NAND4_X2 U14647 ( .A1(n14011), .A2(n18462), .A3(n18992), .A4(n18986), .ZN(
        n14025) );
  NAND2_X2 U14648 ( .A1(DMEM_BUS_OUT[22]), .A2(n18654), .ZN(n14018) );
  NAND2_X2 U14649 ( .A1(ID_EXEC_OUT[54]), .A2(n15712), .ZN(n17842) );
  INV_X4 U14650 ( .A(n14012), .ZN(n14013) );
  AOI21_X4 U14651 ( .B1(n14013), .B2(n13985), .A(n14104), .ZN(n14014) );
  NAND3_X4 U14652 ( .A1(n14016), .A2(n14015), .A3(n14014), .ZN(n17840) );
  NAND2_X2 U14653 ( .A1(n18664), .A2(n17840), .ZN(n14017) );
  NAND3_X4 U14654 ( .A1(n14018), .A2(n17842), .A3(n14017), .ZN(n18980) );
  NAND2_X2 U14655 ( .A1(DMEM_BUS_OUT[17]), .A2(n18654), .ZN(n14024) );
  NAND2_X2 U14656 ( .A1(ID_EXEC_OUT[49]), .A2(n15712), .ZN(n17137) );
  AOI22_X2 U14657 ( .A1(MEM_WB_OUT[17]), .A2(n13878), .B1(MEM_WB_OUT[86]), 
        .B2(n14102), .ZN(n14022) );
  NAND2_X2 U14658 ( .A1(MEM_WB_OUT[54]), .A2(n13224), .ZN(n14021) );
  NAND3_X4 U14659 ( .A1(n14024), .A2(n17137), .A3(n14023), .ZN(n18888) );
  NAND2_X2 U14660 ( .A1(DMEM_BUS_OUT[18]), .A2(n13157), .ZN(n14030) );
  NAND2_X2 U14661 ( .A1(ID_EXEC_OUT[50]), .A2(n13356), .ZN(n18564) );
  NAND2_X2 U14662 ( .A1(MEM_WB_OUT[55]), .A2(n13223), .ZN(n14027) );
  NAND2_X2 U14663 ( .A1(n13405), .A2(n17331), .ZN(n14029) );
  NAND3_X4 U14664 ( .A1(n14030), .A2(n18564), .A3(n14029), .ZN(n18559) );
  NAND2_X2 U14665 ( .A1(DMEM_BUS_OUT[19]), .A2(n18654), .ZN(n14035) );
  NAND2_X2 U14666 ( .A1(ID_EXEC_OUT[51]), .A2(n13356), .ZN(n17904) );
  NAND2_X2 U14667 ( .A1(MEM_WB_OUT[56]), .A2(n13223), .ZN(n14032) );
  NAND2_X2 U14668 ( .A1(n13406), .A2(n17382), .ZN(n14034) );
  NAND3_X4 U14669 ( .A1(n14035), .A2(n17904), .A3(n14034), .ZN(n18911) );
  NAND2_X2 U14670 ( .A1(MEM_WB_OUT[62]), .A2(n13223), .ZN(n14041) );
  NOR2_X4 U14671 ( .A1(n14092), .A2(n12033), .ZN(n14039) );
  NOR2_X4 U14672 ( .A1(n14038), .A2(n14039), .ZN(n14040) );
  AOI21_X4 U14673 ( .B1(DMEM_BUS_OUT[25]), .B2(n18654), .A(n18384), .ZN(n18383) );
  NAND2_X2 U14674 ( .A1(DMEM_BUS_OUT[27]), .A2(n13157), .ZN(n14050) );
  INV_X4 U14675 ( .A(ID_EXEC_OUT[61]), .ZN(n14051) );
  NAND2_X2 U14676 ( .A1(n14052), .A2(n13056), .ZN(n14059) );
  NAND2_X2 U14678 ( .A1(MEM_WB_OUT[66]), .A2(n13223), .ZN(n14056) );
  NAND2_X2 U14679 ( .A1(n14059), .A2(n14058), .ZN(n18457) );
  INV_X4 U14680 ( .A(n18457), .ZN(n14061) );
  NAND2_X2 U14681 ( .A1(DMEM_BUS_OUT[29]), .A2(n13157), .ZN(n14060) );
  NAND2_X2 U14682 ( .A1(ID_EXEC_OUT[55]), .A2(n15712), .ZN(n14072) );
  NOR2_X4 U14683 ( .A1(n13877), .A2(n10940), .ZN(n14064) );
  NAND2_X2 U14684 ( .A1(MEM_WB_OUT[23]), .A2(n13878), .ZN(n14062) );
  INV_X4 U14685 ( .A(n14062), .ZN(n14063) );
  NAND3_X4 U14686 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[23]), .A2(
        n13880), .A3(n13073), .ZN(n14077) );
  NAND2_X2 U14687 ( .A1(DMEM_BUS_OUT[23]), .A2(n13157), .ZN(n14070) );
  NAND3_X4 U14688 ( .A1(n14072), .A2(n14071), .A3(n14070), .ZN(n18922) );
  NOR3_X4 U14689 ( .A1(n13878), .A2(n13073), .A3(n10910), .ZN(n14075) );
  NOR3_X4 U14690 ( .A1(n14076), .A2(n12501), .A3(n14075), .ZN(n14084) );
  INV_X4 U14691 ( .A(n14077), .ZN(n14082) );
  AOI22_X2 U14692 ( .A1(n14082), .A2(n14081), .B1(n14080), .B2(n14079), .ZN(
        n14083) );
  NAND2_X2 U14693 ( .A1(n13157), .A2(DMEM_BUS_OUT[31]), .ZN(n18926) );
  NAND3_X4 U14694 ( .A1(n13156), .A2(n18926), .A3(n13155), .ZN(n19125) );
  AOI22_X2 U14695 ( .A1(MEM_WB_OUT[28]), .A2(n13877), .B1(MEM_WB_OUT[97]), 
        .B2(n14102), .ZN(n14089) );
  NAND2_X2 U14696 ( .A1(MEM_WB_OUT[65]), .A2(n13224), .ZN(n14088) );
  NOR2_X4 U14697 ( .A1(n14086), .A2(n14085), .ZN(n14087) );
  NAND3_X4 U14698 ( .A1(n14089), .A2(n14088), .A3(n14087), .ZN(n15678) );
  NAND2_X2 U14699 ( .A1(DMEM_BUS_OUT[28]), .A2(n13157), .ZN(n14090) );
  NAND2_X2 U14700 ( .A1(MEM_WB_OUT[61]), .A2(n13223), .ZN(n14096) );
  NOR2_X4 U14701 ( .A1(n14103), .A2(n12066), .ZN(n14093) );
  NOR2_X4 U14702 ( .A1(n14094), .A2(n14093), .ZN(n14095) );
  NAND3_X4 U14703 ( .A1(n14097), .A2(n14096), .A3(n14095), .ZN(n15770) );
  NAND2_X2 U14704 ( .A1(n14101), .A2(n14100), .ZN(n18293) );
  NAND2_X2 U14705 ( .A1(MEM_WB_OUT[53]), .A2(n13223), .ZN(n14107) );
  NAND3_X4 U14707 ( .A1(n14111), .A2(n14110), .A3(n14109), .ZN(n18884) );
  NAND4_X2 U14708 ( .A1(n14115), .A2(n14114), .A3(n14113), .A4(n14112), .ZN(
        n6892) );
  NAND2_X2 U14709 ( .A1(MEM_WB_OUT[0]), .A2(n13878), .ZN(n14121) );
  NAND2_X2 U14710 ( .A1(MEM_WB_OUT[37]), .A2(n13223), .ZN(n14120) );
  OAI211_X2 U14711 ( .C1(n14122), .C2(n13165), .A(n14121), .B(n14120), .ZN(
        n18623) );
  INV_X4 U14712 ( .A(n18623), .ZN(n18662) );
  AOI21_X4 U14713 ( .B1(n18654), .B2(DMEM_BUS_OUT[0]), .A(n18653), .ZN(n18587)
         );
  INV_X4 U14714 ( .A(n19068), .ZN(n16791) );
  NAND2_X2 U14715 ( .A1(DMEM_BUS_OUT[6]), .A2(n18654), .ZN(n14128) );
  NAND2_X2 U14716 ( .A1(ID_EXEC_OUT[38]), .A2(n13356), .ZN(n16145) );
  AOI22_X2 U14717 ( .A1(MEM_WB_OUT[43]), .A2(n13222), .B1(MEM_WB_OUT[6]), .B2(
        n13877), .ZN(n14126) );
  NAND2_X2 U14718 ( .A1(n13406), .A2(n16147), .ZN(n14127) );
  NAND3_X4 U14719 ( .A1(n14128), .A2(n16145), .A3(n14127), .ZN(n19038) );
  NAND2_X2 U14720 ( .A1(n16791), .A2(n18534), .ZN(n14135) );
  NAND2_X2 U14721 ( .A1(DMEM_BUS_OUT[3]), .A2(n18654), .ZN(n14131) );
  NAND2_X2 U14722 ( .A1(ID_EXEC_OUT[35]), .A2(n13356), .ZN(n17566) );
  AOI22_X2 U14723 ( .A1(MEM_WB_OUT[40]), .A2(n13222), .B1(MEM_WB_OUT[3]), .B2(
        n13877), .ZN(n14129) );
  NAND2_X2 U14724 ( .A1(n13406), .A2(n16918), .ZN(n14130) );
  NAND3_X4 U14725 ( .A1(n14131), .A2(n17566), .A3(n14130), .ZN(n18872) );
  NAND2_X2 U14726 ( .A1(DMEM_BUS_OUT[2]), .A2(n18654), .ZN(n14134) );
  NAND2_X2 U14727 ( .A1(n13356), .A2(ID_EXEC_OUT[34]), .ZN(n16870) );
  AOI22_X2 U14728 ( .A1(MEM_WB_OUT[39]), .A2(n13222), .B1(MEM_WB_OUT[2]), .B2(
        n13877), .ZN(n14132) );
  NAND2_X2 U14729 ( .A1(n13406), .A2(n16872), .ZN(n14133) );
  NAND3_X4 U14730 ( .A1(n14134), .A2(n16870), .A3(n14133), .ZN(n18873) );
  NAND2_X2 U14731 ( .A1(DMEM_BUS_OUT[10]), .A2(n18654), .ZN(n14138) );
  NAND2_X2 U14732 ( .A1(ID_EXEC_OUT[42]), .A2(n13356), .ZN(n16296) );
  AOI22_X2 U14733 ( .A1(MEM_WB_OUT[47]), .A2(n13222), .B1(MEM_WB_OUT[10]), 
        .B2(n13877), .ZN(n14136) );
  NAND2_X2 U14734 ( .A1(n13406), .A2(n16295), .ZN(n14137) );
  NAND3_X4 U14735 ( .A1(n14138), .A2(n16296), .A3(n14137), .ZN(n19015) );
  NAND2_X2 U14736 ( .A1(DMEM_BUS_OUT[9]), .A2(n18654), .ZN(n14141) );
  NAND2_X2 U14737 ( .A1(ID_EXEC_OUT[41]), .A2(n13356), .ZN(n17046) );
  AOI22_X2 U14738 ( .A1(MEM_WB_OUT[46]), .A2(n13222), .B1(MEM_WB_OUT[9]), .B2(
        n13877), .ZN(n14139) );
  NAND2_X2 U14739 ( .A1(n13406), .A2(n17045), .ZN(n14140) );
  NAND3_X4 U14740 ( .A1(n14141), .A2(n17046), .A3(n14140), .ZN(n19013) );
  NAND2_X2 U14741 ( .A1(DMEM_BUS_OUT[4]), .A2(n18654), .ZN(n14144) );
  NAND2_X2 U14742 ( .A1(ID_EXEC_OUT[36]), .A2(n13356), .ZN(n17309) );
  AOI22_X2 U14743 ( .A1(MEM_WB_OUT[41]), .A2(n13222), .B1(MEM_WB_OUT[4]), .B2(
        n13877), .ZN(n14142) );
  NAND2_X2 U14744 ( .A1(n13406), .A2(n17242), .ZN(n14143) );
  NAND3_X4 U14745 ( .A1(n14144), .A2(n17309), .A3(n14143), .ZN(n18867) );
  NAND2_X2 U14746 ( .A1(DMEM_BUS_OUT[11]), .A2(n18654), .ZN(n14147) );
  NAND2_X2 U14747 ( .A1(ID_EXEC_OUT[43]), .A2(n13356), .ZN(n16409) );
  AOI22_X2 U14748 ( .A1(MEM_WB_OUT[48]), .A2(n13222), .B1(MEM_WB_OUT[11]), 
        .B2(n13877), .ZN(n14145) );
  NAND2_X2 U14749 ( .A1(n13406), .A2(n16350), .ZN(n14146) );
  NAND3_X4 U14750 ( .A1(n14147), .A2(n16409), .A3(n14146), .ZN(n19004) );
  NOR4_X2 U14751 ( .A1(n19015), .A2(n19013), .A3(n18867), .A4(n19004), .ZN(
        n14185) );
  NAND2_X2 U14752 ( .A1(DMEM_BUS_OUT[15]), .A2(n13157), .ZN(n14152) );
  NAND2_X2 U14753 ( .A1(n13164), .A2(
        WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[31]), .ZN(n14150) );
  NAND3_X4 U14754 ( .A1(n14151), .A2(n17871), .A3(n14152), .ZN(n19091) );
  NAND2_X2 U14755 ( .A1(DMEM_BUS_OUT[13]), .A2(n18654), .ZN(n14155) );
  NAND2_X2 U14756 ( .A1(ID_EXEC_OUT[45]), .A2(n13356), .ZN(n17604) );
  AOI22_X2 U14757 ( .A1(MEM_WB_OUT[50]), .A2(n13222), .B1(MEM_WB_OUT[13]), 
        .B2(n13877), .ZN(n14153) );
  NAND2_X2 U14758 ( .A1(n13406), .A2(n16578), .ZN(n14154) );
  NAND3_X4 U14759 ( .A1(n14155), .A2(n17604), .A3(n14154), .ZN(net222497) );
  NAND2_X2 U14760 ( .A1(ID_EXEC_OUT[44]), .A2(n13356), .ZN(n14159) );
  AOI22_X2 U14761 ( .A1(MEM_WB_OUT[49]), .A2(n13223), .B1(MEM_WB_OUT[12]), 
        .B2(n13877), .ZN(n14156) );
  NAND2_X2 U14762 ( .A1(n13406), .A2(n16539), .ZN(n14158) );
  NAND2_X2 U14763 ( .A1(DMEM_BUS_OUT[12]), .A2(n18654), .ZN(n14157) );
  NAND3_X4 U14764 ( .A1(n14159), .A2(n14158), .A3(n14157), .ZN(n19000) );
  NAND2_X2 U14765 ( .A1(ID_EXEC_OUT[40]), .A2(n13356), .ZN(n14163) );
  AOI22_X2 U14766 ( .A1(MEM_WB_OUT[45]), .A2(n13223), .B1(MEM_WB_OUT[8]), .B2(
        n13877), .ZN(n14160) );
  NAND2_X2 U14767 ( .A1(n13406), .A2(n16222), .ZN(n14162) );
  NAND2_X2 U14768 ( .A1(DMEM_BUS_OUT[8]), .A2(n18654), .ZN(n14161) );
  NAND3_X4 U14769 ( .A1(n14163), .A2(n14162), .A3(n14161), .ZN(n19029) );
  NAND2_X2 U14770 ( .A1(ID_EXEC_OUT[39]), .A2(n13356), .ZN(n14167) );
  AOI22_X2 U14771 ( .A1(MEM_WB_OUT[44]), .A2(n13223), .B1(MEM_WB_OUT[7]), .B2(
        n13877), .ZN(n14164) );
  NAND2_X2 U14772 ( .A1(n13406), .A2(n16070), .ZN(n14166) );
  NAND2_X2 U14773 ( .A1(DMEM_BUS_OUT[7]), .A2(n18654), .ZN(n14165) );
  NAND3_X4 U14774 ( .A1(n14167), .A2(n14166), .A3(n14165), .ZN(n16971) );
  NAND2_X2 U14775 ( .A1(ID_EXEC_OUT[37]), .A2(n13356), .ZN(n14171) );
  AOI22_X2 U14776 ( .A1(MEM_WB_OUT[42]), .A2(n13222), .B1(MEM_WB_OUT[5]), .B2(
        n13877), .ZN(n14168) );
  NAND2_X2 U14777 ( .A1(n13406), .A2(n16031), .ZN(n14170) );
  NAND2_X2 U14778 ( .A1(DMEM_BUS_OUT[5]), .A2(n18654), .ZN(n14169) );
  NAND3_X4 U14779 ( .A1(n14171), .A2(n14170), .A3(n14169), .ZN(net225212) );
  NAND2_X2 U14780 ( .A1(ID_EXEC_OUT[46]), .A2(n13356), .ZN(n14175) );
  NAND2_X2 U14781 ( .A1(DMEM_BUS_OUT[14]), .A2(n18654), .ZN(n14173) );
  NAND3_X4 U14782 ( .A1(n14175), .A2(n14174), .A3(n14173), .ZN(n18897) );
  NAND2_X2 U14783 ( .A1(ID_EXEC_OUT[33]), .A2(n13356), .ZN(n14182) );
  AOI22_X2 U14784 ( .A1(n13222), .A2(MEM_WB_OUT[38]), .B1(MEM_WB_OUT[1]), .B2(
        n13877), .ZN(n14177) );
  OAI211_X2 U14785 ( .C1(n13165), .C2(n12033), .A(n13048), .B(n14177), .ZN(
        n15718) );
  NAND2_X2 U14786 ( .A1(n13406), .A2(n15718), .ZN(n14181) );
  NAND2_X2 U14787 ( .A1(n18654), .A2(DMEM_BUS_OUT[1]), .ZN(n14180) );
  NAND3_X4 U14788 ( .A1(n14182), .A2(n14181), .A3(n14180), .ZN(n18870) );
  NOR4_X2 U14789 ( .A1(n16971), .A2(net225212), .A3(n18897), .A4(n18870), .ZN(
        n14183) );
  NAND4_X2 U14790 ( .A1(n14186), .A2(n14185), .A3(n14184), .A4(n14183), .ZN(
        n6893) );
  NAND2_X2 U14791 ( .A1(ID_STAGE_imm16_aluA[16]), .A2(net230387), .ZN(n2564)
         );
  INV_X4 U14792 ( .A(n14187), .ZN(n19163) );
  NOR2_X4 U14793 ( .A1(IF_ID_OUT[32]), .A2(IF_ID_OUT[35]), .ZN(n18768) );
  NOR2_X4 U14794 ( .A1(n12020), .A2(n14208), .ZN(n14209) );
  INV_X4 U14795 ( .A(n14209), .ZN(n5558) );
  INV_X4 U14796 ( .A(n14208), .ZN(n14188) );
  NAND2_X2 U14797 ( .A1(n14188), .A2(net230387), .ZN(n4685) );
  INV_X4 U14798 ( .A(n14233), .ZN(n14238) );
  NOR2_X4 U14799 ( .A1(IF_ID_OUT[37]), .A2(IF_ID_OUT[36]), .ZN(n14255) );
  NOR2_X4 U14800 ( .A1(ID_STAGE_imm16_aluA[31]), .A2(ID_STAGE_imm16_aluA[30]), 
        .ZN(n18771) );
  NAND2_X2 U14801 ( .A1(n14189), .A2(n12300), .ZN(n14190) );
  NOR2_X4 U14802 ( .A1(n14191), .A2(n14190), .ZN(n14204) );
  NOR3_X4 U14803 ( .A1(n14194), .A2(ID_STAGE_imm16_aluA[21]), .A3(n12128), 
        .ZN(n14203) );
  NAND2_X2 U14804 ( .A1(n14196), .A2(n14195), .ZN(n14201) );
  NOR2_X4 U14805 ( .A1(ID_STAGE_imm16_aluA[17]), .A2(ID_STAGE_imm16_aluA[16]), 
        .ZN(n14197) );
  NAND2_X2 U14806 ( .A1(n14197), .A2(n11922), .ZN(n14200) );
  NOR2_X4 U14807 ( .A1(ID_STAGE_imm16_aluA[19]), .A2(ID_STAGE_imm16_aluA[20]), 
        .ZN(n14198) );
  NAND2_X2 U14808 ( .A1(n14198), .A2(n11045), .ZN(n14199) );
  NOR3_X4 U14809 ( .A1(n14201), .A2(n14200), .A3(n14199), .ZN(n14202) );
  NAND3_X4 U14810 ( .A1(n14210), .A2(n12016), .A3(n14205), .ZN(n18781) );
  NAND2_X2 U14811 ( .A1(n18768), .A2(n12020), .ZN(n14206) );
  NOR2_X4 U14812 ( .A1(n18781), .A2(n14206), .ZN(n15631) );
  NAND3_X2 U14813 ( .A1(n5520), .A2(n18780), .A3(n14207), .ZN(n14216) );
  NAND2_X2 U14814 ( .A1(IF_ID_OUT[35]), .A2(n12134), .ZN(n14220) );
  NAND2_X2 U14815 ( .A1(n14211), .A2(n12555), .ZN(n14212) );
  NAND4_X2 U14816 ( .A1(n18769), .A2(net230387), .A3(n14216), .A4(n14215), 
        .ZN(n5555) );
  NAND4_X2 U14817 ( .A1(n18780), .A2(n5520), .A3(n10359), .A4(IF_ID_OUT[34]), 
        .ZN(n5549) );
  INV_X4 U14818 ( .A(n18781), .ZN(n18788) );
  INV_X4 U14819 ( .A(n15393), .ZN(n14217) );
  NAND2_X2 U14820 ( .A1(IF_ID_OUT[34]), .A2(n18768), .ZN(n14221) );
  INV_X4 U14821 ( .A(n14218), .ZN(n18756) );
  NAND2_X2 U14822 ( .A1(n14219), .A2(n18756), .ZN(n14222) );
  OAI22_X2 U14823 ( .A1(n5513), .A2(n14221), .B1(n14233), .B2(n14222), .ZN(
        n5516) );
  INV_X4 U14824 ( .A(n14220), .ZN(n18774) );
  NAND2_X2 U14825 ( .A1(IF_ID_OUT[34]), .A2(n18774), .ZN(n14239) );
  INV_X4 U14826 ( .A(n14239), .ZN(n14254) );
  NAND2_X2 U14827 ( .A1(n14254), .A2(n12555), .ZN(n14224) );
  INV_X4 U14828 ( .A(n14224), .ZN(n14235) );
  INV_X4 U14829 ( .A(n14246), .ZN(n14231) );
  INV_X4 U14830 ( .A(n14221), .ZN(n18754) );
  NAND2_X2 U14831 ( .A1(n18754), .A2(n13221), .ZN(n14266) );
  INV_X4 U14832 ( .A(n14266), .ZN(n14247) );
  INV_X4 U14833 ( .A(n14222), .ZN(n14265) );
  INV_X4 U14834 ( .A(n14241), .ZN(n14256) );
  NAND2_X2 U14835 ( .A1(n14256), .A2(n10840), .ZN(n14232) );
  INV_X4 U14836 ( .A(n14232), .ZN(n14223) );
  AOI22_X2 U14837 ( .A1(n14223), .A2(n14264), .B1(n19301), .B2(n14235), .ZN(
        n14262) );
  NAND2_X2 U14838 ( .A1(n14262), .A2(n14227), .ZN(n14252) );
  INV_X4 U14839 ( .A(n14252), .ZN(n14228) );
  NAND4_X2 U14840 ( .A1(n14230), .A2(n14229), .A3(n14263), .A4(n14228), .ZN(
        n5478) );
  INV_X4 U14841 ( .A(n18766), .ZN(n14264) );
  NAND2_X2 U14842 ( .A1(n14231), .A2(n14264), .ZN(n14237) );
  OAI211_X2 U14843 ( .C1(n5520), .C2(n14242), .A(n14237), .B(n14248), .ZN(
        n5484) );
  NAND2_X2 U14844 ( .A1(ID_STAGE_imm16_aluA[28]), .A2(n14238), .ZN(n14240) );
  INV_X4 U14845 ( .A(n14242), .ZN(n14243) );
  NAND2_X2 U14846 ( .A1(n14243), .A2(n5506), .ZN(n14244) );
  NAND2_X2 U14847 ( .A1(n5506), .A2(n14247), .ZN(n14250) );
  INV_X4 U14848 ( .A(n5516), .ZN(n14249) );
  NAND4_X2 U14849 ( .A1(n14251), .A2(n14250), .A3(n14249), .A4(n14248), .ZN(
        n14253) );
  INV_X4 U14850 ( .A(n14257), .ZN(n14258) );
  INV_X4 U14851 ( .A(n18760), .ZN(n14261) );
  NOR4_X2 U14852 ( .A1(n14268), .A2(n12955), .A3(n5484), .A4(n14267), .ZN(
        n5482) );
  INV_X4 U14853 ( .A(n14269), .ZN(n14272) );
  NAND2_X2 U14854 ( .A1(n14272), .A2(n10368), .ZN(n14278) );
  INV_X4 U14855 ( .A(n14278), .ZN(n14999) );
  INV_X4 U14856 ( .A(n14275), .ZN(n14991) );
  NAND2_X2 U14857 ( .A1(n2531), .A2(net231359), .ZN(n14270) );
  INV_X4 U14858 ( .A(n14270), .ZN(n14293) );
  INV_X4 U14859 ( .A(n14276), .ZN(n14995) );
  INV_X4 U14860 ( .A(n14271), .ZN(n14990) );
  NAND2_X2 U14861 ( .A1(n2533), .A2(net231359), .ZN(n14281) );
  INV_X4 U14862 ( .A(n14281), .ZN(n14273) );
  INV_X4 U14863 ( .A(n14280), .ZN(n14986) );
  NAND2_X2 U14864 ( .A1(n2530), .A2(net231345), .ZN(n14279) );
  INV_X4 U14865 ( .A(n14279), .ZN(n14288) );
  INV_X4 U14866 ( .A(n14274), .ZN(n14997) );
  AOI22_X2 U14867 ( .A1(FP_REG_FILE_reg_out_24__0_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__0_), .B2(n13227), .ZN(n4662) );
  INV_X4 U14868 ( .A(n14277), .ZN(n14982) );
  AOI22_X2 U14869 ( .A1(FP_REG_FILE_reg_out_14__0_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__0_), .B2(n13231), .ZN(n14287) );
  NAND2_X2 U14870 ( .A1(FP_REG_FILE_reg_out_17__0_), .A2(n13234), .ZN(n14286)
         );
  NAND2_X2 U14871 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__0_), .ZN(n14285)
         );
  NAND2_X2 U14872 ( .A1(n14293), .A2(n14986), .ZN(n14283) );
  NAND2_X2 U14873 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__0_), .ZN(n14284)
         );
  NAND4_X2 U14874 ( .A1(n14287), .A2(n14286), .A3(n14285), .A4(n14284), .ZN(
        n4642) );
  NAND2_X2 U14875 ( .A1(FP_REG_FILE_reg_out_1__0_), .A2(n13242), .ZN(n14292)
         );
  NAND2_X2 U14876 ( .A1(FP_REG_FILE_reg_out_12__0_), .A2(n13240), .ZN(n14291)
         );
  NAND2_X2 U14877 ( .A1(n13168), .A2(FP_REG_FILE_reg_out_11__0_), .ZN(n14290)
         );
  NAND2_X2 U14878 ( .A1(n14400), .A2(FP_REG_FILE_reg_out_16__0_), .ZN(n14289)
         );
  NAND4_X2 U14879 ( .A1(n14292), .A2(n14291), .A3(n14290), .A4(n14289), .ZN(
        n4643) );
  OAI22_X2 U14880 ( .A1(n11373), .A2(n13248), .B1(n10400), .B2(n13246), .ZN(
        n14295) );
  AOI22_X2 U14881 ( .A1(FP_REG_FILE_reg_out_24__1_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__1_), .B2(n13227), .ZN(n4629) );
  AOI22_X2 U14882 ( .A1(FP_REG_FILE_reg_out_14__1_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__1_), .B2(n13231), .ZN(n14300) );
  NAND2_X2 U14883 ( .A1(FP_REG_FILE_reg_out_17__1_), .A2(n13235), .ZN(n14299)
         );
  NAND2_X2 U14884 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__1_), .ZN(n14298)
         );
  NAND2_X2 U14885 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__1_), .ZN(n14297)
         );
  NAND4_X2 U14886 ( .A1(n14300), .A2(n14299), .A3(n14298), .A4(n14297), .ZN(
        n4613) );
  NAND2_X2 U14887 ( .A1(FP_REG_FILE_reg_out_1__1_), .A2(n13243), .ZN(n14304)
         );
  NAND2_X2 U14888 ( .A1(FP_REG_FILE_reg_out_12__1_), .A2(n13241), .ZN(n14303)
         );
  NAND2_X2 U14889 ( .A1(n13168), .A2(FP_REG_FILE_reg_out_11__1_), .ZN(n14302)
         );
  NAND2_X2 U14890 ( .A1(n14400), .A2(FP_REG_FILE_reg_out_16__1_), .ZN(n14301)
         );
  NAND4_X2 U14891 ( .A1(n14304), .A2(n14303), .A3(n14302), .A4(n14301), .ZN(
        n4614) );
  OAI22_X2 U14892 ( .A1(n12284), .A2(n13248), .B1(n10913), .B2(n13246), .ZN(
        n14306) );
  AOI22_X2 U14893 ( .A1(FP_REG_FILE_reg_out_24__2_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__2_), .B2(n13227), .ZN(n4600) );
  AOI22_X2 U14894 ( .A1(FP_REG_FILE_reg_out_14__2_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__2_), .B2(n13231), .ZN(n14311) );
  NAND2_X2 U14895 ( .A1(FP_REG_FILE_reg_out_17__2_), .A2(n13234), .ZN(n14310)
         );
  NAND2_X2 U14896 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__2_), .ZN(n14309)
         );
  NAND2_X2 U14897 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__2_), .ZN(n14308)
         );
  NAND4_X2 U14898 ( .A1(n14311), .A2(n14310), .A3(n14309), .A4(n14308), .ZN(
        n4584) );
  NAND2_X2 U14899 ( .A1(FP_REG_FILE_reg_out_1__2_), .A2(n13242), .ZN(n14315)
         );
  NAND2_X2 U14900 ( .A1(FP_REG_FILE_reg_out_12__2_), .A2(n13240), .ZN(n14314)
         );
  NAND2_X2 U14901 ( .A1(n13168), .A2(FP_REG_FILE_reg_out_11__2_), .ZN(n14313)
         );
  NAND2_X2 U14902 ( .A1(n14400), .A2(FP_REG_FILE_reg_out_16__2_), .ZN(n14312)
         );
  NAND4_X2 U14903 ( .A1(n14315), .A2(n14314), .A3(n14313), .A4(n14312), .ZN(
        n4585) );
  OAI22_X2 U14904 ( .A1(n11394), .A2(n13248), .B1(n10401), .B2(n13246), .ZN(
        n14317) );
  AOI22_X2 U14905 ( .A1(FP_REG_FILE_reg_out_24__3_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__3_), .B2(n13227), .ZN(n4571) );
  AOI22_X2 U14906 ( .A1(FP_REG_FILE_reg_out_14__3_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__3_), .B2(n13231), .ZN(n14322) );
  NAND2_X2 U14907 ( .A1(FP_REG_FILE_reg_out_17__3_), .A2(n13235), .ZN(n14321)
         );
  NAND2_X2 U14908 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__3_), .ZN(n14320)
         );
  NAND2_X2 U14909 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__3_), .ZN(n14319)
         );
  NAND4_X2 U14910 ( .A1(n14322), .A2(n14321), .A3(n14320), .A4(n14319), .ZN(
        n4555) );
  NAND2_X2 U14911 ( .A1(FP_REG_FILE_reg_out_1__3_), .A2(n13243), .ZN(n14326)
         );
  NAND2_X2 U14912 ( .A1(FP_REG_FILE_reg_out_12__3_), .A2(n13241), .ZN(n14325)
         );
  NAND2_X2 U14913 ( .A1(n13168), .A2(FP_REG_FILE_reg_out_11__3_), .ZN(n14324)
         );
  NAND2_X2 U14914 ( .A1(n14400), .A2(FP_REG_FILE_reg_out_16__3_), .ZN(n14323)
         );
  NAND4_X2 U14915 ( .A1(n14326), .A2(n14325), .A3(n14324), .A4(n14323), .ZN(
        n4556) );
  OAI22_X2 U14916 ( .A1(n11397), .A2(n13248), .B1(n10402), .B2(n13246), .ZN(
        n14328) );
  AOI22_X2 U14917 ( .A1(FP_REG_FILE_reg_out_24__4_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__4_), .B2(n13227), .ZN(n4542) );
  AOI22_X2 U14918 ( .A1(FP_REG_FILE_reg_out_14__4_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__4_), .B2(n13231), .ZN(n14333) );
  NAND2_X2 U14919 ( .A1(FP_REG_FILE_reg_out_17__4_), .A2(n13234), .ZN(n14332)
         );
  NAND2_X2 U14920 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__4_), .ZN(n14331)
         );
  NAND2_X2 U14921 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__4_), .ZN(n14330)
         );
  NAND4_X2 U14922 ( .A1(n14333), .A2(n14332), .A3(n14331), .A4(n14330), .ZN(
        n4526) );
  NAND2_X2 U14923 ( .A1(FP_REG_FILE_reg_out_1__4_), .A2(n13242), .ZN(n14337)
         );
  NAND2_X2 U14924 ( .A1(FP_REG_FILE_reg_out_12__4_), .A2(n13240), .ZN(n14336)
         );
  NAND2_X2 U14925 ( .A1(n13168), .A2(FP_REG_FILE_reg_out_11__4_), .ZN(n14335)
         );
  NAND2_X2 U14926 ( .A1(n14400), .A2(FP_REG_FILE_reg_out_16__4_), .ZN(n14334)
         );
  NAND4_X2 U14927 ( .A1(n14337), .A2(n14336), .A3(n14335), .A4(n14334), .ZN(
        n4527) );
  OAI22_X2 U14928 ( .A1(n11398), .A2(n13248), .B1(n10403), .B2(n13246), .ZN(
        n14339) );
  AOI22_X2 U14929 ( .A1(FP_REG_FILE_reg_out_24__5_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__5_), .B2(n13227), .ZN(n4513) );
  AOI22_X2 U14930 ( .A1(FP_REG_FILE_reg_out_14__5_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__5_), .B2(n13231), .ZN(n14344) );
  NAND2_X2 U14931 ( .A1(FP_REG_FILE_reg_out_17__5_), .A2(n13235), .ZN(n14343)
         );
  NAND2_X2 U14932 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__5_), .ZN(n14342)
         );
  NAND2_X2 U14933 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__5_), .ZN(n14341)
         );
  NAND4_X2 U14934 ( .A1(n14344), .A2(n14343), .A3(n14342), .A4(n14341), .ZN(
        n4497) );
  NAND2_X2 U14935 ( .A1(FP_REG_FILE_reg_out_1__5_), .A2(n13243), .ZN(n14348)
         );
  NAND2_X2 U14936 ( .A1(FP_REG_FILE_reg_out_12__5_), .A2(n13241), .ZN(n14347)
         );
  NAND2_X2 U14937 ( .A1(n13168), .A2(FP_REG_FILE_reg_out_11__5_), .ZN(n14346)
         );
  NAND2_X2 U14938 ( .A1(n14400), .A2(FP_REG_FILE_reg_out_16__5_), .ZN(n14345)
         );
  NAND4_X2 U14939 ( .A1(n14348), .A2(n14347), .A3(n14346), .A4(n14345), .ZN(
        n4498) );
  OAI22_X2 U14940 ( .A1(n11399), .A2(n13248), .B1(n10404), .B2(n13246), .ZN(
        n14350) );
  AOI22_X2 U14941 ( .A1(FP_REG_FILE_reg_out_24__6_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__6_), .B2(n13227), .ZN(n4483) );
  AOI22_X2 U14942 ( .A1(FP_REG_FILE_reg_out_14__6_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__6_), .B2(n13231), .ZN(n14355) );
  NAND2_X2 U14943 ( .A1(FP_REG_FILE_reg_out_17__6_), .A2(n13234), .ZN(n14354)
         );
  NAND2_X2 U14944 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__6_), .ZN(n14353)
         );
  NAND2_X2 U14945 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__6_), .ZN(n14352)
         );
  NAND4_X2 U14946 ( .A1(n14355), .A2(n14354), .A3(n14353), .A4(n14352), .ZN(
        n4467) );
  NAND2_X2 U14947 ( .A1(FP_REG_FILE_reg_out_1__6_), .A2(n13242), .ZN(n14359)
         );
  NAND2_X2 U14948 ( .A1(FP_REG_FILE_reg_out_12__6_), .A2(n13240), .ZN(n14358)
         );
  NAND2_X2 U14949 ( .A1(n13168), .A2(FP_REG_FILE_reg_out_11__6_), .ZN(n14357)
         );
  NAND2_X2 U14950 ( .A1(n14400), .A2(FP_REG_FILE_reg_out_16__6_), .ZN(n14356)
         );
  NAND4_X2 U14951 ( .A1(n14359), .A2(n14358), .A3(n14357), .A4(n14356), .ZN(
        n4468) );
  OAI22_X2 U14952 ( .A1(n11400), .A2(n13248), .B1(n10405), .B2(n13246), .ZN(
        n14361) );
  AOI22_X2 U14953 ( .A1(FP_REG_FILE_reg_out_24__7_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__7_), .B2(n13227), .ZN(n4454) );
  AOI22_X2 U14954 ( .A1(FP_REG_FILE_reg_out_14__7_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__7_), .B2(n13231), .ZN(n14366) );
  NAND2_X2 U14955 ( .A1(FP_REG_FILE_reg_out_17__7_), .A2(n13235), .ZN(n14365)
         );
  NAND2_X2 U14956 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__7_), .ZN(n14364)
         );
  NAND2_X2 U14957 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__7_), .ZN(n14363)
         );
  NAND4_X2 U14958 ( .A1(n14366), .A2(n14365), .A3(n14364), .A4(n14363), .ZN(
        n4438) );
  NAND2_X2 U14959 ( .A1(FP_REG_FILE_reg_out_1__7_), .A2(n13243), .ZN(n14370)
         );
  NAND2_X2 U14960 ( .A1(FP_REG_FILE_reg_out_12__7_), .A2(n13241), .ZN(n14369)
         );
  NAND2_X2 U14961 ( .A1(n13168), .A2(FP_REG_FILE_reg_out_11__7_), .ZN(n14368)
         );
  NAND2_X2 U14962 ( .A1(n14400), .A2(FP_REG_FILE_reg_out_16__7_), .ZN(n14367)
         );
  NAND4_X2 U14963 ( .A1(n14370), .A2(n14369), .A3(n14368), .A4(n14367), .ZN(
        n4439) );
  OAI22_X2 U14964 ( .A1(n11401), .A2(n13248), .B1(n10406), .B2(n13246), .ZN(
        n14372) );
  AOI22_X2 U14965 ( .A1(FP_REG_FILE_reg_out_24__8_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__8_), .B2(n13227), .ZN(n4425) );
  AOI22_X2 U14966 ( .A1(FP_REG_FILE_reg_out_14__8_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__8_), .B2(n13231), .ZN(n14377) );
  NAND2_X2 U14967 ( .A1(FP_REG_FILE_reg_out_17__8_), .A2(n13234), .ZN(n14376)
         );
  NAND2_X2 U14968 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__8_), .ZN(n14375)
         );
  NAND2_X2 U14969 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__8_), .ZN(n14374)
         );
  NAND4_X2 U14970 ( .A1(n14377), .A2(n14376), .A3(n14375), .A4(n14374), .ZN(
        n4409) );
  NAND2_X2 U14971 ( .A1(FP_REG_FILE_reg_out_1__8_), .A2(n13242), .ZN(n14381)
         );
  NAND2_X2 U14972 ( .A1(FP_REG_FILE_reg_out_12__8_), .A2(n13240), .ZN(n14380)
         );
  NAND2_X2 U14973 ( .A1(n13168), .A2(FP_REG_FILE_reg_out_11__8_), .ZN(n14379)
         );
  NAND2_X2 U14974 ( .A1(n14400), .A2(FP_REG_FILE_reg_out_16__8_), .ZN(n14378)
         );
  NAND4_X2 U14975 ( .A1(n14381), .A2(n14380), .A3(n14379), .A4(n14378), .ZN(
        n4410) );
  OAI22_X2 U14976 ( .A1(n11402), .A2(n13248), .B1(n10407), .B2(n13246), .ZN(
        n14383) );
  AOI22_X2 U14977 ( .A1(FP_REG_FILE_reg_out_24__9_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__9_), .B2(n13227), .ZN(n4396) );
  AOI22_X2 U14978 ( .A1(FP_REG_FILE_reg_out_14__9_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__9_), .B2(n13231), .ZN(n14388) );
  NAND2_X2 U14979 ( .A1(FP_REG_FILE_reg_out_17__9_), .A2(n13235), .ZN(n14387)
         );
  NAND2_X2 U14980 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__9_), .ZN(n14386)
         );
  NAND2_X2 U14981 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__9_), .ZN(n14385)
         );
  NAND4_X2 U14982 ( .A1(n14388), .A2(n14387), .A3(n14386), .A4(n14385), .ZN(
        n4380) );
  NAND2_X2 U14983 ( .A1(FP_REG_FILE_reg_out_1__9_), .A2(n13243), .ZN(n14392)
         );
  NAND2_X2 U14984 ( .A1(FP_REG_FILE_reg_out_12__9_), .A2(n13241), .ZN(n14391)
         );
  NAND2_X2 U14985 ( .A1(n13168), .A2(FP_REG_FILE_reg_out_11__9_), .ZN(n14390)
         );
  NAND2_X2 U14986 ( .A1(n14400), .A2(FP_REG_FILE_reg_out_16__9_), .ZN(n14389)
         );
  NAND4_X2 U14987 ( .A1(n14392), .A2(n14391), .A3(n14390), .A4(n14389), .ZN(
        n4381) );
  OAI22_X2 U14988 ( .A1(n11403), .A2(n13248), .B1(n10408), .B2(n13246), .ZN(
        n14394) );
  AOI22_X2 U14989 ( .A1(FP_REG_FILE_reg_out_24__10_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__10_), .B2(n13226), .ZN(n4367) );
  AOI22_X2 U14990 ( .A1(FP_REG_FILE_reg_out_14__10_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__10_), .B2(n13230), .ZN(n14399) );
  NAND2_X2 U14991 ( .A1(FP_REG_FILE_reg_out_17__10_), .A2(n13235), .ZN(n14398)
         );
  NAND2_X2 U14992 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__10_), .ZN(n14397)
         );
  NAND2_X2 U14993 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__10_), .ZN(n14396)
         );
  NAND4_X2 U14994 ( .A1(n14399), .A2(n14398), .A3(n14397), .A4(n14396), .ZN(
        n4351) );
  NAND2_X2 U14995 ( .A1(FP_REG_FILE_reg_out_1__10_), .A2(n13243), .ZN(n14404)
         );
  NAND2_X2 U14996 ( .A1(FP_REG_FILE_reg_out_12__10_), .A2(n13241), .ZN(n14403)
         );
  NAND2_X2 U14997 ( .A1(n13168), .A2(FP_REG_FILE_reg_out_11__10_), .ZN(n14402)
         );
  NAND2_X2 U14998 ( .A1(n14400), .A2(FP_REG_FILE_reg_out_16__10_), .ZN(n14401)
         );
  NAND4_X2 U14999 ( .A1(n14404), .A2(n14403), .A3(n14402), .A4(n14401), .ZN(
        n4352) );
  OAI22_X2 U15000 ( .A1(n11374), .A2(n13248), .B1(n10409), .B2(n13246), .ZN(
        n14406) );
  AOI22_X2 U15001 ( .A1(FP_REG_FILE_reg_out_24__11_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__11_), .B2(n13226), .ZN(n4338) );
  AOI22_X2 U15002 ( .A1(FP_REG_FILE_reg_out_14__11_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__11_), .B2(n13230), .ZN(n14411) );
  NAND2_X2 U15003 ( .A1(FP_REG_FILE_reg_out_17__11_), .A2(n13235), .ZN(n14410)
         );
  NAND2_X2 U15004 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__11_), .ZN(n14409)
         );
  NAND2_X2 U15005 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__11_), .ZN(n14408)
         );
  NAND4_X2 U15006 ( .A1(n14411), .A2(n14410), .A3(n14409), .A4(n14408), .ZN(
        n4322) );
  AOI22_X2 U15007 ( .A1(FP_REG_FILE_reg_out_1__11_), .A2(n13243), .B1(
        FP_REG_FILE_reg_out_12__11_), .B2(n13241), .ZN(n14415) );
  NAND2_X2 U15008 ( .A1(n14415), .A2(n14414), .ZN(n4323) );
  OAI22_X2 U15009 ( .A1(n11375), .A2(n13249), .B1(n10410), .B2(n13247), .ZN(
        n14417) );
  AOI22_X2 U15010 ( .A1(FP_REG_FILE_reg_out_24__12_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__12_), .B2(n13226), .ZN(n4309) );
  AOI22_X2 U15011 ( .A1(FP_REG_FILE_reg_out_14__12_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__12_), .B2(n13230), .ZN(n14422) );
  NAND2_X2 U15012 ( .A1(FP_REG_FILE_reg_out_17__12_), .A2(n13235), .ZN(n14421)
         );
  NAND2_X2 U15013 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__12_), .ZN(n14420)
         );
  NAND2_X2 U15014 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__12_), .ZN(n14419)
         );
  NAND4_X2 U15015 ( .A1(n14422), .A2(n14421), .A3(n14420), .A4(n14419), .ZN(
        n4293) );
  AOI22_X2 U15016 ( .A1(FP_REG_FILE_reg_out_1__12_), .A2(n13243), .B1(
        FP_REG_FILE_reg_out_12__12_), .B2(n13241), .ZN(n14426) );
  NAND2_X2 U15017 ( .A1(n14426), .A2(n14425), .ZN(n4294) );
  OAI22_X2 U15018 ( .A1(n11376), .A2(n13249), .B1(n10411), .B2(n13246), .ZN(
        n14428) );
  AOI22_X2 U15019 ( .A1(FP_REG_FILE_reg_out_24__13_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__13_), .B2(n13226), .ZN(n4280) );
  AOI22_X2 U15020 ( .A1(FP_REG_FILE_reg_out_14__13_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__13_), .B2(n13230), .ZN(n14433) );
  NAND2_X2 U15021 ( .A1(FP_REG_FILE_reg_out_17__13_), .A2(n13235), .ZN(n14432)
         );
  NAND2_X2 U15022 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__13_), .ZN(n14431)
         );
  NAND2_X2 U15023 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__13_), .ZN(n14430)
         );
  NAND4_X2 U15024 ( .A1(n14433), .A2(n14432), .A3(n14431), .A4(n14430), .ZN(
        n4264) );
  AOI22_X2 U15025 ( .A1(FP_REG_FILE_reg_out_1__13_), .A2(n13243), .B1(
        FP_REG_FILE_reg_out_12__13_), .B2(n13241), .ZN(n14437) );
  NAND2_X2 U15026 ( .A1(n14437), .A2(n14436), .ZN(n4265) );
  OAI22_X2 U15027 ( .A1(n11377), .A2(n13249), .B1(n10412), .B2(n13247), .ZN(
        n14439) );
  AOI22_X2 U15028 ( .A1(FP_REG_FILE_reg_out_24__14_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__14_), .B2(n13226), .ZN(n4251) );
  AOI22_X2 U15029 ( .A1(FP_REG_FILE_reg_out_14__14_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__14_), .B2(n13230), .ZN(n14444) );
  NAND2_X2 U15030 ( .A1(FP_REG_FILE_reg_out_17__14_), .A2(n13235), .ZN(n14443)
         );
  NAND2_X2 U15031 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__14_), .ZN(n14442)
         );
  NAND2_X2 U15032 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__14_), .ZN(n14441)
         );
  NAND4_X2 U15033 ( .A1(n14444), .A2(n14443), .A3(n14442), .A4(n14441), .ZN(
        n4235) );
  AOI22_X2 U15034 ( .A1(FP_REG_FILE_reg_out_1__14_), .A2(n13243), .B1(
        FP_REG_FILE_reg_out_12__14_), .B2(n13241), .ZN(n14448) );
  NAND2_X2 U15035 ( .A1(n14448), .A2(n14447), .ZN(n4236) );
  OAI22_X2 U15036 ( .A1(n11378), .A2(n13249), .B1(n10413), .B2(n13246), .ZN(
        n14450) );
  AOI22_X2 U15037 ( .A1(FP_REG_FILE_reg_out_24__15_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__15_), .B2(n13226), .ZN(n4222) );
  AOI22_X2 U15038 ( .A1(FP_REG_FILE_reg_out_14__15_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__15_), .B2(n13230), .ZN(n14455) );
  NAND2_X2 U15039 ( .A1(FP_REG_FILE_reg_out_17__15_), .A2(n13235), .ZN(n14454)
         );
  NAND2_X2 U15040 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__15_), .ZN(n14453)
         );
  NAND2_X2 U15041 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__15_), .ZN(n14452)
         );
  NAND4_X2 U15042 ( .A1(n14455), .A2(n14454), .A3(n14453), .A4(n14452), .ZN(
        n4206) );
  AOI22_X2 U15043 ( .A1(FP_REG_FILE_reg_out_1__15_), .A2(n13243), .B1(
        FP_REG_FILE_reg_out_12__15_), .B2(n13241), .ZN(n14459) );
  NAND2_X2 U15044 ( .A1(n14459), .A2(n14458), .ZN(n4207) );
  OAI22_X2 U15045 ( .A1(n11379), .A2(n13249), .B1(n10414), .B2(n13247), .ZN(
        n14461) );
  AOI22_X2 U15046 ( .A1(FP_REG_FILE_reg_out_24__16_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__16_), .B2(n13226), .ZN(n4192) );
  AOI22_X2 U15047 ( .A1(FP_REG_FILE_reg_out_14__16_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__16_), .B2(n13230), .ZN(n14466) );
  NAND2_X2 U15048 ( .A1(FP_REG_FILE_reg_out_17__16_), .A2(n13235), .ZN(n14465)
         );
  NAND2_X2 U15049 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__16_), .ZN(n14464)
         );
  NAND2_X2 U15050 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__16_), .ZN(n14463)
         );
  NAND4_X2 U15051 ( .A1(n14466), .A2(n14465), .A3(n14464), .A4(n14463), .ZN(
        n4176) );
  AOI22_X2 U15052 ( .A1(FP_REG_FILE_reg_out_1__16_), .A2(n13243), .B1(
        FP_REG_FILE_reg_out_12__16_), .B2(n13241), .ZN(n14470) );
  NAND2_X2 U15053 ( .A1(n14470), .A2(n14469), .ZN(n4177) );
  OAI22_X2 U15054 ( .A1(n11380), .A2(n13249), .B1(n10415), .B2(n13246), .ZN(
        n14472) );
  AOI22_X2 U15055 ( .A1(FP_REG_FILE_reg_out_24__17_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__17_), .B2(n13226), .ZN(n4163) );
  AOI22_X2 U15056 ( .A1(FP_REG_FILE_reg_out_14__17_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__17_), .B2(n13230), .ZN(n14477) );
  NAND2_X2 U15057 ( .A1(FP_REG_FILE_reg_out_17__17_), .A2(n13235), .ZN(n14476)
         );
  NAND2_X2 U15058 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__17_), .ZN(n14475)
         );
  NAND2_X2 U15059 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__17_), .ZN(n14474)
         );
  NAND4_X2 U15060 ( .A1(n14477), .A2(n14476), .A3(n14475), .A4(n14474), .ZN(
        n4147) );
  AOI22_X2 U15061 ( .A1(FP_REG_FILE_reg_out_1__17_), .A2(n13243), .B1(
        FP_REG_FILE_reg_out_12__17_), .B2(n13241), .ZN(n14481) );
  NAND2_X2 U15062 ( .A1(n14481), .A2(n14480), .ZN(n4148) );
  OAI22_X2 U15063 ( .A1(n11381), .A2(n13249), .B1(n10416), .B2(n13247), .ZN(
        n14483) );
  AOI22_X2 U15064 ( .A1(FP_REG_FILE_reg_out_24__18_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__18_), .B2(n13226), .ZN(n4134) );
  AOI22_X2 U15065 ( .A1(FP_REG_FILE_reg_out_14__18_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__18_), .B2(n13230), .ZN(n14488) );
  NAND2_X2 U15066 ( .A1(FP_REG_FILE_reg_out_17__18_), .A2(n13235), .ZN(n14487)
         );
  NAND2_X2 U15067 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__18_), .ZN(n14486)
         );
  NAND2_X2 U15068 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__18_), .ZN(n14485)
         );
  NAND4_X2 U15069 ( .A1(n14488), .A2(n14487), .A3(n14486), .A4(n14485), .ZN(
        n4118) );
  AOI22_X2 U15070 ( .A1(FP_REG_FILE_reg_out_1__18_), .A2(n13243), .B1(
        FP_REG_FILE_reg_out_12__18_), .B2(n13241), .ZN(n14492) );
  NAND2_X2 U15071 ( .A1(n14492), .A2(n14491), .ZN(n4119) );
  OAI22_X2 U15072 ( .A1(n11382), .A2(n13249), .B1(n10417), .B2(n13246), .ZN(
        n14494) );
  AOI22_X2 U15073 ( .A1(FP_REG_FILE_reg_out_24__19_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__19_), .B2(n13226), .ZN(n4105) );
  AOI22_X2 U15074 ( .A1(FP_REG_FILE_reg_out_14__19_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__19_), .B2(n13230), .ZN(n14499) );
  NAND2_X2 U15075 ( .A1(FP_REG_FILE_reg_out_17__19_), .A2(n13235), .ZN(n14498)
         );
  NAND2_X2 U15076 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__19_), .ZN(n14497)
         );
  NAND2_X2 U15077 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__19_), .ZN(n14496)
         );
  NAND4_X2 U15078 ( .A1(n14499), .A2(n14498), .A3(n14497), .A4(n14496), .ZN(
        n4089) );
  AOI22_X2 U15079 ( .A1(FP_REG_FILE_reg_out_1__19_), .A2(n13243), .B1(
        FP_REG_FILE_reg_out_12__19_), .B2(n13241), .ZN(n14503) );
  NAND2_X2 U15080 ( .A1(n14503), .A2(n14502), .ZN(n4090) );
  OAI22_X2 U15081 ( .A1(n11383), .A2(n13249), .B1(n10418), .B2(n13247), .ZN(
        n14505) );
  AOI22_X2 U15082 ( .A1(FP_REG_FILE_reg_out_24__20_), .A2(n13229), .B1(
        FP_REG_FILE_reg_out_23__20_), .B2(n13226), .ZN(n4076) );
  AOI22_X2 U15083 ( .A1(FP_REG_FILE_reg_out_14__20_), .A2(n13233), .B1(
        FP_REG_FILE_reg_out_13__20_), .B2(n13230), .ZN(n14510) );
  NAND2_X2 U15084 ( .A1(FP_REG_FILE_reg_out_17__20_), .A2(n13235), .ZN(n14509)
         );
  NAND2_X2 U15085 ( .A1(n13237), .A2(FP_REG_FILE_reg_out_0__20_), .ZN(n14508)
         );
  NAND2_X2 U15086 ( .A1(n13239), .A2(FP_REG_FILE_reg_out_10__20_), .ZN(n14507)
         );
  NAND4_X2 U15087 ( .A1(n14510), .A2(n14509), .A3(n14508), .A4(n14507), .ZN(
        n4060) );
  AOI22_X2 U15088 ( .A1(FP_REG_FILE_reg_out_1__20_), .A2(n13243), .B1(
        FP_REG_FILE_reg_out_12__20_), .B2(n13241), .ZN(n14514) );
  NAND2_X2 U15089 ( .A1(n14514), .A2(n14513), .ZN(n4061) );
  OAI22_X2 U15090 ( .A1(n11384), .A2(n13249), .B1(n10419), .B2(n13246), .ZN(
        n14516) );
  AOI22_X2 U15091 ( .A1(FP_REG_FILE_reg_out_24__21_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__21_), .B2(n13227), .ZN(n4047) );
  AOI22_X2 U15092 ( .A1(FP_REG_FILE_reg_out_14__21_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__21_), .B2(n13231), .ZN(n14521) );
  NAND2_X2 U15093 ( .A1(FP_REG_FILE_reg_out_17__21_), .A2(n13234), .ZN(n14520)
         );
  NAND2_X2 U15094 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__21_), .ZN(n14519)
         );
  NAND2_X2 U15095 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__21_), .ZN(n14518)
         );
  NAND4_X2 U15096 ( .A1(n14521), .A2(n14520), .A3(n14519), .A4(n14518), .ZN(
        n4031) );
  AOI22_X2 U15097 ( .A1(FP_REG_FILE_reg_out_1__21_), .A2(n13242), .B1(
        FP_REG_FILE_reg_out_12__21_), .B2(n13240), .ZN(n14525) );
  NAND2_X2 U15098 ( .A1(n14525), .A2(n14524), .ZN(n4032) );
  OAI22_X2 U15099 ( .A1(n11385), .A2(n13249), .B1(n10420), .B2(n13247), .ZN(
        n14527) );
  AOI22_X2 U15100 ( .A1(FP_REG_FILE_reg_out_24__22_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__22_), .B2(n13226), .ZN(n4018) );
  AOI22_X2 U15101 ( .A1(FP_REG_FILE_reg_out_14__22_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__22_), .B2(n13230), .ZN(n14532) );
  NAND2_X2 U15102 ( .A1(FP_REG_FILE_reg_out_17__22_), .A2(n13234), .ZN(n14531)
         );
  NAND2_X2 U15103 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__22_), .ZN(n14530)
         );
  NAND2_X2 U15104 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__22_), .ZN(n14529)
         );
  NAND4_X2 U15105 ( .A1(n14532), .A2(n14531), .A3(n14530), .A4(n14529), .ZN(
        n4002) );
  AOI22_X2 U15106 ( .A1(FP_REG_FILE_reg_out_1__22_), .A2(n13242), .B1(
        FP_REG_FILE_reg_out_12__22_), .B2(n13240), .ZN(n14536) );
  NAND2_X2 U15107 ( .A1(n14536), .A2(n14535), .ZN(n4003) );
  OAI22_X2 U15108 ( .A1(n11386), .A2(n13249), .B1(n10421), .B2(n13247), .ZN(
        n14538) );
  AOI22_X2 U15109 ( .A1(FP_REG_FILE_reg_out_24__23_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__23_), .B2(n13227), .ZN(n3989) );
  AOI22_X2 U15110 ( .A1(FP_REG_FILE_reg_out_14__23_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__23_), .B2(n13231), .ZN(n14543) );
  NAND2_X2 U15111 ( .A1(FP_REG_FILE_reg_out_17__23_), .A2(n13234), .ZN(n14542)
         );
  NAND2_X2 U15112 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__23_), .ZN(n14541)
         );
  NAND2_X2 U15113 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__23_), .ZN(n14540)
         );
  NAND4_X2 U15114 ( .A1(n14543), .A2(n14542), .A3(n14541), .A4(n14540), .ZN(
        n3973) );
  AOI22_X2 U15115 ( .A1(FP_REG_FILE_reg_out_1__23_), .A2(n13242), .B1(
        FP_REG_FILE_reg_out_12__23_), .B2(n13240), .ZN(n14547) );
  NAND2_X2 U15116 ( .A1(n14547), .A2(n14546), .ZN(n3974) );
  OAI22_X2 U15117 ( .A1(n11387), .A2(n13248), .B1(n10422), .B2(n13247), .ZN(
        n14549) );
  AOI22_X2 U15118 ( .A1(FP_REG_FILE_reg_out_24__24_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__24_), .B2(n13226), .ZN(n3960) );
  AOI22_X2 U15119 ( .A1(FP_REG_FILE_reg_out_14__24_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__24_), .B2(n13230), .ZN(n14554) );
  NAND2_X2 U15120 ( .A1(FP_REG_FILE_reg_out_17__24_), .A2(n13234), .ZN(n14553)
         );
  NAND2_X2 U15121 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__24_), .ZN(n14552)
         );
  NAND2_X2 U15122 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__24_), .ZN(n14551)
         );
  NAND4_X2 U15123 ( .A1(n14554), .A2(n14553), .A3(n14552), .A4(n14551), .ZN(
        n3944) );
  AOI22_X2 U15124 ( .A1(FP_REG_FILE_reg_out_1__24_), .A2(n13242), .B1(
        FP_REG_FILE_reg_out_12__24_), .B2(n13240), .ZN(n14558) );
  NAND2_X2 U15125 ( .A1(n14558), .A2(n14557), .ZN(n3945) );
  OAI22_X2 U15126 ( .A1(n11388), .A2(n13249), .B1(n10423), .B2(n13247), .ZN(
        n14560) );
  AOI22_X2 U15127 ( .A1(FP_REG_FILE_reg_out_24__25_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__25_), .B2(n13227), .ZN(n3931) );
  AOI22_X2 U15128 ( .A1(FP_REG_FILE_reg_out_14__25_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__25_), .B2(n13231), .ZN(n14565) );
  NAND2_X2 U15129 ( .A1(FP_REG_FILE_reg_out_17__25_), .A2(n13234), .ZN(n14564)
         );
  NAND2_X2 U15130 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__25_), .ZN(n14563)
         );
  NAND2_X2 U15131 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__25_), .ZN(n14562)
         );
  NAND4_X2 U15132 ( .A1(n14565), .A2(n14564), .A3(n14563), .A4(n14562), .ZN(
        n3915) );
  AOI22_X2 U15133 ( .A1(FP_REG_FILE_reg_out_1__25_), .A2(n13242), .B1(
        FP_REG_FILE_reg_out_12__25_), .B2(n13240), .ZN(n14569) );
  NAND2_X2 U15134 ( .A1(n14569), .A2(n14568), .ZN(n3916) );
  OAI22_X2 U15135 ( .A1(n11389), .A2(n13248), .B1(n10424), .B2(n13247), .ZN(
        n14571) );
  AOI22_X2 U15136 ( .A1(FP_REG_FILE_reg_out_24__26_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__26_), .B2(n13226), .ZN(n3901) );
  AOI22_X2 U15137 ( .A1(FP_REG_FILE_reg_out_14__26_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__26_), .B2(n13230), .ZN(n14576) );
  NAND2_X2 U15138 ( .A1(FP_REG_FILE_reg_out_17__26_), .A2(n13234), .ZN(n14575)
         );
  NAND2_X2 U15139 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__26_), .ZN(n14574)
         );
  NAND2_X2 U15140 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__26_), .ZN(n14573)
         );
  NAND4_X2 U15141 ( .A1(n14576), .A2(n14575), .A3(n14574), .A4(n14573), .ZN(
        n3885) );
  AOI22_X2 U15142 ( .A1(FP_REG_FILE_reg_out_1__26_), .A2(n13242), .B1(
        FP_REG_FILE_reg_out_12__26_), .B2(n13240), .ZN(n14580) );
  NAND2_X2 U15143 ( .A1(n14580), .A2(n14579), .ZN(n3886) );
  OAI22_X2 U15144 ( .A1(n11390), .A2(n13249), .B1(n10425), .B2(n13247), .ZN(
        n14582) );
  AOI22_X2 U15145 ( .A1(FP_REG_FILE_reg_out_24__27_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__27_), .B2(n13227), .ZN(n3872) );
  AOI22_X2 U15146 ( .A1(FP_REG_FILE_reg_out_14__27_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__27_), .B2(n13231), .ZN(n14587) );
  NAND2_X2 U15147 ( .A1(FP_REG_FILE_reg_out_17__27_), .A2(n13234), .ZN(n14586)
         );
  NAND2_X2 U15148 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__27_), .ZN(n14585)
         );
  NAND2_X2 U15149 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__27_), .ZN(n14584)
         );
  NAND4_X2 U15150 ( .A1(n14587), .A2(n14586), .A3(n14585), .A4(n14584), .ZN(
        n3856) );
  AOI22_X2 U15151 ( .A1(FP_REG_FILE_reg_out_1__27_), .A2(n13242), .B1(
        FP_REG_FILE_reg_out_12__27_), .B2(n13240), .ZN(n14591) );
  NAND2_X2 U15152 ( .A1(n14591), .A2(n14590), .ZN(n3857) );
  OAI22_X2 U15153 ( .A1(n11391), .A2(n13248), .B1(n10426), .B2(n13247), .ZN(
        n14593) );
  AOI22_X2 U15154 ( .A1(FP_REG_FILE_reg_out_24__28_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__28_), .B2(n13226), .ZN(n3843) );
  AOI22_X2 U15155 ( .A1(FP_REG_FILE_reg_out_14__28_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__28_), .B2(n13230), .ZN(n14598) );
  NAND2_X2 U15156 ( .A1(FP_REG_FILE_reg_out_17__28_), .A2(n13234), .ZN(n14597)
         );
  NAND2_X2 U15157 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__28_), .ZN(n14596)
         );
  NAND2_X2 U15158 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__28_), .ZN(n14595)
         );
  NAND4_X2 U15159 ( .A1(n14598), .A2(n14597), .A3(n14596), .A4(n14595), .ZN(
        n3827) );
  AOI22_X2 U15160 ( .A1(FP_REG_FILE_reg_out_1__28_), .A2(n13242), .B1(
        FP_REG_FILE_reg_out_12__28_), .B2(n13240), .ZN(n14602) );
  NAND2_X2 U15161 ( .A1(n14602), .A2(n14601), .ZN(n3828) );
  OAI22_X2 U15162 ( .A1(n11392), .A2(n13249), .B1(n10427), .B2(n13247), .ZN(
        n14604) );
  AOI22_X2 U15163 ( .A1(FP_REG_FILE_reg_out_24__29_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__29_), .B2(n13227), .ZN(n3814) );
  AOI22_X2 U15164 ( .A1(FP_REG_FILE_reg_out_14__29_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__29_), .B2(n13231), .ZN(n14609) );
  NAND2_X2 U15165 ( .A1(FP_REG_FILE_reg_out_17__29_), .A2(n13234), .ZN(n14608)
         );
  NAND2_X2 U15166 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__29_), .ZN(n14607)
         );
  NAND2_X2 U15167 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__29_), .ZN(n14606)
         );
  NAND4_X2 U15168 ( .A1(n14609), .A2(n14608), .A3(n14607), .A4(n14606), .ZN(
        n3798) );
  AOI22_X2 U15169 ( .A1(FP_REG_FILE_reg_out_1__29_), .A2(n13242), .B1(
        FP_REG_FILE_reg_out_12__29_), .B2(n13240), .ZN(n14613) );
  NAND2_X2 U15170 ( .A1(n14613), .A2(n14612), .ZN(n3799) );
  OAI22_X2 U15171 ( .A1(n11393), .A2(n13248), .B1(n10428), .B2(n13247), .ZN(
        n14615) );
  AOI22_X2 U15172 ( .A1(FP_REG_FILE_reg_out_24__30_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__30_), .B2(n13226), .ZN(n3785) );
  AOI22_X2 U15173 ( .A1(FP_REG_FILE_reg_out_14__30_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__30_), .B2(n13230), .ZN(n14620) );
  NAND2_X2 U15174 ( .A1(FP_REG_FILE_reg_out_17__30_), .A2(n13234), .ZN(n14619)
         );
  NAND2_X2 U15175 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__30_), .ZN(n14618)
         );
  NAND2_X2 U15176 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__30_), .ZN(n14617)
         );
  NAND4_X2 U15177 ( .A1(n14620), .A2(n14619), .A3(n14618), .A4(n14617), .ZN(
        n3769) );
  AOI22_X2 U15178 ( .A1(FP_REG_FILE_reg_out_1__30_), .A2(n13242), .B1(
        FP_REG_FILE_reg_out_12__30_), .B2(n13240), .ZN(n14624) );
  NAND2_X2 U15179 ( .A1(n14624), .A2(n14623), .ZN(n3770) );
  OAI22_X2 U15180 ( .A1(n11395), .A2(n13249), .B1(n10429), .B2(n13247), .ZN(
        n14626) );
  AOI22_X2 U15181 ( .A1(FP_REG_FILE_reg_out_24__31_), .A2(n13228), .B1(
        FP_REG_FILE_reg_out_23__31_), .B2(n13227), .ZN(n3743) );
  AOI22_X2 U15182 ( .A1(FP_REG_FILE_reg_out_14__31_), .A2(n13232), .B1(
        FP_REG_FILE_reg_out_13__31_), .B2(n13231), .ZN(n14631) );
  NAND2_X2 U15183 ( .A1(FP_REG_FILE_reg_out_17__31_), .A2(n13234), .ZN(n14630)
         );
  NAND2_X2 U15184 ( .A1(n13236), .A2(FP_REG_FILE_reg_out_0__31_), .ZN(n14629)
         );
  NAND2_X2 U15185 ( .A1(n13238), .A2(FP_REG_FILE_reg_out_10__31_), .ZN(n14628)
         );
  NAND4_X2 U15186 ( .A1(n14631), .A2(n14630), .A3(n14629), .A4(n14628), .ZN(
        n3708) );
  AOI22_X2 U15187 ( .A1(FP_REG_FILE_reg_out_1__31_), .A2(n13242), .B1(
        FP_REG_FILE_reg_out_12__31_), .B2(n13240), .ZN(n14637) );
  NAND2_X2 U15188 ( .A1(n14637), .A2(n14636), .ZN(n3709) );
  OAI22_X2 U15189 ( .A1(n11396), .A2(n13248), .B1(n10430), .B2(n13247), .ZN(
        n14639) );
  NAND2_X2 U15191 ( .A1(net230393), .A2(offset_26_id[6]), .ZN(n18752) );
  INV_X4 U15192 ( .A(n18752), .ZN(n14644) );
  INV_X4 U15193 ( .A(n14641), .ZN(n15608) );
  NAND2_X2 U15194 ( .A1(net230393), .A2(n11922), .ZN(n14642) );
  INV_X4 U15195 ( .A(n14642), .ZN(n14647) );
  INV_X4 U15196 ( .A(n10824), .ZN(n18813) );
  NAND2_X2 U15197 ( .A1(n14647), .A2(n18813), .ZN(n14643) );
  INV_X4 U15198 ( .A(n14643), .ZN(n19162) );
  INV_X4 U15199 ( .A(n14645), .ZN(n15616) );
  INV_X4 U15200 ( .A(n14649), .ZN(n15609) );
  OAI221_X2 U15201 ( .B1(n12321), .B2(n13254), .C1(n10650), .C2(n13708), .A(
        n14652), .ZN(n3685) );
  NAND2_X2 U15202 ( .A1(n10161), .A2(n15603), .ZN(n14968) );
  INV_X4 U15203 ( .A(n14656), .ZN(n15621) );
  NAND2_X2 U15204 ( .A1(n19162), .A2(n15621), .ZN(n14657) );
  NAND2_X2 U15205 ( .A1(n10160), .A2(n15621), .ZN(n14658) );
  NAND2_X2 U15206 ( .A1(n10161), .A2(n15621), .ZN(n14659) );
  INV_X4 U15207 ( .A(n14659), .ZN(n19161) );
  NAND2_X2 U15208 ( .A1(FP_REG_FILE_reg_out_11__0_), .A2(n13264), .ZN(n14663)
         );
  NAND2_X2 U15209 ( .A1(FP_REG_FILE_reg_out_25__0_), .A2(n13262), .ZN(n14662)
         );
  NAND2_X2 U15210 ( .A1(n14760), .A2(FP_REG_FILE_reg_out_24__0_), .ZN(n14661)
         );
  NAND2_X2 U15211 ( .A1(n10352), .A2(FP_REG_FILE_reg_out_18__0_), .ZN(n14660)
         );
  NAND4_X2 U15212 ( .A1(n14663), .A2(n14662), .A3(n14661), .A4(n14660), .ZN(
        n3659) );
  OAI221_X2 U15213 ( .B1(n12322), .B2(n13254), .C1(n12271), .C2(n13708), .A(
        n14666), .ZN(n3640) );
  NAND2_X2 U15214 ( .A1(FP_REG_FILE_reg_out_11__1_), .A2(n13265), .ZN(n14673)
         );
  NAND2_X2 U15215 ( .A1(FP_REG_FILE_reg_out_25__1_), .A2(n13263), .ZN(n14672)
         );
  NAND2_X2 U15216 ( .A1(n14760), .A2(FP_REG_FILE_reg_out_24__1_), .ZN(n14671)
         );
  NAND2_X2 U15217 ( .A1(n10352), .A2(FP_REG_FILE_reg_out_18__1_), .ZN(n14670)
         );
  NAND4_X2 U15218 ( .A1(n14673), .A2(n14672), .A3(n14671), .A4(n14670), .ZN(
        n3625) );
  OAI221_X2 U15219 ( .B1(n12323), .B2(n13254), .C1(n10665), .C2(n13708), .A(
        n14676), .ZN(n3606) );
  NAND2_X2 U15220 ( .A1(FP_REG_FILE_reg_out_11__2_), .A2(n13264), .ZN(n14683)
         );
  NAND2_X2 U15221 ( .A1(FP_REG_FILE_reg_out_25__2_), .A2(n13262), .ZN(n14682)
         );
  NAND2_X2 U15222 ( .A1(n14760), .A2(FP_REG_FILE_reg_out_24__2_), .ZN(n14681)
         );
  NAND2_X2 U15223 ( .A1(n10352), .A2(FP_REG_FILE_reg_out_18__2_), .ZN(n14680)
         );
  NAND4_X2 U15224 ( .A1(n14683), .A2(n14682), .A3(n14681), .A4(n14680), .ZN(
        n3591) );
  OAI221_X2 U15225 ( .B1(n12324), .B2(n13254), .C1(n10666), .C2(n13708), .A(
        n14686), .ZN(n3572) );
  NAND2_X2 U15226 ( .A1(FP_REG_FILE_reg_out_11__3_), .A2(n13265), .ZN(n14693)
         );
  NAND2_X2 U15227 ( .A1(FP_REG_FILE_reg_out_25__3_), .A2(n13263), .ZN(n14692)
         );
  NAND2_X2 U15228 ( .A1(n14760), .A2(FP_REG_FILE_reg_out_24__3_), .ZN(n14691)
         );
  NAND2_X2 U15229 ( .A1(n10352), .A2(FP_REG_FILE_reg_out_18__3_), .ZN(n14690)
         );
  NAND4_X2 U15230 ( .A1(n14693), .A2(n14692), .A3(n14691), .A4(n14690), .ZN(
        n3557) );
  OAI221_X2 U15231 ( .B1(n12325), .B2(n13254), .C1(n10667), .C2(n13708), .A(
        n14696), .ZN(n3537) );
  NAND2_X2 U15232 ( .A1(FP_REG_FILE_reg_out_11__4_), .A2(n13264), .ZN(n14703)
         );
  NAND2_X2 U15233 ( .A1(FP_REG_FILE_reg_out_25__4_), .A2(n13262), .ZN(n14702)
         );
  NAND2_X2 U15234 ( .A1(n14760), .A2(FP_REG_FILE_reg_out_24__4_), .ZN(n14701)
         );
  NAND2_X2 U15235 ( .A1(n10352), .A2(FP_REG_FILE_reg_out_18__4_), .ZN(n14700)
         );
  NAND4_X2 U15236 ( .A1(n14703), .A2(n14702), .A3(n14701), .A4(n14700), .ZN(
        n3522) );
  OAI221_X2 U15237 ( .B1(n12326), .B2(n13254), .C1(n10668), .C2(n13708), .A(
        n14706), .ZN(n3503) );
  NAND2_X2 U15238 ( .A1(FP_REG_FILE_reg_out_11__5_), .A2(n13265), .ZN(n14713)
         );
  NAND2_X2 U15239 ( .A1(FP_REG_FILE_reg_out_25__5_), .A2(n13263), .ZN(n14712)
         );
  NAND2_X2 U15240 ( .A1(n14760), .A2(FP_REG_FILE_reg_out_24__5_), .ZN(n14711)
         );
  NAND2_X2 U15241 ( .A1(n10352), .A2(FP_REG_FILE_reg_out_18__5_), .ZN(n14710)
         );
  NAND4_X2 U15242 ( .A1(n14713), .A2(n14712), .A3(n14711), .A4(n14710), .ZN(
        n3488) );
  OAI221_X2 U15243 ( .B1(n12327), .B2(n13254), .C1(n10669), .C2(n13708), .A(
        n14716), .ZN(n3469) );
  NAND2_X2 U15244 ( .A1(FP_REG_FILE_reg_out_11__6_), .A2(n13264), .ZN(n14723)
         );
  NAND2_X2 U15245 ( .A1(FP_REG_FILE_reg_out_25__6_), .A2(n13262), .ZN(n14722)
         );
  NAND2_X2 U15246 ( .A1(n14760), .A2(FP_REG_FILE_reg_out_24__6_), .ZN(n14721)
         );
  NAND2_X2 U15247 ( .A1(n10352), .A2(FP_REG_FILE_reg_out_18__6_), .ZN(n14720)
         );
  NAND4_X2 U15248 ( .A1(n14723), .A2(n14722), .A3(n14721), .A4(n14720), .ZN(
        n3454) );
  OAI221_X2 U15249 ( .B1(n12328), .B2(n13254), .C1(n10670), .C2(n13708), .A(
        n14726), .ZN(n3435) );
  NAND2_X2 U15250 ( .A1(FP_REG_FILE_reg_out_11__7_), .A2(n13265), .ZN(n14733)
         );
  NAND2_X2 U15251 ( .A1(FP_REG_FILE_reg_out_25__7_), .A2(n13263), .ZN(n14732)
         );
  NAND2_X2 U15252 ( .A1(n14760), .A2(FP_REG_FILE_reg_out_24__7_), .ZN(n14731)
         );
  NAND2_X2 U15253 ( .A1(n10352), .A2(FP_REG_FILE_reg_out_18__7_), .ZN(n14730)
         );
  NAND4_X2 U15254 ( .A1(n14733), .A2(n14732), .A3(n14731), .A4(n14730), .ZN(
        n3420) );
  OAI221_X2 U15255 ( .B1(n12329), .B2(n13254), .C1(n10671), .C2(n13708), .A(
        n14736), .ZN(n3401) );
  NAND2_X2 U15256 ( .A1(FP_REG_FILE_reg_out_11__8_), .A2(n13264), .ZN(n14743)
         );
  NAND2_X2 U15257 ( .A1(FP_REG_FILE_reg_out_25__8_), .A2(n13262), .ZN(n14742)
         );
  NAND2_X2 U15258 ( .A1(n14760), .A2(FP_REG_FILE_reg_out_24__8_), .ZN(n14741)
         );
  NAND2_X2 U15259 ( .A1(n10352), .A2(FP_REG_FILE_reg_out_18__8_), .ZN(n14740)
         );
  NAND4_X2 U15260 ( .A1(n14743), .A2(n14742), .A3(n14741), .A4(n14740), .ZN(
        n3386) );
  OAI221_X2 U15261 ( .B1(n12330), .B2(n13254), .C1(n10672), .C2(n13708), .A(
        n14746), .ZN(n3367) );
  NAND2_X2 U15262 ( .A1(FP_REG_FILE_reg_out_11__9_), .A2(n13265), .ZN(n14753)
         );
  NAND2_X2 U15263 ( .A1(FP_REG_FILE_reg_out_25__9_), .A2(n13263), .ZN(n14752)
         );
  NAND2_X2 U15264 ( .A1(n14760), .A2(FP_REG_FILE_reg_out_24__9_), .ZN(n14751)
         );
  NAND2_X2 U15265 ( .A1(n10352), .A2(FP_REG_FILE_reg_out_18__9_), .ZN(n14750)
         );
  NAND4_X2 U15266 ( .A1(n14753), .A2(n14752), .A3(n14751), .A4(n14750), .ZN(
        n3352) );
  OAI221_X2 U15267 ( .B1(n12331), .B2(n13254), .C1(n10651), .C2(n13708), .A(
        n14756), .ZN(n3333) );
  NAND2_X2 U15268 ( .A1(FP_REG_FILE_reg_out_11__10_), .A2(n13265), .ZN(n14764)
         );
  NAND2_X2 U15269 ( .A1(FP_REG_FILE_reg_out_25__10_), .A2(n13263), .ZN(n14763)
         );
  NAND2_X2 U15270 ( .A1(n14760), .A2(FP_REG_FILE_reg_out_24__10_), .ZN(n14762)
         );
  NAND2_X2 U15271 ( .A1(n10352), .A2(FP_REG_FILE_reg_out_18__10_), .ZN(n14761)
         );
  NAND4_X2 U15272 ( .A1(n14764), .A2(n14763), .A3(n14762), .A4(n14761), .ZN(
        n3318) );
  OAI221_X2 U15273 ( .B1(n12332), .B2(n13255), .C1(n10652), .C2(n13709), .A(
        n14767), .ZN(n3299) );
  AOI22_X2 U15274 ( .A1(FP_REG_FILE_reg_out_11__11_), .A2(n13265), .B1(
        FP_REG_FILE_reg_out_25__11_), .B2(n13263), .ZN(n14774) );
  NAND2_X2 U15275 ( .A1(n14774), .A2(n14773), .ZN(n3284) );
  OAI221_X2 U15276 ( .B1(n12333), .B2(n13255), .C1(n10653), .C2(n13708), .A(
        n14777), .ZN(n3265) );
  AOI22_X2 U15277 ( .A1(FP_REG_FILE_reg_out_11__12_), .A2(n13265), .B1(
        FP_REG_FILE_reg_out_25__12_), .B2(n13263), .ZN(n14784) );
  NAND2_X2 U15278 ( .A1(n14784), .A2(n14783), .ZN(n3250) );
  OAI221_X2 U15279 ( .B1(n12334), .B2(n13255), .C1(n10654), .C2(n13709), .A(
        n14787), .ZN(n3231) );
  AOI22_X2 U15280 ( .A1(FP_REG_FILE_reg_out_11__13_), .A2(n13265), .B1(
        FP_REG_FILE_reg_out_25__13_), .B2(n13263), .ZN(n14794) );
  NAND2_X2 U15281 ( .A1(n14794), .A2(n14793), .ZN(n3216) );
  OAI221_X2 U15282 ( .B1(n12335), .B2(n13255), .C1(n10655), .C2(n13708), .A(
        n14797), .ZN(n3196) );
  AOI22_X2 U15283 ( .A1(FP_REG_FILE_reg_out_11__14_), .A2(n13265), .B1(
        FP_REG_FILE_reg_out_25__14_), .B2(n13263), .ZN(n14804) );
  NAND2_X2 U15284 ( .A1(n14804), .A2(n14803), .ZN(n3181) );
  OAI221_X2 U15285 ( .B1(n12336), .B2(n13255), .C1(n10656), .C2(n13709), .A(
        n14807), .ZN(n3162) );
  AOI22_X2 U15286 ( .A1(FP_REG_FILE_reg_out_11__15_), .A2(n13265), .B1(
        FP_REG_FILE_reg_out_25__15_), .B2(n13263), .ZN(n14814) );
  NAND2_X2 U15287 ( .A1(n14814), .A2(n14813), .ZN(n3147) );
  OAI221_X2 U15288 ( .B1(n12337), .B2(n13255), .C1(n10657), .C2(n13708), .A(
        n14817), .ZN(n3128) );
  AOI22_X2 U15289 ( .A1(FP_REG_FILE_reg_out_11__16_), .A2(n13265), .B1(
        FP_REG_FILE_reg_out_25__16_), .B2(n13263), .ZN(n14824) );
  NAND2_X2 U15290 ( .A1(n14824), .A2(n14823), .ZN(n3113) );
  OAI221_X2 U15291 ( .B1(n12338), .B2(n13255), .C1(n10658), .C2(n13709), .A(
        n14827), .ZN(n3094) );
  AOI22_X2 U15292 ( .A1(FP_REG_FILE_reg_out_11__17_), .A2(n13265), .B1(
        FP_REG_FILE_reg_out_25__17_), .B2(n13263), .ZN(n14834) );
  NAND2_X2 U15293 ( .A1(n14834), .A2(n14833), .ZN(n3079) );
  OAI221_X2 U15294 ( .B1(n12339), .B2(n13255), .C1(n10659), .C2(n13708), .A(
        n14837), .ZN(n3060) );
  AOI22_X2 U15295 ( .A1(FP_REG_FILE_reg_out_11__18_), .A2(n13265), .B1(
        FP_REG_FILE_reg_out_25__18_), .B2(n13263), .ZN(n14844) );
  NAND2_X2 U15296 ( .A1(n14844), .A2(n14843), .ZN(n3045) );
  OAI221_X2 U15297 ( .B1(n12340), .B2(n13255), .C1(n10660), .C2(n13709), .A(
        n14847), .ZN(n3026) );
  AOI22_X2 U15298 ( .A1(FP_REG_FILE_reg_out_11__19_), .A2(n13265), .B1(
        FP_REG_FILE_reg_out_25__19_), .B2(n13263), .ZN(n14854) );
  NAND2_X2 U15299 ( .A1(n14854), .A2(n14853), .ZN(n3011) );
  OAI221_X2 U15300 ( .B1(n12341), .B2(n13255), .C1(n10661), .C2(n13708), .A(
        n14857), .ZN(n2992) );
  AOI22_X2 U15301 ( .A1(FP_REG_FILE_reg_out_11__20_), .A2(n13265), .B1(
        FP_REG_FILE_reg_out_25__20_), .B2(n13263), .ZN(n14864) );
  NAND2_X2 U15302 ( .A1(n14864), .A2(n14863), .ZN(n2977) );
  OAI221_X2 U15303 ( .B1(n12342), .B2(n13255), .C1(n10662), .C2(n13709), .A(
        n14867), .ZN(n2958) );
  AOI22_X2 U15304 ( .A1(FP_REG_FILE_reg_out_11__21_), .A2(n13264), .B1(
        FP_REG_FILE_reg_out_25__21_), .B2(n13262), .ZN(n14874) );
  NAND2_X2 U15305 ( .A1(n14874), .A2(n14873), .ZN(n2943) );
  OAI221_X2 U15306 ( .B1(n12343), .B2(n13255), .C1(n10663), .C2(n13709), .A(
        n14877), .ZN(n2924) );
  AOI22_X2 U15307 ( .A1(FP_REG_FILE_reg_out_11__22_), .A2(n13264), .B1(
        FP_REG_FILE_reg_out_25__22_), .B2(n13262), .ZN(n14884) );
  NAND2_X2 U15308 ( .A1(n14884), .A2(n14883), .ZN(n2909) );
  OAI221_X2 U15309 ( .B1(n12344), .B2(n13254), .C1(n10664), .C2(n13709), .A(
        n14887), .ZN(n2890) );
  AOI22_X2 U15310 ( .A1(FP_REG_FILE_reg_out_11__23_), .A2(n13264), .B1(
        FP_REG_FILE_reg_out_25__23_), .B2(n13262), .ZN(n14894) );
  NAND2_X2 U15311 ( .A1(n14894), .A2(n14893), .ZN(n2875) );
  OAI221_X2 U15312 ( .B1(n11479), .B2(n13255), .C1(n11281), .C2(n13709), .A(
        n14897), .ZN(n2855) );
  AOI22_X2 U15313 ( .A1(FP_REG_FILE_reg_out_11__24_), .A2(n13264), .B1(
        FP_REG_FILE_reg_out_25__24_), .B2(n13262), .ZN(n14904) );
  NAND2_X2 U15314 ( .A1(n14904), .A2(n14903), .ZN(n2840) );
  OAI221_X2 U15315 ( .B1(n11480), .B2(n13254), .C1(n11282), .C2(n13709), .A(
        n14907), .ZN(n2821) );
  AOI22_X2 U15316 ( .A1(FP_REG_FILE_reg_out_11__25_), .A2(n13264), .B1(
        FP_REG_FILE_reg_out_25__25_), .B2(n13262), .ZN(n14914) );
  NAND2_X2 U15317 ( .A1(n14914), .A2(n14913), .ZN(n2806) );
  OAI221_X2 U15318 ( .B1(n11481), .B2(n13255), .C1(n11283), .C2(n13709), .A(
        n14917), .ZN(n2787) );
  AOI22_X2 U15319 ( .A1(FP_REG_FILE_reg_out_11__26_), .A2(n13264), .B1(
        FP_REG_FILE_reg_out_25__26_), .B2(n13262), .ZN(n14924) );
  NAND2_X2 U15320 ( .A1(n14924), .A2(n14923), .ZN(n2772) );
  OAI221_X2 U15321 ( .B1(n11482), .B2(n13254), .C1(n11284), .C2(n13709), .A(
        n14927), .ZN(n2753) );
  AOI22_X2 U15322 ( .A1(FP_REG_FILE_reg_out_11__27_), .A2(n13264), .B1(
        FP_REG_FILE_reg_out_25__27_), .B2(n13262), .ZN(n14934) );
  NAND2_X2 U15323 ( .A1(n14934), .A2(n14933), .ZN(n2738) );
  OAI221_X2 U15324 ( .B1(n11483), .B2(n13255), .C1(n11285), .C2(n13709), .A(
        n14937), .ZN(n2719) );
  AOI22_X2 U15325 ( .A1(FP_REG_FILE_reg_out_11__28_), .A2(n13264), .B1(
        FP_REG_FILE_reg_out_25__28_), .B2(n13262), .ZN(n14944) );
  NAND2_X2 U15326 ( .A1(n14944), .A2(n14943), .ZN(n2704) );
  OAI221_X2 U15327 ( .B1(n11484), .B2(n13254), .C1(n11286), .C2(n13709), .A(
        n14947), .ZN(n2685) );
  AOI22_X2 U15328 ( .A1(FP_REG_FILE_reg_out_11__29_), .A2(n13264), .B1(
        FP_REG_FILE_reg_out_25__29_), .B2(n13262), .ZN(n14954) );
  NAND2_X2 U15329 ( .A1(n14954), .A2(n14953), .ZN(n2670) );
  OAI221_X2 U15330 ( .B1(n11485), .B2(n13255), .C1(n11287), .C2(n13709), .A(
        n14957), .ZN(n2651) );
  AOI22_X2 U15331 ( .A1(FP_REG_FILE_reg_out_11__30_), .A2(n13264), .B1(
        FP_REG_FILE_reg_out_25__30_), .B2(n13262), .ZN(n14964) );
  NAND2_X2 U15332 ( .A1(n14964), .A2(n14963), .ZN(n2636) );
  OAI221_X2 U15333 ( .B1(n11486), .B2(n13254), .C1(n11288), .C2(n13709), .A(
        n14967), .ZN(n2602) );
  AOI22_X2 U15334 ( .A1(FP_REG_FILE_reg_out_11__31_), .A2(n13264), .B1(
        FP_REG_FILE_reg_out_25__31_), .B2(n13262), .ZN(n14976) );
  NAND2_X2 U15335 ( .A1(n14976), .A2(n14975), .ZN(n2570) );
  NAND2_X2 U15336 ( .A1(ID_STAGE_imm16_aluA[17]), .A2(net230387), .ZN(n2562)
         );
  NAND2_X2 U15337 ( .A1(ID_STAGE_imm16_aluA[19]), .A2(net230387), .ZN(n2557)
         );
  NAND2_X2 U15338 ( .A1(ID_STAGE_imm16_aluA[20]), .A2(net230387), .ZN(n2555)
         );
  NOR2_X4 U15340 ( .A1(n14977), .A2(n12539), .ZN(n14979) );
  NAND2_X2 U15341 ( .A1(n14979), .A2(n14978), .ZN(n2532) );
  NAND2_X2 U15342 ( .A1(n14990), .A2(n2511), .ZN(n14980) );
  INV_X4 U15343 ( .A(n14980), .ZN(n19158) );
  NAND2_X2 U15344 ( .A1(n14991), .A2(n2508), .ZN(n14981) );
  INV_X4 U15345 ( .A(n14981), .ZN(n19156) );
  NAND2_X2 U15346 ( .A1(n2506), .A2(n14998), .ZN(n15328) );
  OAI22_X2 U15347 ( .A1(n10325), .A2(n13181), .B1(n12721), .B2(n13266), .ZN(
        n2515) );
  NAND2_X2 U15348 ( .A1(n14982), .A2(n2508), .ZN(n2182) );
  NAND2_X2 U15349 ( .A1(n14995), .A2(n2503), .ZN(n15335) );
  NAND2_X2 U15350 ( .A1(n14986), .A2(n2508), .ZN(n15334) );
  NAND2_X2 U15351 ( .A1(n14990), .A2(n2508), .ZN(n1871) );
  NAND2_X2 U15352 ( .A1(n2503), .A2(n14998), .ZN(n15330) );
  NAND2_X2 U15353 ( .A1(n14986), .A2(n2503), .ZN(n15329) );
  INV_X4 U15354 ( .A(n2524), .ZN(n15005) );
  NAND2_X2 U15355 ( .A1(n2506), .A2(n14997), .ZN(n17769) );
  OAI22_X2 U15356 ( .A1(n13184), .A2(n11881), .B1(n13364), .B2(n12828), .ZN(
        n14994) );
  NAND2_X2 U15357 ( .A1(n14997), .A2(n2503), .ZN(n17776) );
  NAND2_X2 U15358 ( .A1(n14995), .A2(n2508), .ZN(n17774) );
  INV_X4 U15359 ( .A(n2532), .ZN(n14996) );
  OAI221_X2 U15360 ( .B1(n12413), .B2(n13382), .C1(n12786), .C2(n13377), .A(
        n12964), .ZN(n15002) );
  NAND2_X2 U15361 ( .A1(n2506), .A2(n14999), .ZN(n17775) );
  NAND2_X2 U15362 ( .A1(n2511), .A2(n14997), .ZN(n17771) );
  OAI22_X2 U15363 ( .A1(n13379), .A2(n12767), .B1(n13368), .B2(n11838), .ZN(
        n15001) );
  NAND2_X2 U15364 ( .A1(n2508), .A2(n14998), .ZN(n17773) );
  NAND2_X2 U15365 ( .A1(n2503), .A2(n14999), .ZN(n17772) );
  OAI22_X2 U15366 ( .A1(n11847), .A2(n13373), .B1(n10861), .B2(n13371), .ZN(
        n15000) );
  NAND4_X2 U15367 ( .A1(n15006), .A2(n15005), .A3(n15004), .A4(n15003), .ZN(
        n2498) );
  OAI22_X2 U15368 ( .A1(n10338), .A2(n13181), .B1(n12735), .B2(n13266), .ZN(
        n2486) );
  INV_X4 U15369 ( .A(n2493), .ZN(n15021) );
  OAI22_X2 U15370 ( .A1(n13184), .A2(n11882), .B1(n13364), .B2(n12888), .ZN(
        n15015) );
  INV_X4 U15371 ( .A(n15718), .ZN(n17168) );
  OAI221_X2 U15372 ( .B1(n12454), .B2(n13383), .C1(n12804), .C2(n13377), .A(
        n12975), .ZN(n15018) );
  OAI22_X2 U15373 ( .A1(n13379), .A2(n12768), .B1(n13368), .B2(n11839), .ZN(
        n15017) );
  OAI22_X2 U15374 ( .A1(n11860), .A2(n13373), .B1(n10868), .B2(n13371), .ZN(
        n15016) );
  NAND4_X2 U15375 ( .A1(n15022), .A2(n15021), .A3(n15020), .A4(n15019), .ZN(
        n2478) );
  OAI22_X2 U15376 ( .A1(n10335), .A2(n13181), .B1(n12732), .B2(n13266), .ZN(
        n2466) );
  INV_X4 U15377 ( .A(n2473), .ZN(n15037) );
  OAI22_X2 U15378 ( .A1(n13184), .A2(n11883), .B1(n13364), .B2(n12874), .ZN(
        n15031) );
  INV_X4 U15379 ( .A(n16872), .ZN(n16844) );
  OAI221_X2 U15380 ( .B1(n12442), .B2(n13383), .C1(n12799), .C2(n13377), .A(
        n12970), .ZN(n15034) );
  OAI22_X2 U15381 ( .A1(n13379), .A2(n12769), .B1(n13368), .B2(n11840), .ZN(
        n15033) );
  OAI22_X2 U15382 ( .A1(n11855), .A2(n13373), .B1(n10867), .B2(n13371), .ZN(
        n15032) );
  NAND4_X2 U15383 ( .A1(n15038), .A2(n15037), .A3(n15036), .A4(n15035), .ZN(
        n2458) );
  OAI22_X2 U15384 ( .A1(n10336), .A2(n13181), .B1(n12733), .B2(n13266), .ZN(
        n2446) );
  NOR2_X4 U15385 ( .A1(n12875), .A2(n13276), .ZN(n15039) );
  NOR3_X4 U15386 ( .A1(n15041), .A2(n15040), .A3(n15039), .ZN(n2443) );
  OAI22_X2 U15387 ( .A1(n10339), .A2(n13181), .B1(n12736), .B2(n13266), .ZN(
        n2426) );
  NOR2_X4 U15388 ( .A1(n12889), .A2(n13276), .ZN(n15044) );
  NOR3_X4 U15389 ( .A1(n15046), .A2(n15045), .A3(n15044), .ZN(n2423) );
  OAI22_X2 U15390 ( .A1(n10326), .A2(n13181), .B1(n12722), .B2(n13266), .ZN(
        n2406) );
  INV_X4 U15391 ( .A(n2413), .ZN(n15063) );
  OAI22_X2 U15392 ( .A1(n13184), .A2(n11884), .B1(n13364), .B2(n12832), .ZN(
        n15057) );
  INV_X4 U15393 ( .A(n16031), .ZN(n15978) );
  OAI221_X2 U15394 ( .B1(n12414), .B2(n13383), .C1(n12787), .C2(n13377), .A(
        n12971), .ZN(n15060) );
  OAI22_X2 U15395 ( .A1(n13379), .A2(n12770), .B1(n13368), .B2(n11841), .ZN(
        n15059) );
  OAI22_X2 U15396 ( .A1(n11848), .A2(n13374), .B1(n10862), .B2(n13370), .ZN(
        n15058) );
  NAND4_X2 U15397 ( .A1(n15064), .A2(n15063), .A3(n15062), .A4(n15061), .ZN(
        n2398) );
  OAI22_X2 U15398 ( .A1(n10327), .A2(n13181), .B1(n12723), .B2(n13266), .ZN(
        n2386) );
  NOR2_X4 U15399 ( .A1(n12833), .A2(n13276), .ZN(n15065) );
  NOR3_X4 U15400 ( .A1(n15067), .A2(n15066), .A3(n15065), .ZN(n2383) );
  OAI22_X2 U15401 ( .A1(n10331), .A2(n13181), .B1(n12727), .B2(n13266), .ZN(
        n2366) );
  INV_X4 U15402 ( .A(n2373), .ZN(n15084) );
  OAI22_X2 U15403 ( .A1(n13184), .A2(n11885), .B1(n13364), .B2(n12852), .ZN(
        n15078) );
  INV_X4 U15404 ( .A(n16070), .ZN(n16441) );
  OAI221_X2 U15405 ( .B1(n12428), .B2(n13383), .C1(n12792), .C2(n13377), .A(
        n12972), .ZN(n15081) );
  OAI22_X2 U15406 ( .A1(n13379), .A2(n12771), .B1(n13368), .B2(n11842), .ZN(
        n15080) );
  OAI22_X2 U15407 ( .A1(n12226), .A2(n13374), .B1(n10864), .B2(n13370), .ZN(
        n15079) );
  NAND4_X2 U15408 ( .A1(n15085), .A2(n15084), .A3(n15083), .A4(n15082), .ZN(
        n2358) );
  OAI22_X2 U15409 ( .A1(n10328), .A2(n13181), .B1(n12724), .B2(n13266), .ZN(
        n2345) );
  INV_X4 U15410 ( .A(n2352), .ZN(n15100) );
  OAI22_X2 U15411 ( .A1(n13184), .A2(n11886), .B1(n13364), .B2(n12840), .ZN(
        n15094) );
  INV_X4 U15412 ( .A(n16222), .ZN(n16176) );
  OAI221_X2 U15413 ( .B1(n12419), .B2(n13383), .C1(n12789), .C2(n13377), .A(
        n12973), .ZN(n15097) );
  OAI22_X2 U15414 ( .A1(n13379), .A2(n12772), .B1(n13368), .B2(n11843), .ZN(
        n15096) );
  OAI22_X2 U15415 ( .A1(n12225), .A2(n13374), .B1(n10863), .B2(n13370), .ZN(
        n15095) );
  NAND4_X2 U15416 ( .A1(n15101), .A2(n15100), .A3(n15099), .A4(n15098), .ZN(
        n2337) );
  OAI22_X2 U15417 ( .A1(n10337), .A2(n13181), .B1(n12734), .B2(n13266), .ZN(
        n2325) );
  NOR2_X4 U15418 ( .A1(n12879), .A2(n13276), .ZN(n15102) );
  NOR3_X4 U15419 ( .A1(n15104), .A2(n15103), .A3(n15102), .ZN(n2322) );
  OAI22_X2 U15420 ( .A1(n10329), .A2(n13181), .B1(n12725), .B2(n13266), .ZN(
        n2305) );
  NOR2_X4 U15421 ( .A1(n12841), .A2(n13276), .ZN(n15107) );
  NOR3_X4 U15422 ( .A1(n15109), .A2(n15108), .A3(n15107), .ZN(n2302) );
  OAI22_X2 U15423 ( .A1(n10330), .A2(n13181), .B1(n12726), .B2(n13267), .ZN(
        n2285) );
  NOR2_X4 U15424 ( .A1(n12845), .A2(n13276), .ZN(n15112) );
  NOR3_X4 U15425 ( .A1(n15114), .A2(n15113), .A3(n15112), .ZN(n2282) );
  OAI22_X2 U15426 ( .A1(n10332), .A2(n13181), .B1(n12728), .B2(n13267), .ZN(
        n2265) );
  INV_X4 U15427 ( .A(n2272), .ZN(n15131) );
  OAI22_X2 U15428 ( .A1(n13184), .A2(n12773), .B1(n13365), .B2(n12856), .ZN(
        n15125) );
  INV_X4 U15429 ( .A(n16539), .ZN(n16494) );
  OAI221_X2 U15430 ( .B1(n12429), .B2(n13383), .C1(n12793), .C2(n13377), .A(
        n12974), .ZN(n15128) );
  OAI22_X2 U15431 ( .A1(n13379), .A2(n12774), .B1(n13368), .B2(n11844), .ZN(
        n15127) );
  OAI22_X2 U15432 ( .A1(n12227), .A2(n13374), .B1(n10865), .B2(n13370), .ZN(
        n15126) );
  NAND4_X2 U15433 ( .A1(n15132), .A2(n15131), .A3(n15130), .A4(n15129), .ZN(
        n2257) );
  OAI22_X2 U15434 ( .A1(n10333), .A2(n13181), .B1(n12729), .B2(n13267), .ZN(
        n2245) );
  NOR2_X4 U15435 ( .A1(n12857), .A2(n13275), .ZN(n15133) );
  NOR3_X4 U15436 ( .A1(n15135), .A2(n15134), .A3(n15133), .ZN(n2242) );
  OAI22_X2 U15437 ( .A1(n10334), .A2(n13181), .B1(n12730), .B2(n13267), .ZN(
        n2225) );
  INV_X4 U15438 ( .A(n2232), .ZN(n15152) );
  OAI22_X2 U15439 ( .A1(n13184), .A2(n11887), .B1(n13364), .B2(n12864), .ZN(
        n15146) );
  INV_X4 U15440 ( .A(n17737), .ZN(n16639) );
  OAI221_X2 U15441 ( .B1(n12434), .B2(n13382), .C1(n12795), .C2(n13377), .A(
        n12976), .ZN(n15149) );
  OAI22_X2 U15442 ( .A1(n13379), .A2(n12775), .B1(n13368), .B2(n11845), .ZN(
        n15148) );
  OAI22_X2 U15443 ( .A1(n12228), .A2(n13374), .B1(n10866), .B2(n13370), .ZN(
        n15147) );
  NAND4_X2 U15444 ( .A1(n15153), .A2(n15152), .A3(n15151), .A4(n15150), .ZN(
        n2217) );
  OAI22_X2 U15445 ( .A1(n12279), .A2(n13181), .B1(n12731), .B2(n13267), .ZN(
        n2204) );
  NOR2_X4 U15446 ( .A1(n12865), .A2(n13275), .ZN(n15154) );
  NOR3_X4 U15447 ( .A1(n15156), .A2(n15155), .A3(n15154), .ZN(n2198) );
  OAI22_X2 U15448 ( .A1(n12441), .A2(n13267), .B1(n10767), .B2(n13180), .ZN(
        n2185) );
  OAI22_X2 U15449 ( .A1(n10751), .A2(n13736), .B1(n12440), .B2(n13270), .ZN(
        n15161) );
  OAI221_X2 U15450 ( .B1(n10705), .B2(n13278), .C1(n12439), .C2(n13275), .A(
        n12959), .ZN(n15164) );
  OAI22_X2 U15451 ( .A1(n13379), .A2(n12776), .B1(n13368), .B2(n11694), .ZN(
        n15167) );
  NAND2_X2 U15452 ( .A1(n15172), .A2(n15171), .ZN(n2168) );
  OAI22_X2 U15453 ( .A1(n12453), .A2(n13267), .B1(n10768), .B2(n13180), .ZN(
        n2163) );
  OAI22_X2 U15454 ( .A1(n10752), .A2(n13736), .B1(n12452), .B2(n13270), .ZN(
        n15175) );
  INV_X4 U15455 ( .A(n1866), .ZN(n15286) );
  NAND2_X2 U15456 ( .A1(n15286), .A2(ID_STAGE_imm16_aluA[17]), .ZN(n15176) );
  OAI221_X2 U15457 ( .B1(n10706), .B2(n13278), .C1(n12451), .C2(n13275), .A(
        n15176), .ZN(n15179) );
  OAI22_X2 U15458 ( .A1(n12461), .A2(n13267), .B1(n10769), .B2(n13180), .ZN(
        n2142) );
  OAI22_X2 U15459 ( .A1(n10753), .A2(n13736), .B1(n12460), .B2(n13270), .ZN(
        n15182) );
  NAND2_X2 U15460 ( .A1(n15286), .A2(ID_STAGE_imm16_aluA[18]), .ZN(n15183) );
  OAI221_X2 U15461 ( .B1(n10707), .B2(n13278), .C1(n12459), .C2(n13275), .A(
        n15183), .ZN(n15186) );
  OAI22_X2 U15462 ( .A1(n12464), .A2(n13267), .B1(n10770), .B2(n13180), .ZN(
        n2122) );
  OAI22_X2 U15463 ( .A1(n10754), .A2(n13736), .B1(n12463), .B2(n13270), .ZN(
        n15189) );
  NAND2_X2 U15464 ( .A1(n15286), .A2(ID_STAGE_imm16_aluA[19]), .ZN(n15190) );
  OAI221_X2 U15465 ( .B1(n10708), .B2(n13278), .C1(n12462), .C2(n13275), .A(
        n15190), .ZN(n15193) );
  OAI22_X2 U15466 ( .A1(n12467), .A2(n13267), .B1(n10771), .B2(n13180), .ZN(
        n2102) );
  OAI22_X2 U15467 ( .A1(n10755), .A2(n13736), .B1(n12466), .B2(n13270), .ZN(
        n15196) );
  OAI221_X2 U15468 ( .B1(n10709), .B2(n13278), .C1(n12465), .C2(n13275), .A(
        n12960), .ZN(n15199) );
  OAI22_X2 U15469 ( .A1(n12470), .A2(n13267), .B1(n10772), .B2(n13180), .ZN(
        n2082) );
  OAI22_X2 U15470 ( .A1(n10756), .A2(n13736), .B1(n12469), .B2(n13270), .ZN(
        n15202) );
  OAI221_X2 U15471 ( .B1(n10710), .B2(n13278), .C1(n12468), .C2(n13275), .A(
        n12961), .ZN(n15205) );
  OAI22_X2 U15472 ( .A1(n12473), .A2(n13266), .B1(n10340), .B2(n13180), .ZN(
        n2062) );
  OAI22_X2 U15473 ( .A1(n10757), .A2(n13736), .B1(n12472), .B2(n13270), .ZN(
        n15208) );
  OAI221_X2 U15474 ( .B1(n10711), .B2(n13278), .C1(n12471), .C2(n13275), .A(
        n12967), .ZN(n15211) );
  OAI22_X2 U15475 ( .A1(n12476), .A2(n13267), .B1(n10341), .B2(n13180), .ZN(
        n2042) );
  OAI22_X2 U15476 ( .A1(n10758), .A2(n13736), .B1(n12475), .B2(n13270), .ZN(
        n15214) );
  OAI221_X2 U15477 ( .B1(n10712), .B2(n13278), .C1(n12474), .C2(n13275), .A(
        n12963), .ZN(n15217) );
  OAI22_X2 U15478 ( .A1(n13379), .A2(n12777), .B1(n13367), .B2(n11715), .ZN(
        n15220) );
  NAND2_X2 U15479 ( .A1(n15225), .A2(n15224), .ZN(n2027) );
  OAI22_X2 U15480 ( .A1(n12479), .A2(n13266), .B1(n10342), .B2(n13180), .ZN(
        n2022) );
  OAI22_X2 U15481 ( .A1(n10759), .A2(n13736), .B1(n12478), .B2(n13270), .ZN(
        n15228) );
  OAI221_X2 U15482 ( .B1(n10713), .B2(n13278), .C1(n12477), .C2(n13275), .A(
        n12968), .ZN(n15231) );
  OAI22_X2 U15483 ( .A1(n13379), .A2(n12778), .B1(n13367), .B2(n11718), .ZN(
        n15234) );
  INV_X4 U15484 ( .A(n15770), .ZN(n18047) );
  NAND2_X2 U15485 ( .A1(n15239), .A2(n15238), .ZN(n2007) );
  OAI22_X2 U15486 ( .A1(n12482), .A2(n13267), .B1(n10343), .B2(n13180), .ZN(
        n2002) );
  OAI22_X2 U15487 ( .A1(n10760), .A2(n13735), .B1(n12481), .B2(n13270), .ZN(
        n15242) );
  OAI221_X2 U15488 ( .B1(n10714), .B2(n13278), .C1(n12480), .C2(n13275), .A(
        n12958), .ZN(n15245) );
  OAI22_X2 U15489 ( .A1(n13380), .A2(n12779), .B1(n13367), .B2(n11721), .ZN(
        n15248) );
  NAND2_X2 U15490 ( .A1(n15253), .A2(n15252), .ZN(n1987) );
  OAI22_X2 U15491 ( .A1(n12485), .A2(n13266), .B1(n10344), .B2(n13180), .ZN(
        n1982) );
  OAI22_X2 U15492 ( .A1(n10761), .A2(n13735), .B1(n12484), .B2(n13270), .ZN(
        n15256) );
  NAND2_X2 U15493 ( .A1(n15286), .A2(ID_STAGE_imm16_aluA[26]), .ZN(n15257) );
  OAI221_X2 U15494 ( .B1(n12277), .B2(n13278), .C1(n12483), .C2(n13275), .A(
        n15257), .ZN(n15260) );
  OAI22_X2 U15495 ( .A1(n13380), .A2(n12780), .B1(n13367), .B2(n11724), .ZN(
        n15263) );
  INV_X4 U15496 ( .A(n15837), .ZN(n18135) );
  NAND2_X2 U15497 ( .A1(n15268), .A2(n15267), .ZN(n1967) );
  OAI22_X2 U15498 ( .A1(n12488), .A2(n13267), .B1(n10345), .B2(n13180), .ZN(
        n1962) );
  OAI22_X2 U15499 ( .A1(n10762), .A2(n13735), .B1(n12487), .B2(n13270), .ZN(
        n15271) );
  OAI221_X2 U15500 ( .B1(n10715), .B2(n13279), .C1(n12486), .C2(n13276), .A(
        n12969), .ZN(n15274) );
  OAI22_X2 U15501 ( .A1(n13380), .A2(n12781), .B1(n13367), .B2(n11727), .ZN(
        n15277) );
  INV_X4 U15502 ( .A(n15682), .ZN(n18176) );
  NAND2_X2 U15503 ( .A1(n15282), .A2(n15281), .ZN(n1947) );
  OAI22_X2 U15504 ( .A1(n12491), .A2(n13266), .B1(n10346), .B2(n13180), .ZN(
        n1941) );
  OAI22_X2 U15505 ( .A1(n10763), .A2(n13735), .B1(n12490), .B2(n13270), .ZN(
        n15285) );
  NAND2_X2 U15506 ( .A1(n15286), .A2(ID_STAGE_imm16_aluA[28]), .ZN(n15287) );
  OAI221_X2 U15507 ( .B1(n12278), .B2(n13279), .C1(n12489), .C2(n13276), .A(
        n15287), .ZN(n15290) );
  OAI22_X2 U15508 ( .A1(n13380), .A2(n12782), .B1(n13367), .B2(n11730), .ZN(
        n15293) );
  INV_X4 U15509 ( .A(n15678), .ZN(n18221) );
  NAND2_X2 U15510 ( .A1(n15298), .A2(n15297), .ZN(n1926) );
  OAI22_X2 U15511 ( .A1(n12494), .A2(n13267), .B1(n10347), .B2(n13180), .ZN(
        n1921) );
  OAI22_X2 U15512 ( .A1(n10764), .A2(n13735), .B1(n12493), .B2(n13269), .ZN(
        n15301) );
  OAI221_X2 U15513 ( .B1(n10716), .B2(n13279), .C1(n12492), .C2(n13276), .A(
        n12966), .ZN(n15304) );
  OAI22_X2 U15514 ( .A1(n13380), .A2(n12783), .B1(n13367), .B2(n11733), .ZN(
        n15307) );
  NAND2_X2 U15515 ( .A1(n15312), .A2(n15311), .ZN(n1906) );
  OAI22_X2 U15516 ( .A1(n12497), .A2(n13266), .B1(n10348), .B2(n13180), .ZN(
        n1901) );
  OAI22_X2 U15517 ( .A1(n10765), .A2(n13735), .B1(n12496), .B2(n13270), .ZN(
        n15315) );
  OAI221_X2 U15518 ( .B1(n10717), .B2(n13279), .C1(n12495), .C2(n13276), .A(
        n12957), .ZN(n15318) );
  OAI22_X2 U15519 ( .A1(n13380), .A2(n12784), .B1(n13367), .B2(n11736), .ZN(
        n15321) );
  NAND2_X2 U15521 ( .A1(n15326), .A2(n15325), .ZN(n1886) );
  OAI22_X2 U15522 ( .A1(n10750), .A2(n13267), .B1(n10257), .B2(n13180), .ZN(
        n1875) );
  OAI22_X2 U15523 ( .A1(n10766), .A2(n13735), .B1(n11469), .B2(n13269), .ZN(
        n15333) );
  OAI221_X2 U15524 ( .B1(n10718), .B2(n13279), .C1(n12766), .C2(n13276), .A(
        n12956), .ZN(n15339) );
  OAI22_X2 U15525 ( .A1(n13380), .A2(n12785), .B1(n13367), .B2(n11846), .ZN(
        n15342) );
  INV_X4 U15526 ( .A(n15671), .ZN(n18930) );
  NAND2_X2 U15527 ( .A1(n15347), .A2(n15346), .ZN(n1832) );
  INV_X4 U15528 ( .A(IMEM_BUS_IN[0]), .ZN(n19164) );
  NAND2_X2 U15529 ( .A1(n10397), .A2(n129), .ZN(n1135) );
  INV_X4 U15530 ( .A(n15348), .ZN(n15349) );
  NAND2_X2 U15531 ( .A1(n10258), .A2(n129), .ZN(n1028) );
  NAND2_X2 U15532 ( .A1(n10258), .A2(n200), .ZN(n959) );
  NAND2_X2 U15533 ( .A1(n10258), .A2(n164), .ZN(n924) );
  INV_X4 U15534 ( .A(n15350), .ZN(n15351) );
  NAND2_X2 U15535 ( .A1(n10322), .A2(n164), .ZN(n787) );
  NAND2_X2 U15536 ( .A1(n12022), .A2(n129), .ZN(n719) );
  NAND2_X2 U15537 ( .A1(n12022), .A2(n94), .ZN(n685) );
  NAND2_X2 U15538 ( .A1(n12022), .A2(n200), .ZN(n651) );
  NAND2_X2 U15539 ( .A1(n12022), .A2(n164), .ZN(n616) );
  INV_X4 U15540 ( .A(n15352), .ZN(n15353) );
  NAND2_X2 U15541 ( .A1(n10531), .A2(n129), .ZN(n581) );
  NAND2_X2 U15542 ( .A1(n10397), .A2(n200), .ZN(n376) );
  NAND2_X2 U15543 ( .A1(n10323), .A2(n200), .ZN(n342) );
  NAND2_X2 U15544 ( .A1(n10397), .A2(n164), .ZN(n272) );
  NAND2_X2 U15545 ( .A1(n10259), .A2(n129), .ZN(n235) );
  NAND2_X2 U15546 ( .A1(n10259), .A2(n94), .ZN(n201) );
  NAND2_X2 U15547 ( .A1(n129), .A2(n10262), .ZN(n95) );
  NAND2_X2 U15548 ( .A1(n94), .A2(n10262), .ZN(n27) );
  INV_X4 U15549 ( .A(n15370), .ZN(n15363) );
  NAND2_X2 U15550 ( .A1(n15363), .A2(n12982), .ZN(n15355) );
  OAI21_X4 U15551 ( .B1(ID_STAGE_imm16_aluA[19]), .B2(n15356), .A(n15355), 
        .ZN(n18775) );
  XNOR2_X2 U15552 ( .A(IMEM_BUS_IN[9]), .B(n15375), .ZN(n15362) );
  NAND2_X2 U15553 ( .A1(n15363), .A2(n10824), .ZN(n15357) );
  OAI21_X4 U15554 ( .B1(ID_STAGE_imm16_aluA[16]), .B2(n15358), .A(n15357), 
        .ZN(n18778) );
  INV_X4 U15555 ( .A(n18778), .ZN(n15374) );
  XNOR2_X2 U15556 ( .A(IMEM_BUS_IN[6]), .B(n15374), .ZN(n15361) );
  NAND2_X2 U15557 ( .A1(n13167), .A2(n12021), .ZN(n15359) );
  INV_X4 U15558 ( .A(n18773), .ZN(n15373) );
  XNOR2_X2 U15559 ( .A(IMEM_BUS_IN[10]), .B(n15373), .ZN(n15360) );
  NAND3_X2 U15560 ( .A1(n15362), .A2(n15361), .A3(n15360), .ZN(n15391) );
  NAND2_X2 U15561 ( .A1(n15363), .A2(n11922), .ZN(n15364) );
  OAI21_X4 U15562 ( .B1(ID_STAGE_imm16_aluA[17]), .B2(n15365), .A(n15364), 
        .ZN(n18777) );
  XNOR2_X2 U15563 ( .A(IMEM_BUS_IN[7]), .B(n15379), .ZN(n15372) );
  NAND2_X2 U15564 ( .A1(IMEM_BUS_IN[2]), .A2(IMEM_BUS_IN[0]), .ZN(n15366) );
  INV_X4 U15565 ( .A(IMEM_BUS_IN[5]), .ZN(n18786) );
  NAND2_X2 U15566 ( .A1(n15368), .A2(n15367), .ZN(n15383) );
  NAND2_X2 U15567 ( .A1(n13167), .A2(n11045), .ZN(n15369) );
  INV_X4 U15568 ( .A(n18776), .ZN(n15384) );
  XNOR2_X2 U15569 ( .A(IMEM_BUS_IN[8]), .B(n15384), .ZN(n15371) );
  NAND3_X2 U15570 ( .A1(n15372), .A2(n15383), .A3(n15371), .ZN(n15390) );
  XNOR2_X2 U15571 ( .A(IMEM_BUS_IN[15]), .B(n15373), .ZN(n15378) );
  XNOR2_X2 U15572 ( .A(IMEM_BUS_IN[11]), .B(n15374), .ZN(n15377) );
  XNOR2_X2 U15573 ( .A(IMEM_BUS_IN[14]), .B(n15375), .ZN(n15376) );
  NAND3_X2 U15574 ( .A1(n15378), .A2(n15377), .A3(n15376), .ZN(n15389) );
  XNOR2_X2 U15575 ( .A(IMEM_BUS_IN[12]), .B(n15379), .ZN(n15387) );
  NAND3_X2 U15576 ( .A1(n15381), .A2(n19170), .A3(n15380), .ZN(n15382) );
  NAND2_X2 U15577 ( .A1(n15383), .A2(n15382), .ZN(n15386) );
  XNOR2_X2 U15578 ( .A(IMEM_BUS_IN[13]), .B(n15384), .ZN(n15385) );
  NAND3_X2 U15579 ( .A1(n15387), .A2(n15386), .A3(n15385), .ZN(n15388) );
  NAND2_X2 U15580 ( .A1(n15392), .A2(n18781), .ZN(n15396) );
  NOR2_X4 U15581 ( .A1(n15394), .A2(n15393), .ZN(n15395) );
  NAND3_X4 U15582 ( .A1(n15397), .A2(n15396), .A3(n15395), .ZN(n15406) );
  NAND2_X2 U15583 ( .A1(n15406), .A2(net231227), .ZN(n15407) );
  NOR2_X4 U15585 ( .A1(n15479), .A2(n15478), .ZN(n15480) );
  NAND3_X4 U15586 ( .A1(IMEM_BUS_OUT[23]), .A2(IMEM_BUS_OUT[24]), .A3(n15398), 
        .ZN(n15469) );
  INV_X4 U15587 ( .A(n15469), .ZN(n15467) );
  NAND3_X4 U15588 ( .A1(IMEM_BUS_OUT[22]), .A2(IMEM_BUS_OUT[21]), .A3(n15467), 
        .ZN(n15464) );
  INV_X4 U15589 ( .A(n15457), .ZN(n15399) );
  NAND3_X4 U15591 ( .A1(IMEM_BUS_OUT[7]), .A2(IMEM_BUS_OUT[8]), .A3(n19352), 
        .ZN(n15431) );
  INV_X4 U15592 ( .A(n15428), .ZN(n15402) );
  INV_X4 U15593 ( .A(n15451), .ZN(n15403) );
  INV_X4 U15594 ( .A(n15447), .ZN(n15404) );
  NOR2_X4 U15595 ( .A1(n15443), .A2(n12034), .ZN(n15405) );
  XNOR2_X2 U15596 ( .A(IMEM_BUS_OUT[0]), .B(n15405), .ZN(n15637) );
  NAND2_X2 U15597 ( .A1(n15406), .A2(net230387), .ZN(n18845) );
  NOR3_X4 U15598 ( .A1(n15407), .A2(n10157), .A3(n13955), .ZN(n15490) );
  NAND2_X2 U15599 ( .A1(n13354), .A2(EXEC_MEM_OUT_109), .ZN(n15408) );
  OAI221_X2 U15600 ( .B1(n13350), .B2(n12715), .C1(n15637), .C2(n13344), .A(
        n15408), .ZN(IF_STAGE_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15601 ( .A1(n13746), .A2(n13284), .B1(n13749), .B2(n11586), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15602 ( .A1(n13753), .A2(n13284), .B1(n12825), .B2(n13750), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15603 ( .A1(n10162), .A2(n13284), .B1(n13755), .B2(n10245), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15604 ( .A1(n13758), .A2(n13284), .B1(n13757), .B2(n11338), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15605 ( .A1(n10163), .A2(n13284), .B1(n13761), .B2(n10949), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15606 ( .A1(n13764), .A2(n13284), .B1(n13763), .B2(n11881), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15607 ( .A1(n13768), .A2(n13284), .B1(n12285), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15608 ( .A1(n10164), .A2(n13284), .B1(n12826), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15609 ( .A1(n13774), .A2(n13284), .B1(n12627), .B2(n13772), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15610 ( .A1(n13779), .A2(n13284), .B1(n12827), .B2(n13776), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15611 ( .A1(n13782), .A2(n13284), .B1(n13781), .B2(n10959), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15612 ( .A1(n13786), .A2(n13285), .B1(n13785), .B2(n10371), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15613 ( .A1(n13790), .A2(n13285), .B1(n13789), .B2(n12937), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15614 ( .A1(n13794), .A2(n13285), .B1(n13793), .B2(n10869), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15615 ( .A1(n13799), .A2(n13285), .B1(n13798), .B2(n10861), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15616 ( .A1(n13804), .A2(n13285), .B1(n13803), .B2(n12413), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15617 ( .A1(n13809), .A2(n13285), .B1(n13807), .B2(n12721), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15618 ( .A1(n13813), .A2(n13285), .B1(n13812), .B2(n10325), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15619 ( .A1(n13817), .A2(n13285), .B1(n10673), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15620 ( .A1(n13821), .A2(n13285), .B1(n13820), .B2(n10871), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15621 ( .A1(n13825), .A2(n13285), .B1(n13824), .B2(n10870), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15622 ( .A1(n13829), .A2(n13285), .B1(n13828), .B2(n12383), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15623 ( .A1(n13833), .A2(n13284), .B1(n13832), .B2(n10505), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15624 ( .A1(n13837), .A2(n13285), .B1(n13836), .B2(n12767), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15625 ( .A1(n10165), .A2(n13285), .B1(n12828), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15626 ( .A1(n13843), .A2(n13285), .B1(n13842), .B2(n10958), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15627 ( .A1(n13847), .A2(n13285), .B1(n13846), .B2(n10690), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15628 ( .A1(n13851), .A2(n13284), .B1(n13850), .B2(n10301), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15629 ( .A1(n10166), .A2(n13285), .B1(n13854), .B2(n12382), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15630 ( .A1(n10167), .A2(n13284), .B1(n13856), .B2(n11838), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15631 ( .A1(n13859), .A2(n13284), .B1(n13858), .B2(n11847), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15632 ( .A1(n13863), .A2(n13284), .B1(n13862), .B2(n12786), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U15633 ( .A(n15443), .B(n12034), .ZN(n17194) );
  NAND2_X2 U15634 ( .A1(n13351), .A2(IMEM_BUS_OUT[1]), .ZN(n15410) );
  NAND2_X2 U15635 ( .A1(n13354), .A2(EXEC_MEM_OUT_110), .ZN(n15409) );
  OAI211_X2 U15636 ( .C1(n17194), .C2(n13345), .A(n15410), .B(n15409), .ZN(
        IF_STAGE_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15637 ( .A1(n13746), .A2(n13286), .B1(n11587), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15638 ( .A1(n13752), .A2(n13286), .B1(n12829), .B2(n13750), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15639 ( .A1(n10162), .A2(n13286), .B1(n10250), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15640 ( .A1(n13758), .A2(n13286), .B1(n11362), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15641 ( .A1(n10163), .A2(n13286), .B1(n10968), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15642 ( .A1(n13764), .A2(n13286), .B1(n11884), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15643 ( .A1(n13768), .A2(n13286), .B1(n12286), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15644 ( .A1(n10164), .A2(n13286), .B1(n12830), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15645 ( .A1(n13774), .A2(n13286), .B1(n12628), .B2(n13772), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15646 ( .A1(n13778), .A2(n13286), .B1(n12831), .B2(n13776), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15647 ( .A1(n13782), .A2(n13286), .B1(n10983), .B2(n13780), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15648 ( .A1(n13786), .A2(n13287), .B1(n10385), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15649 ( .A1(n13790), .A2(n13287), .B1(n12940), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15650 ( .A1(n13794), .A2(n13287), .B1(n10880), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15651 ( .A1(n13799), .A2(n13287), .B1(n13797), .B2(n10862), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15652 ( .A1(n13804), .A2(n13287), .B1(n13802), .B2(n12414), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15653 ( .A1(n13809), .A2(n13287), .B1(n13807), .B2(n12722), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15654 ( .A1(n13813), .A2(n13287), .B1(n13811), .B2(n10326), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15655 ( .A1(n13817), .A2(n13287), .B1(n10678), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15656 ( .A1(n13821), .A2(n13287), .B1(n10882), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15657 ( .A1(n13825), .A2(n13287), .B1(n10881), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15658 ( .A1(n13829), .A2(n13287), .B1(n12393), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15659 ( .A1(n13833), .A2(n13286), .B1(n10510), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15660 ( .A1(n13837), .A2(n13287), .B1(n12770), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15661 ( .A1(n10165), .A2(n13287), .B1(n12832), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15662 ( .A1(n13843), .A2(n13286), .B1(n10982), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15663 ( .A1(n13847), .A2(n13287), .B1(n10691), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15664 ( .A1(n13851), .A2(n13286), .B1(n10306), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15665 ( .A1(n10166), .A2(n13287), .B1(n12392), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15666 ( .A1(n10167), .A2(n13286), .B1(n11841), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15667 ( .A1(n13859), .A2(n13286), .B1(n13857), .B2(n11848), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15668 ( .A1(n13863), .A2(n13287), .B1(n13861), .B2(n12787), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15669 ( .A1(n13746), .A2(n13288), .B1(n11588), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15670 ( .A1(n13753), .A2(n13288), .B1(n12833), .B2(n13750), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15671 ( .A1(n10162), .A2(n13288), .B1(n10372), .B2(n13755), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15672 ( .A1(n13758), .A2(n13289), .B1(n11363), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15673 ( .A1(n10163), .A2(n13289), .B1(n10969), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15674 ( .A1(n13764), .A2(n13289), .B1(n12418), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15675 ( .A1(n13768), .A2(n13288), .B1(n12287), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15676 ( .A1(n10164), .A2(n13289), .B1(n12834), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15677 ( .A1(n13774), .A2(n13289), .B1(n12629), .B2(n13772), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15678 ( .A1(n13779), .A2(n13288), .B1(n12835), .B2(n13776), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15679 ( .A1(n13782), .A2(n13289), .B1(n10985), .B2(n13780), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15680 ( .A1(n13786), .A2(n13288), .B1(n10848), .B2(n13785), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15681 ( .A1(n13790), .A2(n13288), .B1(n12945), .B2(n13789), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15682 ( .A1(n13794), .A2(n13288), .B1(n10883), .B2(n13793), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15683 ( .A1(n13799), .A2(n13288), .B1(n10857), .B2(n13798), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15684 ( .A1(n13804), .A2(n13288), .B1(n12415), .B2(n13803), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15685 ( .A1(n13809), .A2(n13288), .B1(n13807), .B2(n12723), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15686 ( .A1(n13813), .A2(n13288), .B1(n13812), .B2(n10327), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15687 ( .A1(n13817), .A2(n13288), .B1(n10679), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15688 ( .A1(n13821), .A2(n13288), .B1(n10885), .B2(n13820), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15689 ( .A1(n13825), .A2(n13288), .B1(n10884), .B2(n13824), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15690 ( .A1(n13829), .A2(n13288), .B1(n12417), .B2(n13828), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15691 ( .A1(n13833), .A2(n13289), .B1(n10511), .B2(n13832), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15692 ( .A1(n13837), .A2(n13289), .B1(n12746), .B2(n13836), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15693 ( .A1(n10165), .A2(n13289), .B1(n12836), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15694 ( .A1(n13843), .A2(n13289), .B1(n10984), .B2(n13842), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15695 ( .A1(n13847), .A2(n13289), .B1(n10692), .B2(n13846), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15696 ( .A1(n13851), .A2(n13289), .B1(n10307), .B2(n13850), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15697 ( .A1(n10166), .A2(n13289), .B1(n12416), .B2(n13854), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15698 ( .A1(n10167), .A2(n13289), .B1(n12737), .B2(n13856), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15699 ( .A1(n13859), .A2(n13289), .B1(n11849), .B2(n13858), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15700 ( .A1(n13863), .A2(n13289), .B1(n12788), .B2(n13862), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15701 ( .A1(n13746), .A2(n13290), .B1(n11589), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15702 ( .A1(n13752), .A2(n13290), .B1(n12837), .B2(n13750), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15703 ( .A1(n10162), .A2(n13290), .B1(n10374), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15704 ( .A1(n13758), .A2(n13291), .B1(n11365), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15705 ( .A1(n10163), .A2(n13291), .B1(n10970), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15706 ( .A1(n13764), .A2(n13291), .B1(n11886), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15707 ( .A1(n13768), .A2(n13290), .B1(n12289), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15708 ( .A1(n10164), .A2(n13291), .B1(n12838), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15709 ( .A1(n13774), .A2(n13291), .B1(n12630), .B2(n13772), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15710 ( .A1(n13778), .A2(n13290), .B1(n12839), .B2(n13776), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15711 ( .A1(n13782), .A2(n13291), .B1(n10987), .B2(n13780), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15712 ( .A1(n13786), .A2(n13290), .B1(n10850), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15713 ( .A1(n13790), .A2(n13290), .B1(n12942), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15714 ( .A1(n13794), .A2(n13290), .B1(n10889), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15715 ( .A1(n13799), .A2(n13290), .B1(n13798), .B2(n10863), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15716 ( .A1(n13804), .A2(n13290), .B1(n13803), .B2(n12419), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15717 ( .A1(n13809), .A2(n13290), .B1(n13807), .B2(n12724), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15718 ( .A1(n13813), .A2(n13290), .B1(n13811), .B2(n10328), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15719 ( .A1(n13817), .A2(n13290), .B1(n10681), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15720 ( .A1(n13821), .A2(n13290), .B1(n10891), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15721 ( .A1(n13825), .A2(n13290), .B1(n10890), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15722 ( .A1(n13829), .A2(n13290), .B1(n12397), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15723 ( .A1(n13833), .A2(n13291), .B1(n10513), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15724 ( .A1(n13837), .A2(n13291), .B1(n12772), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15725 ( .A1(n10165), .A2(n13291), .B1(n12840), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15726 ( .A1(n13843), .A2(n13291), .B1(n10986), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15727 ( .A1(n13847), .A2(n13291), .B1(n10693), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15728 ( .A1(n13851), .A2(n13291), .B1(n10309), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15729 ( .A1(n10166), .A2(n13291), .B1(n12396), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15730 ( .A1(n10167), .A2(n13291), .B1(n11843), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15731 ( .A1(n13859), .A2(n13291), .B1(n13858), .B2(n12225), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15732 ( .A1(n13863), .A2(n13291), .B1(n13862), .B2(n12789), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15733 ( .A1(n13746), .A2(n13292), .B1(n11590), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15734 ( .A1(n13753), .A2(n13292), .B1(n12841), .B2(n13750), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15735 ( .A1(n10162), .A2(n13292), .B1(n10376), .B2(n13755), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15736 ( .A1(n13758), .A2(n13293), .B1(n11367), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15737 ( .A1(n10163), .A2(n13293), .B1(n10971), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15738 ( .A1(n13764), .A2(n13293), .B1(n12423), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15739 ( .A1(n13768), .A2(n13292), .B1(n11409), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15740 ( .A1(n10164), .A2(n13293), .B1(n12842), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15741 ( .A1(n13774), .A2(n13293), .B1(n12631), .B2(n13772), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15742 ( .A1(n13779), .A2(n13292), .B1(n12843), .B2(n13776), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15743 ( .A1(n13782), .A2(n13293), .B1(n10989), .B2(n13780), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15744 ( .A1(n13786), .A2(n13292), .B1(n10852), .B2(n13785), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15745 ( .A1(n13790), .A2(n13292), .B1(n12946), .B2(n13789), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15746 ( .A1(n13794), .A2(n13292), .B1(n10391), .B2(n13793), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15747 ( .A1(n13799), .A2(n13292), .B1(n10858), .B2(n13798), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15748 ( .A1(n13804), .A2(n13292), .B1(n12420), .B2(n13803), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15749 ( .A1(n13809), .A2(n13292), .B1(n13807), .B2(n12725), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15750 ( .A1(n13813), .A2(n13292), .B1(n13812), .B2(n10329), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15751 ( .A1(n13817), .A2(n13292), .B1(n10683), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15752 ( .A1(n13821), .A2(n13292), .B1(n10895), .B2(n13820), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15753 ( .A1(n13825), .A2(n13292), .B1(n10894), .B2(n13824), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15754 ( .A1(n13829), .A2(n13292), .B1(n12422), .B2(n13828), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15755 ( .A1(n13833), .A2(n13293), .B1(n10515), .B2(n13832), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15756 ( .A1(n13837), .A2(n13293), .B1(n12747), .B2(n13836), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15757 ( .A1(n10165), .A2(n13293), .B1(n12844), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15758 ( .A1(n13843), .A2(n13293), .B1(n10988), .B2(n13842), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15759 ( .A1(n13847), .A2(n13293), .B1(n10694), .B2(n13846), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15760 ( .A1(n13851), .A2(n13293), .B1(n10311), .B2(n13850), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15761 ( .A1(n10166), .A2(n13293), .B1(n12421), .B2(n13854), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15762 ( .A1(n10167), .A2(n13293), .B1(n12738), .B2(n13856), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15763 ( .A1(n13859), .A2(n13293), .B1(n11850), .B2(n13858), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15764 ( .A1(n13863), .A2(n13293), .B1(n12790), .B2(n13862), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15765 ( .A1(n13746), .A2(n13294), .B1(n11591), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15766 ( .A1(n13752), .A2(n13294), .B1(n12845), .B2(n13750), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15767 ( .A1(n10162), .A2(n13294), .B1(n10377), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15768 ( .A1(n13758), .A2(n13295), .B1(n11368), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15769 ( .A1(n10163), .A2(n13295), .B1(n10972), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15770 ( .A1(n13764), .A2(n13295), .B1(n12427), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15771 ( .A1(n13768), .A2(n13294), .B1(n11410), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15772 ( .A1(n10164), .A2(n13295), .B1(n12846), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15773 ( .A1(n13774), .A2(n13295), .B1(n12632), .B2(n13772), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15774 ( .A1(n13778), .A2(n13294), .B1(n12847), .B2(n13776), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15775 ( .A1(n13782), .A2(n13295), .B1(n10991), .B2(n13780), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15776 ( .A1(n13786), .A2(n13294), .B1(n10853), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15777 ( .A1(n13790), .A2(n13294), .B1(n12947), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15778 ( .A1(n13794), .A2(n13294), .B1(n10392), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15779 ( .A1(n13799), .A2(n13294), .B1(n10859), .B2(n13798), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15780 ( .A1(n13804), .A2(n13294), .B1(n12424), .B2(n13803), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15781 ( .A1(n13809), .A2(n13294), .B1(n13807), .B2(n12726), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15782 ( .A1(n13813), .A2(n13294), .B1(n13811), .B2(n10330), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15783 ( .A1(n13817), .A2(n13294), .B1(n10684), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15784 ( .A1(n13821), .A2(n13294), .B1(n10897), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15785 ( .A1(n13825), .A2(n13294), .B1(n10896), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15786 ( .A1(n13829), .A2(n13294), .B1(n12426), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15787 ( .A1(n13833), .A2(n13295), .B1(n10516), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15788 ( .A1(n13837), .A2(n13295), .B1(n12748), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15789 ( .A1(n10165), .A2(n13295), .B1(n12848), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15790 ( .A1(n13843), .A2(n13295), .B1(n10990), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15791 ( .A1(n13847), .A2(n13295), .B1(n10695), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15792 ( .A1(n13851), .A2(n13295), .B1(n10312), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15793 ( .A1(n10166), .A2(n13295), .B1(n12425), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15794 ( .A1(n10167), .A2(n13295), .B1(n12739), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15795 ( .A1(n13859), .A2(n13295), .B1(n11851), .B2(n13858), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15796 ( .A1(n13863), .A2(n13295), .B1(n12791), .B2(n13862), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15797 ( .A1(n13746), .A2(n13296), .B1(n11592), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15798 ( .A1(n13753), .A2(n13296), .B1(n12849), .B2(n13750), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15799 ( .A1(n10162), .A2(n13296), .B1(n10373), .B2(n13755), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15800 ( .A1(n13758), .A2(n13297), .B1(n11364), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15801 ( .A1(n10163), .A2(n13297), .B1(n10973), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15802 ( .A1(n13764), .A2(n13297), .B1(n11885), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15803 ( .A1(n13768), .A2(n13296), .B1(n12288), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15804 ( .A1(n10164), .A2(n13297), .B1(n12850), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15805 ( .A1(n13774), .A2(n13297), .B1(n12633), .B2(n13772), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15806 ( .A1(n13779), .A2(n13296), .B1(n12851), .B2(n13776), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15807 ( .A1(n13782), .A2(n13297), .B1(n10993), .B2(n13780), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15808 ( .A1(n13786), .A2(n13296), .B1(n10849), .B2(n13785), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15809 ( .A1(n13790), .A2(n13296), .B1(n12941), .B2(n13789), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15810 ( .A1(n13794), .A2(n13296), .B1(n10886), .B2(n13793), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15811 ( .A1(n13799), .A2(n13296), .B1(n13798), .B2(n10864), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15812 ( .A1(n13804), .A2(n13296), .B1(n13803), .B2(n12428), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15813 ( .A1(n13809), .A2(n13296), .B1(n13807), .B2(n12727), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15814 ( .A1(n13813), .A2(n13296), .B1(n13812), .B2(n10331), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15815 ( .A1(n13817), .A2(n13296), .B1(n10680), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15816 ( .A1(n13821), .A2(n13296), .B1(n10888), .B2(n13820), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15817 ( .A1(n13825), .A2(n13296), .B1(n10887), .B2(n13824), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15818 ( .A1(n13829), .A2(n13296), .B1(n12395), .B2(n13828), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15819 ( .A1(n13833), .A2(n13297), .B1(n10512), .B2(n13832), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15820 ( .A1(n13837), .A2(n13297), .B1(n12771), .B2(n13836), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15821 ( .A1(n10165), .A2(n13297), .B1(n12852), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15822 ( .A1(n13843), .A2(n13297), .B1(n10992), .B2(n13842), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15823 ( .A1(n13847), .A2(n13297), .B1(n10696), .B2(n13846), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15824 ( .A1(n13851), .A2(n13297), .B1(n10308), .B2(n13850), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15825 ( .A1(n10166), .A2(n13297), .B1(n12394), .B2(n13854), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15826 ( .A1(n10167), .A2(n13297), .B1(n11842), .B2(n13856), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15827 ( .A1(n13859), .A2(n13297), .B1(n13858), .B2(n12226), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15828 ( .A1(n13863), .A2(n13297), .B1(n13862), .B2(n12792), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U15829 ( .A(IMEM_BUS_OUT[10]), .B(n15435), .ZN(n16473) );
  NAND2_X2 U15830 ( .A1(n13354), .A2(EXEC_MEM_OUT_119), .ZN(n15411) );
  OAI221_X2 U15831 ( .B1(n16473), .B2(n13345), .C1(n11097), .C2(n13350), .A(
        n15411), .ZN(IF_STAGE_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U15832 ( .A1(n13354), .A2(EXEC_MEM_OUT_120), .ZN(n15414) );
  OAI221_X2 U15833 ( .B1(n16474), .B2(n13345), .C1(n11470), .C2(n13350), .A(
        n15414), .ZN(IF_STAGE_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15834 ( .A1(n13746), .A2(n13298), .B1(n11593), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15835 ( .A1(n13752), .A2(n13298), .B1(n12853), .B2(n13750), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15836 ( .A1(n10162), .A2(n13298), .B1(n10378), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15837 ( .A1(n13758), .A2(n13299), .B1(n11369), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15838 ( .A1(n10163), .A2(n13299), .B1(n10974), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15839 ( .A1(n13764), .A2(n13299), .B1(n12773), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15840 ( .A1(n13768), .A2(n13298), .B1(n11411), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15841 ( .A1(n10164), .A2(n13299), .B1(n12854), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15842 ( .A1(n13774), .A2(n13299), .B1(n12634), .B2(n13772), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15843 ( .A1(n13778), .A2(n13298), .B1(n12855), .B2(n13776), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15844 ( .A1(n13782), .A2(n13299), .B1(n10995), .B2(n13780), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15845 ( .A1(n13786), .A2(n13298), .B1(n10854), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15846 ( .A1(n13790), .A2(n13298), .B1(n12943), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15847 ( .A1(n13794), .A2(n13298), .B1(n10393), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15848 ( .A1(n13799), .A2(n13298), .B1(n13798), .B2(n10865), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15849 ( .A1(n13804), .A2(n13298), .B1(n13803), .B2(n12429), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15850 ( .A1(n13809), .A2(n13298), .B1(n13807), .B2(n12728), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15851 ( .A1(n13813), .A2(n13298), .B1(n13811), .B2(n10332), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15852 ( .A1(n13817), .A2(n13298), .B1(n10685), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15853 ( .A1(n13821), .A2(n13298), .B1(n10899), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15854 ( .A1(n13825), .A2(n13298), .B1(n10898), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15855 ( .A1(n13829), .A2(n13298), .B1(n12400), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15856 ( .A1(n13833), .A2(n13299), .B1(n10517), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15857 ( .A1(n13837), .A2(n13299), .B1(n12774), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15858 ( .A1(n10165), .A2(n13299), .B1(n12856), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15859 ( .A1(n13843), .A2(n13299), .B1(n10994), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15860 ( .A1(n13847), .A2(n13299), .B1(n10697), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15861 ( .A1(n13851), .A2(n13299), .B1(n10313), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15862 ( .A1(n10166), .A2(n13299), .B1(n12399), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15863 ( .A1(n10167), .A2(n13299), .B1(n11844), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15864 ( .A1(n13859), .A2(n13299), .B1(n13858), .B2(n12227), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15865 ( .A1(n13863), .A2(n13299), .B1(n13862), .B2(n12793), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U15866 ( .A1(n13354), .A2(EXEC_MEM_OUT_121), .ZN(n15415) );
  OAI221_X2 U15867 ( .B1(n16520), .B2(n13345), .C1(n12317), .C2(n13350), .A(
        n15415), .ZN(IF_STAGE_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  INV_X4 U15868 ( .A(n15416), .ZN(n15418) );
  NAND2_X2 U15869 ( .A1(n13354), .A2(EXEC_MEM_OUT_122), .ZN(n15419) );
  OAI221_X2 U15870 ( .B1(n16617), .B2(n13345), .C1(n12989), .C2(n13350), .A(
        n15419), .ZN(IF_STAGE_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15871 ( .A1(n13746), .A2(n13300), .B1(n11594), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15872 ( .A1(n13753), .A2(n13300), .B1(n12857), .B2(n13750), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15873 ( .A1(n10162), .A2(n13300), .B1(n10379), .B2(n13755), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15874 ( .A1(n13758), .A2(n13301), .B1(n11370), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15875 ( .A1(n10163), .A2(n13301), .B1(n10975), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15876 ( .A1(n13764), .A2(n13301), .B1(n12433), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15877 ( .A1(n13768), .A2(n13300), .B1(n11412), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15878 ( .A1(n10164), .A2(n13301), .B1(n12858), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15879 ( .A1(n13774), .A2(n13301), .B1(n12635), .B2(n13772), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15880 ( .A1(n13779), .A2(n13300), .B1(n12859), .B2(n13776), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15881 ( .A1(n13782), .A2(n13301), .B1(n10997), .B2(n13780), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15882 ( .A1(n13786), .A2(n13300), .B1(n10855), .B2(n13785), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15883 ( .A1(n13790), .A2(n13300), .B1(n12948), .B2(n13789), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15884 ( .A1(n13794), .A2(n13300), .B1(n10394), .B2(n13793), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15885 ( .A1(n13799), .A2(n13300), .B1(n10252), .B2(n13797), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15886 ( .A1(n13804), .A2(n13300), .B1(n12430), .B2(n13802), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15887 ( .A1(n13809), .A2(n13300), .B1(n13807), .B2(n12729), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15888 ( .A1(n13813), .A2(n13300), .B1(n13812), .B2(n10333), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15889 ( .A1(n13817), .A2(n13300), .B1(n10686), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15890 ( .A1(n13821), .A2(n13300), .B1(n10901), .B2(n13820), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15891 ( .A1(n13825), .A2(n13300), .B1(n10900), .B2(n13824), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15892 ( .A1(n13829), .A2(n13300), .B1(n12432), .B2(n13828), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15893 ( .A1(n13833), .A2(n13301), .B1(n10518), .B2(n13832), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15894 ( .A1(n13837), .A2(n13301), .B1(n12749), .B2(n13836), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15895 ( .A1(n10165), .A2(n13301), .B1(n12860), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15896 ( .A1(n13843), .A2(n13301), .B1(n10996), .B2(n13842), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15897 ( .A1(n13847), .A2(n13301), .B1(n10698), .B2(n13846), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15898 ( .A1(n13851), .A2(n13301), .B1(n10314), .B2(n13850), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15899 ( .A1(n10166), .A2(n13301), .B1(n12431), .B2(n13854), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15900 ( .A1(n10167), .A2(n13301), .B1(n12740), .B2(n13856), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15901 ( .A1(n13859), .A2(n13301), .B1(n11852), .B2(n13857), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15902 ( .A1(n13863), .A2(n13301), .B1(n12794), .B2(n13861), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U15903 ( .A(IMEM_BUS_OUT[14]), .B(n15420), .ZN(n16665) );
  NAND2_X2 U15904 ( .A1(n13354), .A2(EXEC_MEM_OUT_123), .ZN(n15421) );
  OAI221_X2 U15905 ( .B1(n16665), .B2(n13345), .C1(n12988), .C2(n13350), .A(
        n15421), .ZN(IF_STAGE_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15906 ( .A1(n13746), .A2(n13302), .B1(n11595), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15907 ( .A1(n13752), .A2(n13302), .B1(n12861), .B2(n13750), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15908 ( .A1(n10162), .A2(n13302), .B1(n10380), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15909 ( .A1(n13758), .A2(n13303), .B1(n11371), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15910 ( .A1(n10163), .A2(n13303), .B1(n10976), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15911 ( .A1(n13764), .A2(n13303), .B1(n11887), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15912 ( .A1(n13768), .A2(n13302), .B1(n11413), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15913 ( .A1(n10164), .A2(n13303), .B1(n12862), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15914 ( .A1(n13774), .A2(n13303), .B1(n12636), .B2(n13772), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15915 ( .A1(n13778), .A2(n13302), .B1(n12863), .B2(n13776), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15916 ( .A1(n13782), .A2(n13303), .B1(n10999), .B2(n13780), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15917 ( .A1(n13786), .A2(n13302), .B1(n10856), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15918 ( .A1(n13790), .A2(n13302), .B1(n12944), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15919 ( .A1(n13794), .A2(n13302), .B1(n10395), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15920 ( .A1(n13799), .A2(n13302), .B1(n13798), .B2(n10866), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15921 ( .A1(n13804), .A2(n13302), .B1(n13803), .B2(n12434), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15922 ( .A1(n13809), .A2(n13302), .B1(n13807), .B2(n12730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15923 ( .A1(n13813), .A2(n13302), .B1(n13811), .B2(n10334), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15924 ( .A1(n13817), .A2(n13302), .B1(n10687), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15925 ( .A1(n13821), .A2(n13302), .B1(n10903), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15926 ( .A1(n13825), .A2(n13302), .B1(n10902), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15927 ( .A1(n13829), .A2(n13302), .B1(n12402), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15928 ( .A1(n13833), .A2(n13303), .B1(n10519), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15929 ( .A1(n13837), .A2(n13303), .B1(n12775), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15930 ( .A1(n10165), .A2(n13303), .B1(n12864), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15931 ( .A1(n13843), .A2(n13303), .B1(n10998), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15932 ( .A1(n13847), .A2(n13303), .B1(n10699), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15933 ( .A1(n13851), .A2(n13303), .B1(n10315), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15934 ( .A1(n10166), .A2(n13303), .B1(n12401), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15935 ( .A1(n10167), .A2(n13303), .B1(n11845), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15936 ( .A1(n13859), .A2(n13303), .B1(n13858), .B2(n12228), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15937 ( .A1(n13863), .A2(n13303), .B1(n13862), .B2(n12795), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15938 ( .A1(n13746), .A2(n13305), .B1(n11596), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15939 ( .A1(n13753), .A2(n13305), .B1(n12865), .B2(n13750), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15940 ( .A1(n10162), .A2(n13304), .B1(n10846), .B2(n13755), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15941 ( .A1(n13758), .A2(n13304), .B1(n11372), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15942 ( .A1(n10163), .A2(n13305), .B1(n12080), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15943 ( .A1(n13764), .A2(n13305), .B1(n12438), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15944 ( .A1(n13768), .A2(n13304), .B1(n11414), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15945 ( .A1(n10164), .A2(n13305), .B1(n12866), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15946 ( .A1(n13774), .A2(n13304), .B1(n12637), .B2(n13772), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15947 ( .A1(n13779), .A2(n13305), .B1(n12867), .B2(n13776), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15948 ( .A1(n13782), .A2(n13304), .B1(n11000), .B2(n13780), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15949 ( .A1(n13786), .A2(n13304), .B1(n12024), .B2(n13785), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15950 ( .A1(n13790), .A2(n13304), .B1(n12952), .B2(n13789), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15951 ( .A1(n13794), .A2(n13304), .B1(n10396), .B2(n13793), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15952 ( .A1(n13799), .A2(n13304), .B1(n10253), .B2(n13797), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15953 ( .A1(n13804), .A2(n13304), .B1(n12435), .B2(n13802), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15954 ( .A1(n13809), .A2(n13304), .B1(n13807), .B2(n12731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15955 ( .A1(n13813), .A2(n13304), .B1(n13812), .B2(n12279), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15956 ( .A1(n13817), .A2(n13304), .B1(n10688), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15957 ( .A1(n13821), .A2(n13304), .B1(n10905), .B2(n13820), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15958 ( .A1(n13825), .A2(n13304), .B1(n10904), .B2(n13824), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15959 ( .A1(n13829), .A2(n13304), .B1(n12437), .B2(n13828), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15960 ( .A1(n13833), .A2(n13305), .B1(n12041), .B2(n13832), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15961 ( .A1(n13837), .A2(n13305), .B1(n12750), .B2(n13836), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15962 ( .A1(n10165), .A2(n13305), .B1(n12868), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15963 ( .A1(n13843), .A2(n13305), .B1(n12082), .B2(n13842), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15964 ( .A1(n13847), .A2(n13305), .B1(n12276), .B2(n13846), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15965 ( .A1(n13851), .A2(n13305), .B1(n10504), .B2(n13850), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15966 ( .A1(n10166), .A2(n13305), .B1(n12436), .B2(n13854), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15967 ( .A1(n10167), .A2(n13305), .B1(n12741), .B2(n13856), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15968 ( .A1(n13859), .A2(n13305), .B1(n11853), .B2(n13857), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15969 ( .A1(n13863), .A2(n13305), .B1(n12796), .B2(n13861), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U15970 ( .A1(n13354), .A2(EXEC_MEM_OUT_124), .ZN(n15424) );
  OAI221_X2 U15971 ( .B1(n16722), .B2(n13345), .C1(n12554), .C2(n13350), .A(
        n15424), .ZN(IF_STAGE_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15972 ( .A1(n13746), .A2(n13306), .B1(n12403), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15973 ( .A1(n13752), .A2(n13306), .B1(n13751), .B2(n12439), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15974 ( .A1(n10162), .A2(n13306), .B1(n11692), .B2(n13755), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15975 ( .A1(n13758), .A2(n13306), .B1(n13757), .B2(n10751), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15976 ( .A1(n10163), .A2(n13306), .B1(n11757), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15977 ( .A1(n13764), .A2(n13306), .B1(n11578), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15978 ( .A1(n13768), .A2(n13306), .B1(n12798), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15979 ( .A1(n10164), .A2(n13306), .B1(n12869), .B2(n13771), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15980 ( .A1(n13775), .A2(n13306), .B1(n13773), .B2(n10705), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15981 ( .A1(n13778), .A2(n13306), .B1(n13777), .B2(n12440), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15982 ( .A1(n13782), .A2(n13306), .B1(n13781), .B2(n10767), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15983 ( .A1(n13787), .A2(n13307), .B1(n11693), .B2(n13785), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15984 ( .A1(n719), .A2(n13307), .B1(n12137), .B2(n13789), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15985 ( .A1(n13795), .A2(n13307), .B1(n10493), .B2(n13793), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15986 ( .A1(n13800), .A2(n13307), .B1(n13798), .B2(n10942), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15987 ( .A1(n13805), .A2(n13307), .B1(n13803), .B2(n12751), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15988 ( .A1(n13809), .A2(n13307), .B1(n13808), .B2(n12441), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15989 ( .A1(n13814), .A2(n13307), .B1(n12570), .B2(n13812), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15990 ( .A1(n13818), .A2(n13307), .B1(n12585), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15991 ( .A1(n13822), .A2(n13307), .B1(n12261), .B2(n13820), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15992 ( .A1(n13826), .A2(n13307), .B1(n10492), .B2(n13824), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15993 ( .A1(n13830), .A2(n13307), .B1(n12290), .B2(n13828), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15994 ( .A1(n13833), .A2(n13307), .B1(n10927), .B2(n13832), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15995 ( .A1(n13837), .A2(n13306), .B1(n12776), .B2(n13836), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15996 ( .A1(n10165), .A2(n13306), .B1(n12870), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15997 ( .A1(n13843), .A2(n13307), .B1(n10520), .B2(n13842), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15998 ( .A1(n13847), .A2(n13306), .B1(n11573), .B2(n13846), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U15999 ( .A1(n13851), .A2(n13307), .B1(n11415), .B2(n13850), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16000 ( .A1(n10166), .A2(n13306), .B1(n11806), .B2(n13854), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16001 ( .A1(n10167), .A2(n13307), .B1(n11694), .B2(n13856), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16002 ( .A1(n13859), .A2(n13307), .B1(n13858), .B2(n11854), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16003 ( .A1(n13863), .A2(n13306), .B1(n13862), .B2(n12797), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16004 ( .A1(n13354), .A2(EXEC_MEM_OUT_125), .ZN(n15425) );
  OAI221_X2 U16005 ( .B1(n16768), .B2(n13345), .C1(n12542), .C2(n13350), .A(
        n15425), .ZN(IF_STAGE_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16006 ( .A1(n13746), .A2(n13308), .B1(n12387), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16007 ( .A1(n13752), .A2(n13308), .B1(n12871), .B2(n13751), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16008 ( .A1(n10162), .A2(n13308), .B1(n10247), .B2(n13755), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16009 ( .A1(n13758), .A2(n13308), .B1(n11359), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16010 ( .A1(n10163), .A2(n13308), .B1(n10977), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16011 ( .A1(n13764), .A2(n13308), .B1(n11883), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16012 ( .A1(n13768), .A2(n13308), .B1(n11405), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16013 ( .A1(n10164), .A2(n13308), .B1(n12872), .B2(n13771), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16014 ( .A1(n13775), .A2(n13308), .B1(n12638), .B2(n13773), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16015 ( .A1(n13778), .A2(n13308), .B1(n12873), .B2(n13777), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16016 ( .A1(n13782), .A2(n13308), .B1(n12083), .B2(n13780), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16017 ( .A1(n13787), .A2(n13309), .B1(n10382), .B2(n13785), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16018 ( .A1(n719), .A2(n13308), .B1(n12939), .B2(n13789), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16019 ( .A1(n13795), .A2(n13309), .B1(n10387), .B2(n13793), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16020 ( .A1(n13800), .A2(n13308), .B1(n13798), .B2(n10867), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16021 ( .A1(n13805), .A2(n13309), .B1(n13803), .B2(n12442), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16022 ( .A1(n13809), .A2(n13308), .B1(n13808), .B2(n12732), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16023 ( .A1(n13814), .A2(n13309), .B1(n13812), .B2(n10335), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16024 ( .A1(n13818), .A2(n13308), .B1(n10675), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16025 ( .A1(n13822), .A2(n13309), .B1(n10875), .B2(n13820), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16026 ( .A1(n13826), .A2(n13308), .B1(n10874), .B2(n13824), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16027 ( .A1(n13830), .A2(n13309), .B1(n12389), .B2(n13828), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16028 ( .A1(n13833), .A2(n13309), .B1(n10507), .B2(n13832), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16029 ( .A1(n13837), .A2(n13309), .B1(n12769), .B2(n13836), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16030 ( .A1(n10165), .A2(n13309), .B1(n12874), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16031 ( .A1(n13843), .A2(n13309), .B1(n11001), .B2(n13842), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16032 ( .A1(n13847), .A2(n13309), .B1(n10700), .B2(n13846), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16033 ( .A1(n13851), .A2(n13309), .B1(n10303), .B2(n13850), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16034 ( .A1(n10166), .A2(n13309), .B1(n12388), .B2(n13854), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16035 ( .A1(n10167), .A2(n13309), .B1(n11840), .B2(n13856), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16036 ( .A1(n13859), .A2(n13309), .B1(n13858), .B2(n11855), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16037 ( .A1(n13863), .A2(n13309), .B1(n13862), .B2(n12799), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16038 ( .A1(n13746), .A2(n13310), .B1(n12390), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16039 ( .A1(n13752), .A2(n13310), .B1(n12875), .B2(n13751), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16040 ( .A1(n10162), .A2(n13310), .B1(n10248), .B2(n13755), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16041 ( .A1(n13758), .A2(n13310), .B1(n11360), .B2(n13757), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16042 ( .A1(n10163), .A2(n13310), .B1(n10978), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16043 ( .A1(n13764), .A2(n13310), .B1(n12446), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16044 ( .A1(n13768), .A2(n13310), .B1(n11406), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16045 ( .A1(n10164), .A2(n13310), .B1(n12876), .B2(n13771), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16046 ( .A1(n13775), .A2(n13310), .B1(n12639), .B2(n13773), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16047 ( .A1(n13778), .A2(n13310), .B1(n12877), .B2(n13777), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16048 ( .A1(n13782), .A2(n13310), .B1(n12084), .B2(n13781), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16049 ( .A1(n13787), .A2(n13311), .B1(n10383), .B2(n13785), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16050 ( .A1(n719), .A2(n13310), .B1(n12949), .B2(n13789), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16051 ( .A1(n13795), .A2(n13311), .B1(n10388), .B2(n13793), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16052 ( .A1(n13800), .A2(n13310), .B1(n10254), .B2(n13797), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16053 ( .A1(n13805), .A2(n13311), .B1(n12443), .B2(n13802), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16054 ( .A1(n13809), .A2(n13310), .B1(n13808), .B2(n12733), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16055 ( .A1(n13814), .A2(n13311), .B1(n13812), .B2(n10336), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16056 ( .A1(n13818), .A2(n13310), .B1(n10676), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16057 ( .A1(n13822), .A2(n13311), .B1(n10877), .B2(n13820), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16058 ( .A1(n13826), .A2(n13310), .B1(n10876), .B2(n13824), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16059 ( .A1(n13830), .A2(n13311), .B1(n12445), .B2(n13828), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16060 ( .A1(n13833), .A2(n13311), .B1(n10508), .B2(n13832), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16061 ( .A1(n13837), .A2(n13311), .B1(n12752), .B2(n13836), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16062 ( .A1(n10165), .A2(n13311), .B1(n12878), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16063 ( .A1(n13843), .A2(n13311), .B1(n11002), .B2(n13842), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16064 ( .A1(n13847), .A2(n13311), .B1(n10701), .B2(n13846), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16065 ( .A1(n13851), .A2(n13311), .B1(n10304), .B2(n13850), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16066 ( .A1(n10166), .A2(n13311), .B1(n12444), .B2(n13854), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16067 ( .A1(n10167), .A2(n13311), .B1(n12742), .B2(n13856), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16068 ( .A1(n13859), .A2(n13311), .B1(n11856), .B2(n13857), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16069 ( .A1(n13863), .A2(n13311), .B1(n12800), .B2(n13861), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16070 ( .A1(n13351), .A2(IMEM_BUS_OUT[5]), .ZN(n15427) );
  NAND2_X2 U16071 ( .A1(n13354), .A2(EXEC_MEM_OUT_114), .ZN(n15426) );
  OAI211_X2 U16072 ( .C1(n16958), .C2(n13345), .A(n15427), .B(n15426), .ZN(
        IF_STAGE_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16073 ( .A1(n13354), .A2(EXEC_MEM_OUT_115), .ZN(n15430) );
  OAI221_X2 U16074 ( .B1(n16968), .B2(n13345), .C1(n12559), .C2(n13350), .A(
        n15430), .ZN(IF_STAGE_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16075 ( .A1(n13354), .A2(EXEC_MEM_OUT_116), .ZN(n15433) );
  OAI221_X2 U16076 ( .B1(n16467), .B2(n13345), .C1(n12544), .C2(n13350), .A(
        n15433), .ZN(IF_STAGE_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16077 ( .A1(n13354), .A2(EXEC_MEM_OUT_117), .ZN(n15434) );
  OAI221_X2 U16078 ( .B1(n16974), .B2(n13345), .C1(n12318), .C2(n13350), .A(
        n15434), .ZN(IF_STAGE_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16079 ( .A1(n13746), .A2(n13312), .B1(n12398), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16080 ( .A1(n13752), .A2(n13312), .B1(n12879), .B2(n13751), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16081 ( .A1(n10162), .A2(n13312), .B1(n10375), .B2(n13755), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16082 ( .A1(n13758), .A2(n13312), .B1(n11366), .B2(n13757), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16083 ( .A1(n10163), .A2(n13312), .B1(n10979), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16084 ( .A1(n13764), .A2(n13312), .B1(n12450), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16085 ( .A1(n13768), .A2(n13312), .B1(n11408), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16086 ( .A1(n10164), .A2(n13312), .B1(n12880), .B2(n13771), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16087 ( .A1(n13775), .A2(n13312), .B1(n12640), .B2(n13773), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16088 ( .A1(n13778), .A2(n13312), .B1(n12881), .B2(n13777), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16089 ( .A1(n13782), .A2(n13312), .B1(n12085), .B2(n13781), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16090 ( .A1(n13787), .A2(n13313), .B1(n10851), .B2(n13785), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16091 ( .A1(n719), .A2(n13312), .B1(n12950), .B2(n13789), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16092 ( .A1(n13795), .A2(n13313), .B1(n10390), .B2(n13793), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16093 ( .A1(n13800), .A2(n13312), .B1(n10255), .B2(n13797), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16094 ( .A1(n13805), .A2(n13313), .B1(n12447), .B2(n13802), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16095 ( .A1(n13809), .A2(n13312), .B1(n13808), .B2(n12734), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16096 ( .A1(n13814), .A2(n13313), .B1(n13812), .B2(n10337), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16097 ( .A1(n13818), .A2(n13312), .B1(n10682), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16098 ( .A1(n13822), .A2(n13313), .B1(n10893), .B2(n13820), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16099 ( .A1(n13826), .A2(n13312), .B1(n10892), .B2(n13824), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16100 ( .A1(n13830), .A2(n13313), .B1(n12449), .B2(n13828), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16101 ( .A1(n13833), .A2(n13313), .B1(n10514), .B2(n13832), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16102 ( .A1(n13837), .A2(n13313), .B1(n12753), .B2(n13836), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16103 ( .A1(n10165), .A2(n13313), .B1(n12882), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16104 ( .A1(n13843), .A2(n13313), .B1(n11003), .B2(n13842), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16105 ( .A1(n13847), .A2(n13313), .B1(n10702), .B2(n13846), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16106 ( .A1(n13851), .A2(n13313), .B1(n10310), .B2(n13850), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16107 ( .A1(n10166), .A2(n13313), .B1(n12448), .B2(n13854), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16108 ( .A1(n10167), .A2(n13313), .B1(n12743), .B2(n13856), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16109 ( .A1(n13859), .A2(n13313), .B1(n11857), .B2(n13857), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16110 ( .A1(n13863), .A2(n13313), .B1(n12801), .B2(n13861), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  INV_X4 U16111 ( .A(n15436), .ZN(n15438) );
  NAND2_X2 U16112 ( .A1(n13354), .A2(EXEC_MEM_OUT_118), .ZN(n15439) );
  OAI221_X2 U16113 ( .B1(n17031), .B2(n13345), .C1(n12315), .C2(n13349), .A(
        n15439), .ZN(IF_STAGE_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16114 ( .A1(n13746), .A2(n13314), .B1(n12404), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16115 ( .A1(n13752), .A2(n13314), .B1(n13751), .B2(n12451), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16116 ( .A1(n10162), .A2(n13314), .B1(n11695), .B2(n13755), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16117 ( .A1(n13758), .A2(n13314), .B1(n13756), .B2(n10752), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16118 ( .A1(n10163), .A2(n13314), .B1(n11758), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16119 ( .A1(n13764), .A2(n13314), .B1(n11782), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16120 ( .A1(n13768), .A2(n13314), .B1(n12803), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16121 ( .A1(n10164), .A2(n13314), .B1(n12883), .B2(n13771), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16122 ( .A1(n13775), .A2(n13314), .B1(n13773), .B2(n10706), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16123 ( .A1(n13778), .A2(n13314), .B1(n13777), .B2(n12452), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16124 ( .A1(n13782), .A2(n13314), .B1(n13780), .B2(n10768), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16125 ( .A1(n13787), .A2(n13314), .B1(n11696), .B2(n13785), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16126 ( .A1(n719), .A2(n13315), .B1(n11274), .B2(n13789), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16127 ( .A1(n13795), .A2(n13315), .B1(n10495), .B2(n13793), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16128 ( .A1(n13800), .A2(n13314), .B1(n10230), .B2(n13797), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16129 ( .A1(n13805), .A2(n13315), .B1(n11859), .B2(n13802), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16130 ( .A1(n13809), .A2(n13314), .B1(n13808), .B2(n12453), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16131 ( .A1(n13814), .A2(n13315), .B1(n12571), .B2(n13812), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16132 ( .A1(n13818), .A2(n13314), .B1(n12586), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16133 ( .A1(n13822), .A2(n13315), .B1(n11275), .B2(n13820), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16134 ( .A1(n13826), .A2(n13314), .B1(n10494), .B2(n13824), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16135 ( .A1(n13830), .A2(n13315), .B1(n12291), .B2(n13828), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16136 ( .A1(n13833), .A2(n13315), .B1(n10928), .B2(n13832), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16137 ( .A1(n13837), .A2(n13315), .B1(n12754), .B2(n13836), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16138 ( .A1(n10165), .A2(n13315), .B1(n12884), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16139 ( .A1(n13843), .A2(n13315), .B1(n10316), .B2(n13842), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16140 ( .A1(n13847), .A2(n13315), .B1(n11783), .B2(n13846), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16141 ( .A1(n13851), .A2(n13315), .B1(n11416), .B2(n13850), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16142 ( .A1(n10166), .A2(n13315), .B1(n11807), .B2(n13854), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16143 ( .A1(n10167), .A2(n13315), .B1(n11697), .B2(n13856), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16144 ( .A1(n13859), .A2(n13315), .B1(n11858), .B2(n13857), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16145 ( .A1(n13863), .A2(n13315), .B1(n12802), .B2(n13861), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16146 ( .A1(n13354), .A2(EXEC_MEM_OUT_126), .ZN(n15442) );
  OAI221_X2 U16147 ( .B1(n17116), .B2(n13345), .C1(n12993), .C2(n13349), .A(
        n15442), .ZN(IF_STAGE_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16148 ( .A1(n13746), .A2(n13316), .B1(n12384), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16149 ( .A1(n13752), .A2(n13316), .B1(n12885), .B2(n13751), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16150 ( .A1(n10162), .A2(n13316), .B1(n10246), .B2(n13755), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16151 ( .A1(n13758), .A2(n13316), .B1(n11358), .B2(n13757), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16152 ( .A1(n10163), .A2(n13316), .B1(n10980), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16153 ( .A1(n13764), .A2(n13316), .B1(n11882), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16154 ( .A1(n13768), .A2(n13316), .B1(n11404), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16155 ( .A1(n10164), .A2(n13316), .B1(n12886), .B2(n13771), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16156 ( .A1(n13775), .A2(n13316), .B1(n12641), .B2(n13773), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16157 ( .A1(n13778), .A2(n13316), .B1(n12887), .B2(n13777), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16158 ( .A1(n13782), .A2(n13316), .B1(n12086), .B2(n13781), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16159 ( .A1(n13787), .A2(n13317), .B1(n10381), .B2(n13785), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16160 ( .A1(n719), .A2(n13316), .B1(n12938), .B2(n13789), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16161 ( .A1(n13795), .A2(n13317), .B1(n10386), .B2(n13793), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16162 ( .A1(n13800), .A2(n13316), .B1(n13798), .B2(n10868), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16163 ( .A1(n13805), .A2(n13317), .B1(n13803), .B2(n12454), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16164 ( .A1(n13809), .A2(n13316), .B1(n13808), .B2(n12735), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16165 ( .A1(n13814), .A2(n13317), .B1(n13812), .B2(n10338), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16166 ( .A1(n13818), .A2(n13316), .B1(n10674), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16167 ( .A1(n13822), .A2(n13317), .B1(n10873), .B2(n13820), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16168 ( .A1(n13826), .A2(n13316), .B1(n10872), .B2(n13824), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16169 ( .A1(n13830), .A2(n13317), .B1(n12386), .B2(n13828), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16170 ( .A1(n13833), .A2(n13317), .B1(n10506), .B2(n13832), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16171 ( .A1(n13837), .A2(n13317), .B1(n12768), .B2(n13836), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16172 ( .A1(n10165), .A2(n13317), .B1(n12888), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16173 ( .A1(n13843), .A2(n13317), .B1(n11004), .B2(n13842), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16174 ( .A1(n13847), .A2(n13317), .B1(n10703), .B2(n13846), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16175 ( .A1(n13851), .A2(n13317), .B1(n10302), .B2(n13850), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16176 ( .A1(n10166), .A2(n13317), .B1(n12385), .B2(n13854), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16177 ( .A1(n10167), .A2(n13317), .B1(n11839), .B2(n13856), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16178 ( .A1(n13859), .A2(n13317), .B1(n13858), .B2(n11860), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16179 ( .A1(n13863), .A2(n13317), .B1(n13862), .B2(n12804), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16180 ( .A1(n13351), .A2(IMEM_BUS_OUT[2]), .ZN(n15446) );
  NAND2_X2 U16181 ( .A1(n13354), .A2(EXEC_MEM_OUT_111), .ZN(n15445) );
  OAI211_X2 U16182 ( .C1(n17211), .C2(n13345), .A(n15446), .B(n15445), .ZN(
        IF_STAGE_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  INV_X4 U16183 ( .A(n15452), .ZN(n15448) );
  OAI21_X4 U16184 ( .B1(IMEM_BUS_OUT[3]), .B2(n15448), .A(n15447), .ZN(n16957)
         );
  NAND2_X2 U16185 ( .A1(n13351), .A2(IMEM_BUS_OUT[3]), .ZN(n15450) );
  NAND2_X2 U16186 ( .A1(n13354), .A2(EXEC_MEM_OUT_112), .ZN(n15449) );
  OAI211_X2 U16187 ( .C1(n16957), .C2(n13345), .A(n15450), .B(n15449), .ZN(
        IF_STAGE_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16188 ( .A1(n13746), .A2(n13318), .B1(n12391), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16189 ( .A1(n13752), .A2(n13318), .B1(n12889), .B2(n13751), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16190 ( .A1(n10162), .A2(n13318), .B1(n10249), .B2(n13755), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16191 ( .A1(n13758), .A2(n13318), .B1(n11361), .B2(n13757), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16192 ( .A1(n10163), .A2(n13318), .B1(n10981), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16193 ( .A1(n13764), .A2(n13318), .B1(n12458), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16194 ( .A1(n13768), .A2(n13318), .B1(n11407), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16195 ( .A1(n10164), .A2(n13318), .B1(n12890), .B2(n13771), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16196 ( .A1(n13775), .A2(n13318), .B1(n12642), .B2(n13773), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16197 ( .A1(n13778), .A2(n13318), .B1(n12891), .B2(n13777), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16198 ( .A1(n13782), .A2(n13318), .B1(n12087), .B2(n13781), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16199 ( .A1(n13787), .A2(n13319), .B1(n10384), .B2(n13785), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16200 ( .A1(n719), .A2(n13318), .B1(n12951), .B2(n13789), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16201 ( .A1(n13795), .A2(n13319), .B1(n10389), .B2(n13793), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16202 ( .A1(n13800), .A2(n13318), .B1(n10256), .B2(n13797), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16203 ( .A1(n13805), .A2(n13319), .B1(n12455), .B2(n13802), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16204 ( .A1(n13809), .A2(n13318), .B1(n13808), .B2(n12736), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16205 ( .A1(n13814), .A2(n13319), .B1(n13812), .B2(n10339), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16206 ( .A1(n13818), .A2(n13318), .B1(n10677), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16207 ( .A1(n13822), .A2(n13319), .B1(n10879), .B2(n13820), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16208 ( .A1(n13826), .A2(n13318), .B1(n10878), .B2(n13824), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16209 ( .A1(n13830), .A2(n13319), .B1(n12457), .B2(n13828), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16210 ( .A1(n13833), .A2(n13319), .B1(n10509), .B2(n13832), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16211 ( .A1(n13837), .A2(n13319), .B1(n12755), .B2(n13836), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16212 ( .A1(n10165), .A2(n13319), .B1(n12892), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16213 ( .A1(n13843), .A2(n13319), .B1(n11005), .B2(n13842), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16214 ( .A1(n13847), .A2(n13319), .B1(n10704), .B2(n13846), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16215 ( .A1(n13851), .A2(n13319), .B1(n10305), .B2(n13850), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16216 ( .A1(n10166), .A2(n13319), .B1(n12456), .B2(n13854), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16217 ( .A1(n10167), .A2(n13319), .B1(n12744), .B2(n13856), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16218 ( .A1(n13859), .A2(n13319), .B1(n11861), .B2(n13857), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16219 ( .A1(n13863), .A2(n13319), .B1(n12805), .B2(n13861), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16220 ( .A1(n13351), .A2(IMEM_BUS_OUT[4]), .ZN(n15454) );
  NAND2_X2 U16221 ( .A1(n13354), .A2(EXEC_MEM_OUT_113), .ZN(n15453) );
  OAI211_X2 U16222 ( .C1(n17284), .C2(n13345), .A(n15454), .B(n15453), .ZN(
        IF_STAGE_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16223 ( .A1(n13354), .A2(EXEC_MEM_OUT_127), .ZN(n15456) );
  OAI221_X2 U16224 ( .B1(n17381), .B2(n13344), .C1(n12560), .C2(n13349), .A(
        n15456), .ZN(IF_STAGE_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16225 ( .A1(n13746), .A2(n13320), .B1(n12405), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16226 ( .A1(n13752), .A2(n13320), .B1(n13750), .B2(n12459), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16227 ( .A1(n10162), .A2(n13320), .B1(n11698), .B2(n13755), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16228 ( .A1(n13758), .A2(n13320), .B1(n13757), .B2(n10753), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16229 ( .A1(n10163), .A2(n13320), .B1(n11759), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16230 ( .A1(n13764), .A2(n13320), .B1(n11579), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16231 ( .A1(n13768), .A2(n13320), .B1(n12807), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16232 ( .A1(n10164), .A2(n13320), .B1(n12893), .B2(n13771), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16233 ( .A1(n13775), .A2(n13320), .B1(n13772), .B2(n10707), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16234 ( .A1(n13778), .A2(n13320), .B1(n13776), .B2(n12460), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16235 ( .A1(n13782), .A2(n13320), .B1(n13781), .B2(n10769), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16236 ( .A1(n13787), .A2(n13321), .B1(n11699), .B2(n13785), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16237 ( .A1(n719), .A2(n13321), .B1(n11098), .B2(n13789), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16238 ( .A1(n13795), .A2(n13320), .B1(n10497), .B2(n13793), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16239 ( .A1(n13800), .A2(n13321), .B1(n10231), .B2(n13797), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16240 ( .A1(n13805), .A2(n13320), .B1(n11863), .B2(n13802), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16241 ( .A1(n13809), .A2(n13321), .B1(n13808), .B2(n12461), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16242 ( .A1(n13814), .A2(n13320), .B1(n12572), .B2(n13812), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16243 ( .A1(n13818), .A2(n13321), .B1(n12587), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16244 ( .A1(n13822), .A2(n13320), .B1(n11276), .B2(n13820), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16245 ( .A1(n13826), .A2(n13321), .B1(n10496), .B2(n13824), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16246 ( .A1(n13830), .A2(n13320), .B1(n12292), .B2(n13828), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16247 ( .A1(n13833), .A2(n13321), .B1(n10929), .B2(n13832), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16248 ( .A1(n13837), .A2(n13321), .B1(n12756), .B2(n13836), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16249 ( .A1(n10165), .A2(n13321), .B1(n12894), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16250 ( .A1(n13843), .A2(n13321), .B1(n10317), .B2(n13842), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16251 ( .A1(n13847), .A2(n13321), .B1(n11574), .B2(n13846), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16252 ( .A1(n13851), .A2(n13321), .B1(n11417), .B2(n13850), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16253 ( .A1(n10166), .A2(n13321), .B1(n11808), .B2(n13854), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16254 ( .A1(n10167), .A2(n13321), .B1(n11700), .B2(n13856), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16255 ( .A1(n13859), .A2(n13321), .B1(n11862), .B2(n13857), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16256 ( .A1(n13863), .A2(n13321), .B1(n12806), .B2(n13861), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16257 ( .A1(n13746), .A2(n13322), .B1(n12406), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16258 ( .A1(n13752), .A2(n13322), .B1(n13751), .B2(n12462), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16259 ( .A1(n10162), .A2(n13322), .B1(n11701), .B2(n13755), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16260 ( .A1(n13758), .A2(n13322), .B1(n13756), .B2(n10754), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16261 ( .A1(n10163), .A2(n13322), .B1(n11760), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16262 ( .A1(n13764), .A2(n13322), .B1(n11580), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16263 ( .A1(n13768), .A2(n13322), .B1(n12809), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16264 ( .A1(n10164), .A2(n13322), .B1(n12895), .B2(n13771), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16265 ( .A1(n13775), .A2(n13322), .B1(n13773), .B2(n10708), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16266 ( .A1(n13778), .A2(n13322), .B1(n13777), .B2(n12463), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16267 ( .A1(n13782), .A2(n13322), .B1(n13780), .B2(n10770), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16268 ( .A1(n13787), .A2(n13323), .B1(n11702), .B2(n13785), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16269 ( .A1(n719), .A2(n13323), .B1(n11099), .B2(n13789), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16270 ( .A1(n13795), .A2(n13322), .B1(n10499), .B2(n13793), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16271 ( .A1(n13800), .A2(n13323), .B1(n10232), .B2(n13797), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16272 ( .A1(n13805), .A2(n13322), .B1(n11865), .B2(n13802), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16273 ( .A1(n13809), .A2(n13323), .B1(n13808), .B2(n12464), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16274 ( .A1(n13814), .A2(n13322), .B1(n12573), .B2(n13812), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16275 ( .A1(n13818), .A2(n13323), .B1(n12588), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16276 ( .A1(n13822), .A2(n13322), .B1(n11277), .B2(n13820), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16277 ( .A1(n13826), .A2(n13323), .B1(n10498), .B2(n13824), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16278 ( .A1(n13830), .A2(n13322), .B1(n12293), .B2(n13828), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16279 ( .A1(n13833), .A2(n13323), .B1(n10930), .B2(n13832), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16280 ( .A1(n13837), .A2(n13323), .B1(n12757), .B2(n13836), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16281 ( .A1(n10165), .A2(n13323), .B1(n12896), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16282 ( .A1(n13843), .A2(n13323), .B1(n10318), .B2(n13842), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16283 ( .A1(n13847), .A2(n13323), .B1(n11575), .B2(n13846), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16284 ( .A1(n13851), .A2(n13323), .B1(n11418), .B2(n13850), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16285 ( .A1(n10166), .A2(n13323), .B1(n11809), .B2(n13854), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16286 ( .A1(n10167), .A2(n13323), .B1(n11703), .B2(n13856), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16287 ( .A1(n13859), .A2(n13323), .B1(n11864), .B2(n13857), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16288 ( .A1(n13863), .A2(n13323), .B1(n12808), .B2(n13861), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16289 ( .A1(n13354), .A2(EXEC_MEM_OUT_128), .ZN(n15458) );
  OAI221_X2 U16290 ( .B1(n17432), .B2(n13344), .C1(n12716), .C2(n13349), .A(
        n15458), .ZN(IF_STAGE_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16291 ( .A1(n13746), .A2(n13324), .B1(n12407), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16292 ( .A1(n13752), .A2(n13324), .B1(n13750), .B2(n12465), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16293 ( .A1(n10162), .A2(n13324), .B1(n11704), .B2(n13755), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16294 ( .A1(n13758), .A2(n13324), .B1(n13757), .B2(n10755), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16295 ( .A1(n10163), .A2(n13324), .B1(n11761), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16296 ( .A1(n13764), .A2(n13324), .B1(n11581), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16297 ( .A1(n13768), .A2(n13324), .B1(n12811), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16298 ( .A1(n10164), .A2(n13324), .B1(n12897), .B2(n13771), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16299 ( .A1(n13775), .A2(n13324), .B1(n13772), .B2(n10709), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16300 ( .A1(n13778), .A2(n13324), .B1(n13776), .B2(n12466), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16301 ( .A1(n13782), .A2(n13324), .B1(n13781), .B2(n10771), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16302 ( .A1(n13787), .A2(n13324), .B1(n11705), .B2(n13785), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16303 ( .A1(n719), .A2(n13325), .B1(n11100), .B2(n13789), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16304 ( .A1(n13795), .A2(n13325), .B1(n10501), .B2(n13793), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16305 ( .A1(n13800), .A2(n13324), .B1(n10233), .B2(n13797), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16306 ( .A1(n13805), .A2(n13325), .B1(n11868), .B2(n13802), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16307 ( .A1(n13809), .A2(n13325), .B1(n13808), .B2(n12467), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16308 ( .A1(n13814), .A2(n13324), .B1(n12574), .B2(n13811), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16309 ( .A1(n13818), .A2(n13325), .B1(n12589), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16310 ( .A1(n13822), .A2(n13324), .B1(n11278), .B2(n13820), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16311 ( .A1(n13826), .A2(n13325), .B1(n10500), .B2(n13824), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16312 ( .A1(n13830), .A2(n13324), .B1(n12294), .B2(n13828), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16313 ( .A1(n13833), .A2(n13325), .B1(n10931), .B2(n13832), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16314 ( .A1(n13837), .A2(n13325), .B1(n11866), .B2(n13836), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16315 ( .A1(n10165), .A2(n13325), .B1(n12898), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16316 ( .A1(n13843), .A2(n13325), .B1(n10319), .B2(n13842), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16317 ( .A1(n13847), .A2(n13325), .B1(n11576), .B2(n13846), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16318 ( .A1(n13851), .A2(n13325), .B1(n11419), .B2(n13850), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16319 ( .A1(n10166), .A2(n13325), .B1(n11810), .B2(n13854), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16320 ( .A1(n10167), .A2(n13325), .B1(n11706), .B2(n13856), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16321 ( .A1(n13859), .A2(n13325), .B1(n11867), .B2(n13857), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16322 ( .A1(n13863), .A2(n13325), .B1(n12810), .B2(n13861), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16323 ( .A1(n15464), .A2(n12567), .ZN(n15461) );
  NAND2_X2 U16324 ( .A1(n15461), .A2(n15460), .ZN(n17488) );
  NAND2_X2 U16325 ( .A1(n13354), .A2(EXEC_MEM_OUT_129), .ZN(n15462) );
  OAI221_X2 U16326 ( .B1(n17488), .B2(n13344), .C1(n12567), .C2(n13349), .A(
        n15462), .ZN(IF_STAGE_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16327 ( .A1(n13746), .A2(n13326), .B1(n12408), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16328 ( .A1(n13752), .A2(n13326), .B1(n13751), .B2(n12468), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16329 ( .A1(n10162), .A2(n13326), .B1(n11707), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16330 ( .A1(n13758), .A2(n13326), .B1(n13756), .B2(n10756), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16331 ( .A1(n10163), .A2(n13326), .B1(n11762), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16332 ( .A1(n13764), .A2(n13326), .B1(n11582), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16333 ( .A1(n13768), .A2(n13326), .B1(n12813), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16334 ( .A1(n10164), .A2(n13326), .B1(n12899), .B2(n13771), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16335 ( .A1(n13775), .A2(n13326), .B1(n13773), .B2(n10710), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16336 ( .A1(n13778), .A2(n13326), .B1(n13777), .B2(n12469), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16337 ( .A1(n13782), .A2(n13326), .B1(n13780), .B2(n10772), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16338 ( .A1(n13787), .A2(n13326), .B1(n11708), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16339 ( .A1(n719), .A2(n13327), .B1(n11101), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16340 ( .A1(n13795), .A2(n13327), .B1(n10503), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16341 ( .A1(n13800), .A2(n13326), .B1(n10234), .B2(n13797), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16342 ( .A1(n13805), .A2(n13327), .B1(n11871), .B2(n13802), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16343 ( .A1(n13809), .A2(n13327), .B1(n13808), .B2(n12470), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16344 ( .A1(n13814), .A2(n13326), .B1(n12575), .B2(n13811), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16345 ( .A1(n13818), .A2(n13327), .B1(n12590), .B2(n13815), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16346 ( .A1(n13822), .A2(n13326), .B1(n11279), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16347 ( .A1(n13826), .A2(n13327), .B1(n10502), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16348 ( .A1(n13830), .A2(n13326), .B1(n12295), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16349 ( .A1(n13833), .A2(n13327), .B1(n10932), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16350 ( .A1(n13837), .A2(n13327), .B1(n11869), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16351 ( .A1(n10165), .A2(n13327), .B1(n12900), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16352 ( .A1(n13843), .A2(n13327), .B1(n10320), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16353 ( .A1(n13847), .A2(n13327), .B1(n11577), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16354 ( .A1(n13851), .A2(n13327), .B1(n11420), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16355 ( .A1(n10166), .A2(n13327), .B1(n11811), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16356 ( .A1(n10167), .A2(n13327), .B1(n11709), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16357 ( .A1(n13859), .A2(n13327), .B1(n11870), .B2(n13857), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16358 ( .A1(n13863), .A2(n13327), .B1(n12812), .B2(n13861), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  INV_X4 U16359 ( .A(n15463), .ZN(n15465) );
  NAND2_X2 U16360 ( .A1(n15465), .A2(n15464), .ZN(n17672) );
  NAND2_X2 U16361 ( .A1(n13354), .A2(EXEC_MEM_OUT_130), .ZN(n15466) );
  OAI221_X2 U16362 ( .B1(n17672), .B2(n13344), .C1(n12314), .C2(n13349), .A(
        n15466), .ZN(IF_STAGE_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16363 ( .A1(n13746), .A2(n13328), .B1(n12409), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16364 ( .A1(n13753), .A2(n13328), .B1(n13750), .B2(n12471), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16365 ( .A1(n10162), .A2(n13328), .B1(n11710), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16366 ( .A1(n13758), .A2(n13328), .B1(n13757), .B2(n10757), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16367 ( .A1(n10163), .A2(n13328), .B1(n11763), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16368 ( .A1(n13764), .A2(n13328), .B1(n10792), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16369 ( .A1(n13768), .A2(n13328), .B1(n12815), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16370 ( .A1(n10164), .A2(n13328), .B1(n12901), .B2(n13771), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16371 ( .A1(n13774), .A2(n13328), .B1(n13772), .B2(n10711), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16372 ( .A1(n13779), .A2(n13328), .B1(n13776), .B2(n12472), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16373 ( .A1(n787), .A2(n13328), .B1(n13781), .B2(n10340), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16374 ( .A1(n13786), .A2(n13329), .B1(n11711), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16375 ( .A1(n13790), .A2(n13329), .B1(n12138), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16376 ( .A1(n13794), .A2(n13329), .B1(n10292), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16377 ( .A1(n13799), .A2(n13329), .B1(n10324), .B2(n13797), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16378 ( .A1(n13804), .A2(n13329), .B1(n11872), .B2(n13802), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16379 ( .A1(n13809), .A2(n13329), .B1(n13808), .B2(n12473), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16380 ( .A1(n13813), .A2(n13329), .B1(n12576), .B2(n13811), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16381 ( .A1(n13817), .A2(n13329), .B1(n12591), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16382 ( .A1(n13821), .A2(n13329), .B1(n12262), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16383 ( .A1(n13825), .A2(n13329), .B1(n10918), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16384 ( .A1(n13829), .A2(n13329), .B1(n11421), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16385 ( .A1(n13833), .A2(n13328), .B1(n10521), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16386 ( .A1(n13837), .A2(n13329), .B1(n12250), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16387 ( .A1(n10165), .A2(n13329), .B1(n12902), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16388 ( .A1(n272), .A2(n13328), .B1(n10321), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16389 ( .A1(n13847), .A2(n13329), .B1(n10783), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16390 ( .A1(n13851), .A2(n13328), .B1(n10741), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16391 ( .A1(n10166), .A2(n13329), .B1(n11812), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16392 ( .A1(n10167), .A2(n13328), .B1(n11712), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16393 ( .A1(n13859), .A2(n13328), .B1(n12213), .B2(n13857), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16394 ( .A1(n27), .A2(n13329), .B1(n12814), .B2(n13861), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U16395 ( .A(IMEM_BUS_OUT[22]), .B(n15467), .ZN(n17826) );
  NAND2_X2 U16396 ( .A1(n13354), .A2(EXEC_MEM_OUT_131), .ZN(n15468) );
  OAI221_X2 U16397 ( .B1(n17826), .B2(n13344), .C1(n12181), .C2(n13349), .A(
        n15468), .ZN(IF_STAGE_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16398 ( .A1(n13746), .A2(n13330), .B1(n12410), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16399 ( .A1(n13753), .A2(n13330), .B1(n13751), .B2(n12474), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16400 ( .A1(n10162), .A2(n13330), .B1(n11713), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16401 ( .A1(n13758), .A2(n13330), .B1(n13756), .B2(n10758), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16402 ( .A1(n10163), .A2(n13330), .B1(n11764), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16403 ( .A1(n13764), .A2(n13330), .B1(n10793), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16404 ( .A1(n13768), .A2(n13330), .B1(n11888), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16405 ( .A1(n10164), .A2(n13330), .B1(n12903), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16406 ( .A1(n13774), .A2(n13330), .B1(n13773), .B2(n10712), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16407 ( .A1(n13779), .A2(n13330), .B1(n13777), .B2(n12475), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16408 ( .A1(n787), .A2(n13330), .B1(n13780), .B2(n10341), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16409 ( .A1(n13786), .A2(n13331), .B1(n11714), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16410 ( .A1(n719), .A2(n13331), .B1(n12139), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16411 ( .A1(n13795), .A2(n13331), .B1(n10293), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16412 ( .A1(n13800), .A2(n13331), .B1(n13798), .B2(n10533), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16413 ( .A1(n13805), .A2(n13331), .B1(n13803), .B2(n12758), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16414 ( .A1(n13809), .A2(n13331), .B1(n13807), .B2(n12476), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16415 ( .A1(n13813), .A2(n13331), .B1(n12577), .B2(n13811), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16416 ( .A1(n13817), .A2(n13331), .B1(n12592), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16417 ( .A1(n13821), .A2(n13331), .B1(n12263), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16418 ( .A1(n13825), .A2(n13331), .B1(n10919), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16419 ( .A1(n13829), .A2(n13331), .B1(n11422), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16420 ( .A1(n13833), .A2(n13331), .B1(n10522), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16421 ( .A1(n13837), .A2(n13330), .B1(n12777), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16422 ( .A1(n10165), .A2(n13330), .B1(n12904), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16423 ( .A1(n272), .A2(n13331), .B1(n12042), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16424 ( .A1(n13847), .A2(n13330), .B1(n10784), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16425 ( .A1(n13851), .A2(n13331), .B1(n10742), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16426 ( .A1(n10166), .A2(n13330), .B1(n11813), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16427 ( .A1(n10167), .A2(n13331), .B1(n11715), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16428 ( .A1(n13859), .A2(n13331), .B1(n13858), .B2(n11873), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16429 ( .A1(n27), .A2(n13330), .B1(n13862), .B2(n12816), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16430 ( .A1(n13354), .A2(EXEC_MEM_OUT_132), .ZN(n15471) );
  OAI221_X2 U16431 ( .B1(n17973), .B2(n13345), .C1(n12313), .C2(n13349), .A(
        n15471), .ZN(IF_STAGE_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16432 ( .A1(n13354), .A2(EXEC_MEM_OUT_133), .ZN(n15472) );
  OAI221_X2 U16433 ( .B1(n18063), .B2(n13344), .C1(n12319), .C2(n13349), .A(
        n15472), .ZN(IF_STAGE_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16434 ( .A1(n13746), .A2(n13332), .B1(n11497), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16435 ( .A1(n13753), .A2(n13332), .B1(n13751), .B2(n12477), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16436 ( .A1(n10162), .A2(n13332), .B1(n11716), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16437 ( .A1(n13758), .A2(n13332), .B1(n13756), .B2(n10759), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16438 ( .A1(n10163), .A2(n13332), .B1(n11765), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16439 ( .A1(n13764), .A2(n13332), .B1(n10794), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16440 ( .A1(n13768), .A2(n13332), .B1(n11889), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16441 ( .A1(n10164), .A2(n13332), .B1(n12905), .B2(n13771), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16442 ( .A1(n13774), .A2(n13332), .B1(n13773), .B2(n10713), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16443 ( .A1(n13779), .A2(n13332), .B1(n13777), .B2(n12478), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16444 ( .A1(n13782), .A2(n13332), .B1(n13780), .B2(n10342), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16445 ( .A1(n13786), .A2(n13333), .B1(n11717), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16446 ( .A1(n13790), .A2(n13333), .B1(n12140), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16447 ( .A1(n13794), .A2(n13333), .B1(n10294), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16448 ( .A1(n13799), .A2(n13333), .B1(n13797), .B2(n10534), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16449 ( .A1(n13804), .A2(n13333), .B1(n13802), .B2(n12759), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16450 ( .A1(n13809), .A2(n13333), .B1(n13808), .B2(n12479), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16451 ( .A1(n13813), .A2(n13333), .B1(n12578), .B2(n13811), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16452 ( .A1(n13817), .A2(n13333), .B1(n12593), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16453 ( .A1(n13821), .A2(n13333), .B1(n12264), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16454 ( .A1(n13825), .A2(n13333), .B1(n10920), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16455 ( .A1(n13829), .A2(n13333), .B1(n11423), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16456 ( .A1(n13833), .A2(n13332), .B1(n10523), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16457 ( .A1(n13837), .A2(n13333), .B1(n12778), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16458 ( .A1(n10165), .A2(n13333), .B1(n12906), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16459 ( .A1(n272), .A2(n13332), .B1(n12043), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16460 ( .A1(n13847), .A2(n13333), .B1(n10785), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16461 ( .A1(n13851), .A2(n13332), .B1(n10743), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16462 ( .A1(n10166), .A2(n13333), .B1(n11814), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16463 ( .A1(n10167), .A2(n13332), .B1(n11718), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16464 ( .A1(n13859), .A2(n13332), .B1(n13857), .B2(n11874), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16465 ( .A1(n13863), .A2(n13333), .B1(n13861), .B2(n12817), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  INV_X4 U16466 ( .A(n15473), .ZN(n15475) );
  NAND2_X2 U16467 ( .A1(n13354), .A2(EXEC_MEM_OUT_134), .ZN(n15476) );
  OAI221_X2 U16468 ( .B1(n18106), .B2(n13344), .C1(n12689), .C2(n13349), .A(
        n15476), .ZN(IF_STAGE_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16469 ( .A1(n13746), .A2(n13334), .B1(n11498), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16470 ( .A1(n13753), .A2(n13334), .B1(n13750), .B2(n12480), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16471 ( .A1(n10162), .A2(n13334), .B1(n11719), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16472 ( .A1(n13758), .A2(n13334), .B1(n13757), .B2(n10760), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16473 ( .A1(n10163), .A2(n13334), .B1(n11766), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16474 ( .A1(n13764), .A2(n13334), .B1(n10795), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16475 ( .A1(n13768), .A2(n13334), .B1(n11890), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16476 ( .A1(n10164), .A2(n13334), .B1(n12907), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16477 ( .A1(n13774), .A2(n13334), .B1(n13772), .B2(n10714), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16478 ( .A1(n13779), .A2(n13334), .B1(n13776), .B2(n12481), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16479 ( .A1(n787), .A2(n13334), .B1(n13781), .B2(n10343), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16480 ( .A1(n13786), .A2(n13335), .B1(n11720), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16481 ( .A1(n13790), .A2(n13335), .B1(n12141), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16482 ( .A1(n13795), .A2(n13335), .B1(n10295), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16483 ( .A1(n13799), .A2(n13335), .B1(n13798), .B2(n10535), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16484 ( .A1(n13804), .A2(n13335), .B1(n13803), .B2(n12760), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16485 ( .A1(n13809), .A2(n13335), .B1(n13807), .B2(n12482), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16486 ( .A1(n13813), .A2(n13335), .B1(n12579), .B2(n13811), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16487 ( .A1(n13817), .A2(n13335), .B1(n12594), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16488 ( .A1(n13821), .A2(n13335), .B1(n12265), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16489 ( .A1(n13825), .A2(n13335), .B1(n10921), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16490 ( .A1(n13829), .A2(n13335), .B1(n11424), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16491 ( .A1(n13833), .A2(n13334), .B1(n10524), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16492 ( .A1(n13837), .A2(n13335), .B1(n12779), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16493 ( .A1(n10165), .A2(n13335), .B1(n12908), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16494 ( .A1(n272), .A2(n13334), .B1(n12044), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16495 ( .A1(n13847), .A2(n13335), .B1(n10786), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16496 ( .A1(n13851), .A2(n13334), .B1(n10744), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16497 ( .A1(n10166), .A2(n13335), .B1(n11815), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16498 ( .A1(n10167), .A2(n13334), .B1(n11721), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16499 ( .A1(n13859), .A2(n13334), .B1(n13858), .B2(n11875), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16500 ( .A1(n27), .A2(n13335), .B1(n13862), .B2(n12818), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16501 ( .A1(n13354), .A2(EXEC_MEM_OUT_135), .ZN(n15477) );
  OAI221_X2 U16502 ( .B1(n18151), .B2(n13344), .C1(n12552), .C2(n13349), .A(
        n15477), .ZN(IF_STAGE_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16503 ( .A1(n13746), .A2(n13336), .B1(n11499), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16504 ( .A1(n13753), .A2(n13336), .B1(n13751), .B2(n12483), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16505 ( .A1(n10162), .A2(n13336), .B1(n11722), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16506 ( .A1(n13758), .A2(n13336), .B1(n13757), .B2(n10761), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16507 ( .A1(n10163), .A2(n13336), .B1(n11767), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16508 ( .A1(n13764), .A2(n13336), .B1(n10796), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16509 ( .A1(n13768), .A2(n13336), .B1(n11891), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16510 ( .A1(n10164), .A2(n13336), .B1(n12909), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16511 ( .A1(n13774), .A2(n13336), .B1(n13773), .B2(n12277), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16512 ( .A1(n13779), .A2(n13336), .B1(n13777), .B2(n12484), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16513 ( .A1(n787), .A2(n13336), .B1(n13781), .B2(n10344), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16514 ( .A1(n13786), .A2(n13337), .B1(n11723), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16515 ( .A1(n13790), .A2(n13337), .B1(n12142), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16516 ( .A1(n13794), .A2(n13337), .B1(n10296), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16517 ( .A1(n13800), .A2(n13337), .B1(n13797), .B2(n10536), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16518 ( .A1(n13805), .A2(n13337), .B1(n13802), .B2(n12761), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16519 ( .A1(n13809), .A2(n13337), .B1(n13808), .B2(n12485), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16520 ( .A1(n13813), .A2(n13337), .B1(n12580), .B2(n13811), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16521 ( .A1(n13817), .A2(n13337), .B1(n12595), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16522 ( .A1(n13821), .A2(n13337), .B1(n12266), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16523 ( .A1(n13825), .A2(n13337), .B1(n10922), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16524 ( .A1(n13829), .A2(n13337), .B1(n11425), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16525 ( .A1(n13833), .A2(n13336), .B1(n10525), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16526 ( .A1(n13837), .A2(n13337), .B1(n12780), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16527 ( .A1(n10165), .A2(n13337), .B1(n12910), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16528 ( .A1(n272), .A2(n13336), .B1(n12045), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16529 ( .A1(n13847), .A2(n13337), .B1(n10787), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16530 ( .A1(n13851), .A2(n13336), .B1(n10745), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16531 ( .A1(n10166), .A2(n13337), .B1(n11816), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16532 ( .A1(n10167), .A2(n13336), .B1(n11724), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16533 ( .A1(n13859), .A2(n13336), .B1(n13857), .B2(n11876), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16534 ( .A1(n13863), .A2(n13337), .B1(n13861), .B2(n12819), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16535 ( .A1(n13746), .A2(n13338), .B1(n11500), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16536 ( .A1(n13753), .A2(n13338), .B1(n13751), .B2(n12486), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16537 ( .A1(n10162), .A2(n13338), .B1(n11725), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16538 ( .A1(n13758), .A2(n13338), .B1(n13757), .B2(n10762), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16539 ( .A1(n10163), .A2(n13338), .B1(n11768), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16540 ( .A1(n13764), .A2(n13338), .B1(n10797), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16541 ( .A1(n13768), .A2(n13338), .B1(n11892), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16542 ( .A1(n10164), .A2(n13338), .B1(n12911), .B2(n13771), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16543 ( .A1(n13774), .A2(n13338), .B1(n13773), .B2(n10715), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16544 ( .A1(n13779), .A2(n13338), .B1(n13777), .B2(n12487), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16545 ( .A1(n787), .A2(n13338), .B1(n13781), .B2(n10345), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16546 ( .A1(n13786), .A2(n13339), .B1(n11726), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16547 ( .A1(n13790), .A2(n13339), .B1(n12143), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16548 ( .A1(n13795), .A2(n13339), .B1(n10297), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16549 ( .A1(n13800), .A2(n13339), .B1(n13798), .B2(n10537), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16550 ( .A1(n13805), .A2(n13339), .B1(n13803), .B2(n12762), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16551 ( .A1(n13809), .A2(n13339), .B1(n13807), .B2(n12488), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16552 ( .A1(n13813), .A2(n13339), .B1(n12581), .B2(n13811), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16553 ( .A1(n13817), .A2(n13339), .B1(n12596), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16554 ( .A1(n13821), .A2(n13339), .B1(n12267), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16555 ( .A1(n13825), .A2(n13339), .B1(n10923), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16556 ( .A1(n13829), .A2(n13339), .B1(n11426), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16557 ( .A1(n13833), .A2(n13338), .B1(n10526), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16558 ( .A1(n13837), .A2(n13339), .B1(n12781), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16559 ( .A1(n10165), .A2(n13339), .B1(n12912), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16560 ( .A1(n272), .A2(n13338), .B1(n12046), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16561 ( .A1(n13847), .A2(n13339), .B1(n10788), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16562 ( .A1(n13851), .A2(n13338), .B1(n10746), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16563 ( .A1(n10166), .A2(n13339), .B1(n11817), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16564 ( .A1(n10167), .A2(n13338), .B1(n11727), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16565 ( .A1(n13859), .A2(n13338), .B1(n13858), .B2(n11877), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16566 ( .A1(n13863), .A2(n13339), .B1(n13862), .B2(n12820), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16567 ( .A1(n15479), .A2(n15478), .ZN(n15482) );
  NAND2_X2 U16568 ( .A1(n15482), .A2(n15481), .ZN(n18194) );
  NAND2_X2 U16569 ( .A1(n13354), .A2(EXEC_MEM_OUT_136), .ZN(n15483) );
  OAI221_X2 U16570 ( .B1(n18194), .B2(n13344), .C1(n15478), .C2(n13349), .A(
        n15483), .ZN(IF_STAGE_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16571 ( .A1(n13746), .A2(n13340), .B1(n11501), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16572 ( .A1(n13753), .A2(n13340), .B1(n13751), .B2(n12489), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16573 ( .A1(n10162), .A2(n13340), .B1(n11728), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16574 ( .A1(n13758), .A2(n13340), .B1(n13757), .B2(n10763), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16575 ( .A1(n10163), .A2(n13340), .B1(n11769), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16576 ( .A1(n13764), .A2(n13340), .B1(n10798), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16577 ( .A1(n13768), .A2(n13340), .B1(n11893), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16578 ( .A1(n10164), .A2(n13340), .B1(n12913), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16579 ( .A1(n13774), .A2(n13340), .B1(n13773), .B2(n12278), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16580 ( .A1(n13779), .A2(n13340), .B1(n13777), .B2(n12490), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16581 ( .A1(n787), .A2(n13340), .B1(n13781), .B2(n10346), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16582 ( .A1(n13786), .A2(n13341), .B1(n11729), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16583 ( .A1(n13790), .A2(n13341), .B1(n12144), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16584 ( .A1(n13794), .A2(n13341), .B1(n10298), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16585 ( .A1(n13799), .A2(n13341), .B1(n13797), .B2(n10538), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16586 ( .A1(n13804), .A2(n13341), .B1(n13802), .B2(n12763), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16587 ( .A1(n13809), .A2(n13341), .B1(n13808), .B2(n12491), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16588 ( .A1(n13813), .A2(n13341), .B1(n12582), .B2(n13811), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16589 ( .A1(n13817), .A2(n13341), .B1(n12597), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16590 ( .A1(n13821), .A2(n13341), .B1(n12268), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16591 ( .A1(n13825), .A2(n13341), .B1(n10924), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16592 ( .A1(n13829), .A2(n13341), .B1(n11427), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16593 ( .A1(n13833), .A2(n13340), .B1(n10527), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16594 ( .A1(n13837), .A2(n13341), .B1(n12782), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16595 ( .A1(n10165), .A2(n13341), .B1(n12914), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16596 ( .A1(n13843), .A2(n13340), .B1(n12047), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16597 ( .A1(n13847), .A2(n13341), .B1(n10789), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16598 ( .A1(n13851), .A2(n13340), .B1(n10747), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16599 ( .A1(n10166), .A2(n13341), .B1(n11818), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16600 ( .A1(n10167), .A2(n13340), .B1(n11730), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16601 ( .A1(n13859), .A2(n13340), .B1(n13857), .B2(n11878), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16602 ( .A1(n13863), .A2(n13341), .B1(n13861), .B2(n12821), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16603 ( .A1(n13354), .A2(EXEC_MEM_OUT_137), .ZN(n15484) );
  OAI221_X2 U16604 ( .B1(n18237), .B2(n13344), .C1(n12553), .C2(n13349), .A(
        n15484), .ZN(IF_STAGE_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16605 ( .A1(n13746), .A2(n13342), .B1(n11502), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16606 ( .A1(n13753), .A2(n13342), .B1(n13751), .B2(n12492), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16607 ( .A1(n10162), .A2(n13342), .B1(n11731), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16608 ( .A1(n13758), .A2(n13342), .B1(n13757), .B2(n10764), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16609 ( .A1(n10163), .A2(n13342), .B1(n11770), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16610 ( .A1(n13764), .A2(n13342), .B1(n10799), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16611 ( .A1(n13768), .A2(n13342), .B1(n11894), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16612 ( .A1(n10164), .A2(n13342), .B1(n12915), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16613 ( .A1(n13774), .A2(n13342), .B1(n13773), .B2(n10716), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16614 ( .A1(n13779), .A2(n13342), .B1(n13777), .B2(n12493), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16615 ( .A1(n787), .A2(n13342), .B1(n13781), .B2(n10347), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16616 ( .A1(n13786), .A2(n13343), .B1(n11732), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16617 ( .A1(n13790), .A2(n13343), .B1(n12145), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16618 ( .A1(n13795), .A2(n13343), .B1(n10299), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16619 ( .A1(n13799), .A2(n13343), .B1(n13798), .B2(n10539), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16620 ( .A1(n13804), .A2(n13343), .B1(n13803), .B2(n12764), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16621 ( .A1(n13809), .A2(n13343), .B1(n13807), .B2(n12494), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16622 ( .A1(n13813), .A2(n13343), .B1(n12583), .B2(n13811), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16623 ( .A1(n13817), .A2(n13343), .B1(n12598), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16624 ( .A1(n13821), .A2(n13343), .B1(n12269), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16625 ( .A1(n13825), .A2(n13343), .B1(n10925), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16626 ( .A1(n13829), .A2(n13343), .B1(n11428), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16627 ( .A1(n13833), .A2(n13342), .B1(n10528), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16628 ( .A1(n13837), .A2(n13343), .B1(n12783), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16629 ( .A1(n10165), .A2(n13343), .B1(n12916), .B2(n13839), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16630 ( .A1(n13843), .A2(n13342), .B1(n12048), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16631 ( .A1(n13847), .A2(n13343), .B1(n10790), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16632 ( .A1(n13851), .A2(n13342), .B1(n10748), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16633 ( .A1(n10166), .A2(n13343), .B1(n11819), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16634 ( .A1(n10167), .A2(n13342), .B1(n11733), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16635 ( .A1(n13859), .A2(n13342), .B1(n13858), .B2(n11879), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16636 ( .A1(n13863), .A2(n13343), .B1(n13862), .B2(n12822), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U16637 ( .A1(n13354), .A2(EXEC_MEM_OUT_138), .ZN(n15487) );
  MUX2_X2 U16638 ( .A(n13344), .B(n13350), .S(IMEM_BUS_OUT[29]), .Z(n15486) );
  NAND2_X2 U16639 ( .A1(n15487), .A2(n15486), .ZN(
        IF_STAGE_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16640 ( .A1(n13746), .A2(n13347), .B1(n11503), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16641 ( .A1(n13753), .A2(n13347), .B1(n13751), .B2(n12495), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16642 ( .A1(n10162), .A2(n13347), .B1(n11734), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16643 ( .A1(n13758), .A2(n13347), .B1(n13757), .B2(n10765), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16644 ( .A1(n10163), .A2(n13347), .B1(n11771), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16645 ( .A1(n13764), .A2(n13347), .B1(n10800), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16646 ( .A1(n13768), .A2(n13347), .B1(n11895), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16647 ( .A1(n10164), .A2(n13347), .B1(n12917), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16648 ( .A1(n13774), .A2(n13347), .B1(n13773), .B2(n10717), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16649 ( .A1(n13779), .A2(n13347), .B1(n13777), .B2(n12496), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16650 ( .A1(n787), .A2(n13347), .B1(n13781), .B2(n10348), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16651 ( .A1(n13786), .A2(n13348), .B1(n11735), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16652 ( .A1(n13790), .A2(n13348), .B1(n12146), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16653 ( .A1(n13794), .A2(n13348), .B1(n10300), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16654 ( .A1(n13800), .A2(n13348), .B1(n13797), .B2(n10540), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16655 ( .A1(n13805), .A2(n13348), .B1(n13802), .B2(n12765), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16656 ( .A1(n13809), .A2(n13348), .B1(n13808), .B2(n12497), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16657 ( .A1(n13813), .A2(n13348), .B1(n12584), .B2(n13811), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16658 ( .A1(n13817), .A2(n13348), .B1(n12599), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16659 ( .A1(n13821), .A2(n13348), .B1(n12270), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16660 ( .A1(n13825), .A2(n13348), .B1(n10926), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16661 ( .A1(n13829), .A2(n13348), .B1(n11429), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16662 ( .A1(n13833), .A2(n13347), .B1(n10529), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16663 ( .A1(n13837), .A2(n13348), .B1(n12784), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16664 ( .A1(n10165), .A2(n13348), .B1(n12918), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16665 ( .A1(n13843), .A2(n13347), .B1(n12049), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16666 ( .A1(n13847), .A2(n13348), .B1(n10791), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16667 ( .A1(n13851), .A2(n13347), .B1(n10749), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16668 ( .A1(n10166), .A2(n13348), .B1(n11820), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16669 ( .A1(n10167), .A2(n13347), .B1(n11736), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16670 ( .A1(n13859), .A2(n13347), .B1(n13857), .B2(n11880), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16671 ( .A1(n13863), .A2(n13348), .B1(n13861), .B2(n12823), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI21_X4 U16672 ( .B1(EXEC_MEM_OUT_141), .B2(n13956), .A(n13349), .ZN(n15489) );
  OAI22_X2 U16673 ( .A1(n11504), .A2(n13355), .B1(n12311), .B2(n15491), .ZN(
        n10104) );
  OAI22_X2 U16674 ( .A1(n13746), .A2(n13352), .B1(n12135), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16675 ( .A1(n13753), .A2(n13352), .B1(n13750), .B2(n12766), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16676 ( .A1(n10162), .A2(n13352), .B1(n12412), .B2(n13754), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16677 ( .A1(n13758), .A2(n13352), .B1(n13757), .B2(n10766), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16678 ( .A1(n10163), .A2(n13352), .B1(n12088), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16679 ( .A1(n13764), .A2(n13352), .B1(n12063), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16680 ( .A1(n13768), .A2(n13352), .B1(n10689), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16681 ( .A1(n10164), .A2(n13352), .B1(n12919), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16682 ( .A1(n13774), .A2(n13352), .B1(n13772), .B2(n10718), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16683 ( .A1(n13779), .A2(n13352), .B1(n13776), .B2(n11469), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16684 ( .A1(n787), .A2(n13352), .B1(n13781), .B2(n10257), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16685 ( .A1(n13786), .A2(n13353), .B1(n12411), .B2(n13784), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16686 ( .A1(n13790), .A2(n13353), .B1(n12062), .B2(n13788), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16687 ( .A1(n13795), .A2(n13353), .B1(n10251), .B2(n13792), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16688 ( .A1(n13800), .A2(n13353), .B1(n13798), .B2(n10367), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16689 ( .A1(n13805), .A2(n13353), .B1(n13803), .B2(n12498), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16690 ( .A1(n13809), .A2(n13353), .B1(n13807), .B2(n10750), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16691 ( .A1(n13813), .A2(n13353), .B1(n12643), .B2(n13812), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16692 ( .A1(n13817), .A2(n13353), .B1(n12666), .B2(n13816), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16693 ( .A1(n13821), .A2(n13353), .B1(n12081), .B2(n13819), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16694 ( .A1(n13825), .A2(n13353), .B1(n10847), .B2(n13823), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16695 ( .A1(n13829), .A2(n13353), .B1(n11430), .B2(n13827), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16696 ( .A1(n13833), .A2(n13352), .B1(n10530), .B2(n13831), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16697 ( .A1(n13837), .A2(n13353), .B1(n12785), .B2(n13835), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16698 ( .A1(n10165), .A2(n13353), .B1(n12920), .B2(n13840), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16699 ( .A1(n13843), .A2(n13352), .B1(n12025), .B2(n13841), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16700 ( .A1(n13847), .A2(n13353), .B1(n12177), .B2(n13845), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16701 ( .A1(n13851), .A2(n13352), .B1(n10461), .B2(n13849), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16702 ( .A1(n10166), .A2(n13353), .B1(n12298), .B2(n13853), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16703 ( .A1(n10167), .A2(n13352), .B1(n11846), .B2(n13855), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16704 ( .A1(n13859), .A2(n13352), .B1(n13858), .B2(n12079), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16705 ( .A1(n13863), .A2(n13353), .B1(n13862), .B2(n12824), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U16706 ( .A1(n11505), .A2(n13355), .B1(n12312), .B2(n15491), .ZN(
        n10105) );
  XNOR2_X2 U16707 ( .A(ID_EXEC_OUT[202]), .B(MEM_WB_REG_MEM_WB_REG_N144), .ZN(
        n15496) );
  NAND3_X4 U16708 ( .A1(n15496), .A2(n15495), .A3(n15494), .ZN(n15497) );
  NAND2_X2 U16709 ( .A1(n13411), .A2(ID_EXEC_OUT[160]), .ZN(n15513) );
  NAND2_X2 U16710 ( .A1(DMEM_BUS_OUT[32]), .A2(net231321), .ZN(n15512) );
  INV_X4 U16711 ( .A(n15506), .ZN(n15507) );
  NAND2_X2 U16712 ( .A1(n13414), .A2(DMEM_BUS_OUT[0]), .ZN(n15511) );
  INV_X4 U16713 ( .A(n12040), .ZN(n15509) );
  NAND2_X2 U16714 ( .A1(n13415), .A2(n15509), .ZN(n15510) );
  NAND4_X2 U16715 ( .A1(n15513), .A2(n15512), .A3(n15511), .A4(n15510), .ZN(
        n7294) );
  NAND2_X2 U16716 ( .A1(n13409), .A2(n13149), .ZN(n15514) );
  OAI211_X2 U16717 ( .C1(n12170), .C2(net231227), .A(n15514), .B(n6754), .ZN(
        n7298) );
  NAND2_X2 U16718 ( .A1(n13410), .A2(n18922), .ZN(n15515) );
  OAI211_X2 U16719 ( .C1(n12169), .C2(net231227), .A(n15515), .B(n6756), .ZN(
        n7302) );
  NAND2_X2 U16720 ( .A1(n13410), .A2(n18911), .ZN(n15516) );
  OAI211_X2 U16721 ( .C1(n12165), .C2(net231225), .A(n15516), .B(n6761), .ZN(
        n7306) );
  NAND2_X2 U16722 ( .A1(n13409), .A2(n18980), .ZN(n15517) );
  OAI211_X2 U16723 ( .C1(n12168), .C2(net231223), .A(n15517), .B(n6757), .ZN(
        n7310) );
  NAND2_X2 U16724 ( .A1(n13410), .A2(n17712), .ZN(n15518) );
  OAI211_X2 U16725 ( .C1(n12167), .C2(net231225), .A(n15518), .B(n6759), .ZN(
        n7314) );
  NAND2_X2 U16726 ( .A1(n13412), .A2(ID_EXEC_OUT[163]), .ZN(n15522) );
  NAND2_X2 U16727 ( .A1(DMEM_BUS_OUT[35]), .A2(net231321), .ZN(n15521) );
  NAND2_X2 U16728 ( .A1(n13414), .A2(DMEM_BUS_OUT[3]), .ZN(n15520) );
  NAND2_X2 U16729 ( .A1(n13415), .A2(MEM_WB_OUT[40]), .ZN(n15519) );
  NAND4_X2 U16730 ( .A1(n15522), .A2(n15521), .A3(n15520), .A4(n15519), .ZN(
        n7315) );
  NAND2_X2 U16731 ( .A1(n13409), .A2(n17505), .ZN(n15523) );
  OAI211_X2 U16732 ( .C1(n12166), .C2(net231225), .A(n15523), .B(n6760), .ZN(
        n7319) );
  NAND2_X2 U16733 ( .A1(n13411), .A2(ID_EXEC_OUT[164]), .ZN(n15527) );
  NAND2_X2 U16734 ( .A1(DMEM_BUS_OUT[36]), .A2(net231321), .ZN(n15526) );
  NAND2_X2 U16735 ( .A1(n13413), .A2(DMEM_BUS_OUT[4]), .ZN(n15525) );
  NAND2_X2 U16736 ( .A1(n13415), .A2(MEM_WB_OUT[41]), .ZN(n15524) );
  NAND4_X2 U16737 ( .A1(n15527), .A2(n15526), .A3(n15525), .A4(n15524), .ZN(
        n7320) );
  NAND2_X2 U16738 ( .A1(n13410), .A2(n18867), .ZN(n15528) );
  OAI211_X2 U16739 ( .C1(n12150), .C2(net231225), .A(n15528), .B(n6778), .ZN(
        n7324) );
  INV_X4 U16740 ( .A(net225906), .ZN(net227046) );
  AOI21_X4 U16741 ( .B1(net232881), .B2(n12065), .A(n10369), .ZN(net225529) );
  MUX2_X2 U16742 ( .A(n11565), .B(n12562), .S(net239627), .Z(net223589) );
  OAI21_X4 U16743 ( .B1(net239782), .B2(n13042), .A(n15529), .ZN(net223365) );
  INV_X4 U16744 ( .A(net239527), .ZN(net227269) );
  NAND2_X2 U16745 ( .A1(nextPC_ex_out[24]), .A2(nextPC_ex_out[26]), .ZN(
        net227241) );
  INV_X4 U16746 ( .A(net227241), .ZN(net227240) );
  MUX2_X2 U16747 ( .A(n11566), .B(n12563), .S(net239782), .Z(net223743) );
  INV_X4 U16748 ( .A(net227236), .ZN(net227233) );
  NAND3_X4 U16749 ( .A1(net227213), .A2(n15537), .A3(net227233), .ZN(net227164) );
  NAND3_X4 U16750 ( .A1(net233181), .A2(net227232), .A3(net227233), .ZN(
        net227163) );
  MUX2_X2 U16751 ( .A(n11567), .B(n12564), .S(net239782), .Z(net223985) );
  INV_X4 U16752 ( .A(net223985), .ZN(net227177) );
  NOR2_X4 U16753 ( .A1(nextPC_ex_out[20]), .A2(net227177), .ZN(n15540) );
  INV_X4 U16754 ( .A(n15535), .ZN(n15545) );
  OAI21_X4 U16755 ( .B1(n15539), .B2(n13111), .A(net223743), .ZN(net223797) );
  NAND2_X2 U16756 ( .A1(nextPC_ex_out[21]), .A2(nextPC_ex_out[22]), .ZN(
        net227150) );
  INV_X4 U16757 ( .A(net227187), .ZN(net227182) );
  INV_X4 U16758 ( .A(net223743), .ZN(net227198) );
  NOR3_X4 U16759 ( .A1(n15541), .A2(net227197), .A3(net227198), .ZN(n17673) );
  NAND2_X2 U16760 ( .A1(nextPC_ex_out[21]), .A2(nextPC_ex_out[23]), .ZN(n15542) );
  NOR2_X4 U16761 ( .A1(net227165), .A2(n12558), .ZN(net227183) );
  NOR2_X4 U16762 ( .A1(n13065), .A2(net227170), .ZN(n15546) );
  INV_X4 U16763 ( .A(net227167), .ZN(net227169) );
  AOI21_X4 U16764 ( .B1(n15546), .B2(n17675), .A(net227169), .ZN(net227159) );
  NOR2_X4 U16765 ( .A1(net227165), .A2(net227166), .ZN(net227160) );
  MUX2_X2 U16766 ( .A(n11568), .B(n12565), .S(net239782), .Z(net224493) );
  NAND2_X2 U16767 ( .A1(net224493), .A2(net227135), .ZN(n15547) );
  MUX2_X2 U16768 ( .A(n12072), .B(n12551), .S(net239782), .Z(net227117) );
  NAND3_X4 U16769 ( .A1(n15552), .A2(net227115), .A3(net227116), .ZN(net227108) );
  MUX2_X2 U16770 ( .A(n11569), .B(n12566), .S(net239782), .Z(net227110) );
  NAND2_X2 U16771 ( .A1(n16969), .A2(n10366), .ZN(net225187) );
  INV_X4 U16772 ( .A(n16969), .ZN(n15553) );
  NAND2_X2 U16773 ( .A1(n15553), .A2(nextPC_ex_out[7]), .ZN(net225188) );
  INV_X4 U16774 ( .A(net225187), .ZN(net225191) );
  INV_X4 U16775 ( .A(n15554), .ZN(n15642) );
  NAND2_X2 U16776 ( .A1(net227035), .A2(n17215), .ZN(n15556) );
  INV_X4 U16777 ( .A(n15556), .ZN(n15564) );
  NAND2_X2 U16778 ( .A1(nextPC_ex_out[2]), .A2(nextPC_ex_out[3]), .ZN(n15645)
         );
  NOR2_X4 U16779 ( .A1(n15564), .A2(n15645), .ZN(n15561) );
  INV_X4 U16780 ( .A(net224713), .ZN(net224711) );
  NAND2_X2 U16781 ( .A1(net224711), .A2(nextPC_ex_out[1]), .ZN(n15652) );
  NAND2_X2 U16782 ( .A1(net224704), .A2(n10362), .ZN(n15647) );
  NAND2_X2 U16783 ( .A1(nextPC_ex_out[0]), .A2(net224711), .ZN(n15557) );
  INV_X4 U16784 ( .A(n15563), .ZN(n15558) );
  NAND2_X2 U16785 ( .A1(n15570), .A2(net226995), .ZN(net227020) );
  NOR2_X4 U16786 ( .A1(n10132), .A2(net231915), .ZN(n15578) );
  NAND2_X2 U16787 ( .A1(EXEC_MEM_OUT_109), .A2(net231323), .ZN(n15567) );
  OAI211_X2 U16788 ( .C1(n16791), .C2(net223104), .A(n15568), .B(n15567), .ZN(
        n15569) );
  INV_X4 U16789 ( .A(n15569), .ZN(n15575) );
  INV_X4 U16790 ( .A(n15570), .ZN(n15571) );
  NAND2_X2 U16791 ( .A1(n10361), .A2(n15571), .ZN(n15573) );
  INV_X4 U16792 ( .A(net226995), .ZN(net224848) );
  NAND2_X2 U16793 ( .A1(n10361), .A2(net224848), .ZN(n15572) );
  NAND2_X2 U16794 ( .A1(nextPC_ex_out[0]), .A2(n10362), .ZN(n15574) );
  NAND2_X2 U16795 ( .A1(n15575), .A2(n15574), .ZN(n15576) );
  NOR4_X2 U16796 ( .A1(n15582), .A2(n11583), .A3(n5467), .A4(n5466), .ZN(
        n15597) );
  NOR3_X4 U16797 ( .A1(n15597), .A2(n11922), .A3(n18813), .ZN(n15613) );
  OAI22_X2 U16798 ( .A1(n13419), .A2(n12786), .B1(n13417), .B2(n11847), .ZN(
        n15587) );
  NOR3_X4 U16799 ( .A1(n15597), .A2(n10824), .A3(offset_26_id[6]), .ZN(n15617)
         );
  OAI22_X2 U16800 ( .A1(n13424), .A2(n12826), .B1(n13422), .B2(n12825), .ZN(
        n15586) );
  NOR3_X4 U16801 ( .A1(n15597), .A2(n11922), .A3(n10824), .ZN(n15620) );
  NAND2_X2 U16802 ( .A1(n15609), .A2(n15617), .ZN(n15583) );
  INV_X4 U16803 ( .A(n15583), .ZN(n18690) );
  NAND2_X2 U16804 ( .A1(REG_FILE_reg_out_17__0_), .A2(n13436), .ZN(n15584) );
  OAI221_X2 U16805 ( .B1(n13432), .B2(n12827), .C1(n13427), .C2(n12721), .A(
        n15584), .ZN(n15585) );
  NAND2_X2 U16806 ( .A1(n15620), .A2(n15609), .ZN(n18697) );
  AOI22_X2 U16807 ( .A1(REG_FILE_reg_out_25__0_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__0_), .B2(n13441), .ZN(n15595) );
  NAND2_X2 U16808 ( .A1(n15616), .A2(n15620), .ZN(n18698) );
  NOR3_X4 U16809 ( .A1(n15597), .A2(n18813), .A3(offset_26_id[6]), .ZN(n15610)
         );
  OAI22_X2 U16810 ( .A1(n12383), .A2(n13444), .B1(n10505), .B2(n13442), .ZN(
        n15590) );
  OAI22_X2 U16811 ( .A1(n10301), .A2(n13190), .B1(n10690), .B2(n18699), .ZN(
        n15589) );
  OAI22_X2 U16812 ( .A1(n11838), .A2(n13192), .B1(n12382), .B2(n13193), .ZN(
        n15588) );
  NAND2_X2 U16813 ( .A1(n15621), .A2(n15610), .ZN(n18705) );
  NAND4_X2 U16814 ( .A1(n15596), .A2(n15595), .A3(n15594), .A4(n15593), .ZN(
        n15630) );
  INV_X4 U16815 ( .A(n15597), .ZN(n18713) );
  NAND2_X2 U16816 ( .A1(n13456), .A2(REG_FILE_reg_out_12__0_), .ZN(n15606) );
  NAND2_X2 U16817 ( .A1(n10241), .A2(n15620), .ZN(n18718) );
  NAND2_X2 U16818 ( .A1(n10241), .A2(n15613), .ZN(n18721) );
  AOI22_X2 U16819 ( .A1(n13464), .A2(REG_FILE_reg_out_0__0_), .B1(
        REG_FILE_reg_out_15__0_), .B2(n13466), .ZN(n15604) );
  NAND4_X2 U16820 ( .A1(n15607), .A2(n15606), .A3(n15605), .A4(n15604), .ZN(
        n15629) );
  NAND2_X2 U16821 ( .A1(n15616), .A2(n15617), .ZN(n18733) );
  NAND4_X2 U16822 ( .A1(n15627), .A2(n15626), .A3(n15625), .A4(n15624), .ZN(
        n15628) );
  NOR3_X4 U16823 ( .A1(n15630), .A2(n15629), .A3(n15628), .ZN(n15636) );
  OAI22_X2 U16824 ( .A1(n11506), .A2(net231253), .B1(net230381), .B2(n15636), 
        .ZN(n7326) );
  NAND2_X2 U16825 ( .A1(n13166), .A2(net230387), .ZN(n18188) );
  INV_X4 U16826 ( .A(n18188), .ZN(n15632) );
  NAND2_X2 U16827 ( .A1(n13205), .A2(ID_STAGE_imm16_aluA[16]), .ZN(n16766) );
  NAND2_X2 U16828 ( .A1(ID_EXEC_OUT[64]), .A2(net231319), .ZN(n15635) );
  OAI211_X2 U16829 ( .C1(n15636), .C2(n13476), .A(n17267), .B(n15635), .ZN(
        n7327) );
  OAI22_X2 U16831 ( .A1(n15638), .A2(net231253), .B1(n13481), .B2(n15637), 
        .ZN(n7332) );
  NAND2_X2 U16832 ( .A1(net224711), .A2(n10362), .ZN(n15640) );
  NAND2_X2 U16833 ( .A1(net224704), .A2(nextPC_ex_out[1]), .ZN(n15639) );
  NAND2_X2 U16834 ( .A1(n15640), .A2(n15639), .ZN(n15643) );
  INV_X4 U16835 ( .A(n15652), .ZN(n15646) );
  NAND2_X2 U16836 ( .A1(n15646), .A2(n15645), .ZN(n15656) );
  NAND2_X2 U16837 ( .A1(n13412), .A2(ID_EXEC_OUT[161]), .ZN(n15661) );
  NAND2_X2 U16838 ( .A1(DMEM_BUS_OUT[33]), .A2(net231321), .ZN(n15660) );
  NAND2_X2 U16839 ( .A1(n13413), .A2(DMEM_BUS_OUT[1]), .ZN(n15659) );
  NAND2_X2 U16840 ( .A1(n13415), .A2(MEM_WB_OUT[38]), .ZN(n15658) );
  NAND4_X2 U16841 ( .A1(n15661), .A2(n15660), .A3(n15659), .A4(n15658), .ZN(
        n7334) );
  INV_X4 U16842 ( .A(n15665), .ZN(n15666) );
  NOR2_X4 U16843 ( .A1(n15668), .A2(n15667), .ZN(n15670) );
  NAND2_X2 U16844 ( .A1(DMEM_BUS_OUT[31]), .A2(n13485), .ZN(n18931) );
  NAND3_X4 U16845 ( .A1(n15673), .A2(n18931), .A3(n15672), .ZN(n19105) );
  NAND2_X2 U16846 ( .A1(n19105), .A2(n11913), .ZN(n17874) );
  INV_X4 U16847 ( .A(n17874), .ZN(n19124) );
  NAND2_X2 U16848 ( .A1(net230393), .A2(n12017), .ZN(n19138) );
  INV_X4 U16849 ( .A(n19138), .ZN(n18669) );
  MUX2_X2 U16850 ( .A(n15675), .B(n15674), .S(ID_EXEC_OUT[157]), .Z(n15676) );
  NAND2_X2 U16851 ( .A1(n18669), .A2(n15676), .ZN(n19104) );
  NAND2_X2 U16852 ( .A1(n13401), .A2(n15678), .ZN(n15679) );
  NAND3_X4 U16853 ( .A1(n15681), .A2(n15680), .A3(n15679), .ZN(n18860) );
  INV_X4 U16854 ( .A(n18860), .ZN(n18945) );
  NAND2_X2 U16855 ( .A1(n18945), .A2(n18373), .ZN(n16007) );
  NAND2_X2 U16856 ( .A1(DMEM_BUS_OUT[29]), .A2(n13484), .ZN(n15688) );
  NAND3_X4 U16857 ( .A1(n15689), .A2(n15688), .A3(n15687), .ZN(n18862) );
  NAND2_X2 U16858 ( .A1(n18271), .A2(n18943), .ZN(n18469) );
  INV_X4 U16859 ( .A(n18469), .ZN(n18309) );
  NAND2_X2 U16860 ( .A1(n18309), .A2(n18873), .ZN(n15699) );
  NAND2_X2 U16861 ( .A1(net232816), .A2(n18980), .ZN(n15692) );
  NAND2_X2 U16862 ( .A1(n13385), .A2(n19038), .ZN(n15691) );
  NAND2_X2 U16863 ( .A1(n18373), .A2(n18860), .ZN(n16797) );
  INV_X4 U16864 ( .A(n16797), .ZN(n16816) );
  NAND2_X2 U16865 ( .A1(n13358), .A2(n18897), .ZN(n17843) );
  NAND2_X2 U16866 ( .A1(net223324), .A2(n13159), .ZN(n15690) );
  NAND4_X2 U16867 ( .A1(n15692), .A2(n15691), .A3(n17843), .A4(n15690), .ZN(
        n17298) );
  INV_X4 U16868 ( .A(n17298), .ZN(n15697) );
  NAND2_X2 U16869 ( .A1(n13358), .A2(n19015), .ZN(n15693) );
  INV_X4 U16870 ( .A(n15693), .ZN(n17517) );
  INV_X4 U16871 ( .A(n18559), .ZN(n18902) );
  MUX2_X2 U16872 ( .A(n15697), .B(n15696), .S(n18943), .Z(n15698) );
  NAND2_X2 U16873 ( .A1(n15699), .A2(n15698), .ZN(n18642) );
  INV_X4 U16874 ( .A(n18642), .ZN(n15709) );
  NAND3_X2 U16875 ( .A1(n18929), .A2(n15700), .A3(n13098), .ZN(n15701) );
  NAND3_X4 U16876 ( .A1(n15703), .A2(n15702), .A3(n15701), .ZN(n18641) );
  NAND2_X2 U16877 ( .A1(n13385), .A2(n19029), .ZN(n16208) );
  NAND2_X2 U16878 ( .A1(net232816), .A2(n13149), .ZN(n15704) );
  NAND3_X4 U16879 ( .A1(n16208), .A2(n18245), .A3(n15704), .ZN(n17299) );
  NAND2_X2 U16880 ( .A1(n13392), .A2(n17299), .ZN(n15708) );
  NAND2_X2 U16881 ( .A1(n18943), .A2(n18641), .ZN(n16060) );
  INV_X4 U16882 ( .A(n16060), .ZN(n18540) );
  NAND2_X2 U16883 ( .A1(net232816), .A2(n17505), .ZN(n15706) );
  NAND2_X2 U16884 ( .A1(n13385), .A2(n18867), .ZN(n16024) );
  NAND2_X2 U16885 ( .A1(n13358), .A2(n19000), .ZN(n17509) );
  NAND2_X2 U16886 ( .A1(net223324), .A2(n13163), .ZN(n15705) );
  NAND4_X2 U16887 ( .A1(n15706), .A2(n16024), .A3(n17509), .A4(n15705), .ZN(
        n18636) );
  NAND2_X2 U16888 ( .A1(n13396), .A2(n18636), .ZN(n15707) );
  NAND2_X2 U16889 ( .A1(n18644), .A2(n16876), .ZN(n15754) );
  NAND2_X2 U16890 ( .A1(n6625), .A2(ID_EXEC_OUT[157]), .ZN(n15711) );
  NAND2_X2 U16891 ( .A1(n15710), .A2(n12030), .ZN(n18668) );
  NAND2_X2 U16892 ( .A1(n15711), .A2(n18668), .ZN(n15714) );
  NAND2_X2 U16893 ( .A1(n17982), .A2(n15718), .ZN(n15717) );
  NAND2_X2 U16894 ( .A1(n13208), .A2(n13356), .ZN(n15713) );
  INV_X4 U16895 ( .A(n15713), .ZN(n17983) );
  NAND2_X2 U16896 ( .A1(n17983), .A2(ID_EXEC_OUT[33]), .ZN(n15716) );
  NAND2_X2 U16897 ( .A1(n12540), .A2(n15714), .ZN(n17870) );
  NAND2_X2 U16898 ( .A1(n18566), .A2(DMEM_BUS_OUT[1]), .ZN(n15715) );
  NAND3_X2 U16899 ( .A1(n15717), .A2(n15716), .A3(n15715), .ZN(n15722) );
  NAND2_X2 U16900 ( .A1(n13484), .A2(DMEM_BUS_OUT[1]), .ZN(n15721) );
  NAND2_X2 U16901 ( .A1(ID_EXEC_OUT[65]), .A2(n13403), .ZN(n15720) );
  NAND2_X2 U16902 ( .A1(n13400), .A2(n15718), .ZN(n15719) );
  NAND3_X4 U16903 ( .A1(n15721), .A2(n15720), .A3(n15719), .ZN(n18869) );
  NAND2_X2 U16904 ( .A1(n15722), .A2(n18869), .ZN(n15753) );
  INV_X4 U16905 ( .A(n19105), .ZN(n15728) );
  NAND2_X2 U16906 ( .A1(n15728), .A2(ID_EXEC_OUT[158]), .ZN(n18003) );
  INV_X4 U16907 ( .A(n18003), .ZN(n15723) );
  NAND2_X2 U16908 ( .A1(n13385), .A2(n18870), .ZN(n15724) );
  NAND2_X2 U16909 ( .A1(n15724), .A2(n16064), .ZN(n17304) );
  INV_X4 U16910 ( .A(n18641), .ZN(n19100) );
  NAND2_X2 U16911 ( .A1(n18943), .A2(n19100), .ZN(n19101) );
  INV_X4 U16912 ( .A(n19101), .ZN(n18340) );
  MUX2_X2 U16913 ( .A(n16879), .B(n17304), .S(n13388), .Z(n16882) );
  INV_X4 U16914 ( .A(n16877), .ZN(n15725) );
  INV_X4 U16915 ( .A(n15726), .ZN(n18678) );
  NAND2_X2 U16916 ( .A1(n19105), .A2(ID_EXEC_OUT[158]), .ZN(n18008) );
  INV_X4 U16917 ( .A(n18008), .ZN(n19088) );
  NAND2_X2 U16918 ( .A1(n13385), .A2(n16971), .ZN(n15731) );
  NAND2_X2 U16919 ( .A1(net223324), .A2(n13151), .ZN(n15730) );
  NAND2_X2 U16920 ( .A1(net232816), .A2(n18922), .ZN(n15729) );
  NAND4_X2 U16921 ( .A1(n15731), .A2(n17992), .A3(n15730), .A4(n15729), .ZN(
        n16883) );
  NAND2_X2 U16922 ( .A1(n13392), .A2(n16883), .ZN(n15747) );
  NAND2_X2 U16924 ( .A1(n13358), .A2(n19013), .ZN(n17125) );
  INV_X4 U16925 ( .A(n19101), .ZN(n15733) );
  NAND2_X2 U16926 ( .A1(n13385), .A2(n18872), .ZN(n15738) );
  NAND2_X2 U16927 ( .A1(n13358), .A2(n19004), .ZN(n17525) );
  NAND2_X2 U16928 ( .A1(net232816), .A2(n18911), .ZN(n15736) );
  NAND4_X2 U16929 ( .A1(n15738), .A2(n17525), .A3(n15737), .A4(n15736), .ZN(
        n16886) );
  INV_X4 U16930 ( .A(n16886), .ZN(n15739) );
  NAND2_X2 U16931 ( .A1(net223324), .A2(n13161), .ZN(n15741) );
  NAND2_X2 U16932 ( .A1(n13359), .A2(net222497), .ZN(n17696) );
  NAND2_X2 U16933 ( .A1(n13385), .A2(net225212), .ZN(n16009) );
  NAND2_X2 U16934 ( .A1(net232816), .A2(n17712), .ZN(n15740) );
  NAND4_X2 U16935 ( .A1(n15741), .A2(n17696), .A3(n16009), .A4(n15740), .ZN(
        n16885) );
  INV_X4 U16936 ( .A(n16885), .ZN(n15742) );
  NAND2_X2 U16937 ( .A1(n19100), .A2(n18862), .ZN(n18637) );
  INV_X4 U16938 ( .A(n18870), .ZN(n17121) );
  NAND2_X2 U16939 ( .A1(n13385), .A2(n15733), .ZN(n18284) );
  OAI22_X2 U16940 ( .A1(n15742), .A2(n18637), .B1(n17121), .B2(n18284), .ZN(
        n15743) );
  NAND3_X4 U16941 ( .A1(n15747), .A2(n15746), .A3(n15745), .ZN(n18643) );
  XNOR2_X2 U16942 ( .A(n18869), .B(n18870), .ZN(n19076) );
  NAND2_X2 U16943 ( .A1(n10398), .A2(n18669), .ZN(n19110) );
  NAND2_X2 U16944 ( .A1(net231319), .A2(DMEM_BUS_OUT[1]), .ZN(n15748) );
  AOI211_X4 U16945 ( .C1(n18360), .C2(n18643), .A(n15750), .B(n15749), .ZN(
        n15751) );
  NAND4_X2 U16946 ( .A1(n15754), .A2(n15753), .A3(n15752), .A4(n15751), .ZN(
        n15932) );
  INV_X4 U16947 ( .A(n15932), .ZN(n15935) );
  NAND2_X2 U16948 ( .A1(ID_EXEC_OUT[69]), .A2(n13403), .ZN(n15757) );
  NAND2_X2 U16949 ( .A1(DMEM_BUS_OUT[5]), .A2(n13484), .ZN(n15756) );
  NAND2_X2 U16950 ( .A1(n13400), .A2(n16031), .ZN(n15755) );
  NAND3_X4 U16951 ( .A1(n15757), .A2(n15756), .A3(n15755), .ZN(net222531) );
  XNOR2_X2 U16952 ( .A(net222531), .B(n13494), .ZN(n15758) );
  XNOR2_X2 U16953 ( .A(n15758), .B(net225212), .ZN(n18611) );
  NAND2_X2 U16954 ( .A1(n15758), .A2(net225212), .ZN(n18601) );
  NAND2_X2 U16955 ( .A1(ID_EXEC_OUT[68]), .A2(n13403), .ZN(n15761) );
  NAND2_X2 U16956 ( .A1(DMEM_BUS_OUT[4]), .A2(n13485), .ZN(n15760) );
  NAND2_X2 U16957 ( .A1(n13400), .A2(n17242), .ZN(n15759) );
  NAND3_X4 U16958 ( .A1(n15761), .A2(n15760), .A3(n15759), .ZN(n18866) );
  XNOR2_X2 U16959 ( .A(n18866), .B(n13493), .ZN(n15923) );
  XNOR2_X2 U16960 ( .A(n15923), .B(n18867), .ZN(n18612) );
  NAND3_X2 U16961 ( .A1(n18929), .A2(n17981), .A3(n13098), .ZN(n15762) );
  NAND3_X4 U16962 ( .A1(n15764), .A2(n15763), .A3(n15762), .ZN(n18921) );
  XNOR2_X2 U16963 ( .A(n18921), .B(n13493), .ZN(n15765) );
  XNOR2_X2 U16964 ( .A(n15765), .B(n18922), .ZN(n17978) );
  NAND3_X4 U16965 ( .A1(n15767), .A2(n15768), .A3(n15766), .ZN(n18979) );
  XNOR2_X2 U16966 ( .A(n18979), .B(n13493), .ZN(n15776) );
  XNOR2_X2 U16967 ( .A(n15776), .B(n18980), .ZN(n17837) );
  INV_X4 U16968 ( .A(n17837), .ZN(n15769) );
  XNOR2_X2 U16969 ( .A(n18924), .B(n13493), .ZN(n15778) );
  NAND2_X2 U16970 ( .A1(n15778), .A2(n13149), .ZN(n17834) );
  NAND2_X2 U16971 ( .A1(n17834), .A2(n17835), .ZN(n15774) );
  XNOR2_X2 U16972 ( .A(n15778), .B(n13149), .ZN(n18306) );
  NAND2_X2 U16973 ( .A1(ID_EXEC_OUT[85]), .A2(n13403), .ZN(n15784) );
  NAND2_X2 U16974 ( .A1(DMEM_BUS_OUT[21]), .A2(n13484), .ZN(n15783) );
  NAND2_X2 U16975 ( .A1(n13400), .A2(n17622), .ZN(n15782) );
  NAND3_X4 U16976 ( .A1(n15784), .A2(n15783), .A3(n15782), .ZN(n18985) );
  XNOR2_X2 U16977 ( .A(n18985), .B(n13493), .ZN(n15794) );
  XNOR2_X2 U16978 ( .A(n15794), .B(n17712), .ZN(n17711) );
  INV_X4 U16979 ( .A(n17711), .ZN(n15793) );
  XNOR2_X2 U16981 ( .A(n18385), .B(n13493), .ZN(n15792) );
  INV_X4 U16982 ( .A(n18395), .ZN(n17499) );
  NAND2_X2 U16983 ( .A1(n17499), .A2(n15793), .ZN(n15795) );
  NAND2_X2 U16984 ( .A1(n15794), .A2(n17712), .ZN(n17895) );
  NAND2_X2 U16985 ( .A1(ID_EXEC_OUT[84]), .A2(n13403), .ZN(n15799) );
  NAND2_X2 U16986 ( .A1(DMEM_BUS_OUT[20]), .A2(n13484), .ZN(n15798) );
  NAND2_X2 U16987 ( .A1(n13400), .A2(n17546), .ZN(n15797) );
  NAND3_X4 U16988 ( .A1(n15799), .A2(n15798), .A3(n15797), .ZN(n18991) );
  XNOR2_X2 U16989 ( .A(n18991), .B(n13493), .ZN(n15802) );
  XNOR2_X2 U16990 ( .A(n15802), .B(n17505), .ZN(n17503) );
  INV_X4 U16991 ( .A(n17503), .ZN(n15800) );
  NAND2_X2 U16992 ( .A1(n15802), .A2(n17505), .ZN(n17897) );
  NAND2_X2 U16993 ( .A1(ID_EXEC_OUT[83]), .A2(n13403), .ZN(n15805) );
  NAND2_X2 U16994 ( .A1(DMEM_BUS_OUT[19]), .A2(n13484), .ZN(n15804) );
  NAND2_X2 U16995 ( .A1(n13400), .A2(n17382), .ZN(n15803) );
  XNOR2_X2 U16996 ( .A(n18914), .B(n13494), .ZN(n15851) );
  XNOR2_X2 U16997 ( .A(n15851), .B(n18911), .ZN(n17901) );
  INV_X4 U16998 ( .A(n17901), .ZN(n16780) );
  NAND2_X2 U16999 ( .A1(ID_EXEC_OUT[82]), .A2(n13403), .ZN(n15808) );
  NAND2_X2 U17000 ( .A1(DMEM_BUS_OUT[18]), .A2(n13484), .ZN(n15807) );
  NAND2_X2 U17001 ( .A1(n13400), .A2(n17331), .ZN(n15806) );
  NAND3_X4 U17002 ( .A1(n15808), .A2(n15807), .A3(n15806), .ZN(n18901) );
  XNOR2_X2 U17003 ( .A(n18901), .B(n13493), .ZN(n15853) );
  XNOR2_X2 U17004 ( .A(n15853), .B(n18559), .ZN(n18561) );
  INV_X4 U17005 ( .A(n18561), .ZN(n16785) );
  NAND2_X2 U17006 ( .A1(n16780), .A2(n16785), .ZN(n15809) );
  INV_X4 U17007 ( .A(n15809), .ZN(n17720) );
  INV_X4 U17008 ( .A(n16787), .ZN(n15855) );
  NAND2_X2 U17009 ( .A1(n17720), .A2(n15855), .ZN(n15826) );
  NAND2_X2 U17010 ( .A1(ID_EXEC_OUT[81]), .A2(n13403), .ZN(n15814) );
  NAND2_X2 U17011 ( .A1(DMEM_BUS_OUT[17]), .A2(n13484), .ZN(n15813) );
  NAND2_X2 U17012 ( .A1(n13400), .A2(n17094), .ZN(n15812) );
  NAND3_X4 U17013 ( .A1(n15814), .A2(n15813), .A3(n15812), .ZN(n18890) );
  XNOR2_X2 U17014 ( .A(n18890), .B(n13493), .ZN(n15815) );
  XNOR2_X2 U17015 ( .A(n15815), .B(n18888), .ZN(n17130) );
  NAND2_X2 U17016 ( .A1(n15815), .A2(n18888), .ZN(n16786) );
  NAND2_X2 U17017 ( .A1(n17130), .A2(n16786), .ZN(n15856) );
  INV_X4 U17018 ( .A(n15856), .ZN(n15825) );
  NAND2_X2 U17019 ( .A1(ID_EXEC_OUT[79]), .A2(n18625), .ZN(n15818) );
  NAND2_X2 U17020 ( .A1(DMEM_BUS_OUT[15]), .A2(n18927), .ZN(n15817) );
  XNOR2_X2 U17021 ( .A(n10129), .B(n13493), .ZN(n15819) );
  INV_X4 U17022 ( .A(n17732), .ZN(n15824) );
  INV_X4 U17023 ( .A(n17733), .ZN(n17884) );
  NAND2_X2 U17024 ( .A1(ID_EXEC_OUT[78]), .A2(n13403), .ZN(n15822) );
  NAND2_X2 U17025 ( .A1(DMEM_BUS_OUT[14]), .A2(n13484), .ZN(n15821) );
  NAND2_X2 U17026 ( .A1(n13400), .A2(n17737), .ZN(n15820) );
  NAND3_X4 U17027 ( .A1(n15822), .A2(n15821), .A3(n15820), .ZN(n18896) );
  XNOR2_X2 U17028 ( .A(n18896), .B(n13493), .ZN(n15857) );
  XNOR2_X2 U17029 ( .A(n15857), .B(n18897), .ZN(n17734) );
  INV_X4 U17030 ( .A(n17734), .ZN(n15823) );
  OAI21_X4 U17031 ( .B1(n15824), .B2(n17884), .A(n15823), .ZN(n15864) );
  NOR3_X4 U17032 ( .A1(n15826), .A2(n15825), .A3(n15864), .ZN(n15850) );
  XNOR2_X2 U17033 ( .A(n13159), .B(n13494), .ZN(n15827) );
  XNOR2_X2 U17035 ( .A(n15828), .B(n19105), .ZN(n19108) );
  OAI21_X4 U17036 ( .B1(n19108), .B2(n13493), .A(n15829), .ZN(n18548) );
  OAI21_X4 U17039 ( .B1(n15832), .B2(n18547), .A(n15831), .ZN(n18466) );
  XNOR2_X2 U17040 ( .A(n13161), .B(n13218), .ZN(n15833) );
  XNOR2_X2 U17041 ( .A(n15833), .B(n18862), .ZN(n18467) );
  NAND2_X2 U17042 ( .A1(n15834), .A2(n13161), .ZN(n17492) );
  XNOR2_X2 U17043 ( .A(n18860), .B(n13494), .ZN(n15835) );
  NAND2_X2 U17044 ( .A1(n15835), .A2(n13163), .ZN(n17495) );
  NAND2_X2 U17045 ( .A1(n17492), .A2(n17495), .ZN(n15842) );
  XNOR2_X2 U17046 ( .A(n15835), .B(n13163), .ZN(n18279) );
  XNOR2_X2 U17047 ( .A(n18958), .B(n13494), .ZN(n15845) );
  XNOR2_X2 U17048 ( .A(n15845), .B(n18345), .ZN(n17498) );
  XNOR2_X2 U17049 ( .A(n15844), .B(n13041), .ZN(n18361) );
  AOI211_X4 U17050 ( .C1(n18279), .C2(n17495), .A(n17498), .B(n18361), .ZN(
        n15841) );
  OAI21_X4 U17051 ( .B1(n15843), .B2(n15842), .A(n15841), .ZN(n15849) );
  NAND2_X2 U17052 ( .A1(n15845), .A2(n18345), .ZN(n17894) );
  NAND2_X2 U17053 ( .A1(n17894), .A2(n17895), .ZN(n15846) );
  NOR2_X4 U17054 ( .A1(n15847), .A2(n15846), .ZN(n15848) );
  NAND2_X2 U17055 ( .A1(n15851), .A2(n18911), .ZN(n16781) );
  INV_X4 U17056 ( .A(n16781), .ZN(n15852) );
  NAND2_X2 U17057 ( .A1(n15852), .A2(n16785), .ZN(n17725) );
  INV_X4 U17058 ( .A(n17725), .ZN(n15854) );
  NAND2_X2 U17059 ( .A1(n15853), .A2(n18559), .ZN(n16783) );
  NAND2_X2 U17060 ( .A1(n16783), .A2(n16786), .ZN(n17723) );
  NOR2_X4 U17061 ( .A1(n15854), .A2(n17723), .ZN(n15862) );
  NAND2_X2 U17062 ( .A1(n15856), .A2(n15855), .ZN(n17729) );
  NAND2_X2 U17063 ( .A1(n15857), .A2(n18897), .ZN(n15863) );
  INV_X4 U17064 ( .A(n15863), .ZN(n15860) );
  INV_X4 U17065 ( .A(n17728), .ZN(n15859) );
  OAI211_X2 U17066 ( .C1(n15862), .C2(n17729), .A(n17732), .B(n15861), .ZN(
        n15866) );
  NAND2_X2 U17067 ( .A1(n15864), .A2(n15863), .ZN(n15865) );
  NAND2_X2 U17068 ( .A1(n15866), .A2(n15865), .ZN(n15867) );
  OAI21_X4 U17069 ( .B1(n15869), .B2(n15868), .A(n15867), .ZN(n17591) );
  NAND2_X2 U17070 ( .A1(ID_EXEC_OUT[77]), .A2(n13403), .ZN(n15872) );
  NAND2_X2 U17071 ( .A1(DMEM_BUS_OUT[13]), .A2(n13484), .ZN(n15871) );
  NAND2_X2 U17072 ( .A1(n13399), .A2(n16578), .ZN(n15870) );
  NAND3_X4 U17073 ( .A1(n15872), .A2(n15871), .A3(n15870), .ZN(n18907) );
  XNOR2_X2 U17074 ( .A(n18907), .B(n13494), .ZN(n15874) );
  XNOR2_X2 U17075 ( .A(n15874), .B(net222497), .ZN(n15873) );
  INV_X4 U17076 ( .A(n15873), .ZN(n17593) );
  NAND2_X2 U17077 ( .A1(ID_EXEC_OUT[76]), .A2(n13403), .ZN(n15877) );
  NAND2_X2 U17078 ( .A1(DMEM_BUS_OUT[12]), .A2(n13484), .ZN(n15876) );
  NAND2_X2 U17079 ( .A1(n13399), .A2(n16539), .ZN(n15875) );
  NAND3_X4 U17080 ( .A1(n15877), .A2(n15876), .A3(n15875), .ZN(n18999) );
  XNOR2_X2 U17081 ( .A(n18999), .B(n13494), .ZN(n15878) );
  NAND2_X2 U17082 ( .A1(n15878), .A2(n19000), .ZN(n16397) );
  XNOR2_X2 U17083 ( .A(n15878), .B(n19000), .ZN(n16537) );
  NAND2_X2 U17084 ( .A1(ID_EXEC_OUT[75]), .A2(n13403), .ZN(n15881) );
  NAND2_X2 U17085 ( .A1(DMEM_BUS_OUT[11]), .A2(n13484), .ZN(n15880) );
  NAND2_X2 U17086 ( .A1(n13399), .A2(n16350), .ZN(n15879) );
  NAND3_X4 U17087 ( .A1(n15881), .A2(n15880), .A3(n15879), .ZN(n19003) );
  XNOR2_X2 U17088 ( .A(n19003), .B(n13494), .ZN(n15883) );
  XNOR2_X2 U17089 ( .A(n15883), .B(n19004), .ZN(n16398) );
  AOI21_X4 U17090 ( .B1(n16537), .B2(n16397), .A(n16398), .ZN(n15882) );
  NAND2_X2 U17091 ( .A1(n15883), .A2(n19004), .ZN(n16324) );
  NAND2_X2 U17092 ( .A1(ID_EXEC_OUT[74]), .A2(n13403), .ZN(n15886) );
  NAND2_X2 U17093 ( .A1(DMEM_BUS_OUT[10]), .A2(n13484), .ZN(n15885) );
  NAND2_X2 U17094 ( .A1(n13399), .A2(n16295), .ZN(n15884) );
  NAND3_X4 U17095 ( .A1(n15886), .A2(n15885), .A3(n15884), .ZN(n19016) );
  XNOR2_X2 U17096 ( .A(n19016), .B(n13494), .ZN(n15887) );
  NAND2_X2 U17097 ( .A1(n15887), .A2(n19015), .ZN(n17037) );
  NAND2_X2 U17098 ( .A1(n16324), .A2(n17037), .ZN(n15892) );
  XNOR2_X2 U17099 ( .A(n15887), .B(n19015), .ZN(n17036) );
  NAND2_X2 U17100 ( .A1(ID_EXEC_OUT[73]), .A2(n13403), .ZN(n15890) );
  NAND2_X2 U17101 ( .A1(DMEM_BUS_OUT[9]), .A2(n13484), .ZN(n15889) );
  NAND2_X2 U17102 ( .A1(n13399), .A2(n17045), .ZN(n15888) );
  NAND3_X4 U17103 ( .A1(n15890), .A2(n15889), .A3(n15888), .ZN(n19012) );
  XNOR2_X2 U17104 ( .A(n19012), .B(n13494), .ZN(n15896) );
  XNOR2_X2 U17105 ( .A(n15896), .B(n19013), .ZN(n17041) );
  AOI21_X4 U17106 ( .B1(n17036), .B2(n17037), .A(n17041), .ZN(n15891) );
  OAI21_X4 U17107 ( .B1(n12994), .B2(n15892), .A(n15891), .ZN(n16077) );
  NAND2_X2 U17108 ( .A1(ID_EXEC_OUT[72]), .A2(n13403), .ZN(n15895) );
  NAND2_X2 U17109 ( .A1(DMEM_BUS_OUT[8]), .A2(n13484), .ZN(n15894) );
  NAND2_X2 U17110 ( .A1(n13399), .A2(n16222), .ZN(n15893) );
  NAND3_X4 U17111 ( .A1(n15895), .A2(n15894), .A3(n15893), .ZN(n19028) );
  XNOR2_X2 U17112 ( .A(n19028), .B(n13494), .ZN(n15898) );
  NAND2_X2 U17113 ( .A1(n15898), .A2(n19029), .ZN(n16080) );
  NAND2_X2 U17114 ( .A1(n15896), .A2(n19013), .ZN(n16078) );
  INV_X4 U17115 ( .A(n16080), .ZN(n15903) );
  XNOR2_X2 U17116 ( .A(n15898), .B(n19029), .ZN(n16081) );
  INV_X4 U17117 ( .A(n16081), .ZN(n16220) );
  NAND2_X2 U17118 ( .A1(DMEM_BUS_OUT[7]), .A2(n13485), .ZN(n15901) );
  NAND2_X2 U17119 ( .A1(ID_EXEC_OUT[71]), .A2(n13403), .ZN(n15900) );
  NAND2_X2 U17120 ( .A1(n13399), .A2(n16070), .ZN(n15899) );
  NAND3_X4 U17121 ( .A1(n15901), .A2(n15900), .A3(n15899), .ZN(n18878) );
  XNOR2_X2 U17122 ( .A(n18878), .B(n13494), .ZN(n15904) );
  XNOR2_X2 U17123 ( .A(n15904), .B(n16971), .ZN(n16083) );
  INV_X4 U17124 ( .A(n16083), .ZN(n15902) );
  OAI21_X4 U17125 ( .B1(n15903), .B2(n16220), .A(n15902), .ZN(n15906) );
  NAND2_X2 U17126 ( .A1(n15904), .A2(n16971), .ZN(n15905) );
  OAI21_X4 U17127 ( .B1(n15907), .B2(n15906), .A(n15905), .ZN(n16142) );
  NAND2_X2 U17128 ( .A1(ID_EXEC_OUT[70]), .A2(n13403), .ZN(n15910) );
  NAND2_X2 U17129 ( .A1(DMEM_BUS_OUT[6]), .A2(n13485), .ZN(n15909) );
  NAND2_X2 U17130 ( .A1(n13399), .A2(n16147), .ZN(n15908) );
  NAND3_X4 U17131 ( .A1(n15910), .A2(n15909), .A3(n15908), .ZN(n16154) );
  XNOR2_X2 U17132 ( .A(n16154), .B(n13494), .ZN(n15912) );
  XNOR2_X2 U17133 ( .A(n15912), .B(n19038), .ZN(n16141) );
  INV_X4 U17134 ( .A(n16141), .ZN(n15911) );
  NAND2_X2 U17135 ( .A1(n15912), .A2(n19038), .ZN(n18610) );
  NAND2_X2 U17136 ( .A1(ID_EXEC_OUT[67]), .A2(n13403), .ZN(n15917) );
  NAND2_X2 U17137 ( .A1(DMEM_BUS_OUT[3]), .A2(n13484), .ZN(n15916) );
  NAND2_X2 U17138 ( .A1(n13399), .A2(n16918), .ZN(n15915) );
  NAND3_X4 U17139 ( .A1(n15917), .A2(n15916), .A3(n15915), .ZN(n18877) );
  XNOR2_X2 U17140 ( .A(n18877), .B(n13494), .ZN(n15924) );
  NAND2_X2 U17141 ( .A1(n15924), .A2(n18872), .ZN(n18595) );
  NAND2_X2 U17142 ( .A1(ID_EXEC_OUT[66]), .A2(n13403), .ZN(n15920) );
  NAND2_X2 U17143 ( .A1(DMEM_BUS_OUT[2]), .A2(n13484), .ZN(n15919) );
  NAND2_X2 U17144 ( .A1(n13399), .A2(n16872), .ZN(n15918) );
  NAND3_X4 U17145 ( .A1(n15920), .A2(n15919), .A3(n15918), .ZN(n16892) );
  XNOR2_X2 U17146 ( .A(n16892), .B(n13494), .ZN(n15921) );
  NAND2_X2 U17147 ( .A1(n15921), .A2(n18873), .ZN(n18590) );
  NAND2_X2 U17148 ( .A1(n18595), .A2(n18590), .ZN(n15922) );
  XNOR2_X2 U17149 ( .A(n15921), .B(n18873), .ZN(n18597) );
  NAND2_X2 U17150 ( .A1(n18597), .A2(n18590), .ZN(n15925) );
  NAND2_X2 U17151 ( .A1(n15922), .A2(n15925), .ZN(n15926) );
  NAND2_X2 U17152 ( .A1(n15923), .A2(n18867), .ZN(n17557) );
  NAND2_X2 U17153 ( .A1(n15926), .A2(n17557), .ZN(n15929) );
  XNOR2_X2 U17154 ( .A(n15924), .B(n18872), .ZN(n18594) );
  INV_X4 U17155 ( .A(n18594), .ZN(n17560) );
  NAND2_X2 U17156 ( .A1(n15925), .A2(n17560), .ZN(n15927) );
  NAND2_X2 U17157 ( .A1(n15927), .A2(n15926), .ZN(n15928) );
  OAI21_X4 U17158 ( .B1(n16899), .B2(n15929), .A(n15928), .ZN(n15930) );
  XNOR2_X2 U17159 ( .A(n18869), .B(n11041), .ZN(n18589) );
  XNOR2_X2 U17160 ( .A(n18589), .B(n18870), .ZN(n18592) );
  XNOR2_X2 U17161 ( .A(n15930), .B(n18592), .ZN(n15934) );
  NAND2_X2 U17162 ( .A1(n13409), .A2(n18888), .ZN(n15936) );
  OAI211_X2 U17163 ( .C1(n12163), .C2(net231225), .A(n15936), .B(n6763), .ZN(
        n7340) );
  NAND2_X2 U17164 ( .A1(n13411), .A2(ID_EXEC_OUT[169]), .ZN(n15940) );
  NAND2_X2 U17165 ( .A1(DMEM_BUS_OUT[41]), .A2(net231321), .ZN(n15939) );
  NAND2_X2 U17166 ( .A1(n13413), .A2(DMEM_BUS_OUT[9]), .ZN(n15938) );
  NAND2_X2 U17167 ( .A1(n13415), .A2(MEM_WB_OUT[46]), .ZN(n15937) );
  NAND4_X2 U17168 ( .A1(n15940), .A2(n15939), .A3(n15938), .A4(n15937), .ZN(
        n7341) );
  NAND2_X2 U17169 ( .A1(n13410), .A2(n19013), .ZN(n15941) );
  OAI211_X2 U17170 ( .C1(n12155), .C2(net231227), .A(n15941), .B(n6773), .ZN(
        n7345) );
  NAND2_X2 U17171 ( .A1(n13412), .A2(ID_EXEC_OUT[162]), .ZN(n15945) );
  NAND2_X2 U17172 ( .A1(DMEM_BUS_OUT[34]), .A2(net231321), .ZN(n15944) );
  NAND2_X2 U17173 ( .A1(n13414), .A2(DMEM_BUS_OUT[2]), .ZN(n15943) );
  NAND2_X2 U17174 ( .A1(n13415), .A2(MEM_WB_OUT[39]), .ZN(n15942) );
  NAND4_X2 U17175 ( .A1(n15945), .A2(n15944), .A3(n15943), .A4(n15942), .ZN(
        n7346) );
  NAND2_X2 U17176 ( .A1(n13410), .A2(n19000), .ZN(n15946) );
  OAI211_X2 U17177 ( .C1(n12158), .C2(net231225), .A(n15946), .B(n6770), .ZN(
        n7350) );
  NAND2_X2 U17178 ( .A1(n13411), .A2(ID_EXEC_OUT[168]), .ZN(n15950) );
  NAND2_X2 U17179 ( .A1(DMEM_BUS_OUT[40]), .A2(net231321), .ZN(n15949) );
  NAND2_X2 U17180 ( .A1(n13413), .A2(DMEM_BUS_OUT[8]), .ZN(n15948) );
  NAND2_X2 U17181 ( .A1(n13415), .A2(MEM_WB_OUT[45]), .ZN(n15947) );
  NAND4_X2 U17182 ( .A1(n15950), .A2(n15949), .A3(n15948), .A4(n15947), .ZN(
        n7351) );
  NAND2_X2 U17183 ( .A1(n13412), .A2(ID_EXEC_OUT[166]), .ZN(n15954) );
  NAND2_X2 U17184 ( .A1(DMEM_BUS_OUT[38]), .A2(net231321), .ZN(n15953) );
  NAND2_X2 U17185 ( .A1(n13413), .A2(DMEM_BUS_OUT[6]), .ZN(n15952) );
  NAND2_X2 U17186 ( .A1(n13415), .A2(MEM_WB_OUT[43]), .ZN(n15951) );
  NAND4_X2 U17187 ( .A1(n15954), .A2(n15953), .A3(n15952), .A4(n15951), .ZN(
        n7352) );
  NAND2_X2 U17188 ( .A1(n13410), .A2(n19038), .ZN(n15955) );
  OAI211_X2 U17189 ( .C1(n12152), .C2(net231225), .A(n15955), .B(n6776), .ZN(
        n7356) );
  NAND2_X2 U17190 ( .A1(n13411), .A2(ID_EXEC_OUT[167]), .ZN(n15959) );
  NAND2_X2 U17191 ( .A1(DMEM_BUS_OUT[39]), .A2(net231321), .ZN(n15958) );
  NAND2_X2 U17192 ( .A1(n13414), .A2(DMEM_BUS_OUT[7]), .ZN(n15957) );
  NAND2_X2 U17193 ( .A1(n13415), .A2(MEM_WB_OUT[44]), .ZN(n15956) );
  NAND4_X2 U17194 ( .A1(n15959), .A2(n15958), .A3(n15957), .A4(n15956), .ZN(
        n7357) );
  NAND2_X2 U17195 ( .A1(n13412), .A2(ID_EXEC_OUT[165]), .ZN(n15963) );
  NAND2_X2 U17196 ( .A1(DMEM_BUS_OUT[37]), .A2(net231321), .ZN(n15962) );
  NAND2_X2 U17197 ( .A1(n13414), .A2(DMEM_BUS_OUT[5]), .ZN(n15961) );
  NAND2_X2 U17198 ( .A1(n13415), .A2(MEM_WB_OUT[42]), .ZN(n15960) );
  NAND4_X2 U17199 ( .A1(n15963), .A2(n15962), .A3(n15961), .A4(n15960), .ZN(
        n7358) );
  NAND2_X2 U17200 ( .A1(n13410), .A2(net225212), .ZN(n15964) );
  OAI211_X2 U17201 ( .C1(n12151), .C2(net231223), .A(n15964), .B(n6777), .ZN(
        n7362) );
  OAI22_X2 U17202 ( .A1(n13419), .A2(n12787), .B1(n13417), .B2(n11848), .ZN(
        n15968) );
  OAI22_X2 U17203 ( .A1(n13424), .A2(n12830), .B1(n13422), .B2(n12829), .ZN(
        n15967) );
  NAND2_X2 U17204 ( .A1(REG_FILE_reg_out_17__5_), .A2(n13436), .ZN(n15965) );
  OAI221_X2 U17205 ( .B1(n13432), .B2(n12831), .C1(n13427), .C2(n12722), .A(
        n15965), .ZN(n15966) );
  AOI22_X2 U17206 ( .A1(REG_FILE_reg_out_25__5_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__5_), .B2(n10350), .ZN(n15976) );
  OAI22_X2 U17207 ( .A1(n12393), .A2(n13444), .B1(n10510), .B2(n13442), .ZN(
        n15971) );
  OAI22_X2 U17208 ( .A1(n10306), .A2(n13190), .B1(n10691), .B2(n18699), .ZN(
        n15970) );
  OAI22_X2 U17209 ( .A1(n11841), .A2(n13192), .B1(n12392), .B2(n13193), .ZN(
        n15969) );
  NAND4_X2 U17210 ( .A1(n15977), .A2(n15976), .A3(n15975), .A4(n15974), .ZN(
        n16002) );
  NAND2_X2 U17211 ( .A1(n13456), .A2(REG_FILE_reg_out_12__5_), .ZN(n15986) );
  AOI22_X2 U17212 ( .A1(n13464), .A2(REG_FILE_reg_out_0__5_), .B1(
        REG_FILE_reg_out_15__5_), .B2(n13466), .ZN(n15984) );
  NAND4_X2 U17213 ( .A1(n15987), .A2(n15986), .A3(n15985), .A4(n15984), .ZN(
        n16001) );
  NAND4_X2 U17214 ( .A1(n15999), .A2(n15998), .A3(n15997), .A4(n15996), .ZN(
        n16000) );
  NOR3_X4 U17215 ( .A1(n16002), .A2(n16001), .A3(n16000), .ZN(n16003) );
  OAI22_X2 U17216 ( .A1(n11507), .A2(net231251), .B1(net230383), .B2(n16003), 
        .ZN(n7363) );
  OAI221_X2 U17217 ( .B1(n12502), .B2(net231221), .C1(n16003), .C2(n13477), 
        .A(n17267), .ZN(n7364) );
  MUX2_X2 U17218 ( .A(DMEM_BUS_OUT[5]), .B(MEM_WB_OUT[42]), .S(net231297), .Z(
        n7366) );
  XNOR2_X2 U17219 ( .A(n17294), .B(n18611), .ZN(n16005) );
  XNOR2_X2 U17220 ( .A(net222531), .B(net225212), .ZN(n19040) );
  INV_X4 U17221 ( .A(n18872), .ZN(n17526) );
  NAND2_X2 U17222 ( .A1(n17526), .A2(n16064), .ZN(n16008) );
  NAND2_X2 U17223 ( .A1(n16064), .A2(n16007), .ZN(n16062) );
  NAND2_X2 U17224 ( .A1(n16008), .A2(n16062), .ZN(n17307) );
  NAND2_X2 U17225 ( .A1(n16009), .A2(n16064), .ZN(n16389) );
  NAND2_X2 U17226 ( .A1(n13388), .A2(n16389), .ZN(n16012) );
  INV_X4 U17227 ( .A(n18637), .ZN(n19097) );
  NAND2_X2 U17228 ( .A1(n13392), .A2(n16879), .ZN(n16010) );
  INV_X4 U17229 ( .A(n16010), .ZN(n16026) );
  AOI21_X4 U17230 ( .B1(n13487), .B2(n17304), .A(n16026), .ZN(n16011) );
  OAI211_X2 U17231 ( .C1(n16060), .C2(n17307), .A(n16012), .B(n16011), .ZN(
        n16151) );
  INV_X4 U17232 ( .A(n16151), .ZN(n16018) );
  NAND2_X2 U17233 ( .A1(n13389), .A2(n16885), .ZN(n16016) );
  NAND2_X2 U17234 ( .A1(n13397), .A2(n16883), .ZN(n16015) );
  NAND2_X2 U17236 ( .A1(n13385), .A2(n19013), .ZN(n16301) );
  NAND2_X2 U17237 ( .A1(n13385), .A2(n19004), .ZN(n16390) );
  NAND2_X2 U17238 ( .A1(n13359), .A2(n18911), .ZN(n18269) );
  NAND3_X4 U17239 ( .A1(n16390), .A2(n18269), .A3(n16013), .ZN(n16290) );
  AOI22_X2 U17240 ( .A1(n13487), .A2(n16884), .B1(n13392), .B2(n16290), .ZN(
        n16014) );
  NAND3_X4 U17241 ( .A1(n16016), .A2(n16015), .A3(n16014), .ZN(n17322) );
  INV_X4 U17242 ( .A(n17322), .ZN(n16017) );
  OAI22_X2 U17243 ( .A1(n16018), .A2(n13211), .B1(n16017), .B2(n13214), .ZN(
        n16039) );
  NAND2_X2 U17244 ( .A1(n13386), .A2(n19015), .ZN(n16311) );
  NAND2_X2 U17245 ( .A1(n13359), .A2(n18559), .ZN(n18252) );
  NAND2_X2 U17246 ( .A1(net232816), .A2(n18345), .ZN(n16019) );
  NAND2_X2 U17247 ( .A1(n13386), .A2(n19000), .ZN(n16524) );
  NAND2_X2 U17248 ( .A1(n13359), .A2(n17505), .ZN(n18247) );
  NAND2_X2 U17249 ( .A1(net232816), .A2(n13163), .ZN(n16020) );
  NAND3_X4 U17250 ( .A1(n16524), .A2(n18247), .A3(n16020), .ZN(n16402) );
  AOI22_X2 U17251 ( .A1(n13487), .A2(n17300), .B1(n13392), .B2(n16402), .ZN(
        n16022) );
  AOI22_X2 U17252 ( .A1(n13388), .A2(n17298), .B1(n13397), .B2(n17299), .ZN(
        n16021) );
  NAND2_X2 U17253 ( .A1(n16022), .A2(n16021), .ZN(n16144) );
  INV_X4 U17254 ( .A(n16144), .ZN(n16023) );
  NAND2_X2 U17255 ( .A1(n16024), .A2(n16064), .ZN(n16310) );
  NAND2_X2 U17256 ( .A1(n13389), .A2(n16310), .ZN(n16029) );
  NAND2_X2 U17257 ( .A1(n13386), .A2(n18873), .ZN(n16025) );
  NAND2_X2 U17258 ( .A1(n16025), .A2(n16064), .ZN(n16878) );
  NAND2_X2 U17259 ( .A1(n13396), .A2(n16878), .ZN(n16028) );
  AOI21_X4 U17260 ( .B1(n13487), .B2(n16877), .A(n16026), .ZN(n16027) );
  INV_X4 U17261 ( .A(n16030), .ZN(n17316) );
  NAND2_X2 U17262 ( .A1(n17982), .A2(n16031), .ZN(n16034) );
  NAND2_X2 U17263 ( .A1(n17983), .A2(ID_EXEC_OUT[37]), .ZN(n16033) );
  NAND2_X2 U17264 ( .A1(n18566), .A2(DMEM_BUS_OUT[5]), .ZN(n16032) );
  NAND3_X2 U17265 ( .A1(n16034), .A2(n16033), .A3(n16032), .ZN(n16035) );
  NAND2_X2 U17266 ( .A1(n16035), .A2(net222531), .ZN(n16036) );
  MUX2_X2 U17267 ( .A(DMEM_BUS_OUT[7]), .B(MEM_WB_OUT[44]), .S(net231297), .Z(
        n7368) );
  AOI22_X2 U17268 ( .A1(DMEM_BUS_OUT[7]), .A2(net231307), .B1(ID_EXEC_OUT[211]), .B2(n13216), .ZN(n16088) );
  NAND2_X2 U17269 ( .A1(n13385), .A2(net222497), .ZN(n16774) );
  NAND2_X2 U17270 ( .A1(net232816), .A2(n13161), .ZN(n16043) );
  NAND3_X4 U17271 ( .A1(n16774), .A2(net223079), .A3(n16043), .ZN(n16544) );
  NAND2_X2 U17272 ( .A1(n13392), .A2(n16544), .ZN(n16046) );
  NAND2_X2 U17273 ( .A1(n13389), .A2(n16883), .ZN(n16045) );
  NAND2_X2 U17274 ( .A1(n13487), .A2(n16290), .ZN(n16044) );
  NAND4_X2 U17275 ( .A1(n16047), .A2(n16046), .A3(n16045), .A4(n16044), .ZN(
        n16152) );
  NAND2_X2 U17276 ( .A1(n16152), .A2(n18360), .ZN(n16058) );
  NAND2_X2 U17277 ( .A1(n13397), .A2(n17300), .ZN(n16052) );
  NAND2_X2 U17278 ( .A1(n13385), .A2(n18897), .ZN(n16796) );
  NAND2_X2 U17279 ( .A1(n13359), .A2(n18980), .ZN(n18535) );
  NAND3_X4 U17281 ( .A1(n16796), .A2(n18535), .A3(n16048), .ZN(n17597) );
  NAND2_X2 U17282 ( .A1(n13392), .A2(n17597), .ZN(n16051) );
  NAND2_X2 U17283 ( .A1(n13389), .A2(n17299), .ZN(n16050) );
  NAND2_X2 U17284 ( .A1(n13488), .A2(n16402), .ZN(n16049) );
  NAND4_X2 U17285 ( .A1(n16052), .A2(n16051), .A3(n16050), .A4(n16049), .ZN(
        n16214) );
  NAND2_X2 U17286 ( .A1(n16214), .A2(n17908), .ZN(n16057) );
  NAND2_X2 U17287 ( .A1(n18534), .A2(n16064), .ZN(n16053) );
  NAND2_X2 U17288 ( .A1(n16053), .A2(n16062), .ZN(n16209) );
  NAND2_X2 U17289 ( .A1(n13487), .A2(n16878), .ZN(n16055) );
  AOI22_X2 U17290 ( .A1(n13397), .A2(n16310), .B1(n13392), .B2(n16877), .ZN(
        n16054) );
  OAI211_X2 U17291 ( .C1(n19101), .C2(n16209), .A(n16055), .B(n16054), .ZN(
        n16157) );
  NAND2_X2 U17292 ( .A1(n16157), .A2(n18302), .ZN(n16056) );
  NAND2_X2 U17293 ( .A1(n17304), .A2(n16059), .ZN(n16068) );
  INV_X4 U17294 ( .A(n16060), .ZN(n16061) );
  NAND2_X2 U17295 ( .A1(n16389), .A2(n16061), .ZN(n16067) );
  INV_X4 U17296 ( .A(n16971), .ZN(n19089) );
  INV_X4 U17297 ( .A(n16062), .ZN(n16063) );
  AOI21_X4 U17298 ( .B1(n19089), .B2(n16064), .A(n16063), .ZN(n17584) );
  NAND2_X2 U17299 ( .A1(n17584), .A2(n15733), .ZN(n16066) );
  INV_X4 U17300 ( .A(n17307), .ZN(n16299) );
  NAND2_X2 U17301 ( .A1(n16299), .A2(n13488), .ZN(n16065) );
  NAND4_X2 U17302 ( .A1(n16068), .A2(n16067), .A3(n16066), .A4(n16065), .ZN(
        n16069) );
  INV_X4 U17303 ( .A(n16069), .ZN(n16226) );
  NOR2_X4 U17304 ( .A1(n16226), .A2(n13211), .ZN(n16075) );
  AOI22_X2 U17305 ( .A1(n17983), .A2(ID_EXEC_OUT[39]), .B1(n18566), .B2(
        DMEM_BUS_OUT[7]), .ZN(n16073) );
  NAND2_X2 U17306 ( .A1(n17982), .A2(n16070), .ZN(n16072) );
  INV_X4 U17307 ( .A(n18878), .ZN(n16071) );
  NOR3_X4 U17308 ( .A1(n16076), .A2(n16075), .A3(n16074), .ZN(n16087) );
  INV_X4 U17309 ( .A(n16079), .ZN(n16219) );
  OAI21_X4 U17310 ( .B1(n16081), .B2(n16219), .A(n16080), .ZN(n16082) );
  XNOR2_X2 U17311 ( .A(n16082), .B(n16083), .ZN(n16085) );
  XNOR2_X2 U17312 ( .A(n18878), .B(n16971), .ZN(n19031) );
  NAND3_X4 U17314 ( .A1(n16086), .A2(n16087), .A3(n16088), .ZN(n7369) );
  OAI22_X2 U17315 ( .A1(n13419), .A2(n12788), .B1(n13417), .B2(n11849), .ZN(
        n16092) );
  OAI22_X2 U17316 ( .A1(n13424), .A2(n12834), .B1(n13421), .B2(n12833), .ZN(
        n16091) );
  NAND2_X2 U17317 ( .A1(REG_FILE_reg_out_17__6_), .A2(n13436), .ZN(n16089) );
  OAI221_X2 U17318 ( .B1(n13432), .B2(n12835), .C1(n13427), .C2(n12723), .A(
        n16089), .ZN(n16090) );
  AOI22_X2 U17319 ( .A1(REG_FILE_reg_out_25__6_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__6_), .B2(n10350), .ZN(n16100) );
  OAI22_X2 U17320 ( .A1(n12417), .A2(n13444), .B1(n10511), .B2(n13442), .ZN(
        n16095) );
  OAI22_X2 U17321 ( .A1(n10307), .A2(n13190), .B1(n10692), .B2(n18699), .ZN(
        n16094) );
  OAI22_X2 U17322 ( .A1(n12737), .A2(n13192), .B1(n12416), .B2(n13193), .ZN(
        n16093) );
  NAND4_X2 U17323 ( .A1(n16101), .A2(n16100), .A3(n16099), .A4(n16098), .ZN(
        n16125) );
  INV_X4 U17324 ( .A(n16147), .ZN(n16130) );
  NAND2_X2 U17325 ( .A1(n13456), .A2(REG_FILE_reg_out_12__6_), .ZN(n16109) );
  AOI22_X2 U17326 ( .A1(n13464), .A2(REG_FILE_reg_out_0__6_), .B1(
        REG_FILE_reg_out_15__6_), .B2(n13466), .ZN(n16107) );
  NAND4_X2 U17327 ( .A1(n16110), .A2(n16109), .A3(n16108), .A4(n16107), .ZN(
        n16124) );
  NAND4_X2 U17328 ( .A1(n16122), .A2(n16121), .A3(n16120), .A4(n16119), .ZN(
        n16123) );
  NOR3_X4 U17329 ( .A1(n16125), .A2(n16124), .A3(n16123), .ZN(n16126) );
  OAI22_X2 U17330 ( .A1(n11508), .A2(net231253), .B1(net230383), .B2(n16126), 
        .ZN(n7370) );
  OAI221_X2 U17331 ( .B1(n12503), .B2(net231221), .C1(n16126), .C2(n13477), 
        .A(n17267), .ZN(n7371) );
  NOR2_X4 U17332 ( .A1(n2379), .A2(n2380), .ZN(n16139) );
  NOR4_X2 U17333 ( .A1(n2381), .A2(n16129), .A3(n16128), .A4(n16127), .ZN(
        n16137) );
  OAI22_X2 U17334 ( .A1(n12415), .A2(n13383), .B1(n13380), .B2(n12746), .ZN(
        n16134) );
  OAI222_X2 U17335 ( .A1(n11849), .A2(n13374), .B1(n10857), .B2(n13370), .C1(
        n13367), .C2(n12737), .ZN(n16133) );
  NAND4_X2 U17336 ( .A1(n16139), .A2(n16138), .A3(n16137), .A4(n16136), .ZN(
        n16140) );
  MUX2_X2 U17337 ( .A(n16140), .B(ID_EXEC_OUT[38]), .S(net231295), .Z(n7372)
         );
  NAND2_X2 U17338 ( .A1(n18360), .A2(n16144), .ZN(n16160) );
  NAND2_X2 U17339 ( .A1(n18566), .A2(DMEM_BUS_OUT[6]), .ZN(n16148) );
  INV_X4 U17340 ( .A(n16154), .ZN(n19039) );
  AOI221_X2 U17341 ( .B1(n18644), .B2(n16152), .C1(n19118), .C2(n16151), .A(
        n16150), .ZN(n16159) );
  NAND2_X2 U17342 ( .A1(DMEM_BUS_OUT[6]), .A2(net231321), .ZN(n16153) );
  XNOR2_X2 U17343 ( .A(n16154), .B(n19038), .ZN(n19035) );
  NAND2_X2 U17345 ( .A1(n13410), .A2(n19029), .ZN(n16162) );
  OAI211_X2 U17346 ( .C1(n12154), .C2(net231225), .A(n16162), .B(n6774), .ZN(
        n7378) );
  OAI22_X2 U17347 ( .A1(n13419), .A2(n12789), .B1(n13417), .B2(n12225), .ZN(
        n16166) );
  OAI22_X2 U17348 ( .A1(n13424), .A2(n12838), .B1(n13422), .B2(n12837), .ZN(
        n16165) );
  NAND2_X2 U17349 ( .A1(REG_FILE_reg_out_17__8_), .A2(n13436), .ZN(n16163) );
  OAI221_X2 U17350 ( .B1(n13432), .B2(n12839), .C1(n13427), .C2(n12724), .A(
        n16163), .ZN(n16164) );
  AOI22_X2 U17351 ( .A1(REG_FILE_reg_out_25__8_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__8_), .B2(n10350), .ZN(n16174) );
  OAI22_X2 U17352 ( .A1(n12397), .A2(n13444), .B1(n10513), .B2(n13442), .ZN(
        n16169) );
  OAI22_X2 U17353 ( .A1(n10309), .A2(n13190), .B1(n10693), .B2(n18699), .ZN(
        n16168) );
  OAI22_X2 U17354 ( .A1(n11843), .A2(n13192), .B1(n12396), .B2(n13193), .ZN(
        n16167) );
  NAND4_X2 U17355 ( .A1(n16175), .A2(n16174), .A3(n16173), .A4(n16172), .ZN(
        n16200) );
  NAND2_X2 U17356 ( .A1(n13456), .A2(REG_FILE_reg_out_12__8_), .ZN(n16184) );
  AOI22_X2 U17357 ( .A1(n13464), .A2(REG_FILE_reg_out_0__8_), .B1(
        REG_FILE_reg_out_15__8_), .B2(n13466), .ZN(n16182) );
  NAND4_X2 U17358 ( .A1(n16185), .A2(n16184), .A3(n16183), .A4(n16182), .ZN(
        n16199) );
  NAND4_X2 U17359 ( .A1(n16197), .A2(n16196), .A3(n16195), .A4(n16194), .ZN(
        n16198) );
  NOR3_X4 U17360 ( .A1(n16200), .A2(n16199), .A3(n16198), .ZN(n16201) );
  OAI22_X2 U17361 ( .A1(n11509), .A2(net231251), .B1(net230381), .B2(n16201), 
        .ZN(n7379) );
  OAI221_X2 U17362 ( .B1(n12504), .B2(net231221), .C1(n16201), .C2(n13476), 
        .A(n17267), .ZN(n7380) );
  MUX2_X2 U17363 ( .A(DMEM_BUS_OUT[8]), .B(MEM_WB_OUT[45]), .S(net231295), .Z(
        n7382) );
  NAND2_X2 U17364 ( .A1(n13487), .A2(n16544), .ZN(n16206) );
  NAND2_X2 U17365 ( .A1(n13359), .A2(n18922), .ZN(n19090) );
  NAND2_X2 U17366 ( .A1(net232816), .A2(n13151), .ZN(n16202) );
  NAND3_X4 U17367 ( .A1(n16772), .A2(n19090), .A3(n16202), .ZN(n17753) );
  NAND2_X2 U17368 ( .A1(n13392), .A2(n17753), .ZN(n16205) );
  NAND2_X2 U17369 ( .A1(n13396), .A2(n16290), .ZN(n16204) );
  NAND4_X2 U17370 ( .A1(n16206), .A2(n16205), .A3(n16204), .A4(n16203), .ZN(
        n17050) );
  NAND2_X2 U17371 ( .A1(n16310), .A2(n16300), .ZN(n16213) );
  NAND2_X2 U17372 ( .A1(n16878), .A2(n16207), .ZN(n16212) );
  OAI211_X2 U17373 ( .C1(n19354), .C2(n16797), .A(n16795), .B(n16208), .ZN(
        n17746) );
  NAND2_X2 U17374 ( .A1(n13389), .A2(n17746), .ZN(n16211) );
  INV_X4 U17375 ( .A(n16209), .ZN(n16523) );
  NAND2_X2 U17376 ( .A1(n16523), .A2(n16061), .ZN(n16210) );
  NAND4_X2 U17377 ( .A1(n16213), .A2(n16212), .A3(n16211), .A4(n16210), .ZN(
        n17051) );
  AOI22_X2 U17378 ( .A1(n17050), .A2(n10559), .B1(n17924), .B2(n17051), .ZN(
        n16232) );
  INV_X4 U17379 ( .A(n16214), .ZN(n16215) );
  NOR2_X4 U17380 ( .A1(n16215), .A2(n13215), .ZN(n16218) );
  OAI22_X2 U17381 ( .A1(net231249), .A2(n11986), .B1(n13217), .B2(n10820), 
        .ZN(n16217) );
  XNOR2_X2 U17382 ( .A(n19028), .B(n19029), .ZN(n19025) );
  XNOR2_X2 U17383 ( .A(n16220), .B(n16219), .ZN(n16221) );
  NAND2_X2 U17384 ( .A1(n13492), .A2(n16221), .ZN(n16230) );
  NAND2_X2 U17385 ( .A1(n18566), .A2(DMEM_BUS_OUT[8]), .ZN(n16225) );
  NAND2_X2 U17386 ( .A1(n17983), .A2(ID_EXEC_OUT[40]), .ZN(n16224) );
  NAND2_X2 U17387 ( .A1(n17982), .A2(n16222), .ZN(n16223) );
  AOI21_X4 U17388 ( .B1(n16228), .B2(n19028), .A(n16227), .ZN(n16229) );
  NAND4_X2 U17389 ( .A1(n16232), .A2(n16231), .A3(n16230), .A4(n16229), .ZN(
        n7383) );
  NAND2_X2 U17390 ( .A1(n13410), .A2(n19015), .ZN(n16233) );
  OAI211_X2 U17391 ( .C1(n12156), .C2(net231225), .A(n16233), .B(n6772), .ZN(
        n7387) );
  NAND2_X2 U17392 ( .A1(n13412), .A2(ID_EXEC_OUT[170]), .ZN(n16237) );
  NAND2_X2 U17393 ( .A1(DMEM_BUS_OUT[42]), .A2(net231321), .ZN(n16236) );
  NAND2_X2 U17394 ( .A1(n13414), .A2(DMEM_BUS_OUT[10]), .ZN(n16235) );
  NAND2_X2 U17395 ( .A1(n13415), .A2(MEM_WB_OUT[47]), .ZN(n16234) );
  NAND4_X2 U17396 ( .A1(n16237), .A2(n16236), .A3(n16235), .A4(n16234), .ZN(
        n7388) );
  OAI22_X2 U17397 ( .A1(n13419), .A2(n12790), .B1(n13417), .B2(n11850), .ZN(
        n16241) );
  OAI22_X2 U17398 ( .A1(n13424), .A2(n12842), .B1(n13421), .B2(n12841), .ZN(
        n16240) );
  NAND2_X2 U17399 ( .A1(REG_FILE_reg_out_17__10_), .A2(n13436), .ZN(n16238) );
  OAI221_X2 U17400 ( .B1(n13432), .B2(n12843), .C1(n13427), .C2(n12725), .A(
        n16238), .ZN(n16239) );
  AOI22_X2 U17401 ( .A1(REG_FILE_reg_out_25__10_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__10_), .B2(n10350), .ZN(n16249) );
  OAI22_X2 U17402 ( .A1(n12422), .A2(n13444), .B1(n10515), .B2(n13442), .ZN(
        n16244) );
  OAI22_X2 U17403 ( .A1(n10311), .A2(n13190), .B1(n10694), .B2(n18699), .ZN(
        n16243) );
  OAI22_X2 U17404 ( .A1(n12738), .A2(n13192), .B1(n12421), .B2(n13193), .ZN(
        n16242) );
  NAND4_X2 U17405 ( .A1(n16250), .A2(n16249), .A3(n16248), .A4(n16247), .ZN(
        n16274) );
  NAND2_X2 U17406 ( .A1(n13456), .A2(REG_FILE_reg_out_12__10_), .ZN(n16258) );
  AOI22_X2 U17407 ( .A1(n13464), .A2(REG_FILE_reg_out_0__10_), .B1(
        REG_FILE_reg_out_15__10_), .B2(n13466), .ZN(n16256) );
  NAND4_X2 U17408 ( .A1(n16259), .A2(n16258), .A3(n16257), .A4(n16256), .ZN(
        n16273) );
  NAND4_X2 U17409 ( .A1(n16271), .A2(n16270), .A3(n16269), .A4(n16268), .ZN(
        n16272) );
  NOR3_X4 U17410 ( .A1(n16274), .A2(n16273), .A3(n16272), .ZN(n16275) );
  OAI22_X2 U17411 ( .A1(n11510), .A2(net231253), .B1(net230381), .B2(n16275), 
        .ZN(n7389) );
  OAI221_X2 U17412 ( .B1(n12505), .B2(net231221), .C1(n16275), .C2(n13477), 
        .A(n17267), .ZN(n7390) );
  NOR2_X4 U17413 ( .A1(n2298), .A2(n2299), .ZN(n16288) );
  NOR4_X2 U17414 ( .A1(n2300), .A2(n16278), .A3(n16277), .A4(n16276), .ZN(
        n16286) );
  OAI22_X2 U17415 ( .A1(n12420), .A2(n13383), .B1(n13380), .B2(n12747), .ZN(
        n16283) );
  OAI222_X2 U17416 ( .A1(n11850), .A2(n13374), .B1(n10858), .B2(n13370), .C1(
        n13367), .C2(n12738), .ZN(n16282) );
  NAND4_X2 U17417 ( .A1(n16288), .A2(n16287), .A3(n16286), .A4(n16285), .ZN(
        n16289) );
  MUX2_X2 U17418 ( .A(n16289), .B(ID_EXEC_OUT[42]), .S(net231297), .Z(n7391)
         );
  NAND2_X2 U17419 ( .A1(n13487), .A2(n17753), .ZN(n16294) );
  NAND2_X2 U17420 ( .A1(n13386), .A2(n18888), .ZN(n17120) );
  NAND2_X2 U17421 ( .A1(n13389), .A2(n16290), .ZN(n16292) );
  NAND2_X2 U17422 ( .A1(n13396), .A2(n16544), .ZN(n16291) );
  NAND4_X2 U17423 ( .A1(n16294), .A2(n16293), .A3(n16292), .A4(n16291), .ZN(
        n16408) );
  NAND2_X2 U17424 ( .A1(n18644), .A2(n16408), .ZN(n16309) );
  OAI22_X2 U17425 ( .A1(n16279), .A2(n18569), .B1(n13209), .B2(n16296), .ZN(
        n16297) );
  NAND2_X2 U17426 ( .A1(n16299), .A2(n16059), .ZN(n16306) );
  NAND2_X2 U17427 ( .A1(n16300), .A2(n16389), .ZN(n16305) );
  NAND2_X2 U17428 ( .A1(n13359), .A2(n18870), .ZN(n16302) );
  NAND2_X2 U17429 ( .A1(n13389), .A2(n17585), .ZN(n16304) );
  NAND2_X2 U17430 ( .A1(n17584), .A2(n16061), .ZN(n16303) );
  NAND4_X2 U17431 ( .A1(n16306), .A2(n16305), .A3(n16304), .A4(n16303), .ZN(
        n17056) );
  NAND2_X2 U17432 ( .A1(n17056), .A2(n18302), .ZN(n16307) );
  NAND2_X2 U17433 ( .A1(n13392), .A2(n16310), .ZN(n16315) );
  NAND2_X2 U17434 ( .A1(n16523), .A2(n13488), .ZN(n16314) );
  NAND2_X2 U17435 ( .A1(n13359), .A2(n18873), .ZN(n16312) );
  AOI22_X2 U17436 ( .A1(n13388), .A2(n17747), .B1(n13397), .B2(n17746), .ZN(
        n16313) );
  INV_X4 U17437 ( .A(n16422), .ZN(n16316) );
  NOR2_X4 U17438 ( .A1(n16318), .A2(n16317), .ZN(n16331) );
  NAND2_X2 U17439 ( .A1(n13487), .A2(n17597), .ZN(n16323) );
  NAND2_X2 U17440 ( .A1(n13359), .A2(n13149), .ZN(n16319) );
  NAND2_X2 U17441 ( .A1(n16319), .A2(n16790), .ZN(n17598) );
  NAND2_X2 U17442 ( .A1(n13392), .A2(n17598), .ZN(n16322) );
  NAND2_X2 U17443 ( .A1(n13396), .A2(n16402), .ZN(n16321) );
  NAND2_X2 U17444 ( .A1(n13389), .A2(n17300), .ZN(n16320) );
  NAND4_X2 U17445 ( .A1(n16323), .A2(n16322), .A3(n16321), .A4(n16320), .ZN(
        n17057) );
  NAND2_X2 U17446 ( .A1(n18360), .A2(n17057), .ZN(n16330) );
  AOI22_X2 U17447 ( .A1(DMEM_BUS_OUT[10]), .A2(net231307), .B1(
        ID_EXEC_OUT[214]), .B2(n13216), .ZN(n16329) );
  XNOR2_X2 U17448 ( .A(n17040), .B(n17036), .ZN(n16327) );
  XNOR2_X2 U17449 ( .A(n19016), .B(n19015), .ZN(n19011) );
  NAND4_X2 U17450 ( .A1(n16328), .A2(n16330), .A3(n16329), .A4(n16331), .ZN(
        n7393) );
  NAND2_X2 U17451 ( .A1(n13410), .A2(n19004), .ZN(n16332) );
  OAI211_X2 U17452 ( .C1(n12157), .C2(net231225), .A(n16332), .B(n6771), .ZN(
        n7397) );
  NAND2_X2 U17453 ( .A1(n13412), .A2(ID_EXEC_OUT[171]), .ZN(n16336) );
  NAND2_X2 U17454 ( .A1(DMEM_BUS_OUT[43]), .A2(net231321), .ZN(n16335) );
  NAND2_X2 U17455 ( .A1(n13414), .A2(DMEM_BUS_OUT[11]), .ZN(n16334) );
  NAND2_X2 U17456 ( .A1(n13416), .A2(MEM_WB_OUT[48]), .ZN(n16333) );
  NAND4_X2 U17457 ( .A1(n16336), .A2(n16335), .A3(n16334), .A4(n16333), .ZN(
        n7398) );
  OAI22_X2 U17458 ( .A1(n13419), .A2(n12791), .B1(n13417), .B2(n11851), .ZN(
        n16340) );
  OAI22_X2 U17459 ( .A1(n13423), .A2(n12846), .B1(n13422), .B2(n12845), .ZN(
        n16339) );
  NAND2_X2 U17460 ( .A1(REG_FILE_reg_out_17__11_), .A2(n13436), .ZN(n16337) );
  OAI221_X2 U17461 ( .B1(n13432), .B2(n12847), .C1(n13427), .C2(n12726), .A(
        n16337), .ZN(n16338) );
  AOI22_X2 U17462 ( .A1(REG_FILE_reg_out_25__11_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__11_), .B2(n10350), .ZN(n16348) );
  OAI22_X2 U17463 ( .A1(n12426), .A2(n13444), .B1(n10516), .B2(n13442), .ZN(
        n16343) );
  OAI22_X2 U17464 ( .A1(n10312), .A2(n13190), .B1(n10695), .B2(n18699), .ZN(
        n16342) );
  OAI22_X2 U17465 ( .A1(n12739), .A2(n13192), .B1(n12425), .B2(n13193), .ZN(
        n16341) );
  NAND4_X2 U17466 ( .A1(n16349), .A2(n16348), .A3(n16347), .A4(n16346), .ZN(
        n16374) );
  INV_X4 U17467 ( .A(n16350), .ZN(n16413) );
  NAND2_X2 U17468 ( .A1(n13456), .A2(REG_FILE_reg_out_12__11_), .ZN(n16358) );
  AOI22_X2 U17469 ( .A1(n13464), .A2(REG_FILE_reg_out_0__11_), .B1(
        REG_FILE_reg_out_15__11_), .B2(n13466), .ZN(n16356) );
  NAND4_X2 U17470 ( .A1(n16359), .A2(n16358), .A3(n16357), .A4(n16356), .ZN(
        n16373) );
  NAND4_X2 U17471 ( .A1(n16371), .A2(n16370), .A3(n16369), .A4(n16368), .ZN(
        n16372) );
  NOR3_X4 U17472 ( .A1(n16374), .A2(n16373), .A3(n16372), .ZN(n16375) );
  OAI22_X2 U17473 ( .A1(n11511), .A2(net231255), .B1(net230381), .B2(n16375), 
        .ZN(n7399) );
  OAI221_X2 U17474 ( .B1(n12506), .B2(net231221), .C1(n16375), .C2(n13477), 
        .A(n17267), .ZN(n7400) );
  NOR2_X4 U17475 ( .A1(n2278), .A2(n2279), .ZN(n16387) );
  NOR4_X2 U17476 ( .A1(n2280), .A2(n16378), .A3(n16377), .A4(n16376), .ZN(
        n16385) );
  OAI22_X2 U17477 ( .A1(n12424), .A2(n13383), .B1(n13380), .B2(n12748), .ZN(
        n16382) );
  OAI222_X2 U17478 ( .A1(n11851), .A2(n13374), .B1(n10859), .B2(n13370), .C1(
        n13367), .C2(n12739), .ZN(n16381) );
  NAND4_X2 U17479 ( .A1(n16387), .A2(n16386), .A3(n16385), .A4(n16384), .ZN(
        n16388) );
  MUX2_X2 U17480 ( .A(n16388), .B(ID_EXEC_OUT[43]), .S(net231295), .Z(n7401)
         );
  NAND2_X2 U17481 ( .A1(n13393), .A2(n16389), .ZN(n16394) );
  NAND2_X2 U17482 ( .A1(n17584), .A2(n13488), .ZN(n16393) );
  NAND2_X2 U17483 ( .A1(n13358), .A2(n18872), .ZN(n16391) );
  AOI22_X2 U17484 ( .A1(n13388), .A2(n17586), .B1(n13397), .B2(n17585), .ZN(
        n16392) );
  NAND2_X2 U17485 ( .A1(n17924), .A2(n16530), .ZN(n16426) );
  OAI21_X4 U17486 ( .B1(n16537), .B2(n12990), .A(n16397), .ZN(n16399) );
  XNOR2_X2 U17487 ( .A(n16399), .B(n16398), .ZN(n16400) );
  NAND2_X2 U17488 ( .A1(n16400), .A2(n13492), .ZN(n16425) );
  NAND2_X2 U17489 ( .A1(n13487), .A2(n17598), .ZN(n16406) );
  NAND2_X2 U17490 ( .A1(n13358), .A2(n18345), .ZN(n16401) );
  NAND2_X2 U17491 ( .A1(n13386), .A2(n18559), .ZN(n17515) );
  NAND2_X2 U17492 ( .A1(n16401), .A2(n17515), .ZN(n17595) );
  NAND2_X2 U17493 ( .A1(n13392), .A2(n17595), .ZN(n16405) );
  NAND2_X2 U17494 ( .A1(n13389), .A2(n16402), .ZN(n16404) );
  NAND2_X2 U17495 ( .A1(n13396), .A2(n17597), .ZN(n16403) );
  NAND4_X2 U17496 ( .A1(n16406), .A2(n16405), .A3(n16404), .A4(n16403), .ZN(
        n16407) );
  INV_X4 U17497 ( .A(n16407), .ZN(n16532) );
  NOR2_X4 U17498 ( .A1(n16532), .A2(n13207), .ZN(n16418) );
  INV_X4 U17499 ( .A(n16408), .ZN(n16416) );
  INV_X4 U17500 ( .A(n16409), .ZN(n16410) );
  NAND2_X2 U17501 ( .A1(n16410), .A2(n13208), .ZN(n16412) );
  NAND2_X2 U17502 ( .A1(n18566), .A2(DMEM_BUS_OUT[11]), .ZN(n16411) );
  OAI211_X2 U17503 ( .C1(n16413), .C2(n18569), .A(n16412), .B(n16411), .ZN(
        n16414) );
  NAND2_X2 U17504 ( .A1(n16414), .A2(n19003), .ZN(n16415) );
  OAI21_X4 U17505 ( .B1(n16416), .B2(n13214), .A(n16415), .ZN(n16417) );
  NAND2_X2 U17506 ( .A1(DMEM_BUS_OUT[11]), .A2(net231321), .ZN(n16419) );
  XNOR2_X2 U17507 ( .A(n19003), .B(n19004), .ZN(n19001) );
  NAND4_X2 U17508 ( .A1(n16425), .A2(n16426), .A3(n16424), .A4(n16423), .ZN(
        n7403) );
  NAND2_X2 U17509 ( .A1(n13410), .A2(n16971), .ZN(n16427) );
  OAI211_X2 U17510 ( .C1(n12153), .C2(net231227), .A(n16427), .B(n6775), .ZN(
        n7407) );
  OAI22_X2 U17511 ( .A1(n13419), .A2(n12792), .B1(n13417), .B2(n12226), .ZN(
        n16431) );
  OAI22_X2 U17512 ( .A1(n13423), .A2(n12850), .B1(n13422), .B2(n12849), .ZN(
        n16430) );
  NAND2_X2 U17513 ( .A1(REG_FILE_reg_out_17__7_), .A2(n13436), .ZN(n16428) );
  OAI221_X2 U17514 ( .B1(n13432), .B2(n12851), .C1(n13427), .C2(n12727), .A(
        n16428), .ZN(n16429) );
  AOI22_X2 U17515 ( .A1(REG_FILE_reg_out_25__7_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__7_), .B2(n10350), .ZN(n16439) );
  OAI22_X2 U17516 ( .A1(n12395), .A2(n13444), .B1(n10512), .B2(n13442), .ZN(
        n16434) );
  OAI22_X2 U17517 ( .A1(n10308), .A2(n13190), .B1(n10696), .B2(n18699), .ZN(
        n16433) );
  OAI22_X2 U17518 ( .A1(n11842), .A2(n13192), .B1(n12394), .B2(n13193), .ZN(
        n16432) );
  NAND4_X2 U17519 ( .A1(n16440), .A2(n16439), .A3(n16438), .A4(n16437), .ZN(
        n16465) );
  NAND2_X2 U17520 ( .A1(n13456), .A2(REG_FILE_reg_out_12__7_), .ZN(n16449) );
  AOI22_X2 U17521 ( .A1(n13464), .A2(REG_FILE_reg_out_0__7_), .B1(
        REG_FILE_reg_out_15__7_), .B2(n13466), .ZN(n16447) );
  NAND4_X2 U17522 ( .A1(n16450), .A2(n16449), .A3(n16448), .A4(n16447), .ZN(
        n16464) );
  NAND4_X2 U17523 ( .A1(n16462), .A2(n16461), .A3(n16460), .A4(n16459), .ZN(
        n16463) );
  NOR3_X4 U17524 ( .A1(n16465), .A2(n16464), .A3(n16463), .ZN(n16466) );
  OAI22_X2 U17525 ( .A1(n11512), .A2(net231251), .B1(net230381), .B2(n16466), 
        .ZN(n7408) );
  OAI221_X2 U17526 ( .B1(n12507), .B2(net231221), .C1(n16466), .C2(n13476), 
        .A(n17267), .ZN(n7409) );
  MUX2_X2 U17527 ( .A(MEM_WB_REG_MEM_WB_REG_N173), .B(MEM_WB_OUT[7]), .S(
        net231295), .Z(n7411) );
  OAI22_X2 U17528 ( .A1(n12195), .A2(net231253), .B1(n13481), .B2(n16467), 
        .ZN(n7414) );
  XNOR2_X2 U17529 ( .A(net225906), .B(n11919), .ZN(n16468) );
  XNOR2_X2 U17530 ( .A(n16469), .B(n16468), .ZN(n16472) );
  NAND2_X2 U17531 ( .A1(net231615), .A2(n19015), .ZN(n16471) );
  NAND2_X2 U17532 ( .A1(EXEC_MEM_OUT_119), .A2(net231321), .ZN(n16470) );
  OAI211_X2 U17533 ( .C1(n16472), .C2(net231915), .A(n16471), .B(n16470), .ZN(
        n7415) );
  MUX2_X2 U17534 ( .A(MEM_WB_REG_MEM_WB_REG_N170), .B(MEM_WB_OUT[10]), .S(
        net231295), .Z(n7416) );
  OAI22_X2 U17535 ( .A1(n19331), .A2(net231251), .B1(n13481), .B2(n16473), 
        .ZN(n7419) );
  MUX2_X2 U17536 ( .A(MEM_WB_REG_MEM_WB_REG_N169), .B(MEM_WB_OUT[11]), .S(
        net231295), .Z(n7420) );
  OAI22_X2 U17537 ( .A1(net231247), .A2(n12018), .B1(n19330), .B2(net230381), 
        .ZN(n7422) );
  OAI22_X2 U17538 ( .A1(n19330), .A2(net231251), .B1(n13481), .B2(n16474), 
        .ZN(n7423) );
  XNOR2_X2 U17539 ( .A(net225890), .B(net225889), .ZN(n16476) );
  NAND2_X2 U17540 ( .A1(net231615), .A2(n19004), .ZN(n16475) );
  OAI221_X2 U17541 ( .B1(net231227), .B2(n11473), .C1(n16476), .C2(net231915), 
        .A(n16475), .ZN(n7424) );
  NAND2_X2 U17542 ( .A1(n13412), .A2(ID_EXEC_OUT[172]), .ZN(n16480) );
  NAND2_X2 U17543 ( .A1(DMEM_BUS_OUT[44]), .A2(net231321), .ZN(n16479) );
  NAND2_X2 U17544 ( .A1(n13414), .A2(DMEM_BUS_OUT[12]), .ZN(n16478) );
  NAND2_X2 U17545 ( .A1(n13416), .A2(MEM_WB_OUT[49]), .ZN(n16477) );
  NAND4_X2 U17546 ( .A1(n16480), .A2(n16479), .A3(n16478), .A4(n16477), .ZN(
        n7425) );
  OAI22_X2 U17547 ( .A1(n13419), .A2(n12793), .B1(n13417), .B2(n12227), .ZN(
        n16484) );
  OAI22_X2 U17548 ( .A1(n13423), .A2(n12854), .B1(n13422), .B2(n12853), .ZN(
        n16483) );
  NAND2_X2 U17549 ( .A1(REG_FILE_reg_out_17__12_), .A2(n13436), .ZN(n16481) );
  OAI221_X2 U17550 ( .B1(n13432), .B2(n12855), .C1(n13427), .C2(n12728), .A(
        n16481), .ZN(n16482) );
  AOI22_X2 U17551 ( .A1(REG_FILE_reg_out_25__12_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__12_), .B2(n10350), .ZN(n16492) );
  OAI22_X2 U17552 ( .A1(n12400), .A2(n13444), .B1(n10517), .B2(n13442), .ZN(
        n16487) );
  OAI22_X2 U17553 ( .A1(n10313), .A2(n13190), .B1(n10697), .B2(n18699), .ZN(
        n16486) );
  OAI22_X2 U17554 ( .A1(n11844), .A2(n13192), .B1(n12399), .B2(n13193), .ZN(
        n16485) );
  NAND4_X2 U17555 ( .A1(n16493), .A2(n16492), .A3(n16491), .A4(n16490), .ZN(
        n16518) );
  NAND2_X2 U17556 ( .A1(n13456), .A2(REG_FILE_reg_out_12__12_), .ZN(n16502) );
  AOI22_X2 U17557 ( .A1(n13464), .A2(REG_FILE_reg_out_0__12_), .B1(
        REG_FILE_reg_out_15__12_), .B2(n13466), .ZN(n16500) );
  NAND4_X2 U17558 ( .A1(n16503), .A2(n16502), .A3(n16501), .A4(n16500), .ZN(
        n16517) );
  NAND4_X2 U17559 ( .A1(n16515), .A2(n16514), .A3(n16513), .A4(n16512), .ZN(
        n16516) );
  NOR3_X4 U17560 ( .A1(n16518), .A2(n16517), .A3(n16516), .ZN(n16519) );
  OAI22_X2 U17561 ( .A1(n11513), .A2(net231251), .B1(net230381), .B2(n16519), 
        .ZN(n7426) );
  OAI221_X2 U17562 ( .B1(n12508), .B2(net231221), .C1(n16519), .C2(n13476), 
        .A(n17267), .ZN(n7427) );
  MUX2_X2 U17563 ( .A(MEM_WB_REG_MEM_WB_REG_N168), .B(MEM_WB_OUT[12]), .S(
        net231295), .Z(n7429) );
  OAI22_X2 U17564 ( .A1(n12188), .A2(net231255), .B1(n13481), .B2(n16520), 
        .ZN(n7432) );
  MUX2_X2 U17567 ( .A(DMEM_BUS_OUT[12]), .B(MEM_WB_OUT[49]), .S(net231295), 
        .Z(n7434) );
  XNOR2_X2 U17568 ( .A(n18999), .B(n19000), .ZN(n18851) );
  INV_X4 U17569 ( .A(n18851), .ZN(n16529) );
  NAND2_X2 U17570 ( .A1(n16523), .A2(n16059), .ZN(n16528) );
  NAND2_X2 U17571 ( .A1(n13487), .A2(n17746), .ZN(n16527) );
  NAND2_X2 U17572 ( .A1(n13358), .A2(n18867), .ZN(n16525) );
  AOI22_X2 U17573 ( .A1(n13388), .A2(n17910), .B1(n13397), .B2(n17747), .ZN(
        n16526) );
  AOI22_X2 U17574 ( .A1(n13490), .A2(n16529), .B1(n17924), .B2(n17617), .ZN(
        n16555) );
  INV_X4 U17575 ( .A(n16530), .ZN(n16531) );
  NOR2_X4 U17576 ( .A1(n16531), .A2(n13213), .ZN(n16535) );
  OAI22_X2 U17577 ( .A1(net231249), .A2(n11987), .B1(n13217), .B2(n10821), 
        .ZN(n16534) );
  NOR2_X4 U17578 ( .A1(n16532), .A2(n13215), .ZN(n16533) );
  NOR3_X4 U17579 ( .A1(n16535), .A2(n16534), .A3(n16533), .ZN(n16554) );
  NAND2_X2 U17580 ( .A1(n13492), .A2(n16538), .ZN(n16553) );
  NAND2_X2 U17581 ( .A1(n18566), .A2(DMEM_BUS_OUT[12]), .ZN(n16542) );
  NAND2_X2 U17582 ( .A1(n17983), .A2(ID_EXEC_OUT[44]), .ZN(n16541) );
  NAND2_X2 U17583 ( .A1(n17982), .A2(n16539), .ZN(n16540) );
  NAND2_X2 U17584 ( .A1(n13386), .A2(n18911), .ZN(n17530) );
  NAND2_X2 U17585 ( .A1(n16543), .A2(n17530), .ZN(n17917) );
  NAND2_X2 U17586 ( .A1(n13393), .A2(n17917), .ZN(n16547) );
  NAND2_X2 U17587 ( .A1(n13389), .A2(n16544), .ZN(n16546) );
  NAND2_X2 U17588 ( .A1(n13396), .A2(n17753), .ZN(n16545) );
  NAND4_X2 U17589 ( .A1(n16548), .A2(n16547), .A3(n16546), .A4(n16545), .ZN(
        n16549) );
  INV_X4 U17590 ( .A(n16549), .ZN(n17611) );
  NOR2_X4 U17591 ( .A1(n17611), .A2(n13207), .ZN(n16550) );
  AOI21_X4 U17592 ( .B1(n16551), .B2(n18999), .A(n16550), .ZN(n16552) );
  NAND4_X2 U17593 ( .A1(n16555), .A2(n16554), .A3(n16553), .A4(n16552), .ZN(
        n7435) );
  OAI211_X2 U17594 ( .C1(n12162), .C2(net231225), .A(n16556), .B(n6764), .ZN(
        n7439) );
  XNOR2_X2 U17595 ( .A(n16557), .B(net225777), .ZN(n16560) );
  NAND2_X2 U17596 ( .A1(net231615), .A2(net222497), .ZN(n16559) );
  NAND2_X2 U17597 ( .A1(EXEC_MEM_OUT_122), .A2(net231321), .ZN(n16558) );
  OAI211_X2 U17598 ( .C1(n16560), .C2(net231915), .A(n16559), .B(n16558), .ZN(
        n7440) );
  NAND2_X2 U17599 ( .A1(n13412), .A2(ID_EXEC_OUT[173]), .ZN(n16564) );
  NAND2_X2 U17600 ( .A1(DMEM_BUS_OUT[45]), .A2(net231321), .ZN(n16563) );
  NAND2_X2 U17601 ( .A1(n13414), .A2(DMEM_BUS_OUT[13]), .ZN(n16562) );
  NAND2_X2 U17602 ( .A1(n13416), .A2(MEM_WB_OUT[50]), .ZN(n16561) );
  NAND4_X2 U17603 ( .A1(n16564), .A2(n16563), .A3(n16562), .A4(n16561), .ZN(
        n7441) );
  OAI22_X2 U17604 ( .A1(n13419), .A2(n12794), .B1(n13417), .B2(n11852), .ZN(
        n16568) );
  OAI22_X2 U17605 ( .A1(n13423), .A2(n12858), .B1(n13422), .B2(n12857), .ZN(
        n16567) );
  NAND2_X2 U17606 ( .A1(REG_FILE_reg_out_17__13_), .A2(n13436), .ZN(n16565) );
  OAI221_X2 U17607 ( .B1(n13432), .B2(n12859), .C1(n13427), .C2(n12729), .A(
        n16565), .ZN(n16566) );
  AOI22_X2 U17608 ( .A1(REG_FILE_reg_out_25__13_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__13_), .B2(n10350), .ZN(n16576) );
  OAI22_X2 U17609 ( .A1(n12432), .A2(n13444), .B1(n10518), .B2(n13442), .ZN(
        n16571) );
  OAI22_X2 U17610 ( .A1(n10314), .A2(n13190), .B1(n10698), .B2(n18699), .ZN(
        n16570) );
  OAI22_X2 U17611 ( .A1(n12740), .A2(n13192), .B1(n12431), .B2(n13193), .ZN(
        n16569) );
  NAND4_X2 U17612 ( .A1(n16577), .A2(n16576), .A3(n16575), .A4(n16574), .ZN(
        n16602) );
  INV_X4 U17613 ( .A(n16578), .ZN(n17608) );
  NAND2_X2 U17614 ( .A1(n13456), .A2(REG_FILE_reg_out_12__13_), .ZN(n16586) );
  AOI22_X2 U17615 ( .A1(n13464), .A2(REG_FILE_reg_out_0__13_), .B1(
        REG_FILE_reg_out_15__13_), .B2(n13466), .ZN(n16584) );
  NAND4_X2 U17616 ( .A1(n16587), .A2(n16586), .A3(n16585), .A4(n16584), .ZN(
        n16601) );
  NAND4_X2 U17617 ( .A1(n16599), .A2(n16598), .A3(n16597), .A4(n16596), .ZN(
        n16600) );
  NOR3_X4 U17618 ( .A1(n16602), .A2(n16601), .A3(n16600), .ZN(n16603) );
  OAI22_X2 U17619 ( .A1(n11514), .A2(net231253), .B1(net230381), .B2(n16603), 
        .ZN(n7442) );
  OAI221_X2 U17620 ( .B1(n12509), .B2(net231221), .C1(n16603), .C2(n13476), 
        .A(n17267), .ZN(n7443) );
  NOR2_X4 U17621 ( .A1(n2238), .A2(n2239), .ZN(n16615) );
  NOR4_X2 U17622 ( .A1(n2240), .A2(n16606), .A3(n16605), .A4(n16604), .ZN(
        n16613) );
  OAI22_X2 U17623 ( .A1(n12430), .A2(n13383), .B1(n13380), .B2(n12749), .ZN(
        n16610) );
  OAI222_X2 U17624 ( .A1(n11852), .A2(n13374), .B1(n10252), .B2(n13370), .C1(
        n13368), .C2(n12740), .ZN(n16609) );
  NAND4_X2 U17625 ( .A1(n16615), .A2(n16614), .A3(n16613), .A4(n16612), .ZN(
        n16616) );
  MUX2_X2 U17626 ( .A(n16616), .B(ID_EXEC_OUT[45]), .S(net231295), .Z(n7444)
         );
  MUX2_X2 U17627 ( .A(MEM_WB_REG_MEM_WB_REG_N167), .B(MEM_WB_OUT[13]), .S(
        net231295), .Z(n7445) );
  OAI22_X2 U17628 ( .A1(net231249), .A2(n11934), .B1(n19329), .B2(net230383), 
        .ZN(n7447) );
  OAI22_X2 U17629 ( .A1(n19329), .A2(net231253), .B1(n13481), .B2(n16617), 
        .ZN(n7448) );
  XNOR2_X2 U17630 ( .A(n16618), .B(net225681), .ZN(n16621) );
  NAND2_X2 U17631 ( .A1(net231615), .A2(n18897), .ZN(n16620) );
  NAND2_X2 U17632 ( .A1(EXEC_MEM_OUT_123), .A2(net231321), .ZN(n16619) );
  OAI211_X2 U17633 ( .C1(n16621), .C2(net231915), .A(n16620), .B(n16619), .ZN(
        n7449) );
  NAND2_X2 U17634 ( .A1(n13412), .A2(ID_EXEC_OUT[174]), .ZN(n16625) );
  NAND2_X2 U17635 ( .A1(DMEM_BUS_OUT[46]), .A2(net231319), .ZN(n16624) );
  NAND2_X2 U17636 ( .A1(n13414), .A2(DMEM_BUS_OUT[14]), .ZN(n16623) );
  NAND2_X2 U17637 ( .A1(n13416), .A2(MEM_WB_OUT[51]), .ZN(n16622) );
  NAND4_X2 U17638 ( .A1(n16625), .A2(n16624), .A3(n16623), .A4(n16622), .ZN(
        n7450) );
  OAI22_X2 U17639 ( .A1(n13419), .A2(n12795), .B1(n13417), .B2(n12228), .ZN(
        n16629) );
  OAI22_X2 U17640 ( .A1(n13423), .A2(n12862), .B1(n13422), .B2(n12861), .ZN(
        n16628) );
  NAND2_X2 U17641 ( .A1(REG_FILE_reg_out_17__14_), .A2(n13436), .ZN(n16626) );
  OAI221_X2 U17642 ( .B1(n13432), .B2(n12863), .C1(n13427), .C2(n12730), .A(
        n16626), .ZN(n16627) );
  AOI22_X2 U17643 ( .A1(REG_FILE_reg_out_25__14_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__14_), .B2(n10350), .ZN(n16637) );
  OAI22_X2 U17644 ( .A1(n12402), .A2(n13444), .B1(n10519), .B2(n13442), .ZN(
        n16632) );
  OAI22_X2 U17645 ( .A1(n10315), .A2(n13190), .B1(n10699), .B2(n18699), .ZN(
        n16631) );
  OAI22_X2 U17646 ( .A1(n11845), .A2(n13192), .B1(n12401), .B2(n13193), .ZN(
        n16630) );
  NAND4_X2 U17647 ( .A1(n16638), .A2(n16637), .A3(n16636), .A4(n16635), .ZN(
        n16663) );
  NAND2_X2 U17648 ( .A1(n13456), .A2(REG_FILE_reg_out_12__14_), .ZN(n16647) );
  AOI22_X2 U17649 ( .A1(n13464), .A2(REG_FILE_reg_out_0__14_), .B1(
        REG_FILE_reg_out_15__14_), .B2(n13466), .ZN(n16645) );
  NAND4_X2 U17650 ( .A1(n16648), .A2(n16647), .A3(n16646), .A4(n16645), .ZN(
        n16662) );
  NAND4_X2 U17651 ( .A1(n16660), .A2(n16659), .A3(n16658), .A4(n16657), .ZN(
        n16661) );
  NOR3_X4 U17652 ( .A1(n16663), .A2(n16662), .A3(n16661), .ZN(n16664) );
  OAI22_X2 U17653 ( .A1(n11515), .A2(net231253), .B1(net230379), .B2(n16664), 
        .ZN(n7451) );
  OAI221_X2 U17654 ( .B1(n12510), .B2(net231221), .C1(n16664), .C2(n13476), 
        .A(n17267), .ZN(n7452) );
  MUX2_X2 U17655 ( .A(MEM_WB_REG_MEM_WB_REG_N166), .B(MEM_WB_OUT[14]), .S(
        net231295), .Z(n7454) );
  OAI22_X2 U17656 ( .A1(n11541), .A2(net231253), .B1(net230379), .B2(n11993), 
        .ZN(n7455) );
  OAI22_X2 U17657 ( .A1(net231249), .A2(n11993), .B1(n19328), .B2(net230381), 
        .ZN(n7456) );
  OAI22_X2 U17658 ( .A1(n19328), .A2(net231253), .B1(n13481), .B2(n16665), 
        .ZN(n7457) );
  NAND2_X2 U17659 ( .A1(n13412), .A2(ID_EXEC_OUT[175]), .ZN(n16669) );
  NAND2_X2 U17660 ( .A1(DMEM_BUS_OUT[47]), .A2(net231319), .ZN(n16668) );
  NAND2_X2 U17661 ( .A1(n13414), .A2(DMEM_BUS_OUT[15]), .ZN(n16667) );
  NAND2_X2 U17662 ( .A1(n13416), .A2(MEM_WB_OUT[52]), .ZN(n16666) );
  NAND4_X2 U17663 ( .A1(n16669), .A2(n16668), .A3(n16667), .A4(n16666), .ZN(
        n7458) );
  OAI22_X2 U17664 ( .A1(n13419), .A2(n12796), .B1(n13417), .B2(n11853), .ZN(
        n16673) );
  OAI22_X2 U17665 ( .A1(n13423), .A2(n12866), .B1(n13422), .B2(n12865), .ZN(
        n16672) );
  NAND2_X2 U17666 ( .A1(REG_FILE_reg_out_17__15_), .A2(n13435), .ZN(n16670) );
  OAI221_X2 U17667 ( .B1(n13432), .B2(n12867), .C1(n13427), .C2(n12731), .A(
        n16670), .ZN(n16671) );
  AOI22_X2 U17668 ( .A1(REG_FILE_reg_out_25__15_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__15_), .B2(n10350), .ZN(n16681) );
  OAI22_X2 U17669 ( .A1(n12437), .A2(n13444), .B1(n12041), .B2(n13442), .ZN(
        n16676) );
  OAI22_X2 U17670 ( .A1(n10504), .A2(n13190), .B1(n12276), .B2(n18699), .ZN(
        n16675) );
  OAI22_X2 U17671 ( .A1(n12741), .A2(n13192), .B1(n12436), .B2(n13193), .ZN(
        n16674) );
  NAND4_X2 U17672 ( .A1(n16682), .A2(n16681), .A3(n16680), .A4(n16679), .ZN(
        n16706) );
  NAND2_X2 U17673 ( .A1(n13456), .A2(REG_FILE_reg_out_12__15_), .ZN(n16690) );
  AOI22_X2 U17674 ( .A1(n13464), .A2(REG_FILE_reg_out_0__15_), .B1(
        REG_FILE_reg_out_15__15_), .B2(n13466), .ZN(n16688) );
  NAND4_X2 U17675 ( .A1(n16691), .A2(n16690), .A3(n16689), .A4(n16688), .ZN(
        n16705) );
  NAND4_X2 U17676 ( .A1(n16703), .A2(n16702), .A3(n16701), .A4(n16700), .ZN(
        n16704) );
  NOR3_X4 U17677 ( .A1(n16706), .A2(n16705), .A3(n16704), .ZN(n16707) );
  OAI22_X2 U17678 ( .A1(n11516), .A2(net231253), .B1(net230379), .B2(n16707), 
        .ZN(n7459) );
  OAI221_X2 U17679 ( .B1(n12511), .B2(net231221), .C1(n16707), .C2(n13476), 
        .A(n17267), .ZN(n7460) );
  NOR2_X4 U17680 ( .A1(n2193), .A2(n2194), .ZN(n16720) );
  NOR4_X2 U17681 ( .A1(n2195), .A2(n16710), .A3(n16709), .A4(n16708), .ZN(
        n16718) );
  OAI22_X2 U17682 ( .A1(n12435), .A2(n13383), .B1(n13380), .B2(n12750), .ZN(
        n16715) );
  OAI222_X2 U17683 ( .A1(n11853), .A2(n13374), .B1(n10253), .B2(n13370), .C1(
        n13368), .C2(n12741), .ZN(n16714) );
  NAND4_X2 U17684 ( .A1(n16720), .A2(n16719), .A3(n16718), .A4(n16717), .ZN(
        n16721) );
  MUX2_X2 U17685 ( .A(n16721), .B(ID_EXEC_OUT[47]), .S(net231295), .Z(n7461)
         );
  MUX2_X2 U17686 ( .A(MEM_WB_REG_MEM_WB_REG_N165), .B(MEM_WB_OUT[15]), .S(
        net231293), .Z(n7462) );
  OAI22_X2 U17687 ( .A1(n12189), .A2(net231253), .B1(n13481), .B2(n16722), 
        .ZN(n7465) );
  XNOR2_X2 U17688 ( .A(net225527), .B(net225526), .ZN(n16724) );
  OAI221_X2 U17689 ( .B1(net231229), .B2(n11474), .C1(n16724), .C2(net231915), 
        .A(n16723), .ZN(n7466) );
  NAND2_X2 U17690 ( .A1(n13412), .A2(ID_EXEC_OUT[176]), .ZN(n16728) );
  NAND2_X2 U17691 ( .A1(DMEM_BUS_OUT[48]), .A2(net231321), .ZN(n16727) );
  NAND2_X2 U17692 ( .A1(n13414), .A2(DMEM_BUS_OUT[16]), .ZN(n16726) );
  NAND2_X2 U17693 ( .A1(n13416), .A2(MEM_WB_OUT[53]), .ZN(n16725) );
  NAND4_X2 U17694 ( .A1(n16728), .A2(n16727), .A3(n16726), .A4(n16725), .ZN(
        n7467) );
  NAND2_X2 U17695 ( .A1(REG_FILE_reg_out_17__16_), .A2(n13435), .ZN(n16734) );
  OAI22_X2 U17696 ( .A1(n13419), .A2(n12797), .B1(n13418), .B2(n11854), .ZN(
        n16737) );
  OAI22_X2 U17697 ( .A1(n13440), .A2(n12585), .B1(n13438), .B2(n12570), .ZN(
        n16736) );
  NAND2_X2 U17698 ( .A1(n18493), .A2(REG_FILE_reg_out_6__16_), .ZN(n16742) );
  NAND2_X2 U17699 ( .A1(n13191), .A2(REG_FILE_reg_out_7__16_), .ZN(n16741) );
  NAND2_X2 U17700 ( .A1(n18494), .A2(REG_FILE_reg_out_4__16_), .ZN(n16740) );
  NAND2_X2 U17701 ( .A1(n13189), .A2(REG_FILE_reg_out_5__16_), .ZN(n16739) );
  NAND4_X2 U17702 ( .A1(n16742), .A2(n16741), .A3(n16740), .A4(n16739), .ZN(
        n16745) );
  OAI22_X2 U17703 ( .A1(n12290), .A2(n13445), .B1(n10927), .B2(n13443), .ZN(
        n16744) );
  OAI22_X2 U17704 ( .A1(n12776), .A2(n13451), .B1(n10520), .B2(n13448), .ZN(
        n16743) );
  NOR3_X4 U17705 ( .A1(n16745), .A2(n16744), .A3(n16743), .ZN(n16763) );
  NAND2_X2 U17706 ( .A1(n13198), .A2(REG_FILE_reg_out_14__16_), .ZN(n16749) );
  NAND2_X2 U17707 ( .A1(n13200), .A2(REG_FILE_reg_out_1__16_), .ZN(n16748) );
  NAND2_X2 U17708 ( .A1(n18502), .A2(REG_FILE_reg_out_11__16_), .ZN(n16747) );
  NAND2_X2 U17709 ( .A1(n13203), .A2(REG_FILE_reg_out_13__16_), .ZN(n16746) );
  NAND4_X2 U17710 ( .A1(n16749), .A2(n16748), .A3(n16747), .A4(n16746), .ZN(
        n16752) );
  OAI22_X2 U17711 ( .A1(n12137), .A2(n13471), .B1(n10493), .B2(n13467), .ZN(
        n16751) );
  OAI22_X2 U17712 ( .A1(n12261), .A2(n13475), .B1(n10492), .B2(n13472), .ZN(
        n16750) );
  NOR3_X4 U17713 ( .A1(n16752), .A2(n16751), .A3(n16750), .ZN(n16762) );
  NAND2_X2 U17714 ( .A1(n13456), .A2(REG_FILE_reg_out_12__16_), .ZN(n16757) );
  NAND2_X2 U17715 ( .A1(n13194), .A2(REG_FILE_reg_out_19__16_), .ZN(n16756) );
  NAND3_X4 U17716 ( .A1(n16757), .A2(n16756), .A3(n16755), .ZN(n16760) );
  OAI22_X2 U17717 ( .A1(n13460), .A2(n12870), .B1(n13459), .B2(n12751), .ZN(
        n16759) );
  OAI22_X2 U17718 ( .A1(n13465), .A2(n12798), .B1(n12403), .B2(n13463), .ZN(
        n16758) );
  NOR3_X4 U17719 ( .A1(n16760), .A2(n16759), .A3(n16758), .ZN(n16761) );
  NAND4_X2 U17720 ( .A1(n16764), .A2(n16763), .A3(n16762), .A4(n16761), .ZN(
        n16765) );
  INV_X4 U17721 ( .A(n16765), .ZN(n16767) );
  OAI22_X2 U17722 ( .A1(n11517), .A2(net231255), .B1(net230379), .B2(n16767), 
        .ZN(n7468) );
  OAI221_X2 U17723 ( .B1(n12320), .B2(net231221), .C1(n16767), .C2(n13476), 
        .A(n16766), .ZN(n7469) );
  OAI22_X2 U17724 ( .A1(n11103), .A2(net231253), .B1(net230379), .B2(n11928), 
        .ZN(n7472) );
  OAI22_X2 U17725 ( .A1(net231249), .A2(n11928), .B1(n12185), .B2(net230381), 
        .ZN(n7473) );
  OAI22_X2 U17726 ( .A1(n12185), .A2(net231255), .B1(n13481), .B2(n16768), 
        .ZN(n7474) );
  XNOR2_X2 U17727 ( .A(net225448), .B(net225449), .ZN(n16771) );
  NAND2_X2 U17728 ( .A1(EXEC_MEM_OUT_125), .A2(net231323), .ZN(n16769) );
  OAI211_X2 U17729 ( .C1(n16771), .C2(net231915), .A(n16770), .B(n16769), .ZN(
        n7475) );
  MUX2_X2 U17730 ( .A(DMEM_BUS_OUT[16]), .B(MEM_WB_OUT[53]), .S(net231295), 
        .Z(n7476) );
  NAND2_X2 U17731 ( .A1(n13358), .A2(n16971), .ZN(n16773) );
  NAND2_X2 U17732 ( .A1(n13389), .A2(n17697), .ZN(n16779) );
  NAND2_X2 U17733 ( .A1(n13358), .A2(net225212), .ZN(n16775) );
  NAND2_X2 U17734 ( .A1(n13396), .A2(n17587), .ZN(n16778) );
  NAND2_X2 U17735 ( .A1(n13393), .A2(n17585), .ZN(n16777) );
  NAND2_X2 U17736 ( .A1(n13488), .A2(n17586), .ZN(n16776) );
  NAND4_X2 U17737 ( .A1(n16779), .A2(n16778), .A3(n16777), .A4(n16776), .ZN(
        n17878) );
  NAND2_X2 U17738 ( .A1(n19118), .A2(n17878), .ZN(n16829) );
  INV_X4 U17739 ( .A(n16783), .ZN(n16784) );
  AOI21_X4 U17740 ( .B1(n18562), .B2(n16785), .A(n16784), .ZN(n17131) );
  XNOR2_X2 U17741 ( .A(n16788), .B(n16787), .ZN(n16789) );
  NAND2_X2 U17742 ( .A1(n13358), .A2(n19029), .ZN(n18629) );
  INV_X4 U17743 ( .A(n16790), .ZN(n16793) );
  NOR2_X4 U17744 ( .A1(n16793), .A2(n16792), .ZN(n16794) );
  OAI211_X2 U17747 ( .C1(n18534), .C2(n16797), .A(n16796), .B(n16795), .ZN(
        n17909) );
  NAND2_X2 U17748 ( .A1(n13396), .A2(n17909), .ZN(n16800) );
  NAND2_X2 U17749 ( .A1(n13392), .A2(n17747), .ZN(n16799) );
  NAND2_X2 U17750 ( .A1(n13488), .A2(n17910), .ZN(n16798) );
  NAND4_X2 U17751 ( .A1(n16801), .A2(n16800), .A3(n16799), .A4(n16798), .ZN(
        n17145) );
  INV_X4 U17752 ( .A(n17145), .ZN(n16809) );
  NAND2_X2 U17753 ( .A1(n13386), .A2(n18980), .ZN(n17844) );
  NAND2_X2 U17754 ( .A1(n13358), .A2(n13159), .ZN(n16802) );
  NAND2_X2 U17755 ( .A1(n17844), .A2(n16802), .ZN(n17686) );
  NAND2_X2 U17756 ( .A1(n13392), .A2(n17686), .ZN(n16807) );
  NAND2_X2 U17757 ( .A1(n13358), .A2(n13163), .ZN(n16803) );
  NAND2_X2 U17758 ( .A1(n13386), .A2(n17505), .ZN(n17510) );
  NAND2_X2 U17759 ( .A1(n16803), .A2(n17510), .ZN(n17596) );
  NAND2_X2 U17760 ( .A1(n13488), .A2(n17596), .ZN(n16806) );
  NAND2_X2 U17761 ( .A1(n13389), .A2(n17598), .ZN(n16805) );
  NAND2_X2 U17762 ( .A1(n13396), .A2(n17595), .ZN(n16804) );
  NAND4_X2 U17763 ( .A1(n16807), .A2(n16806), .A3(n16805), .A4(n16804), .ZN(
        n17872) );
  NAND2_X2 U17764 ( .A1(n10199), .A2(n17872), .ZN(n16808) );
  OAI21_X4 U17765 ( .B1(n16809), .B2(n18003), .A(n16808), .ZN(n16814) );
  NAND2_X2 U17766 ( .A1(n18566), .A2(DMEM_BUS_OUT[16]), .ZN(n16811) );
  AOI21_X4 U17767 ( .B1(n18651), .B2(n16814), .A(n16813), .ZN(n16827) );
  NAND2_X2 U17768 ( .A1(n13386), .A2(n18922), .ZN(n17988) );
  NAND2_X2 U17769 ( .A1(n17988), .A2(n16815), .ZN(n17918) );
  NAND2_X2 U17770 ( .A1(n13392), .A2(n17918), .ZN(n16821) );
  NAND2_X2 U17771 ( .A1(n13358), .A2(n13161), .ZN(n16817) );
  NAND2_X2 U17772 ( .A1(n13386), .A2(n17712), .ZN(n17693) );
  NAND2_X2 U17773 ( .A1(n16817), .A2(n17693), .ZN(n17916) );
  NAND2_X2 U17774 ( .A1(n13488), .A2(n17916), .ZN(n16820) );
  NAND2_X2 U17775 ( .A1(n13396), .A2(n17917), .ZN(n16818) );
  NAND4_X2 U17776 ( .A1(n16821), .A2(n16820), .A3(n16819), .A4(n16818), .ZN(
        n17149) );
  NAND2_X2 U17777 ( .A1(DMEM_BUS_OUT[16]), .A2(net231323), .ZN(n16822) );
  NAND4_X2 U17778 ( .A1(n16829), .A2(n16828), .A3(n16827), .A4(n16826), .ZN(
        n7477) );
  NAND2_X2 U17779 ( .A1(n13410), .A2(n18873), .ZN(n16830) );
  OAI211_X2 U17780 ( .C1(n12148), .C2(net231225), .A(n16830), .B(n6780), .ZN(
        n7481) );
  OAI22_X2 U17781 ( .A1(n13419), .A2(n12799), .B1(n13418), .B2(n11855), .ZN(
        n16834) );
  OAI22_X2 U17782 ( .A1(n13423), .A2(n12872), .B1(n13422), .B2(n12871), .ZN(
        n16833) );
  NAND2_X2 U17783 ( .A1(REG_FILE_reg_out_17__2_), .A2(n13435), .ZN(n16831) );
  OAI221_X2 U17784 ( .B1(n13432), .B2(n12873), .C1(n13427), .C2(n12732), .A(
        n16831), .ZN(n16832) );
  AOI22_X2 U17785 ( .A1(REG_FILE_reg_out_25__2_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__2_), .B2(n13441), .ZN(n16842) );
  OAI22_X2 U17786 ( .A1(n12389), .A2(n13445), .B1(n10507), .B2(n13443), .ZN(
        n16837) );
  OAI22_X2 U17787 ( .A1(n10303), .A2(n13190), .B1(n10700), .B2(n18699), .ZN(
        n16836) );
  OAI22_X2 U17788 ( .A1(n11840), .A2(n13192), .B1(n12388), .B2(n13193), .ZN(
        n16835) );
  NAND4_X2 U17789 ( .A1(n16843), .A2(n16842), .A3(n16841), .A4(n16840), .ZN(
        n16868) );
  NAND2_X2 U17790 ( .A1(n13456), .A2(REG_FILE_reg_out_12__2_), .ZN(n16852) );
  AOI22_X2 U17791 ( .A1(n13464), .A2(REG_FILE_reg_out_0__2_), .B1(
        REG_FILE_reg_out_15__2_), .B2(n13466), .ZN(n16850) );
  NAND4_X2 U17792 ( .A1(n16853), .A2(n16852), .A3(n16851), .A4(n16850), .ZN(
        n16867) );
  NAND4_X2 U17793 ( .A1(n16865), .A2(n16864), .A3(n16863), .A4(n16862), .ZN(
        n16866) );
  NOR3_X4 U17794 ( .A1(n16868), .A2(n16867), .A3(n16866), .ZN(n16869) );
  OAI22_X2 U17795 ( .A1(n11518), .A2(net231253), .B1(net230379), .B2(n16869), 
        .ZN(n7482) );
  OAI221_X2 U17796 ( .B1(n12512), .B2(net231221), .C1(n16869), .C2(n13476), 
        .A(n17267), .ZN(n7483) );
  NAND2_X2 U17797 ( .A1(n18566), .A2(DMEM_BUS_OUT[2]), .ZN(n16873) );
  INV_X4 U17798 ( .A(n16892), .ZN(n18874) );
  NAND2_X2 U17799 ( .A1(n13397), .A2(n16877), .ZN(n16881) );
  NAND2_X2 U17800 ( .A1(n13390), .A2(n16878), .ZN(n16880) );
  NAND2_X2 U17801 ( .A1(n16879), .A2(n18862), .ZN(n17305) );
  AOI22_X2 U17802 ( .A1(n19118), .A2(n16882), .B1(n17924), .B2(n17565), .ZN(
        n16896) );
  NAND2_X2 U17803 ( .A1(n16300), .A2(n16883), .ZN(n16890) );
  NAND2_X2 U17804 ( .A1(n13397), .A2(n16885), .ZN(n16888) );
  NAND2_X2 U17805 ( .A1(n13390), .A2(n16886), .ZN(n16887) );
  NAND4_X2 U17806 ( .A1(n16890), .A2(n16889), .A3(n16888), .A4(n16887), .ZN(
        n17561) );
  NAND2_X2 U17807 ( .A1(DMEM_BUS_OUT[2]), .A2(net231323), .ZN(n16891) );
  XNOR2_X2 U17808 ( .A(n16892), .B(n18873), .ZN(n19047) );
  NAND3_X4 U17809 ( .A1(n16897), .A2(n16896), .A3(n16895), .ZN(n16901) );
  INV_X4 U17810 ( .A(n16901), .ZN(n16904) );
  NAND2_X2 U17811 ( .A1(n17557), .A2(n18595), .ZN(n18602) );
  NAND2_X2 U17812 ( .A1(n18594), .A2(n18595), .ZN(n16898) );
  OAI21_X4 U17813 ( .B1(n16899), .B2(n18602), .A(n16898), .ZN(n16900) );
  XNOR2_X2 U17814 ( .A(n16900), .B(n18597), .ZN(n16903) );
  NOR2_X4 U17815 ( .A1(n13492), .A2(n16901), .ZN(n16902) );
  OAI22_X2 U17816 ( .A1(n13420), .A2(n12800), .B1(n13418), .B2(n11856), .ZN(
        n16908) );
  OAI22_X2 U17817 ( .A1(n13423), .A2(n12876), .B1(n13422), .B2(n12875), .ZN(
        n16907) );
  NAND2_X2 U17818 ( .A1(REG_FILE_reg_out_17__3_), .A2(n13435), .ZN(n16905) );
  OAI221_X2 U17819 ( .B1(n13432), .B2(n12877), .C1(n13427), .C2(n12733), .A(
        n16905), .ZN(n16906) );
  AOI22_X2 U17820 ( .A1(REG_FILE_reg_out_25__3_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__3_), .B2(n13441), .ZN(n16916) );
  OAI22_X2 U17821 ( .A1(n12445), .A2(n13445), .B1(n10508), .B2(n13443), .ZN(
        n16911) );
  OAI22_X2 U17822 ( .A1(n10304), .A2(n13190), .B1(n10701), .B2(n18699), .ZN(
        n16910) );
  OAI22_X2 U17823 ( .A1(n12742), .A2(n13192), .B1(n12444), .B2(n13193), .ZN(
        n16909) );
  NAND4_X2 U17824 ( .A1(n16917), .A2(n16916), .A3(n16915), .A4(n16914), .ZN(
        n16942) );
  INV_X4 U17825 ( .A(n16918), .ZN(n17570) );
  NAND2_X2 U17826 ( .A1(n13456), .A2(REG_FILE_reg_out_12__3_), .ZN(n16926) );
  AOI22_X2 U17827 ( .A1(n13464), .A2(REG_FILE_reg_out_0__3_), .B1(
        REG_FILE_reg_out_15__3_), .B2(n13466), .ZN(n16924) );
  NAND4_X2 U17828 ( .A1(n16927), .A2(n16926), .A3(n16925), .A4(n16924), .ZN(
        n16941) );
  NAND4_X2 U17829 ( .A1(n16939), .A2(n16938), .A3(n16937), .A4(n16936), .ZN(
        n16940) );
  NOR3_X4 U17830 ( .A1(n16942), .A2(n16941), .A3(n16940), .ZN(n16943) );
  OAI22_X2 U17831 ( .A1(n11519), .A2(net231253), .B1(net230379), .B2(n16943), 
        .ZN(n7487) );
  OAI221_X2 U17832 ( .B1(n12513), .B2(net231221), .C1(n16943), .C2(n13476), 
        .A(n17267), .ZN(n7488) );
  NOR2_X4 U17833 ( .A1(n2439), .A2(n2440), .ZN(n16955) );
  NOR4_X2 U17834 ( .A1(n2441), .A2(n16946), .A3(n16945), .A4(n16944), .ZN(
        n16953) );
  OAI22_X2 U17835 ( .A1(n12443), .A2(n13383), .B1(n13380), .B2(n12752), .ZN(
        n16950) );
  OAI222_X2 U17836 ( .A1(n11856), .A2(n13374), .B1(n10254), .B2(n13370), .C1(
        n13368), .C2(n12742), .ZN(n16949) );
  NAND4_X2 U17837 ( .A1(n16955), .A2(n16954), .A3(n16953), .A4(n16952), .ZN(
        n16956) );
  MUX2_X2 U17838 ( .A(n16956), .B(ID_EXEC_OUT[35]), .S(net231295), .Z(n7489)
         );
  MUX2_X2 U17839 ( .A(MEM_WB_REG_MEM_WB_REG_N177), .B(MEM_WB_OUT[3]), .S(
        net231295), .Z(n7490) );
  OAI22_X2 U17840 ( .A1(n12305), .A2(net231255), .B1(n13481), .B2(n16957), 
        .ZN(n7493) );
  MUX2_X2 U17841 ( .A(MEM_WB_REG_MEM_WB_REG_N175), .B(MEM_WB_OUT[5]), .S(
        net231295), .Z(n7495) );
  OAI22_X2 U17842 ( .A1(n12193), .A2(net231257), .B1(n13481), .B2(n16958), 
        .ZN(n7498) );
  NOR2_X4 U17843 ( .A1(n19349), .A2(n10357), .ZN(n16959) );
  NAND2_X2 U17844 ( .A1(net224704), .A2(nextPC_ex_out[6]), .ZN(n16961) );
  NAND2_X2 U17845 ( .A1(n16962), .A2(n16961), .ZN(n16963) );
  OAI22_X2 U17846 ( .A1(nextPC_ex_out[6]), .A2(net225187), .B1(n10356), .B2(
        net225188), .ZN(net225184) );
  OAI22_X2 U17847 ( .A1(n10356), .A2(net225187), .B1(nextPC_ex_out[6]), .B2(
        net225188), .ZN(net225186) );
  MUX2_X2 U17848 ( .A(MEM_WB_REG_MEM_WB_REG_N174), .B(MEM_WB_OUT[6]), .S(
        net231293), .Z(n7500) );
  OAI22_X2 U17849 ( .A1(n12194), .A2(net231253), .B1(n13481), .B2(n16968), 
        .ZN(n7503) );
  XNOR2_X2 U17850 ( .A(n16969), .B(nextPC_ex_out[7]), .ZN(n16970) );
  AOI22_X2 U17851 ( .A1(EXEC_MEM_OUT_116), .A2(net231307), .B1(net231615), 
        .B2(n16971), .ZN(n16972) );
  MUX2_X2 U17852 ( .A(MEM_WB_REG_MEM_WB_REG_N172), .B(MEM_WB_OUT[8]), .S(
        net231295), .Z(n7505) );
  OAI22_X2 U17853 ( .A1(n12196), .A2(net231255), .B1(n13481), .B2(n16974), 
        .ZN(n7508) );
  XNOR2_X2 U17854 ( .A(net227019), .B(net225160), .ZN(n16978) );
  NAND2_X2 U17855 ( .A1(net231615), .A2(n19029), .ZN(n16977) );
  NAND2_X2 U17856 ( .A1(EXEC_MEM_OUT_117), .A2(net231319), .ZN(n16976) );
  OAI211_X2 U17857 ( .C1(n16978), .C2(net231915), .A(n16977), .B(n16976), .ZN(
        n7509) );
  OAI22_X2 U17858 ( .A1(n13419), .A2(n12801), .B1(n13418), .B2(n11857), .ZN(
        n16982) );
  OAI22_X2 U17859 ( .A1(n13423), .A2(n12880), .B1(n13422), .B2(n12879), .ZN(
        n16981) );
  NAND2_X2 U17860 ( .A1(REG_FILE_reg_out_17__9_), .A2(n13435), .ZN(n16979) );
  OAI221_X2 U17861 ( .B1(n13431), .B2(n12881), .C1(n13427), .C2(n12734), .A(
        n16979), .ZN(n16980) );
  AOI22_X2 U17862 ( .A1(REG_FILE_reg_out_25__9_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__9_), .B2(n13441), .ZN(n16990) );
  OAI22_X2 U17863 ( .A1(n12449), .A2(n13445), .B1(n10514), .B2(n13443), .ZN(
        n16985) );
  OAI22_X2 U17864 ( .A1(n10310), .A2(n13190), .B1(n10702), .B2(n18699), .ZN(
        n16984) );
  OAI22_X2 U17865 ( .A1(n12743), .A2(n13192), .B1(n12448), .B2(n13193), .ZN(
        n16983) );
  NAND4_X2 U17866 ( .A1(n16991), .A2(n16990), .A3(n16989), .A4(n16988), .ZN(
        n17015) );
  NAND2_X2 U17867 ( .A1(n13456), .A2(REG_FILE_reg_out_12__9_), .ZN(n16999) );
  AOI22_X2 U17868 ( .A1(n13464), .A2(REG_FILE_reg_out_0__9_), .B1(
        REG_FILE_reg_out_15__9_), .B2(n13466), .ZN(n16997) );
  NAND4_X2 U17869 ( .A1(n17000), .A2(n16999), .A3(n16998), .A4(n16997), .ZN(
        n17014) );
  NAND4_X2 U17870 ( .A1(n17012), .A2(n17011), .A3(n17010), .A4(n17009), .ZN(
        n17013) );
  NOR3_X4 U17871 ( .A1(n17015), .A2(n17014), .A3(n17013), .ZN(n17016) );
  OAI22_X2 U17872 ( .A1(n11520), .A2(net231255), .B1(net230379), .B2(n17016), 
        .ZN(n7510) );
  OAI221_X2 U17873 ( .B1(n12514), .B2(net231221), .C1(n17016), .C2(n13476), 
        .A(n17267), .ZN(n7511) );
  NOR2_X4 U17874 ( .A1(n2318), .A2(n2319), .ZN(n17029) );
  NOR4_X2 U17875 ( .A1(n2320), .A2(n17019), .A3(n17018), .A4(n17017), .ZN(
        n17027) );
  OAI22_X2 U17876 ( .A1(n12447), .A2(n13383), .B1(n13380), .B2(n12753), .ZN(
        n17024) );
  OAI222_X2 U17877 ( .A1(n11857), .A2(n13374), .B1(n10255), .B2(n13370), .C1(
        n13368), .C2(n12743), .ZN(n17023) );
  NAND4_X2 U17878 ( .A1(n17029), .A2(n17028), .A3(n17027), .A4(n17026), .ZN(
        n17030) );
  MUX2_X2 U17879 ( .A(n17030), .B(ID_EXEC_OUT[41]), .S(net231293), .Z(n7512)
         );
  MUX2_X2 U17880 ( .A(MEM_WB_REG_MEM_WB_REG_N171), .B(MEM_WB_OUT[9]), .S(
        net231295), .Z(n7513) );
  OAI22_X2 U17881 ( .A1(net137185), .A2(net231255), .B1(n13481), .B2(n17031), 
        .ZN(n7516) );
  XNOR2_X2 U17882 ( .A(net225077), .B(nextPC_ex_out[9]), .ZN(n17033) );
  XNOR2_X2 U17883 ( .A(n17032), .B(n17033), .ZN(n17035) );
  NAND2_X2 U17884 ( .A1(net231615), .A2(n19013), .ZN(n17034) );
  INV_X4 U17885 ( .A(n17036), .ZN(n17039) );
  INV_X4 U17886 ( .A(n17037), .ZN(n17038) );
  INV_X4 U17887 ( .A(n17041), .ZN(n17042) );
  XNOR2_X2 U17888 ( .A(n17043), .B(n17042), .ZN(n17044) );
  OAI22_X2 U17889 ( .A1(n17020), .A2(n18569), .B1(n13209), .B2(n17046), .ZN(
        n17047) );
  XNOR2_X2 U17890 ( .A(n19012), .B(n19013), .ZN(n17049) );
  INV_X4 U17891 ( .A(n17049), .ZN(n19023) );
  NAND2_X2 U17892 ( .A1(n13490), .A2(n19023), .ZN(n17063) );
  NAND2_X2 U17893 ( .A1(DMEM_BUS_OUT[9]), .A2(net231323), .ZN(n17055) );
  NAND2_X2 U17894 ( .A1(ID_EXEC_OUT[213]), .A2(n13216), .ZN(n17054) );
  NAND2_X2 U17895 ( .A1(n18360), .A2(n17050), .ZN(n17053) );
  NAND2_X2 U17896 ( .A1(n19118), .A2(n17051), .ZN(n17052) );
  NAND4_X2 U17897 ( .A1(n17055), .A2(n17054), .A3(n17053), .A4(n17052), .ZN(
        n17061) );
  INV_X4 U17898 ( .A(n17056), .ZN(n17059) );
  INV_X4 U17899 ( .A(n17057), .ZN(n17058) );
  OAI22_X2 U17900 ( .A1(n17059), .A2(n13211), .B1(n17058), .B2(n13207), .ZN(
        n17060) );
  NOR2_X4 U17901 ( .A1(n17061), .A2(n17060), .ZN(n17062) );
  NAND4_X2 U17902 ( .A1(n17065), .A2(n17064), .A3(n17063), .A4(n17062), .ZN(
        n7519) );
  NAND2_X2 U17903 ( .A1(n13412), .A2(ID_EXEC_OUT[177]), .ZN(n17069) );
  NAND2_X2 U17904 ( .A1(DMEM_BUS_OUT[49]), .A2(net231319), .ZN(n17068) );
  NAND2_X2 U17905 ( .A1(n13414), .A2(DMEM_BUS_OUT[17]), .ZN(n17067) );
  NAND2_X2 U17906 ( .A1(n13416), .A2(MEM_WB_OUT[54]), .ZN(n17066) );
  NAND4_X2 U17907 ( .A1(n17069), .A2(n17068), .A3(n17067), .A4(n17066), .ZN(
        n7520) );
  NAND2_X2 U17908 ( .A1(REG_FILE_reg_out_17__17_), .A2(n13435), .ZN(n17075) );
  OAI22_X2 U17909 ( .A1(n13420), .A2(n12802), .B1(n13418), .B2(n11858), .ZN(
        n17078) );
  OAI22_X2 U17910 ( .A1(n13440), .A2(n12586), .B1(n13438), .B2(n12571), .ZN(
        n17077) );
  NAND2_X2 U17911 ( .A1(n18493), .A2(REG_FILE_reg_out_6__17_), .ZN(n17083) );
  NAND2_X2 U17912 ( .A1(n13191), .A2(REG_FILE_reg_out_7__17_), .ZN(n17082) );
  NAND2_X2 U17913 ( .A1(n18494), .A2(REG_FILE_reg_out_4__17_), .ZN(n17081) );
  NAND2_X2 U17914 ( .A1(n13189), .A2(REG_FILE_reg_out_5__17_), .ZN(n17080) );
  NAND4_X2 U17915 ( .A1(n17083), .A2(n17082), .A3(n17081), .A4(n17080), .ZN(
        n17086) );
  OAI22_X2 U17916 ( .A1(n12291), .A2(n13445), .B1(n10928), .B2(n13443), .ZN(
        n17085) );
  OAI22_X2 U17917 ( .A1(n12754), .A2(n13450), .B1(n10316), .B2(n13447), .ZN(
        n17084) );
  NOR3_X4 U17918 ( .A1(n17086), .A2(n17085), .A3(n17084), .ZN(n17104) );
  NAND2_X2 U17919 ( .A1(n13198), .A2(REG_FILE_reg_out_14__17_), .ZN(n17090) );
  NAND2_X2 U17920 ( .A1(n13200), .A2(REG_FILE_reg_out_1__17_), .ZN(n17089) );
  NAND2_X2 U17921 ( .A1(n18502), .A2(REG_FILE_reg_out_11__17_), .ZN(n17088) );
  NAND2_X2 U17922 ( .A1(n13203), .A2(REG_FILE_reg_out_13__17_), .ZN(n17087) );
  NAND4_X2 U17923 ( .A1(n17090), .A2(n17089), .A3(n17088), .A4(n17087), .ZN(
        n17093) );
  OAI22_X2 U17924 ( .A1(n11274), .A2(n13470), .B1(n10495), .B2(n13468), .ZN(
        n17092) );
  OAI22_X2 U17925 ( .A1(n11275), .A2(n13474), .B1(n10494), .B2(n13473), .ZN(
        n17091) );
  NOR3_X4 U17926 ( .A1(n17093), .A2(n17092), .A3(n17091), .ZN(n17103) );
  NAND2_X2 U17927 ( .A1(n13456), .A2(REG_FILE_reg_out_12__17_), .ZN(n17098) );
  NAND2_X2 U17928 ( .A1(n13194), .A2(REG_FILE_reg_out_19__17_), .ZN(n17097) );
  INV_X4 U17929 ( .A(n17094), .ZN(n17141) );
  NAND3_X4 U17930 ( .A1(n17098), .A2(n17097), .A3(n17096), .ZN(n17101) );
  OAI22_X2 U17931 ( .A1(n13461), .A2(n12884), .B1(n13458), .B2(n11859), .ZN(
        n17100) );
  OAI22_X2 U17932 ( .A1(n13465), .A2(n12803), .B1(n12404), .B2(n13463), .ZN(
        n17099) );
  NOR3_X4 U17933 ( .A1(n17101), .A2(n17100), .A3(n17099), .ZN(n17102) );
  NAND4_X2 U17934 ( .A1(n17105), .A2(n17104), .A3(n17103), .A4(n17102), .ZN(
        n17106) );
  INV_X4 U17935 ( .A(n17106), .ZN(n17107) );
  OAI22_X2 U17936 ( .A1(n11521), .A2(net231255), .B1(net230379), .B2(n17107), 
        .ZN(n7521) );
  OAI222_X2 U17937 ( .A1(n17107), .A2(n13477), .B1(n12517), .B2(net231223), 
        .C1(n10807), .C2(n13206), .ZN(n7522) );
  NOR2_X4 U17938 ( .A1(n2150), .A2(n17108), .ZN(n17114) );
  NOR2_X4 U17939 ( .A1(n2147), .A2(n2149), .ZN(n17113) );
  OAI222_X2 U17940 ( .A1(n11858), .A2(n13374), .B1(n10230), .B2(n13370), .C1(
        n13368), .C2(n11697), .ZN(n17111) );
  OAI22_X2 U17941 ( .A1(n11859), .A2(n13383), .B1(n13380), .B2(n12754), .ZN(
        n17109) );
  NOR3_X4 U17942 ( .A1(n17111), .A2(n17110), .A3(n17109), .ZN(n17112) );
  NAND3_X2 U17943 ( .A1(n17114), .A2(n17113), .A3(n17112), .ZN(n17115) );
  MUX2_X2 U17944 ( .A(n17115), .B(ID_EXEC_OUT[49]), .S(net231293), .Z(n7523)
         );
  OAI22_X2 U17945 ( .A1(n12186), .A2(net231257), .B1(n13481), .B2(n17116), 
        .ZN(n7527) );
  XNOR2_X2 U17946 ( .A(net224953), .B(net224952), .ZN(n17119) );
  NAND2_X2 U17947 ( .A1(net231615), .A2(n18888), .ZN(n17118) );
  NAND2_X2 U17948 ( .A1(EXEC_MEM_OUT_126), .A2(net231323), .ZN(n17117) );
  OAI211_X2 U17949 ( .C1(n17119), .C2(net231915), .A(n17118), .B(n17117), .ZN(
        n7528) );
  NAND2_X2 U17950 ( .A1(n13488), .A2(n17587), .ZN(n17129) );
  INV_X4 U17951 ( .A(n17120), .ZN(n17123) );
  NOR2_X4 U17952 ( .A1(n17121), .A2(net232817), .ZN(n17122) );
  NAND2_X2 U17953 ( .A1(n13390), .A2(n17994), .ZN(n17128) );
  NAND2_X2 U17954 ( .A1(n13392), .A2(n17586), .ZN(n17127) );
  NAND2_X2 U17955 ( .A1(n13397), .A2(n17697), .ZN(n17126) );
  NAND4_X2 U17956 ( .A1(n17129), .A2(n17128), .A3(n17127), .A4(n17126), .ZN(
        n18581) );
  NAND2_X2 U17957 ( .A1(n17924), .A2(n18581), .ZN(n17153) );
  INV_X4 U17958 ( .A(n17130), .ZN(n17132) );
  XNOR2_X2 U17959 ( .A(n17131), .B(n17132), .ZN(n17133) );
  NAND2_X2 U17960 ( .A1(n13492), .A2(n17133), .ZN(n17152) );
  INV_X4 U17961 ( .A(n17540), .ZN(n17683) );
  AOI22_X2 U17962 ( .A1(n17596), .A2(n18943), .B1(n17683), .B2(n13149), .ZN(
        n17537) );
  NAND2_X2 U17963 ( .A1(n16300), .A2(n17686), .ZN(n17135) );
  NAND2_X2 U17964 ( .A1(n13390), .A2(n17595), .ZN(n17134) );
  OAI211_X2 U17965 ( .C1(n19100), .C2(n17537), .A(n17135), .B(n17134), .ZN(
        n17136) );
  INV_X4 U17966 ( .A(n17136), .ZN(n18573) );
  NAND2_X2 U17967 ( .A1(n17138), .A2(n13208), .ZN(n17140) );
  NAND2_X2 U17968 ( .A1(n18566), .A2(DMEM_BUS_OUT[17]), .ZN(n17139) );
  OAI211_X2 U17969 ( .C1(n17141), .C2(n18569), .A(n17140), .B(n17139), .ZN(
        n17142) );
  OAI21_X4 U17970 ( .B1(n18573), .B2(n13207), .A(n17143), .ZN(n17144) );
  NAND2_X2 U17971 ( .A1(DMEM_BUS_OUT[17]), .A2(net231323), .ZN(n17146) );
  XNOR2_X2 U17972 ( .A(n18890), .B(n18888), .ZN(n18887) );
  NAND4_X2 U17973 ( .A1(n17153), .A2(n17152), .A3(n17151), .A4(n17150), .ZN(
        n7530) );
  NAND2_X2 U17974 ( .A1(n13410), .A2(n18870), .ZN(n17154) );
  OAI211_X2 U17975 ( .C1(n12147), .C2(net231225), .A(n17154), .B(n6781), .ZN(
        n7534) );
  OAI22_X2 U17976 ( .A1(n13419), .A2(n12804), .B1(n13418), .B2(n11860), .ZN(
        n17158) );
  OAI22_X2 U17977 ( .A1(n13423), .A2(n12886), .B1(n13422), .B2(n12885), .ZN(
        n17157) );
  NAND2_X2 U17978 ( .A1(REG_FILE_reg_out_17__1_), .A2(n13435), .ZN(n17155) );
  OAI221_X2 U17979 ( .B1(n13431), .B2(n12887), .C1(n13427), .C2(n12735), .A(
        n17155), .ZN(n17156) );
  AOI22_X2 U17980 ( .A1(REG_FILE_reg_out_25__1_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__1_), .B2(n13441), .ZN(n17166) );
  OAI22_X2 U17981 ( .A1(n12386), .A2(n13445), .B1(n10506), .B2(n13443), .ZN(
        n17161) );
  OAI22_X2 U17982 ( .A1(n10302), .A2(n13190), .B1(n10703), .B2(n18699), .ZN(
        n17160) );
  OAI22_X2 U17983 ( .A1(n11839), .A2(n13192), .B1(n12385), .B2(n13193), .ZN(
        n17159) );
  NAND4_X2 U17984 ( .A1(n17167), .A2(n17166), .A3(n17165), .A4(n17164), .ZN(
        n17192) );
  NAND2_X2 U17985 ( .A1(n13456), .A2(REG_FILE_reg_out_12__1_), .ZN(n17176) );
  AOI22_X2 U17986 ( .A1(n13464), .A2(REG_FILE_reg_out_0__1_), .B1(
        REG_FILE_reg_out_15__1_), .B2(n13466), .ZN(n17174) );
  NAND4_X2 U17987 ( .A1(n17177), .A2(n17176), .A3(n17175), .A4(n17174), .ZN(
        n17191) );
  NAND4_X2 U17988 ( .A1(n17189), .A2(n17188), .A3(n17187), .A4(n17186), .ZN(
        n17190) );
  NOR3_X4 U17989 ( .A1(n17192), .A2(n17191), .A3(n17190), .ZN(n17193) );
  OAI22_X2 U17990 ( .A1(n11522), .A2(net231255), .B1(net230379), .B2(n17193), 
        .ZN(n7535) );
  OAI221_X2 U17991 ( .B1(n12515), .B2(net231221), .C1(n17193), .C2(n13476), 
        .A(n17267), .ZN(n7536) );
  MUX2_X2 U17992 ( .A(MEM_WB_REG_MEM_WB_REG_N179), .B(MEM_WB_OUT[1]), .S(
        net231293), .Z(n7538) );
  OAI22_X2 U17993 ( .A1(n12303), .A2(net231255), .B1(n13480), .B2(n17194), 
        .ZN(n7541) );
  NAND3_X4 U17994 ( .A1(n17215), .A2(n17197), .A3(net224816), .ZN(n17222) );
  NAND2_X2 U17995 ( .A1(nextPC_ex_out[3]), .A2(n10358), .ZN(n17198) );
  NOR3_X4 U17996 ( .A1(n17213), .A2(net224713), .A3(n17198), .ZN(n17199) );
  NAND2_X2 U17997 ( .A1(net224704), .A2(n10364), .ZN(n17212) );
  NAND2_X2 U17998 ( .A1(net224711), .A2(nextPC_ex_out[2]), .ZN(n17200) );
  OAI211_X2 U17999 ( .C1(nextPC_ex_out[2]), .C2(n17212), .A(n17201), .B(n17200), .ZN(n17206) );
  NAND2_X2 U18000 ( .A1(n17202), .A2(n10361), .ZN(n17203) );
  MUX2_X2 U18001 ( .A(MEM_WB_REG_MEM_WB_REG_N178), .B(MEM_WB_OUT[2]), .S(
        net231293), .Z(n7543) );
  OAI22_X2 U18002 ( .A1(n12304), .A2(net231255), .B1(n13480), .B2(n17211), 
        .ZN(n7546) );
  INV_X4 U18003 ( .A(n17212), .ZN(n17214) );
  NAND2_X2 U18004 ( .A1(net224711), .A2(nextPC_ex_out[3]), .ZN(n17223) );
  OAI22_X2 U18005 ( .A1(n13419), .A2(n12805), .B1(n13418), .B2(n11861), .ZN(
        n17232) );
  OAI22_X2 U18006 ( .A1(n13423), .A2(n12890), .B1(n13422), .B2(n12889), .ZN(
        n17231) );
  NAND2_X2 U18007 ( .A1(REG_FILE_reg_out_17__4_), .A2(n13435), .ZN(n17229) );
  OAI221_X2 U18008 ( .B1(n13432), .B2(n12891), .C1(n13427), .C2(n12736), .A(
        n17229), .ZN(n17230) );
  AOI22_X2 U18009 ( .A1(REG_FILE_reg_out_25__4_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__4_), .B2(n13441), .ZN(n17240) );
  OAI22_X2 U18010 ( .A1(n12457), .A2(n13445), .B1(n10509), .B2(n13443), .ZN(
        n17235) );
  OAI22_X2 U18011 ( .A1(n10305), .A2(n13190), .B1(n10704), .B2(n18699), .ZN(
        n17234) );
  OAI22_X2 U18012 ( .A1(n12744), .A2(n13192), .B1(n12456), .B2(n13193), .ZN(
        n17233) );
  NOR3_X4 U18013 ( .A1(n17235), .A2(n17234), .A3(n17233), .ZN(n17239) );
  NAND4_X2 U18014 ( .A1(n17241), .A2(n17240), .A3(n17239), .A4(n17238), .ZN(
        n17266) );
  INV_X4 U18015 ( .A(n17242), .ZN(n17313) );
  NAND2_X2 U18016 ( .A1(n13456), .A2(REG_FILE_reg_out_12__4_), .ZN(n17250) );
  AOI22_X2 U18017 ( .A1(n13464), .A2(REG_FILE_reg_out_0__4_), .B1(
        REG_FILE_reg_out_15__4_), .B2(n13466), .ZN(n17248) );
  NAND4_X2 U18018 ( .A1(n17251), .A2(n17250), .A3(n17249), .A4(n17248), .ZN(
        n17265) );
  NOR2_X4 U18019 ( .A1(n10981), .A2(n13204), .ZN(n17254) );
  NAND4_X2 U18020 ( .A1(n17263), .A2(n17262), .A3(n17261), .A4(n17260), .ZN(
        n17264) );
  NOR3_X4 U18021 ( .A1(n17266), .A2(n17265), .A3(n17264), .ZN(n17268) );
  OAI22_X2 U18022 ( .A1(n11523), .A2(net231255), .B1(net230379), .B2(n17268), 
        .ZN(n7548) );
  OAI221_X2 U18023 ( .B1(n17268), .B2(n13477), .C1(n12516), .C2(net231245), 
        .A(n17267), .ZN(n7549) );
  NOR2_X4 U18024 ( .A1(n2419), .A2(n2420), .ZN(n17282) );
  NOR4_X2 U18025 ( .A1(n2421), .A2(n17273), .A3(n17272), .A4(n17271), .ZN(
        n17280) );
  OAI22_X2 U18026 ( .A1(n12455), .A2(n13383), .B1(n13380), .B2(n12755), .ZN(
        n17277) );
  OAI222_X2 U18027 ( .A1(n11861), .A2(n13374), .B1(n10256), .B2(n13370), .C1(
        n13367), .C2(n12744), .ZN(n17276) );
  NAND4_X2 U18028 ( .A1(n17282), .A2(n17281), .A3(n17280), .A4(n17279), .ZN(
        n17283) );
  MUX2_X2 U18029 ( .A(n17283), .B(ID_EXEC_OUT[36]), .S(net231293), .Z(n7550)
         );
  MUX2_X2 U18030 ( .A(MEM_WB_REG_MEM_WB_REG_N176), .B(MEM_WB_OUT[4]), .S(
        net231293), .Z(n7551) );
  OAI22_X2 U18031 ( .A1(n19327), .A2(net231255), .B1(n13481), .B2(n17284), 
        .ZN(n7554) );
  NAND2_X2 U18032 ( .A1(net224711), .A2(nextPC_ex_out[4]), .ZN(net224710) );
  NAND2_X2 U18033 ( .A1(n17288), .A2(n17287), .ZN(n17289) );
  INV_X4 U18034 ( .A(n17294), .ZN(n17295) );
  OAI21_X4 U18035 ( .B1(n17295), .B2(n18611), .A(n18601), .ZN(n17296) );
  XNOR2_X2 U18036 ( .A(n17296), .B(n18612), .ZN(n17297) );
  NAND2_X2 U18037 ( .A1(n17297), .A2(n13492), .ZN(n17326) );
  NAND2_X2 U18038 ( .A1(n13397), .A2(n17298), .ZN(n17303) );
  NAND2_X2 U18039 ( .A1(n13390), .A2(n18636), .ZN(n17302) );
  AOI22_X2 U18040 ( .A1(n13392), .A2(n17300), .B1(n13487), .B2(n17299), .ZN(
        n17301) );
  NAND2_X2 U18041 ( .A1(n18360), .A2(n17575), .ZN(n17325) );
  NAND2_X2 U18042 ( .A1(n13397), .A2(n17304), .ZN(n17306) );
  OAI211_X2 U18043 ( .C1(n19101), .C2(n17307), .A(n17306), .B(n17305), .ZN(
        n17308) );
  INV_X4 U18044 ( .A(n17308), .ZN(n17574) );
  INV_X4 U18045 ( .A(n17309), .ZN(n17310) );
  NAND2_X2 U18046 ( .A1(n17310), .A2(n13208), .ZN(n17312) );
  NAND2_X2 U18047 ( .A1(n18566), .A2(DMEM_BUS_OUT[4]), .ZN(n17311) );
  OAI211_X2 U18048 ( .C1(n17313), .C2(n18569), .A(n17312), .B(n17311), .ZN(
        n17314) );
  NAND2_X2 U18049 ( .A1(n17314), .A2(n18866), .ZN(n17315) );
  NOR2_X4 U18050 ( .A1(n17318), .A2(n17317), .ZN(n17324) );
  NAND2_X2 U18051 ( .A1(DMEM_BUS_OUT[4]), .A2(net231323), .ZN(n17319) );
  XNOR2_X2 U18052 ( .A(n18866), .B(n18867), .ZN(n19044) );
  NAND4_X2 U18053 ( .A1(n17326), .A2(n17325), .A3(n17324), .A4(n17323), .ZN(
        n7557) );
  XNOR2_X2 U18054 ( .A(n17327), .B(net224658), .ZN(n17330) );
  NAND2_X2 U18055 ( .A1(net231615), .A2(n18559), .ZN(n17329) );
  NAND2_X2 U18056 ( .A1(EXEC_MEM_OUT_127), .A2(net231323), .ZN(n17328) );
  OAI211_X2 U18057 ( .C1(n17330), .C2(net231915), .A(n17329), .B(n17328), .ZN(
        n7558) );
  INV_X4 U18058 ( .A(n17331), .ZN(n18570) );
  NOR2_X4 U18059 ( .A1(n2129), .A2(n17332), .ZN(n17338) );
  NOR2_X4 U18060 ( .A1(n2126), .A2(n2128), .ZN(n17337) );
  OAI222_X2 U18061 ( .A1(n11862), .A2(n13374), .B1(n10231), .B2(n13370), .C1(
        n13367), .C2(n11700), .ZN(n17335) );
  OAI22_X2 U18062 ( .A1(n11863), .A2(n13383), .B1(n13380), .B2(n12756), .ZN(
        n17333) );
  NOR3_X4 U18063 ( .A1(n17335), .A2(n17334), .A3(n17333), .ZN(n17336) );
  NAND3_X2 U18064 ( .A1(n17338), .A2(n17337), .A3(n17336), .ZN(n17339) );
  MUX2_X2 U18065 ( .A(n17339), .B(ID_EXEC_OUT[50]), .S(net231293), .Z(n7559)
         );
  NAND2_X2 U18066 ( .A1(REG_FILE_reg_out_17__18_), .A2(n13435), .ZN(n17345) );
  OAI22_X2 U18067 ( .A1(n13419), .A2(n12806), .B1(n13418), .B2(n11862), .ZN(
        n17348) );
  OAI22_X2 U18068 ( .A1(n13440), .A2(n12587), .B1(n13438), .B2(n12572), .ZN(
        n17347) );
  NAND2_X2 U18069 ( .A1(n18493), .A2(REG_FILE_reg_out_6__18_), .ZN(n17353) );
  NAND2_X2 U18070 ( .A1(n13191), .A2(REG_FILE_reg_out_7__18_), .ZN(n17352) );
  NAND2_X2 U18071 ( .A1(n18494), .A2(REG_FILE_reg_out_4__18_), .ZN(n17351) );
  NAND2_X2 U18072 ( .A1(n13189), .A2(REG_FILE_reg_out_5__18_), .ZN(n17350) );
  NAND4_X2 U18073 ( .A1(n17353), .A2(n17352), .A3(n17351), .A4(n17350), .ZN(
        n17356) );
  OAI22_X2 U18074 ( .A1(n12292), .A2(n13445), .B1(n10929), .B2(n13443), .ZN(
        n17355) );
  OAI22_X2 U18075 ( .A1(n12756), .A2(n13450), .B1(n10317), .B2(n13447), .ZN(
        n17354) );
  NOR3_X4 U18076 ( .A1(n17356), .A2(n17355), .A3(n17354), .ZN(n17373) );
  NAND2_X2 U18077 ( .A1(n13198), .A2(REG_FILE_reg_out_14__18_), .ZN(n17360) );
  NAND2_X2 U18078 ( .A1(n13200), .A2(REG_FILE_reg_out_1__18_), .ZN(n17359) );
  NAND2_X2 U18079 ( .A1(n18502), .A2(REG_FILE_reg_out_11__18_), .ZN(n17358) );
  NAND2_X2 U18080 ( .A1(n13203), .A2(REG_FILE_reg_out_13__18_), .ZN(n17357) );
  NAND4_X2 U18081 ( .A1(n17360), .A2(n17359), .A3(n17358), .A4(n17357), .ZN(
        n17363) );
  OAI22_X2 U18082 ( .A1(n11098), .A2(n13470), .B1(n10497), .B2(n13468), .ZN(
        n17362) );
  OAI22_X2 U18083 ( .A1(n11276), .A2(n13474), .B1(n10496), .B2(n13473), .ZN(
        n17361) );
  NOR3_X4 U18084 ( .A1(n17363), .A2(n17362), .A3(n17361), .ZN(n17372) );
  NAND2_X2 U18085 ( .A1(n13456), .A2(REG_FILE_reg_out_12__18_), .ZN(n17367) );
  NAND2_X2 U18086 ( .A1(n13194), .A2(REG_FILE_reg_out_19__18_), .ZN(n17366) );
  NAND3_X4 U18087 ( .A1(n17367), .A2(n17366), .A3(n17365), .ZN(n17370) );
  OAI22_X2 U18088 ( .A1(n13461), .A2(n12894), .B1(n13458), .B2(n11863), .ZN(
        n17369) );
  OAI22_X2 U18089 ( .A1(n13465), .A2(n12807), .B1(n12405), .B2(n13463), .ZN(
        n17368) );
  NOR3_X4 U18090 ( .A1(n17370), .A2(n17369), .A3(n17368), .ZN(n17371) );
  NAND4_X2 U18091 ( .A1(n17374), .A2(n17373), .A3(n17372), .A4(n17371), .ZN(
        n17375) );
  INV_X4 U18092 ( .A(n17375), .ZN(n17380) );
  OAI222_X2 U18093 ( .A1(n17380), .A2(n13477), .B1(n12518), .B2(net231223), 
        .C1(n11045), .C2(n13206), .ZN(n7560) );
  NAND2_X2 U18094 ( .A1(n13412), .A2(ID_EXEC_OUT[178]), .ZN(n17379) );
  NAND2_X2 U18095 ( .A1(DMEM_BUS_OUT[50]), .A2(net231319), .ZN(n17378) );
  NAND2_X2 U18096 ( .A1(n13414), .A2(DMEM_BUS_OUT[18]), .ZN(n17377) );
  NAND2_X2 U18097 ( .A1(n13416), .A2(MEM_WB_OUT[55]), .ZN(n17376) );
  NAND4_X2 U18098 ( .A1(n17379), .A2(n17378), .A3(n17377), .A4(n17376), .ZN(
        n7561) );
  OAI22_X2 U18099 ( .A1(n11524), .A2(net231255), .B1(net230379), .B2(n17380), 
        .ZN(n7562) );
  OAI22_X2 U18100 ( .A1(n11104), .A2(net231255), .B1(net230379), .B2(n11917), 
        .ZN(n7564) );
  OAI22_X2 U18101 ( .A1(net231251), .A2(n11917), .B1(n12187), .B2(net230383), 
        .ZN(n7565) );
  OAI22_X2 U18102 ( .A1(n12187), .A2(net231255), .B1(n13481), .B2(n17381), 
        .ZN(n7566) );
  INV_X4 U18103 ( .A(n17382), .ZN(n17905) );
  NOR2_X4 U18104 ( .A1(n2109), .A2(n17383), .ZN(n17389) );
  NOR2_X4 U18105 ( .A1(n2106), .A2(n2108), .ZN(n17388) );
  OAI222_X2 U18106 ( .A1(n11864), .A2(n13373), .B1(n10232), .B2(n13371), .C1(
        n13368), .C2(n11703), .ZN(n17386) );
  OAI22_X2 U18107 ( .A1(n11865), .A2(n13383), .B1(n13380), .B2(n12757), .ZN(
        n17384) );
  NOR3_X4 U18108 ( .A1(n17386), .A2(n17385), .A3(n17384), .ZN(n17387) );
  NAND3_X2 U18109 ( .A1(n17389), .A2(n17388), .A3(n17387), .ZN(n17390) );
  MUX2_X2 U18110 ( .A(n17390), .B(ID_EXEC_OUT[51]), .S(net231293), .Z(n7567)
         );
  NAND2_X2 U18111 ( .A1(REG_FILE_reg_out_17__19_), .A2(n13435), .ZN(n17396) );
  OAI22_X2 U18112 ( .A1(n13420), .A2(n12808), .B1(n13418), .B2(n11864), .ZN(
        n17399) );
  OAI22_X2 U18113 ( .A1(n13440), .A2(n12588), .B1(n13438), .B2(n12573), .ZN(
        n17398) );
  NAND2_X2 U18114 ( .A1(n18493), .A2(REG_FILE_reg_out_6__19_), .ZN(n17404) );
  NAND2_X2 U18115 ( .A1(n13191), .A2(REG_FILE_reg_out_7__19_), .ZN(n17403) );
  NAND2_X2 U18116 ( .A1(n18494), .A2(REG_FILE_reg_out_4__19_), .ZN(n17402) );
  NAND2_X2 U18117 ( .A1(n13189), .A2(REG_FILE_reg_out_5__19_), .ZN(n17401) );
  NAND4_X2 U18118 ( .A1(n17404), .A2(n17403), .A3(n17402), .A4(n17401), .ZN(
        n17407) );
  OAI22_X2 U18119 ( .A1(n12293), .A2(n13445), .B1(n10930), .B2(n13443), .ZN(
        n17406) );
  OAI22_X2 U18120 ( .A1(n12757), .A2(n13450), .B1(n10318), .B2(n13447), .ZN(
        n17405) );
  NOR3_X4 U18121 ( .A1(n17407), .A2(n17406), .A3(n17405), .ZN(n17424) );
  NAND2_X2 U18122 ( .A1(n13198), .A2(REG_FILE_reg_out_14__19_), .ZN(n17411) );
  NAND2_X2 U18123 ( .A1(n13200), .A2(REG_FILE_reg_out_1__19_), .ZN(n17410) );
  NAND2_X2 U18124 ( .A1(n18502), .A2(REG_FILE_reg_out_11__19_), .ZN(n17409) );
  NAND2_X2 U18125 ( .A1(n13203), .A2(REG_FILE_reg_out_13__19_), .ZN(n17408) );
  NAND4_X2 U18126 ( .A1(n17411), .A2(n17410), .A3(n17409), .A4(n17408), .ZN(
        n17414) );
  OAI22_X2 U18127 ( .A1(n11099), .A2(n13471), .B1(n10499), .B2(n13468), .ZN(
        n17413) );
  OAI22_X2 U18128 ( .A1(n11277), .A2(n13475), .B1(n10498), .B2(n13473), .ZN(
        n17412) );
  NOR3_X4 U18129 ( .A1(n17414), .A2(n17413), .A3(n17412), .ZN(n17423) );
  NAND2_X2 U18130 ( .A1(n13456), .A2(REG_FILE_reg_out_12__19_), .ZN(n17418) );
  NAND2_X2 U18131 ( .A1(n13194), .A2(REG_FILE_reg_out_19__19_), .ZN(n17417) );
  NAND3_X4 U18132 ( .A1(n17418), .A2(n17417), .A3(n17416), .ZN(n17421) );
  OAI22_X2 U18133 ( .A1(n13461), .A2(n12896), .B1(n13458), .B2(n11865), .ZN(
        n17420) );
  OAI22_X2 U18134 ( .A1(n13465), .A2(n12809), .B1(n12406), .B2(n13463), .ZN(
        n17419) );
  NOR3_X4 U18135 ( .A1(n17421), .A2(n17420), .A3(n17419), .ZN(n17422) );
  NAND4_X2 U18136 ( .A1(n17425), .A2(n17424), .A3(n17423), .A4(n17422), .ZN(
        n17426) );
  INV_X4 U18137 ( .A(n17426), .ZN(n17431) );
  OAI222_X2 U18138 ( .A1(n17431), .A2(n13477), .B1(n12519), .B2(net231223), 
        .C1(n10806), .C2(n13206), .ZN(n7568) );
  NAND2_X2 U18139 ( .A1(n13412), .A2(ID_EXEC_OUT[179]), .ZN(n17430) );
  NAND2_X2 U18140 ( .A1(DMEM_BUS_OUT[51]), .A2(net231321), .ZN(n17429) );
  NAND2_X2 U18141 ( .A1(n13414), .A2(DMEM_BUS_OUT[19]), .ZN(n17428) );
  NAND2_X2 U18142 ( .A1(n13416), .A2(MEM_WB_OUT[56]), .ZN(n17427) );
  NAND4_X2 U18143 ( .A1(n17430), .A2(n17429), .A3(n17428), .A4(n17427), .ZN(
        n7569) );
  OAI22_X2 U18144 ( .A1(n11525), .A2(net231257), .B1(net230379), .B2(n17431), 
        .ZN(n7570) );
  OAI22_X2 U18145 ( .A1(n12190), .A2(net231255), .B1(n13481), .B2(n17432), 
        .ZN(n7574) );
  INV_X4 U18146 ( .A(net224493), .ZN(net224492) );
  XNOR2_X2 U18147 ( .A(net224492), .B(n10242), .ZN(n17434) );
  XNOR2_X2 U18148 ( .A(n17434), .B(n17433), .ZN(n17437) );
  NAND2_X2 U18149 ( .A1(net231615), .A2(n18911), .ZN(n17436) );
  NAND2_X2 U18150 ( .A1(EXEC_MEM_OUT_128), .A2(net231323), .ZN(n17435) );
  OAI211_X2 U18151 ( .C1(n17437), .C2(net231915), .A(n17436), .B(n17435), .ZN(
        n7575) );
  INV_X4 U18152 ( .A(n17546), .ZN(n17470) );
  NOR2_X4 U18153 ( .A1(n2089), .A2(n17438), .ZN(n17444) );
  NOR2_X4 U18154 ( .A1(n2086), .A2(n2088), .ZN(n17443) );
  OAI222_X2 U18155 ( .A1(n11867), .A2(n13374), .B1(n10233), .B2(n13370), .C1(
        n13367), .C2(n11706), .ZN(n17441) );
  OAI22_X2 U18156 ( .A1(n11868), .A2(n13383), .B1(n13380), .B2(n11866), .ZN(
        n17439) );
  NOR3_X4 U18157 ( .A1(n17441), .A2(n17440), .A3(n17439), .ZN(n17442) );
  NAND3_X2 U18158 ( .A1(n17444), .A2(n17443), .A3(n17442), .ZN(n17445) );
  MUX2_X2 U18159 ( .A(n17445), .B(ID_EXEC_OUT[52]), .S(net231293), .Z(n7576)
         );
  NAND2_X2 U18160 ( .A1(REG_FILE_reg_out_17__20_), .A2(n13435), .ZN(n17451) );
  OAI22_X2 U18161 ( .A1(n13419), .A2(n12810), .B1(n13418), .B2(n11867), .ZN(
        n17454) );
  OAI22_X2 U18162 ( .A1(n13440), .A2(n12589), .B1(n13438), .B2(n12574), .ZN(
        n17453) );
  NAND2_X2 U18163 ( .A1(n18493), .A2(REG_FILE_reg_out_6__20_), .ZN(n17459) );
  NAND2_X2 U18164 ( .A1(n13191), .A2(REG_FILE_reg_out_7__20_), .ZN(n17458) );
  NAND2_X2 U18165 ( .A1(n18494), .A2(REG_FILE_reg_out_4__20_), .ZN(n17457) );
  NAND2_X2 U18166 ( .A1(n13189), .A2(REG_FILE_reg_out_5__20_), .ZN(n17456) );
  NAND4_X2 U18167 ( .A1(n17459), .A2(n17458), .A3(n17457), .A4(n17456), .ZN(
        n17462) );
  OAI22_X2 U18168 ( .A1(n12294), .A2(n13445), .B1(n10931), .B2(n13443), .ZN(
        n17461) );
  OAI22_X2 U18169 ( .A1(n11866), .A2(n13450), .B1(n10319), .B2(n13447), .ZN(
        n17460) );
  NOR3_X4 U18170 ( .A1(n17462), .A2(n17461), .A3(n17460), .ZN(n17480) );
  NAND2_X2 U18171 ( .A1(n13198), .A2(REG_FILE_reg_out_14__20_), .ZN(n17466) );
  NAND2_X2 U18172 ( .A1(n13200), .A2(REG_FILE_reg_out_1__20_), .ZN(n17465) );
  NAND2_X2 U18173 ( .A1(n18502), .A2(REG_FILE_reg_out_11__20_), .ZN(n17464) );
  NAND2_X2 U18174 ( .A1(n13203), .A2(REG_FILE_reg_out_13__20_), .ZN(n17463) );
  NAND4_X2 U18175 ( .A1(n17466), .A2(n17465), .A3(n17464), .A4(n17463), .ZN(
        n17469) );
  OAI22_X2 U18176 ( .A1(n11100), .A2(n13470), .B1(n10501), .B2(n13468), .ZN(
        n17468) );
  OAI22_X2 U18177 ( .A1(n11278), .A2(n13474), .B1(n10500), .B2(n13473), .ZN(
        n17467) );
  NOR3_X4 U18178 ( .A1(n17469), .A2(n17468), .A3(n17467), .ZN(n17479) );
  NAND2_X2 U18179 ( .A1(n13456), .A2(REG_FILE_reg_out_12__20_), .ZN(n17474) );
  NAND2_X2 U18180 ( .A1(n13194), .A2(REG_FILE_reg_out_19__20_), .ZN(n17473) );
  OAI22_X2 U18181 ( .A1(n13461), .A2(n12898), .B1(n13458), .B2(n11868), .ZN(
        n17476) );
  OAI22_X2 U18182 ( .A1(n13465), .A2(n12811), .B1(n12407), .B2(n13463), .ZN(
        n17475) );
  NOR3_X4 U18183 ( .A1(n17477), .A2(n17476), .A3(n17475), .ZN(n17478) );
  NAND4_X2 U18184 ( .A1(n17481), .A2(n17480), .A3(n17479), .A4(n17478), .ZN(
        n17482) );
  INV_X4 U18185 ( .A(n17482), .ZN(n17487) );
  OAI222_X2 U18186 ( .A1(n17487), .A2(n13477), .B1(n12520), .B2(net231223), 
        .C1(n12021), .C2(n13206), .ZN(n7577) );
  NAND2_X2 U18187 ( .A1(n13412), .A2(ID_EXEC_OUT[180]), .ZN(n17486) );
  NAND2_X2 U18188 ( .A1(DMEM_BUS_OUT[52]), .A2(net231319), .ZN(n17485) );
  NAND2_X2 U18189 ( .A1(n13414), .A2(DMEM_BUS_OUT[20]), .ZN(n17484) );
  NAND2_X2 U18190 ( .A1(n13416), .A2(MEM_WB_OUT[57]), .ZN(n17483) );
  NAND4_X2 U18191 ( .A1(n17486), .A2(n17485), .A3(n17484), .A4(n17483), .ZN(
        n7578) );
  OAI22_X2 U18192 ( .A1(n11526), .A2(net231257), .B1(net230379), .B2(n17487), 
        .ZN(n7579) );
  OAI22_X2 U18193 ( .A1(n19326), .A2(net231257), .B1(n13480), .B2(n17488), 
        .ZN(n7583) );
  XNOR2_X2 U18194 ( .A(net224402), .B(net233124), .ZN(n17491) );
  NAND2_X2 U18195 ( .A1(net231615), .A2(n17505), .ZN(n17490) );
  NAND2_X2 U18196 ( .A1(EXEC_MEM_OUT_129), .A2(net231323), .ZN(n17489) );
  OAI211_X2 U18197 ( .C1(n17491), .C2(net231915), .A(n17490), .B(n17489), .ZN(
        n7584) );
  INV_X4 U18198 ( .A(n18279), .ZN(n17494) );
  INV_X4 U18199 ( .A(n18362), .ZN(n17497) );
  OAI21_X4 U18200 ( .B1(n17497), .B2(n18361), .A(n17496), .ZN(n18322) );
  INV_X4 U18201 ( .A(n17498), .ZN(n18324) );
  INV_X4 U18202 ( .A(n17895), .ZN(n17500) );
  XNOR2_X2 U18203 ( .A(n17504), .B(n17503), .ZN(n17507) );
  XNOR2_X2 U18204 ( .A(n18991), .B(n17505), .ZN(n18990) );
  NAND2_X2 U18205 ( .A1(net232816), .A2(n18867), .ZN(n17514) );
  INV_X4 U18206 ( .A(n17509), .ZN(n17512) );
  INV_X4 U18207 ( .A(n17510), .ZN(n17511) );
  NOR2_X4 U18208 ( .A1(n17512), .A2(n17511), .ZN(n17513) );
  NAND2_X2 U18209 ( .A1(n13390), .A2(n18338), .ZN(n17523) );
  NAND2_X2 U18210 ( .A1(net232816), .A2(n18873), .ZN(n17519) );
  INV_X4 U18211 ( .A(n17515), .ZN(n17516) );
  NAND2_X2 U18212 ( .A1(n13397), .A2(n18296), .ZN(n17522) );
  NAND2_X2 U18214 ( .A1(n13393), .A2(n17909), .ZN(n17520) );
  NAND4_X2 U18215 ( .A1(n17523), .A2(n17522), .A3(n17521), .A4(n17520), .ZN(
        n17524) );
  INV_X4 U18216 ( .A(n17524), .ZN(n17702) );
  NAND2_X2 U18217 ( .A1(n13397), .A2(n17994), .ZN(n17534) );
  INV_X4 U18218 ( .A(n17525), .ZN(n17528) );
  NOR2_X4 U18219 ( .A1(n17526), .A2(net232817), .ZN(n17527) );
  NOR2_X4 U18220 ( .A1(n17528), .A2(n17527), .ZN(n17529) );
  NAND2_X2 U18221 ( .A1(n13390), .A2(n18328), .ZN(n17533) );
  NAND2_X2 U18222 ( .A1(n16300), .A2(n17697), .ZN(n17532) );
  NAND2_X2 U18223 ( .A1(n13393), .A2(n17587), .ZN(n17531) );
  NAND4_X2 U18224 ( .A1(n17534), .A2(n17533), .A3(n17532), .A4(n17531), .ZN(
        n17923) );
  INV_X4 U18225 ( .A(n17923), .ZN(n17535) );
  OAI22_X2 U18226 ( .A1(n17702), .A2(n18003), .B1(n17535), .B2(n18008), .ZN(
        n17552) );
  NAND2_X2 U18227 ( .A1(n13397), .A2(n17686), .ZN(n17536) );
  INV_X4 U18228 ( .A(n17907), .ZN(n17543) );
  MUX2_X2 U18229 ( .A(n13041), .B(n18966), .S(n19100), .Z(n18308) );
  INV_X4 U18230 ( .A(n18308), .ZN(n17541) );
  NAND2_X2 U18231 ( .A1(n13390), .A2(n17916), .ZN(n17539) );
  NAND2_X2 U18232 ( .A1(n13397), .A2(n17918), .ZN(n17538) );
  INV_X4 U18233 ( .A(n17542), .ZN(n17682) );
  OAI22_X2 U18234 ( .A1(n17543), .A2(n13214), .B1(n17682), .B2(n13207), .ZN(
        n17551) );
  NAND2_X2 U18235 ( .A1(n18566), .A2(DMEM_BUS_OUT[20]), .ZN(n17548) );
  INV_X4 U18236 ( .A(n18991), .ZN(n17547) );
  AOI211_X4 U18237 ( .C1(n18651), .C2(n17552), .A(n17551), .B(n17550), .ZN(
        n17553) );
  NAND3_X4 U18238 ( .A1(n17555), .A2(n17554), .A3(n17553), .ZN(n7586) );
  NAND2_X2 U18239 ( .A1(n13409), .A2(n18872), .ZN(n17556) );
  OAI211_X2 U18240 ( .C1(n12149), .C2(net231227), .A(n17556), .B(n6779), .ZN(
        n7590) );
  NAND2_X2 U18241 ( .A1(n17558), .A2(n17557), .ZN(n17559) );
  XNOR2_X2 U18242 ( .A(n17559), .B(n17560), .ZN(n17582) );
  XNOR2_X2 U18243 ( .A(n18877), .B(n18872), .ZN(n19048) );
  INV_X4 U18244 ( .A(n17561), .ZN(n17564) );
  OAI221_X2 U18245 ( .B1(n19048), .B2(n13491), .C1(n17564), .C2(n13214), .A(
        n17563), .ZN(n17580) );
  INV_X4 U18246 ( .A(n17565), .ZN(n17573) );
  INV_X4 U18247 ( .A(n17566), .ZN(n17567) );
  NAND2_X2 U18248 ( .A1(n17567), .A2(n13208), .ZN(n17569) );
  NAND2_X2 U18249 ( .A1(n18566), .A2(DMEM_BUS_OUT[3]), .ZN(n17568) );
  OAI211_X2 U18250 ( .C1(n17570), .C2(n18569), .A(n17569), .B(n17568), .ZN(
        n17571) );
  NAND2_X2 U18251 ( .A1(n17571), .A2(n18877), .ZN(n17572) );
  NOR2_X4 U18252 ( .A1(n17574), .A2(n13211), .ZN(n17578) );
  INV_X4 U18253 ( .A(n17575), .ZN(n17576) );
  NOR4_X2 U18254 ( .A1(n17580), .A2(n17579), .A3(n17578), .A4(n17577), .ZN(
        n17581) );
  NAND2_X2 U18255 ( .A1(n13409), .A2(net222497), .ZN(n17583) );
  OAI211_X2 U18256 ( .C1(n12159), .C2(net231227), .A(n17583), .B(n6768), .ZN(
        n7596) );
  NAND2_X2 U18257 ( .A1(n17584), .A2(n16059), .ZN(n17590) );
  NAND2_X2 U18258 ( .A1(n13488), .A2(n17585), .ZN(n17589) );
  AOI22_X2 U18259 ( .A1(n13388), .A2(n17587), .B1(n13397), .B2(n17586), .ZN(
        n17588) );
  NAND2_X2 U18260 ( .A1(n17924), .A2(n17742), .ZN(n17621) );
  XNOR2_X2 U18261 ( .A(n17593), .B(n17592), .ZN(n17594) );
  NAND2_X2 U18262 ( .A1(n13492), .A2(n17594), .ZN(n17620) );
  NAND2_X2 U18263 ( .A1(n13488), .A2(n17595), .ZN(n17602) );
  NAND2_X2 U18264 ( .A1(n13393), .A2(n17596), .ZN(n17601) );
  NAND2_X2 U18265 ( .A1(n13390), .A2(n17597), .ZN(n17600) );
  NAND2_X2 U18266 ( .A1(n13397), .A2(n17598), .ZN(n17599) );
  NAND4_X2 U18267 ( .A1(n17602), .A2(n17601), .A3(n17600), .A4(n17599), .ZN(
        n17743) );
  INV_X4 U18268 ( .A(n17743), .ZN(n17603) );
  NOR2_X4 U18269 ( .A1(n17603), .A2(n13207), .ZN(n17613) );
  INV_X4 U18270 ( .A(n17604), .ZN(n17605) );
  NAND2_X2 U18271 ( .A1(n17605), .A2(n13208), .ZN(n17607) );
  NAND2_X2 U18272 ( .A1(n18566), .A2(DMEM_BUS_OUT[13]), .ZN(n17606) );
  OAI211_X2 U18273 ( .C1(n17608), .C2(n18569), .A(n17607), .B(n17606), .ZN(
        n17609) );
  NAND2_X2 U18274 ( .A1(n17609), .A2(n18907), .ZN(n17610) );
  OAI21_X4 U18275 ( .B1(n17611), .B2(n13215), .A(n17610), .ZN(n17612) );
  NOR2_X4 U18276 ( .A1(n17613), .A2(n17612), .ZN(n17619) );
  NAND2_X2 U18277 ( .A1(DMEM_BUS_OUT[13]), .A2(net231323), .ZN(n17614) );
  XNOR2_X2 U18278 ( .A(n18907), .B(net222497), .ZN(n18917) );
  NAND4_X2 U18279 ( .A1(n17621), .A2(n17620), .A3(n17619), .A4(n17618), .ZN(
        n7598) );
  INV_X4 U18280 ( .A(n17622), .ZN(n17681) );
  NOR2_X4 U18281 ( .A1(n2069), .A2(n17623), .ZN(n17629) );
  NOR2_X4 U18282 ( .A1(n2066), .A2(n2068), .ZN(n17628) );
  OAI222_X2 U18283 ( .A1(n11870), .A2(n13373), .B1(n10234), .B2(n13371), .C1(
        n13368), .C2(n11709), .ZN(n17626) );
  OAI22_X2 U18284 ( .A1(n11871), .A2(n13382), .B1(n13380), .B2(n11869), .ZN(
        n17624) );
  NOR3_X4 U18285 ( .A1(n17626), .A2(n17625), .A3(n17624), .ZN(n17627) );
  NAND3_X2 U18286 ( .A1(n17629), .A2(n17628), .A3(n17627), .ZN(n17630) );
  MUX2_X2 U18287 ( .A(n17630), .B(ID_EXEC_OUT[53]), .S(net231293), .Z(n7599)
         );
  NAND2_X2 U18288 ( .A1(REG_FILE_reg_out_17__21_), .A2(n13434), .ZN(n17636) );
  OAI22_X2 U18289 ( .A1(n13420), .A2(n12812), .B1(n13418), .B2(n11870), .ZN(
        n17639) );
  OAI22_X2 U18290 ( .A1(n13440), .A2(n12590), .B1(n13438), .B2(n12575), .ZN(
        n17638) );
  NAND2_X2 U18291 ( .A1(n18493), .A2(REG_FILE_reg_out_6__21_), .ZN(n17644) );
  NAND2_X2 U18292 ( .A1(n13191), .A2(REG_FILE_reg_out_7__21_), .ZN(n17643) );
  NAND2_X2 U18293 ( .A1(n18494), .A2(REG_FILE_reg_out_4__21_), .ZN(n17642) );
  NAND2_X2 U18294 ( .A1(n13189), .A2(REG_FILE_reg_out_5__21_), .ZN(n17641) );
  NAND4_X2 U18295 ( .A1(n17644), .A2(n17643), .A3(n17642), .A4(n17641), .ZN(
        n17647) );
  OAI22_X2 U18296 ( .A1(n12295), .A2(n13445), .B1(n10932), .B2(n13443), .ZN(
        n17646) );
  OAI22_X2 U18297 ( .A1(n11869), .A2(n13450), .B1(n10320), .B2(n13447), .ZN(
        n17645) );
  NAND2_X2 U18298 ( .A1(n13198), .A2(REG_FILE_reg_out_14__21_), .ZN(n17651) );
  NAND2_X2 U18299 ( .A1(n13200), .A2(REG_FILE_reg_out_1__21_), .ZN(n17650) );
  NAND2_X2 U18300 ( .A1(n18502), .A2(REG_FILE_reg_out_11__21_), .ZN(n17649) );
  NAND2_X2 U18301 ( .A1(n13203), .A2(REG_FILE_reg_out_13__21_), .ZN(n17648) );
  NAND4_X2 U18302 ( .A1(n17651), .A2(n17650), .A3(n17649), .A4(n17648), .ZN(
        n17654) );
  OAI22_X2 U18303 ( .A1(n11101), .A2(n13471), .B1(n10503), .B2(n13468), .ZN(
        n17653) );
  OAI22_X2 U18304 ( .A1(n11279), .A2(n13475), .B1(n10502), .B2(n13473), .ZN(
        n17652) );
  NAND2_X2 U18305 ( .A1(n13455), .A2(REG_FILE_reg_out_12__21_), .ZN(n17658) );
  NAND2_X2 U18306 ( .A1(n13194), .A2(REG_FILE_reg_out_19__21_), .ZN(n17657) );
  OAI22_X2 U18307 ( .A1(n13461), .A2(n12900), .B1(n13458), .B2(n11871), .ZN(
        n17660) );
  OAI22_X2 U18308 ( .A1(n13465), .A2(n12813), .B1(n12408), .B2(n13463), .ZN(
        n17659) );
  NAND4_X2 U18309 ( .A1(n17665), .A2(n17664), .A3(n17663), .A4(n17662), .ZN(
        n17666) );
  INV_X4 U18310 ( .A(n17666), .ZN(n17671) );
  OAI222_X2 U18311 ( .A1(n17671), .A2(n13477), .B1(n12521), .B2(net231223), 
        .C1(n11983), .C2(n13206), .ZN(n7600) );
  NAND2_X2 U18312 ( .A1(n13411), .A2(ID_EXEC_OUT[181]), .ZN(n17670) );
  NAND2_X2 U18313 ( .A1(DMEM_BUS_OUT[53]), .A2(net231319), .ZN(n17669) );
  NAND2_X2 U18314 ( .A1(n13413), .A2(DMEM_BUS_OUT[21]), .ZN(n17668) );
  NAND2_X2 U18315 ( .A1(n13416), .A2(MEM_WB_OUT[58]), .ZN(n17667) );
  NAND4_X2 U18316 ( .A1(n17670), .A2(n17669), .A3(n17668), .A4(n17667), .ZN(
        n7601) );
  OAI22_X2 U18317 ( .A1(n11527), .A2(net231257), .B1(net230379), .B2(n17671), 
        .ZN(n7602) );
  OAI22_X2 U18318 ( .A1(n11105), .A2(net231257), .B1(net230377), .B2(n11918), 
        .ZN(n7604) );
  OAI22_X2 U18319 ( .A1(net231249), .A2(n11918), .B1(n19325), .B2(net230381), 
        .ZN(n7605) );
  OAI22_X2 U18320 ( .A1(n19325), .A2(net231257), .B1(n13481), .B2(n17672), 
        .ZN(n7606) );
  XNOR2_X2 U18321 ( .A(net224170), .B(net224171), .ZN(n17678) );
  NAND2_X2 U18322 ( .A1(net231615), .A2(n17712), .ZN(n17677) );
  NAND2_X2 U18323 ( .A1(EXEC_MEM_OUT_130), .A2(net231323), .ZN(n17676) );
  OAI211_X2 U18324 ( .C1(n17678), .C2(net231915), .A(n17677), .B(n17676), .ZN(
        n7607) );
  NAND2_X2 U18325 ( .A1(n18566), .A2(DMEM_BUS_OUT[21]), .ZN(n17679) );
  OAI221_X2 U18326 ( .B1(n17681), .B2(n18569), .C1(n13209), .C2(n17680), .A(
        n17679), .ZN(n17692) );
  NOR2_X4 U18327 ( .A1(n17682), .A2(n13215), .ZN(n17691) );
  NAND2_X2 U18328 ( .A1(n17683), .A2(n19100), .ZN(n17684) );
  INV_X4 U18329 ( .A(n17684), .ZN(n18347) );
  AOI22_X2 U18330 ( .A1(n10843), .A2(n13149), .B1(n18347), .B2(n18345), .ZN(
        n17688) );
  AOI22_X2 U18331 ( .A1(n18310), .A2(n13163), .B1(n13388), .B2(n17686), .ZN(
        n17687) );
  NAND2_X2 U18332 ( .A1(n17688), .A2(n17687), .ZN(n17859) );
  INV_X4 U18333 ( .A(n17859), .ZN(n17689) );
  NAND2_X2 U18334 ( .A1(n13397), .A2(n18328), .ZN(n17701) );
  INV_X4 U18335 ( .A(n17693), .ZN(n17694) );
  NAND2_X2 U18336 ( .A1(n13390), .A2(n18329), .ZN(n17700) );
  NAND2_X2 U18337 ( .A1(n13393), .A2(n17697), .ZN(n17699) );
  NAND2_X2 U18338 ( .A1(n13488), .A2(n17994), .ZN(n17698) );
  NAND4_X2 U18339 ( .A1(n17701), .A2(n17700), .A3(n17699), .A4(n17698), .ZN(
        n17833) );
  INV_X4 U18340 ( .A(n17833), .ZN(n17703) );
  OAI22_X2 U18341 ( .A1(n18003), .A2(n17703), .B1(n17702), .B2(n18008), .ZN(
        n17704) );
  NAND2_X2 U18342 ( .A1(n18651), .A2(n17704), .ZN(n17717) );
  AOI22_X2 U18343 ( .A1(DMEM_BUS_OUT[21]), .A2(net231307), .B1(
        ID_EXEC_OUT[225]), .B2(n13216), .ZN(n17716) );
  XNOR2_X2 U18344 ( .A(n17710), .B(n17711), .ZN(n17714) );
  XNOR2_X2 U18345 ( .A(n18985), .B(n17712), .ZN(n18989) );
  NAND4_X2 U18346 ( .A1(n17715), .A2(n17717), .A3(n17716), .A4(n17718), .ZN(
        n7609) );
  NAND2_X2 U18347 ( .A1(n13409), .A2(n18897), .ZN(n17719) );
  OAI211_X2 U18348 ( .C1(n12160), .C2(net231227), .A(n17719), .B(n6766), .ZN(
        n7613) );
  MUX2_X2 U18349 ( .A(DMEM_BUS_OUT[14]), .B(MEM_WB_OUT[51]), .S(net231293), 
        .Z(n7614) );
  INV_X4 U18350 ( .A(n17723), .ZN(n17724) );
  NAND3_X2 U18351 ( .A1(n17726), .A2(n17725), .A3(n17724), .ZN(n17727) );
  INV_X4 U18352 ( .A(n17727), .ZN(n17730) );
  INV_X4 U18353 ( .A(n17731), .ZN(n17883) );
  XNOR2_X2 U18354 ( .A(n17735), .B(n17734), .ZN(n17736) );
  NAND2_X2 U18355 ( .A1(n13492), .A2(n17736), .ZN(n17767) );
  NAND2_X2 U18356 ( .A1(n17982), .A2(n17737), .ZN(n17740) );
  NAND2_X2 U18357 ( .A1(n17983), .A2(ID_EXEC_OUT[46]), .ZN(n17739) );
  NAND2_X2 U18358 ( .A1(n18566), .A2(DMEM_BUS_OUT[14]), .ZN(n17738) );
  NAND3_X2 U18359 ( .A1(n17740), .A2(n17739), .A3(n17738), .ZN(n17741) );
  NAND2_X2 U18360 ( .A1(n17741), .A2(n18896), .ZN(n17766) );
  INV_X4 U18361 ( .A(n17742), .ZN(n17745) );
  NAND2_X2 U18362 ( .A1(n10199), .A2(n17743), .ZN(n17744) );
  OAI21_X4 U18363 ( .B1(n17745), .B2(n18008), .A(n17744), .ZN(n17761) );
  NAND2_X2 U18364 ( .A1(n16061), .A2(n17910), .ZN(n17751) );
  NAND2_X2 U18365 ( .A1(n13390), .A2(n17909), .ZN(n17750) );
  NAND2_X2 U18366 ( .A1(n13393), .A2(n17746), .ZN(n17749) );
  NAND2_X2 U18367 ( .A1(n16300), .A2(n17747), .ZN(n17748) );
  NAND4_X2 U18368 ( .A1(n17749), .A2(n17750), .A3(n17751), .A4(n17748), .ZN(
        n17752) );
  INV_X4 U18369 ( .A(n17752), .ZN(n17873) );
  NAND2_X2 U18370 ( .A1(n16300), .A2(n17917), .ZN(n17758) );
  NAND2_X2 U18371 ( .A1(n13393), .A2(n17916), .ZN(n17757) );
  NAND2_X2 U18372 ( .A1(n13390), .A2(n17753), .ZN(n17756) );
  NAND4_X2 U18373 ( .A1(n17758), .A2(n17757), .A3(n17756), .A4(n17755), .ZN(
        n17885) );
  NAND2_X2 U18374 ( .A1(n19124), .A2(n17885), .ZN(n17759) );
  OAI21_X4 U18375 ( .B1(n17761), .B2(n17760), .A(n18651), .ZN(n17765) );
  XNOR2_X2 U18376 ( .A(n18896), .B(n18897), .ZN(n18903) );
  INV_X4 U18377 ( .A(n18903), .ZN(n18852) );
  NAND4_X2 U18378 ( .A1(n17767), .A2(n17766), .A3(n17765), .A4(n17764), .ZN(
        n7615) );
  INV_X4 U18379 ( .A(n17840), .ZN(n17808) );
  NOR2_X4 U18380 ( .A1(n2049), .A2(n17770), .ZN(n17782) );
  NOR2_X4 U18381 ( .A1(n2046), .A2(n2048), .ZN(n17781) );
  OAI222_X2 U18382 ( .A1(n12213), .A2(n13374), .B1(n10324), .B2(n13370), .C1(
        n13367), .C2(n11712), .ZN(n17779) );
  OAI22_X2 U18383 ( .A1(n11872), .A2(n13383), .B1(n13380), .B2(n12250), .ZN(
        n17777) );
  NOR3_X4 U18384 ( .A1(n17779), .A2(n17778), .A3(n17777), .ZN(n17780) );
  NAND3_X2 U18385 ( .A1(n17782), .A2(n17781), .A3(n17780), .ZN(n17783) );
  MUX2_X2 U18386 ( .A(n17783), .B(ID_EXEC_OUT[54]), .S(net231293), .Z(n7616)
         );
  NAND2_X2 U18387 ( .A1(REG_FILE_reg_out_17__22_), .A2(n13434), .ZN(n17789) );
  OAI22_X2 U18388 ( .A1(n13420), .A2(n12814), .B1(n13417), .B2(n12213), .ZN(
        n17792) );
  OAI22_X2 U18389 ( .A1(n13440), .A2(n12591), .B1(n13438), .B2(n12576), .ZN(
        n17791) );
  NAND2_X2 U18390 ( .A1(n18493), .A2(REG_FILE_reg_out_6__22_), .ZN(n17797) );
  NAND2_X2 U18391 ( .A1(n13191), .A2(REG_FILE_reg_out_7__22_), .ZN(n17796) );
  NAND2_X2 U18392 ( .A1(n18494), .A2(REG_FILE_reg_out_4__22_), .ZN(n17795) );
  NAND2_X2 U18393 ( .A1(n13189), .A2(REG_FILE_reg_out_5__22_), .ZN(n17794) );
  NAND4_X2 U18394 ( .A1(n17797), .A2(n17796), .A3(n17795), .A4(n17794), .ZN(
        n17800) );
  OAI22_X2 U18395 ( .A1(n11421), .A2(n13445), .B1(n10521), .B2(n13442), .ZN(
        n17799) );
  OAI22_X2 U18396 ( .A1(n12250), .A2(n13451), .B1(n10321), .B2(n13448), .ZN(
        n17798) );
  NAND2_X2 U18397 ( .A1(n13198), .A2(REG_FILE_reg_out_14__22_), .ZN(n17804) );
  NAND2_X2 U18398 ( .A1(n13200), .A2(REG_FILE_reg_out_1__22_), .ZN(n17803) );
  NAND2_X2 U18399 ( .A1(n18502), .A2(REG_FILE_reg_out_11__22_), .ZN(n17802) );
  NAND2_X2 U18400 ( .A1(n13203), .A2(REG_FILE_reg_out_13__22_), .ZN(n17801) );
  NAND4_X2 U18401 ( .A1(n17804), .A2(n17803), .A3(n17802), .A4(n17801), .ZN(
        n17807) );
  OAI22_X2 U18402 ( .A1(n12138), .A2(n13471), .B1(n10292), .B2(n13467), .ZN(
        n17806) );
  OAI22_X2 U18403 ( .A1(n12262), .A2(n13475), .B1(n10918), .B2(n13472), .ZN(
        n17805) );
  NAND2_X2 U18404 ( .A1(n13455), .A2(REG_FILE_reg_out_12__22_), .ZN(n17812) );
  NAND2_X2 U18405 ( .A1(n13194), .A2(REG_FILE_reg_out_19__22_), .ZN(n17811) );
  OAI22_X2 U18406 ( .A1(n13461), .A2(n12902), .B1(n13458), .B2(n11872), .ZN(
        n17814) );
  OAI22_X2 U18407 ( .A1(n18721), .A2(n12815), .B1(n12409), .B2(n13463), .ZN(
        n17813) );
  NAND4_X2 U18408 ( .A1(n17819), .A2(n17818), .A3(n17817), .A4(n17816), .ZN(
        n17820) );
  INV_X4 U18409 ( .A(n17820), .ZN(n17825) );
  OAI222_X2 U18410 ( .A1(n17825), .A2(n13477), .B1(n11478), .B2(net231223), 
        .C1(n18794), .C2(n13206), .ZN(n7617) );
  NAND2_X2 U18411 ( .A1(n13411), .A2(ID_EXEC_OUT[182]), .ZN(n17824) );
  NAND2_X2 U18412 ( .A1(DMEM_BUS_OUT[54]), .A2(net231319), .ZN(n17823) );
  NAND2_X2 U18413 ( .A1(n13413), .A2(DMEM_BUS_OUT[22]), .ZN(n17822) );
  NAND2_X2 U18414 ( .A1(n13416), .A2(MEM_WB_OUT[59]), .ZN(n17821) );
  NAND4_X2 U18415 ( .A1(n17824), .A2(n17823), .A3(n17822), .A4(n17821), .ZN(
        n7618) );
  OAI22_X2 U18416 ( .A1(n11528), .A2(net231257), .B1(net230377), .B2(n17825), 
        .ZN(n7619) );
  OAI22_X2 U18417 ( .A1(n19324), .A2(net231257), .B1(n13480), .B2(n17826), 
        .ZN(n7623) );
  NAND2_X2 U18418 ( .A1(n17828), .A2(n17827), .ZN(n17829) );
  XNOR2_X2 U18419 ( .A(n17830), .B(n17829), .ZN(n17832) );
  NAND2_X2 U18420 ( .A1(net231615), .A2(n18980), .ZN(n17831) );
  OAI221_X2 U18421 ( .B1(net231227), .B2(n11475), .C1(net231915), .C2(n17832), 
        .A(n17831), .ZN(n7624) );
  NAND2_X2 U18422 ( .A1(n19118), .A2(n17833), .ZN(n17866) );
  NAND2_X2 U18423 ( .A1(n17982), .A2(n17840), .ZN(n17841) );
  OAI221_X2 U18424 ( .B1(n13209), .B2(n17842), .C1(n11982), .C2(n17870), .A(
        n17841), .ZN(n17858) );
  NAND2_X2 U18425 ( .A1(n16300), .A2(n18296), .ZN(n17852) );
  NAND2_X2 U18426 ( .A1(net232816), .A2(n19038), .ZN(n17848) );
  INV_X4 U18427 ( .A(n17843), .ZN(n17846) );
  INV_X4 U18428 ( .A(n17844), .ZN(n17845) );
  NOR2_X4 U18429 ( .A1(n17846), .A2(n17845), .ZN(n17847) );
  NAND3_X4 U18430 ( .A1(n17848), .A2(n17993), .A3(n17847), .ZN(n18339) );
  NAND2_X2 U18431 ( .A1(n15733), .A2(n18339), .ZN(n17851) );
  NAND2_X2 U18433 ( .A1(n16061), .A2(n18338), .ZN(n17849) );
  NAND4_X2 U18434 ( .A1(n17852), .A2(n17851), .A3(n17850), .A4(n17849), .ZN(
        n18005) );
  AOI22_X2 U18435 ( .A1(n18310), .A2(n13161), .B1(n13388), .B2(n17918), .ZN(
        n17853) );
  NAND2_X2 U18436 ( .A1(n17854), .A2(n17853), .ZN(n18006) );
  INV_X4 U18437 ( .A(n18006), .ZN(n17855) );
  NOR2_X4 U18438 ( .A1(n17689), .A2(n13214), .ZN(n17862) );
  OAI22_X2 U18439 ( .A1(net231251), .A2(n11982), .B1(n13217), .B2(n10818), 
        .ZN(n17861) );
  NAND4_X2 U18440 ( .A1(n17865), .A2(n17866), .A3(n17864), .A4(n17863), .ZN(
        n7626) );
  OAI211_X2 U18441 ( .C1(n12161), .C2(net231227), .A(n17867), .B(n6765), .ZN(
        n7630) );
  OAI221_X2 U18442 ( .B1(n13209), .B2(n17871), .C1(n12130), .C2(n17870), .A(
        n17869), .ZN(n17877) );
  INV_X4 U18443 ( .A(n17872), .ZN(n17875) );
  AOI22_X2 U18444 ( .A1(n17877), .A2(n13141), .B1(n17876), .B2(n18651), .ZN(
        n17891) );
  INV_X4 U18445 ( .A(n17878), .ZN(n17879) );
  NOR2_X4 U18446 ( .A1(n17879), .A2(n13211), .ZN(n17882) );
  OAI22_X2 U18447 ( .A1(net231251), .A2(n12130), .B1(n13217), .B2(n10822), 
        .ZN(n17881) );
  XNOR2_X2 U18448 ( .A(n18882), .B(n19091), .ZN(n18891) );
  NOR3_X4 U18449 ( .A1(n17882), .A2(n17881), .A3(n17880), .ZN(n17890) );
  XNOR2_X2 U18450 ( .A(n17883), .B(n17884), .ZN(n17888) );
  INV_X4 U18451 ( .A(n17885), .ZN(n17886) );
  NOR2_X4 U18452 ( .A1(n17886), .A2(n13214), .ZN(n17887) );
  XNOR2_X2 U18453 ( .A(n18914), .B(n18911), .ZN(n18879) );
  INV_X4 U18454 ( .A(n17897), .ZN(n17898) );
  XNOR2_X2 U18455 ( .A(n17902), .B(n17901), .ZN(n17932) );
  NAND2_X2 U18456 ( .A1(n18566), .A2(DMEM_BUS_OUT[19]), .ZN(n17903) );
  OAI221_X2 U18457 ( .B1(n17905), .B2(n18569), .C1(n13209), .C2(n17904), .A(
        n17903), .ZN(n17906) );
  NAND2_X2 U18458 ( .A1(n17906), .A2(n18914), .ZN(n17927) );
  NAND2_X2 U18459 ( .A1(n17908), .A2(n17907), .ZN(n17926) );
  INV_X4 U18460 ( .A(n13211), .ZN(n17924) );
  NAND2_X2 U18461 ( .A1(n16300), .A2(n17909), .ZN(n17915) );
  NAND2_X2 U18462 ( .A1(n13390), .A2(n18296), .ZN(n17914) );
  NAND2_X2 U18463 ( .A1(n13393), .A2(n17910), .ZN(n17913) );
  NAND2_X2 U18465 ( .A1(n16061), .A2(n17916), .ZN(n17922) );
  NAND2_X2 U18466 ( .A1(n15733), .A2(n17917), .ZN(n17920) );
  NAND2_X2 U18467 ( .A1(n16300), .A2(n17918), .ZN(n17919) );
  NAND4_X2 U18468 ( .A1(n17922), .A2(n17921), .A3(n17920), .A4(n17919), .ZN(
        n18577) );
  NAND2_X2 U18469 ( .A1(ID_EXEC_OUT[223]), .A2(n13216), .ZN(n17928) );
  NOR2_X4 U18470 ( .A1(n17930), .A2(n17929), .ZN(n17931) );
  OAI221_X2 U18471 ( .B1(n18879), .B2(n13491), .C1(n17932), .C2(n18550), .A(
        n17931), .ZN(n7634) );
  NAND2_X2 U18472 ( .A1(REG_FILE_reg_out_17__23_), .A2(n13434), .ZN(n17938) );
  OAI22_X2 U18473 ( .A1(n13420), .A2(n12816), .B1(n13417), .B2(n11873), .ZN(
        n17941) );
  OAI22_X2 U18474 ( .A1(n13440), .A2(n12592), .B1(n13438), .B2(n12577), .ZN(
        n17940) );
  NOR3_X4 U18475 ( .A1(n17942), .A2(n17941), .A3(n17940), .ZN(n17968) );
  NAND2_X2 U18476 ( .A1(n18493), .A2(REG_FILE_reg_out_6__23_), .ZN(n17946) );
  NAND2_X2 U18477 ( .A1(n13191), .A2(REG_FILE_reg_out_7__23_), .ZN(n17945) );
  NAND2_X2 U18478 ( .A1(n18494), .A2(REG_FILE_reg_out_4__23_), .ZN(n17944) );
  NAND2_X2 U18479 ( .A1(n13189), .A2(REG_FILE_reg_out_5__23_), .ZN(n17943) );
  NAND4_X2 U18480 ( .A1(n17946), .A2(n17945), .A3(n17944), .A4(n17943), .ZN(
        n17949) );
  OAI22_X2 U18481 ( .A1(n11422), .A2(n13444), .B1(n10522), .B2(n13443), .ZN(
        n17948) );
  OAI22_X2 U18482 ( .A1(n12777), .A2(n13451), .B1(n12042), .B2(n13448), .ZN(
        n17947) );
  NAND2_X2 U18483 ( .A1(n13198), .A2(REG_FILE_reg_out_14__23_), .ZN(n17953) );
  NAND2_X2 U18484 ( .A1(n13200), .A2(REG_FILE_reg_out_1__23_), .ZN(n17952) );
  NAND2_X2 U18485 ( .A1(n18502), .A2(REG_FILE_reg_out_11__23_), .ZN(n17951) );
  NAND2_X2 U18486 ( .A1(n13203), .A2(REG_FILE_reg_out_13__23_), .ZN(n17950) );
  NAND4_X2 U18487 ( .A1(n17953), .A2(n17952), .A3(n17951), .A4(n17950), .ZN(
        n17956) );
  OAI22_X2 U18488 ( .A1(n12139), .A2(n13471), .B1(n10293), .B2(n13467), .ZN(
        n17955) );
  OAI22_X2 U18489 ( .A1(n12263), .A2(n13475), .B1(n10919), .B2(n13472), .ZN(
        n17954) );
  NAND2_X2 U18490 ( .A1(n13455), .A2(REG_FILE_reg_out_12__23_), .ZN(n17961) );
  NAND2_X2 U18491 ( .A1(n13194), .A2(REG_FILE_reg_out_19__23_), .ZN(n17960) );
  OAI22_X2 U18492 ( .A1(n13460), .A2(n12904), .B1(n13459), .B2(n12758), .ZN(
        n17963) );
  OAI22_X2 U18493 ( .A1(n13465), .A2(n11888), .B1(n12410), .B2(n13463), .ZN(
        n17962) );
  OAI222_X2 U18494 ( .A1(n10773), .A2(n13477), .B1(n12543), .B2(net231223), 
        .C1(n18790), .C2(n13206), .ZN(n7636) );
  NAND2_X2 U18495 ( .A1(n13411), .A2(ID_EXEC_OUT[183]), .ZN(n17972) );
  NAND2_X2 U18496 ( .A1(DMEM_BUS_OUT[55]), .A2(net231319), .ZN(n17971) );
  NAND2_X2 U18497 ( .A1(n13413), .A2(DMEM_BUS_OUT[23]), .ZN(n17970) );
  NAND2_X2 U18498 ( .A1(n13415), .A2(MEM_WB_OUT[60]), .ZN(n17969) );
  NAND4_X2 U18499 ( .A1(n17972), .A2(n17971), .A3(n17970), .A4(n17969), .ZN(
        n7637) );
  OAI22_X2 U18500 ( .A1(n11529), .A2(net231257), .B1(net230377), .B2(n10773), 
        .ZN(n7638) );
  OAI22_X2 U18501 ( .A1(net231251), .A2(n11985), .B1(n19323), .B2(net230383), 
        .ZN(n7641) );
  OAI22_X2 U18502 ( .A1(n19323), .A2(net231257), .B1(n13481), .B2(n17973), 
        .ZN(n7642) );
  XNOR2_X2 U18503 ( .A(n17974), .B(net223794), .ZN(n17977) );
  NAND2_X2 U18504 ( .A1(net231615), .A2(n18922), .ZN(n17976) );
  NAND2_X2 U18505 ( .A1(EXEC_MEM_OUT_132), .A2(net231323), .ZN(n17975) );
  OAI211_X2 U18506 ( .C1(n17977), .C2(net231915), .A(n17976), .B(n17975), .ZN(
        n7643) );
  MUX2_X2 U18507 ( .A(DMEM_BUS_OUT[23]), .B(MEM_WB_OUT[60]), .S(net231293), 
        .Z(n7644) );
  NAND2_X2 U18509 ( .A1(n17982), .A2(n17981), .ZN(n17986) );
  NAND2_X2 U18510 ( .A1(n17983), .A2(ID_EXEC_OUT[55]), .ZN(n17985) );
  NAND2_X2 U18511 ( .A1(n18566), .A2(DMEM_BUS_OUT[23]), .ZN(n17984) );
  NAND3_X2 U18512 ( .A1(n17986), .A2(n17985), .A3(n17984), .ZN(n17987) );
  INV_X4 U18513 ( .A(n17988), .ZN(n17990) );
  NOR2_X4 U18514 ( .A1(n17990), .A2(n17989), .ZN(n17991) );
  NAND3_X4 U18515 ( .A1(n17993), .A2(n17992), .A3(n17991), .ZN(n18472) );
  AOI22_X2 U18516 ( .A1(n13388), .A2(n18472), .B1(n13397), .B2(n18329), .ZN(
        n17996) );
  AOI22_X2 U18517 ( .A1(n13487), .A2(n18328), .B1(n13392), .B2(n17994), .ZN(
        n17995) );
  NAND2_X2 U18518 ( .A1(n17996), .A2(n17995), .ZN(n18301) );
  INV_X4 U18519 ( .A(n18301), .ZN(n18004) );
  NAND2_X2 U18520 ( .A1(n10843), .A2(n18345), .ZN(n18001) );
  NAND2_X2 U18521 ( .A1(n18309), .A2(n19100), .ZN(n17997) );
  INV_X4 U18522 ( .A(n17997), .ZN(n18346) );
  NAND2_X2 U18523 ( .A1(n18346), .A2(n13149), .ZN(n18000) );
  NAND2_X2 U18524 ( .A1(n18310), .A2(n13159), .ZN(n17999) );
  NAND2_X2 U18525 ( .A1(n18347), .A2(n13163), .ZN(n17998) );
  NAND4_X2 U18526 ( .A1(n18001), .A2(n18000), .A3(n17999), .A4(n17998), .ZN(
        n18292) );
  NAND2_X2 U18527 ( .A1(n19124), .A2(n18292), .ZN(n18002) );
  OAI21_X4 U18528 ( .B1(n18004), .B2(n18003), .A(n18002), .ZN(n18011) );
  INV_X4 U18529 ( .A(n18005), .ZN(n18009) );
  NAND2_X2 U18530 ( .A1(n10199), .A2(n18006), .ZN(n18007) );
  OAI21_X4 U18531 ( .B1(n18011), .B2(n18010), .A(n18651), .ZN(n18016) );
  INV_X4 U18532 ( .A(n18978), .ZN(n18014) );
  NAND4_X2 U18533 ( .A1(n18018), .A2(n18017), .A3(n18016), .A4(n18015), .ZN(
        n7645) );
  OAI211_X2 U18534 ( .C1(n12173), .C2(net231225), .A(n18019), .B(n6750), .ZN(
        n7649) );
  XNOR2_X2 U18535 ( .A(n18020), .B(net223740), .ZN(n18022) );
  NAND2_X2 U18536 ( .A1(net231615), .A2(n13149), .ZN(n18021) );
  OAI221_X2 U18537 ( .B1(net231227), .B2(n11476), .C1(net231915), .C2(n18022), 
        .A(n18021), .ZN(n7650) );
  NAND2_X2 U18538 ( .A1(REG_FILE_reg_out_17__24_), .A2(n13434), .ZN(n18028) );
  OAI22_X2 U18539 ( .A1(n13420), .A2(n12817), .B1(n13417), .B2(n11874), .ZN(
        n18031) );
  OAI22_X2 U18540 ( .A1(n13440), .A2(n12593), .B1(n13438), .B2(n12578), .ZN(
        n18030) );
  NOR3_X4 U18541 ( .A1(n18032), .A2(n18031), .A3(n18030), .ZN(n18058) );
  NAND2_X2 U18542 ( .A1(n18493), .A2(REG_FILE_reg_out_6__24_), .ZN(n18036) );
  NAND2_X2 U18543 ( .A1(n13191), .A2(REG_FILE_reg_out_7__24_), .ZN(n18035) );
  NAND2_X2 U18544 ( .A1(n18494), .A2(REG_FILE_reg_out_4__24_), .ZN(n18034) );
  NAND2_X2 U18545 ( .A1(n13189), .A2(REG_FILE_reg_out_5__24_), .ZN(n18033) );
  NAND4_X2 U18546 ( .A1(n18036), .A2(n18035), .A3(n18034), .A4(n18033), .ZN(
        n18039) );
  OAI22_X2 U18547 ( .A1(n11423), .A2(n13445), .B1(n10523), .B2(n13442), .ZN(
        n18038) );
  OAI22_X2 U18548 ( .A1(n12778), .A2(n13451), .B1(n12043), .B2(n13448), .ZN(
        n18037) );
  NAND2_X2 U18549 ( .A1(n13198), .A2(REG_FILE_reg_out_14__24_), .ZN(n18043) );
  NAND2_X2 U18550 ( .A1(n13200), .A2(REG_FILE_reg_out_1__24_), .ZN(n18042) );
  NAND2_X2 U18551 ( .A1(n18502), .A2(REG_FILE_reg_out_11__24_), .ZN(n18041) );
  NAND2_X2 U18552 ( .A1(n13203), .A2(REG_FILE_reg_out_13__24_), .ZN(n18040) );
  NAND4_X2 U18553 ( .A1(n18043), .A2(n18042), .A3(n18041), .A4(n18040), .ZN(
        n18046) );
  OAI22_X2 U18554 ( .A1(n12140), .A2(n13471), .B1(n10294), .B2(n13467), .ZN(
        n18045) );
  OAI22_X2 U18555 ( .A1(n12264), .A2(n13475), .B1(n10920), .B2(n13472), .ZN(
        n18044) );
  NAND2_X2 U18556 ( .A1(n13455), .A2(REG_FILE_reg_out_12__24_), .ZN(n18051) );
  NAND2_X2 U18557 ( .A1(n13194), .A2(REG_FILE_reg_out_19__24_), .ZN(n18050) );
  OAI22_X2 U18558 ( .A1(n13460), .A2(n12906), .B1(n13459), .B2(n12759), .ZN(
        n18053) );
  OAI22_X2 U18559 ( .A1(n13465), .A2(n11889), .B1(n11497), .B2(n13463), .ZN(
        n18052) );
  OAI222_X2 U18560 ( .A1(n10774), .A2(n13476), .B1(n11560), .B2(net231223), 
        .C1(n12028), .C2(n13206), .ZN(n7652) );
  NAND2_X2 U18561 ( .A1(n13411), .A2(ID_EXEC_OUT[184]), .ZN(n18062) );
  NAND2_X2 U18562 ( .A1(DMEM_BUS_OUT[56]), .A2(net231323), .ZN(n18061) );
  NAND2_X2 U18563 ( .A1(n13413), .A2(DMEM_BUS_OUT[24]), .ZN(n18060) );
  NAND2_X2 U18564 ( .A1(n13416), .A2(MEM_WB_OUT[61]), .ZN(n18059) );
  NAND4_X2 U18565 ( .A1(n18062), .A2(n18061), .A3(n18060), .A4(n18059), .ZN(
        n7653) );
  OAI22_X2 U18566 ( .A1(n11530), .A2(net231257), .B1(net230377), .B2(n10774), 
        .ZN(n7654) );
  OAI22_X2 U18567 ( .A1(n12500), .A2(net231257), .B1(n13481), .B2(n18063), 
        .ZN(n7658) );
  OAI221_X2 U18568 ( .B1(net231227), .B2(n11477), .C1(net231915), .C2(n18065), 
        .A(n18064), .ZN(n7659) );
  NAND2_X2 U18569 ( .A1(REG_FILE_reg_out_17__25_), .A2(n13434), .ZN(n18071) );
  OAI22_X2 U18570 ( .A1(n13420), .A2(n12818), .B1(n13418), .B2(n11875), .ZN(
        n18074) );
  OAI22_X2 U18571 ( .A1(n13440), .A2(n12594), .B1(n13438), .B2(n12579), .ZN(
        n18073) );
  NOR3_X4 U18572 ( .A1(n18075), .A2(n18074), .A3(n18073), .ZN(n18101) );
  NAND2_X2 U18573 ( .A1(n18493), .A2(REG_FILE_reg_out_6__25_), .ZN(n18079) );
  NAND2_X2 U18574 ( .A1(n13191), .A2(REG_FILE_reg_out_7__25_), .ZN(n18078) );
  NAND2_X2 U18575 ( .A1(n18494), .A2(REG_FILE_reg_out_4__25_), .ZN(n18077) );
  NAND2_X2 U18576 ( .A1(n13189), .A2(REG_FILE_reg_out_5__25_), .ZN(n18076) );
  NAND4_X2 U18577 ( .A1(n18079), .A2(n18078), .A3(n18077), .A4(n18076), .ZN(
        n18082) );
  OAI22_X2 U18578 ( .A1(n11424), .A2(n13444), .B1(n10524), .B2(n13443), .ZN(
        n18081) );
  OAI22_X2 U18579 ( .A1(n12779), .A2(n13451), .B1(n12044), .B2(n13448), .ZN(
        n18080) );
  NAND2_X2 U18580 ( .A1(n13198), .A2(REG_FILE_reg_out_14__25_), .ZN(n18086) );
  NAND2_X2 U18581 ( .A1(n13200), .A2(REG_FILE_reg_out_1__25_), .ZN(n18085) );
  NAND2_X2 U18582 ( .A1(n18502), .A2(REG_FILE_reg_out_11__25_), .ZN(n18084) );
  NAND2_X2 U18583 ( .A1(n13203), .A2(REG_FILE_reg_out_13__25_), .ZN(n18083) );
  NAND4_X2 U18584 ( .A1(n18086), .A2(n18085), .A3(n18084), .A4(n18083), .ZN(
        n18089) );
  OAI22_X2 U18585 ( .A1(n12141), .A2(n13471), .B1(n10295), .B2(n13467), .ZN(
        n18088) );
  OAI22_X2 U18586 ( .A1(n12265), .A2(n13475), .B1(n10921), .B2(n13472), .ZN(
        n18087) );
  NAND2_X2 U18587 ( .A1(n13455), .A2(REG_FILE_reg_out_12__25_), .ZN(n18094) );
  NAND2_X2 U18588 ( .A1(n13194), .A2(REG_FILE_reg_out_19__25_), .ZN(n18093) );
  OAI22_X2 U18589 ( .A1(n13460), .A2(n12908), .B1(n13459), .B2(n12760), .ZN(
        n18096) );
  OAI22_X2 U18590 ( .A1(n13465), .A2(n11890), .B1(n11498), .B2(n13463), .ZN(
        n18095) );
  OAI222_X2 U18591 ( .A1(n10775), .A2(n13476), .B1(n11570), .B2(net231223), 
        .C1(n12300), .C2(n13206), .ZN(n7661) );
  NAND2_X2 U18592 ( .A1(n13411), .A2(ID_EXEC_OUT[185]), .ZN(n18105) );
  NAND2_X2 U18593 ( .A1(DMEM_BUS_OUT[57]), .A2(net231319), .ZN(n18104) );
  NAND2_X2 U18594 ( .A1(n13413), .A2(DMEM_BUS_OUT[25]), .ZN(n18103) );
  NAND2_X2 U18595 ( .A1(n13415), .A2(MEM_WB_OUT[62]), .ZN(n18102) );
  NAND4_X2 U18596 ( .A1(n18105), .A2(n18104), .A3(n18103), .A4(n18102), .ZN(
        n7662) );
  OAI22_X2 U18597 ( .A1(n11531), .A2(net231257), .B1(net230377), .B2(n10775), 
        .ZN(n7663) );
  OAI22_X2 U18598 ( .A1(net231249), .A2(net223591), .B1(n19322), .B2(net230383), .ZN(n7666) );
  OAI22_X2 U18599 ( .A1(n19322), .A2(net231257), .B1(n13480), .B2(n18106), 
        .ZN(n7667) );
  INV_X4 U18600 ( .A(n18107), .ZN(n18108) );
  XNOR2_X2 U18601 ( .A(net223586), .B(n18108), .ZN(n18110) );
  NAND2_X2 U18602 ( .A1(net231615), .A2(n18345), .ZN(n18109) );
  OAI221_X2 U18603 ( .B1(net231227), .B2(n12316), .C1(n18110), .C2(net231915), 
        .A(n18109), .ZN(n7668) );
  NAND2_X2 U18604 ( .A1(REG_FILE_reg_out_17__26_), .A2(n13434), .ZN(n18116) );
  OAI22_X2 U18605 ( .A1(n13420), .A2(n12819), .B1(n13417), .B2(n11876), .ZN(
        n18119) );
  OAI22_X2 U18606 ( .A1(n13440), .A2(n12595), .B1(n13438), .B2(n12580), .ZN(
        n18118) );
  NOR3_X4 U18607 ( .A1(n18120), .A2(n18119), .A3(n18118), .ZN(n18146) );
  NAND2_X2 U18608 ( .A1(n18493), .A2(REG_FILE_reg_out_6__26_), .ZN(n18124) );
  NAND2_X2 U18609 ( .A1(n13191), .A2(REG_FILE_reg_out_7__26_), .ZN(n18123) );
  NAND2_X2 U18610 ( .A1(n18494), .A2(REG_FILE_reg_out_4__26_), .ZN(n18122) );
  NAND2_X2 U18611 ( .A1(n13189), .A2(REG_FILE_reg_out_5__26_), .ZN(n18121) );
  NAND4_X2 U18612 ( .A1(n18124), .A2(n18123), .A3(n18122), .A4(n18121), .ZN(
        n18127) );
  OAI22_X2 U18613 ( .A1(n11425), .A2(n13445), .B1(n10525), .B2(n13442), .ZN(
        n18126) );
  OAI22_X2 U18614 ( .A1(n12780), .A2(n13451), .B1(n12045), .B2(n13448), .ZN(
        n18125) );
  NAND2_X2 U18615 ( .A1(n13198), .A2(REG_FILE_reg_out_14__26_), .ZN(n18131) );
  NAND2_X2 U18616 ( .A1(n13200), .A2(REG_FILE_reg_out_1__26_), .ZN(n18130) );
  NAND2_X2 U18617 ( .A1(n18502), .A2(REG_FILE_reg_out_11__26_), .ZN(n18129) );
  NAND2_X2 U18618 ( .A1(n13203), .A2(REG_FILE_reg_out_13__26_), .ZN(n18128) );
  NAND4_X2 U18619 ( .A1(n18131), .A2(n18130), .A3(n18129), .A4(n18128), .ZN(
        n18134) );
  OAI22_X2 U18620 ( .A1(n12142), .A2(n13471), .B1(n10296), .B2(n13467), .ZN(
        n18133) );
  OAI22_X2 U18621 ( .A1(n12266), .A2(n13475), .B1(n10922), .B2(n13472), .ZN(
        n18132) );
  NAND2_X2 U18622 ( .A1(n13455), .A2(REG_FILE_reg_out_12__26_), .ZN(n18139) );
  NAND2_X2 U18623 ( .A1(n13194), .A2(REG_FILE_reg_out_19__26_), .ZN(n18138) );
  OAI22_X2 U18624 ( .A1(n13460), .A2(n12910), .B1(n13459), .B2(n12761), .ZN(
        n18141) );
  OAI22_X2 U18625 ( .A1(n13465), .A2(n11891), .B1(n11499), .B2(n13463), .ZN(
        n18140) );
  OAI222_X2 U18626 ( .A1(n10776), .A2(n13476), .B1(n11561), .B2(net231223), 
        .C1(n10240), .C2(n13206), .ZN(n7670) );
  NAND2_X2 U18627 ( .A1(n13411), .A2(ID_EXEC_OUT[186]), .ZN(n18150) );
  NAND2_X2 U18628 ( .A1(DMEM_BUS_OUT[58]), .A2(net231319), .ZN(n18149) );
  NAND2_X2 U18629 ( .A1(n13413), .A2(DMEM_BUS_OUT[26]), .ZN(n18148) );
  NAND2_X2 U18630 ( .A1(n13416), .A2(MEM_WB_OUT[63]), .ZN(n18147) );
  NAND4_X2 U18631 ( .A1(n18150), .A2(n18149), .A3(n18148), .A4(n18147), .ZN(
        n7671) );
  OAI22_X2 U18632 ( .A1(n11532), .A2(net231259), .B1(net230383), .B2(n10776), 
        .ZN(n7672) );
  OAI22_X2 U18633 ( .A1(n12191), .A2(net231259), .B1(n13480), .B2(n18151), 
        .ZN(n7676) );
  NAND2_X2 U18634 ( .A1(REG_FILE_reg_out_17__27_), .A2(n13434), .ZN(n18157) );
  OAI22_X2 U18635 ( .A1(n13420), .A2(n12820), .B1(n13417), .B2(n11877), .ZN(
        n18160) );
  OAI22_X2 U18636 ( .A1(n13440), .A2(n12596), .B1(n13438), .B2(n12581), .ZN(
        n18159) );
  NOR3_X4 U18637 ( .A1(n18161), .A2(n18160), .A3(n18159), .ZN(n18187) );
  NAND2_X2 U18638 ( .A1(n18493), .A2(REG_FILE_reg_out_6__27_), .ZN(n18165) );
  NAND2_X2 U18639 ( .A1(n13191), .A2(REG_FILE_reg_out_7__27_), .ZN(n18164) );
  NAND2_X2 U18640 ( .A1(n18494), .A2(REG_FILE_reg_out_4__27_), .ZN(n18163) );
  NAND2_X2 U18641 ( .A1(n13189), .A2(REG_FILE_reg_out_5__27_), .ZN(n18162) );
  NAND4_X2 U18642 ( .A1(n18165), .A2(n18164), .A3(n18163), .A4(n18162), .ZN(
        n18168) );
  OAI22_X2 U18643 ( .A1(n11426), .A2(n13444), .B1(n10526), .B2(n13442), .ZN(
        n18167) );
  OAI22_X2 U18644 ( .A1(n12781), .A2(n13451), .B1(n12046), .B2(n13448), .ZN(
        n18166) );
  NAND2_X2 U18645 ( .A1(n13198), .A2(REG_FILE_reg_out_14__27_), .ZN(n18172) );
  NAND2_X2 U18646 ( .A1(n13200), .A2(REG_FILE_reg_out_1__27_), .ZN(n18171) );
  NAND2_X2 U18647 ( .A1(n18502), .A2(REG_FILE_reg_out_11__27_), .ZN(n18170) );
  NAND2_X2 U18648 ( .A1(n13203), .A2(REG_FILE_reg_out_13__27_), .ZN(n18169) );
  NAND4_X2 U18649 ( .A1(n18172), .A2(n18171), .A3(n18170), .A4(n18169), .ZN(
        n18175) );
  OAI22_X2 U18650 ( .A1(n12143), .A2(n13471), .B1(n10297), .B2(n13467), .ZN(
        n18174) );
  OAI22_X2 U18651 ( .A1(n12267), .A2(n13475), .B1(n10923), .B2(n13472), .ZN(
        n18173) );
  NAND2_X2 U18652 ( .A1(n13455), .A2(REG_FILE_reg_out_12__27_), .ZN(n18180) );
  NAND2_X2 U18653 ( .A1(n13194), .A2(REG_FILE_reg_out_19__27_), .ZN(n18179) );
  OAI22_X2 U18654 ( .A1(n13460), .A2(n12912), .B1(n13459), .B2(n12762), .ZN(
        n18182) );
  OAI22_X2 U18655 ( .A1(n13465), .A2(n11892), .B1(n11500), .B2(n13463), .ZN(
        n18181) );
  OAI222_X2 U18656 ( .A1(n18189), .A2(n18188), .B1(n10780), .B2(n13476), .C1(
        n11563), .C2(net231221), .ZN(n7678) );
  NAND2_X2 U18657 ( .A1(n13411), .A2(ID_EXEC_OUT[187]), .ZN(n18193) );
  NAND2_X2 U18658 ( .A1(DMEM_BUS_OUT[59]), .A2(net231319), .ZN(n18192) );
  NAND2_X2 U18659 ( .A1(n13413), .A2(DMEM_BUS_OUT[27]), .ZN(n18191) );
  NAND2_X2 U18660 ( .A1(n13415), .A2(MEM_WB_OUT[64]), .ZN(n18190) );
  NAND4_X2 U18661 ( .A1(n18193), .A2(n18192), .A3(n18191), .A4(n18190), .ZN(
        n7679) );
  OAI22_X2 U18662 ( .A1(n11533), .A2(net231259), .B1(net230381), .B2(n10780), 
        .ZN(n7680) );
  OAI22_X2 U18663 ( .A1(net231251), .A2(net239554), .B1(n19321), .B2(net230381), .ZN(n7683) );
  OAI22_X2 U18664 ( .A1(n19321), .A2(net231259), .B1(n13480), .B2(n18194), 
        .ZN(n7684) );
  XNOR2_X2 U18665 ( .A(net223439), .B(net223440), .ZN(n18196) );
  NAND2_X2 U18666 ( .A1(EXEC_MEM_OUT_136), .A2(net231323), .ZN(n18195) );
  OAI221_X2 U18667 ( .B1(n18196), .B2(net231915), .C1(n18962), .C2(net223104), 
        .A(n18195), .ZN(n7685) );
  NAND2_X2 U18668 ( .A1(REG_FILE_reg_out_17__28_), .A2(n13434), .ZN(n18202) );
  OAI22_X2 U18669 ( .A1(n13420), .A2(n12821), .B1(n13418), .B2(n11878), .ZN(
        n18205) );
  OAI22_X2 U18670 ( .A1(n13440), .A2(n12597), .B1(n13438), .B2(n12582), .ZN(
        n18204) );
  NOR3_X4 U18671 ( .A1(n18206), .A2(n18205), .A3(n18204), .ZN(n18232) );
  NAND2_X2 U18672 ( .A1(n18493), .A2(REG_FILE_reg_out_6__28_), .ZN(n18210) );
  NAND2_X2 U18673 ( .A1(n13191), .A2(REG_FILE_reg_out_7__28_), .ZN(n18209) );
  NAND2_X2 U18674 ( .A1(n18494), .A2(REG_FILE_reg_out_4__28_), .ZN(n18208) );
  NAND2_X2 U18675 ( .A1(n13189), .A2(REG_FILE_reg_out_5__28_), .ZN(n18207) );
  NAND4_X2 U18676 ( .A1(n18210), .A2(n18209), .A3(n18208), .A4(n18207), .ZN(
        n18213) );
  OAI22_X2 U18677 ( .A1(n11427), .A2(n13444), .B1(n10527), .B2(n13443), .ZN(
        n18212) );
  OAI22_X2 U18678 ( .A1(n12782), .A2(n13451), .B1(n12047), .B2(n13448), .ZN(
        n18211) );
  NAND2_X2 U18679 ( .A1(n13198), .A2(REG_FILE_reg_out_14__28_), .ZN(n18217) );
  NAND2_X2 U18680 ( .A1(n13200), .A2(REG_FILE_reg_out_1__28_), .ZN(n18216) );
  NAND2_X2 U18681 ( .A1(n18502), .A2(REG_FILE_reg_out_11__28_), .ZN(n18215) );
  NAND2_X2 U18682 ( .A1(n13203), .A2(REG_FILE_reg_out_13__28_), .ZN(n18214) );
  NAND4_X2 U18683 ( .A1(n18217), .A2(n18216), .A3(n18215), .A4(n18214), .ZN(
        n18220) );
  OAI22_X2 U18684 ( .A1(n12144), .A2(n13471), .B1(n10298), .B2(n13467), .ZN(
        n18219) );
  OAI22_X2 U18685 ( .A1(n12268), .A2(n13475), .B1(n10924), .B2(n13472), .ZN(
        n18218) );
  NAND2_X2 U18686 ( .A1(n13455), .A2(REG_FILE_reg_out_12__28_), .ZN(n18225) );
  NAND2_X2 U18687 ( .A1(n13194), .A2(REG_FILE_reg_out_19__28_), .ZN(n18224) );
  OAI22_X2 U18688 ( .A1(n13460), .A2(n12914), .B1(n13459), .B2(n12763), .ZN(
        n18227) );
  OAI22_X2 U18689 ( .A1(n13465), .A2(n11893), .B1(n11501), .B2(n13463), .ZN(
        n18226) );
  OAI222_X2 U18690 ( .A1(n10777), .A2(n13476), .B1(n11280), .B2(net231223), 
        .C1(n10840), .C2(n13206), .ZN(n7687) );
  NAND2_X2 U18691 ( .A1(n13411), .A2(ID_EXEC_OUT[188]), .ZN(n18236) );
  NAND2_X2 U18692 ( .A1(DMEM_BUS_OUT[60]), .A2(net231319), .ZN(n18235) );
  NAND2_X2 U18693 ( .A1(n13413), .A2(DMEM_BUS_OUT[28]), .ZN(n18234) );
  NAND2_X2 U18694 ( .A1(n13416), .A2(MEM_WB_OUT[65]), .ZN(n18233) );
  NAND4_X2 U18695 ( .A1(n18236), .A2(n18235), .A3(n18234), .A4(n18233), .ZN(
        n7688) );
  OAI22_X2 U18696 ( .A1(n11534), .A2(net231259), .B1(net230377), .B2(n10777), 
        .ZN(n7689) );
  OAI22_X2 U18697 ( .A1(n12192), .A2(net231259), .B1(n18237), .B2(n13481), 
        .ZN(n7693) );
  XNOR2_X2 U18698 ( .A(n18239), .B(n18238), .ZN(n18242) );
  NAND2_X2 U18699 ( .A1(EXEC_MEM_OUT_137), .A2(net231323), .ZN(n18240) );
  OAI211_X2 U18700 ( .C1(n18242), .C2(net231915), .A(n18241), .B(n18240), .ZN(
        n7694) );
  MUX2_X2 U18701 ( .A(DMEM_BUS_OUT[28]), .B(MEM_WB_OUT[65]), .S(net231293), 
        .Z(n7695) );
  NAND2_X2 U18702 ( .A1(n13386), .A2(n13149), .ZN(n18246) );
  NAND2_X2 U18703 ( .A1(net232816), .A2(n19029), .ZN(n18243) );
  NAND4_X2 U18704 ( .A1(n18246), .A2(n18245), .A3(n18244), .A4(n18243), .ZN(
        n18533) );
  AOI22_X2 U18705 ( .A1(n18346), .A2(n13163), .B1(n13487), .B2(n18533), .ZN(
        n18257) );
  NAND2_X2 U18706 ( .A1(net223324), .A2(n18867), .ZN(n18249) );
  NAND2_X2 U18707 ( .A1(net232816), .A2(n19000), .ZN(n18248) );
  NAND2_X2 U18708 ( .A1(n15733), .A2(n18539), .ZN(n18256) );
  NAND2_X2 U18709 ( .A1(n13393), .A2(n18339), .ZN(n18255) );
  NAND2_X2 U18710 ( .A1(n13386), .A2(n18345), .ZN(n18253) );
  NAND2_X2 U18711 ( .A1(net223324), .A2(n18873), .ZN(n18251) );
  NAND2_X2 U18712 ( .A1(net232816), .A2(n19015), .ZN(n18250) );
  NAND4_X2 U18713 ( .A1(n18253), .A2(n18252), .A3(n18251), .A4(n18250), .ZN(
        n18541) );
  NAND2_X2 U18714 ( .A1(n16061), .A2(n18541), .ZN(n18254) );
  NAND4_X2 U18715 ( .A1(n18257), .A2(n18256), .A3(n18255), .A4(n18254), .ZN(
        n18258) );
  INV_X4 U18716 ( .A(n18258), .ZN(n18452) );
  OAI22_X2 U18717 ( .A1(n13217), .A2(n11981), .B1(n18452), .B2(n13211), .ZN(
        n18260) );
  NOR2_X4 U18718 ( .A1(n18260), .A2(n18259), .ZN(n18291) );
  MUX2_X2 U18719 ( .A(n13209), .B(n13491), .S(n18365), .Z(n18264) );
  AOI22_X2 U18720 ( .A1(n13490), .A2(n18262), .B1(n10829), .B2(
        DMEM_BUS_OUT[28]), .ZN(n18263) );
  MUX2_X2 U18721 ( .A(n18264), .B(n18263), .S(n18945), .Z(n18290) );
  NAND2_X2 U18723 ( .A1(n18266), .A2(n18265), .ZN(n18531) );
  NAND2_X2 U18724 ( .A1(n13393), .A2(n18329), .ZN(n18278) );
  NAND2_X2 U18725 ( .A1(n13488), .A2(n18472), .ZN(n18277) );
  NAND2_X2 U18726 ( .A1(net223324), .A2(n18872), .ZN(n18268) );
  NAND2_X2 U18727 ( .A1(net232816), .A2(n19004), .ZN(n18267) );
  NAND4_X2 U18728 ( .A1(n18270), .A2(n18269), .A3(n18268), .A4(n18267), .ZN(
        n19096) );
  NAND2_X2 U18729 ( .A1(net223324), .A2(n18870), .ZN(n18273) );
  NAND2_X2 U18730 ( .A1(net232816), .A2(n19013), .ZN(n18272) );
  NAND4_X2 U18731 ( .A1(n18275), .A2(n18274), .A3(n18273), .A4(n18272), .ZN(
        n18468) );
  AOI22_X2 U18732 ( .A1(n13388), .A2(n19096), .B1(n13397), .B2(n18468), .ZN(
        n18276) );
  AOI22_X2 U18733 ( .A1(n18531), .A2(n10363), .B1(n19118), .B2(n18367), .ZN(
        n18289) );
  NOR3_X4 U18734 ( .A1(n18283), .A2(n18550), .A3(n18282), .ZN(n18287) );
  INV_X4 U18735 ( .A(n13161), .ZN(n18455) );
  INV_X4 U18736 ( .A(n18284), .ZN(n19107) );
  NAND2_X2 U18737 ( .A1(n18644), .A2(n19107), .ZN(n18463) );
  NAND4_X2 U18738 ( .A1(n18291), .A2(n18290), .A3(n18289), .A4(n18288), .ZN(
        n7696) );
  MUX2_X2 U18739 ( .A(DMEM_BUS_OUT[24]), .B(MEM_WB_OUT[61]), .S(net231293), 
        .Z(n7697) );
  MUX2_X2 U18740 ( .A(n13209), .B(n13491), .S(n18925), .Z(n18295) );
  INV_X4 U18741 ( .A(n18924), .ZN(n18859) );
  MUX2_X2 U18742 ( .A(n18295), .B(n18294), .S(n18859), .Z(n18319) );
  NAND2_X2 U18743 ( .A1(n16061), .A2(n18339), .ZN(n18300) );
  NAND2_X2 U18744 ( .A1(n15733), .A2(n18533), .ZN(n18299) );
  NAND2_X2 U18745 ( .A1(n13488), .A2(n18338), .ZN(n18298) );
  NAND2_X2 U18746 ( .A1(n13393), .A2(n18296), .ZN(n18297) );
  NAND4_X2 U18747 ( .A1(n18300), .A2(n18299), .A3(n18298), .A4(n18297), .ZN(
        n18392) );
  AOI22_X2 U18748 ( .A1(n18302), .A2(n18301), .B1(n18392), .B2(n17924), .ZN(
        n18318) );
  NAND2_X2 U18749 ( .A1(n18309), .A2(n18308), .ZN(n18313) );
  NAND2_X2 U18750 ( .A1(n18347), .A2(n13161), .ZN(n18312) );
  NAND2_X2 U18751 ( .A1(n18310), .A2(n13151), .ZN(n18311) );
  NAND3_X4 U18752 ( .A1(n18313), .A2(n18312), .A3(n18311), .ZN(n18394) );
  INV_X4 U18753 ( .A(n18394), .ZN(n18314) );
  NAND4_X2 U18754 ( .A1(n18320), .A2(n18319), .A3(n18318), .A4(n18317), .ZN(
        n7698) );
  NAND2_X2 U18755 ( .A1(n13409), .A2(n18345), .ZN(n18321) );
  OAI211_X2 U18756 ( .C1(n12171), .C2(net231227), .A(n18321), .B(n6752), .ZN(
        n7702) );
  MUX2_X2 U18757 ( .A(DMEM_BUS_OUT[26]), .B(MEM_WB_OUT[63]), .S(net231291), 
        .Z(n7703) );
  XNOR2_X2 U18758 ( .A(n18324), .B(n18323), .ZN(n18327) );
  INV_X4 U18759 ( .A(n18958), .ZN(n18325) );
  AOI21_X4 U18760 ( .B1(n13492), .B2(n18327), .A(n18326), .ZN(n18357) );
  NAND2_X2 U18761 ( .A1(n16061), .A2(n18472), .ZN(n18333) );
  NAND2_X2 U18762 ( .A1(n13388), .A2(n18468), .ZN(n18332) );
  NAND2_X2 U18763 ( .A1(n16207), .A2(n18328), .ZN(n18331) );
  NAND2_X2 U18764 ( .A1(n13488), .A2(n18329), .ZN(n18330) );
  NAND4_X2 U18765 ( .A1(n18333), .A2(n18332), .A3(n18331), .A4(n18330), .ZN(
        n18393) );
  NAND2_X2 U18766 ( .A1(n19118), .A2(n18393), .ZN(n18356) );
  NAND2_X2 U18767 ( .A1(n10363), .A2(n13161), .ZN(n18336) );
  NAND2_X2 U18768 ( .A1(n18347), .A2(n13151), .ZN(n18334) );
  NAND3_X4 U18769 ( .A1(n18336), .A2(n18335), .A3(n18334), .ZN(n18359) );
  XNOR2_X2 U18770 ( .A(n18958), .B(n18345), .ZN(n18959) );
  AOI21_X4 U18771 ( .B1(n18644), .B2(n18359), .A(n18337), .ZN(n18355) );
  NAND2_X2 U18772 ( .A1(n13393), .A2(n18338), .ZN(n18343) );
  NAND2_X2 U18773 ( .A1(n13488), .A2(n18339), .ZN(n18342) );
  AOI22_X2 U18774 ( .A1(n13397), .A2(n18533), .B1(n13388), .B2(n18541), .ZN(
        n18341) );
  NAND3_X4 U18775 ( .A1(n18343), .A2(n18342), .A3(n18341), .ZN(n18368) );
  NAND2_X2 U18776 ( .A1(DMEM_BUS_OUT[26]), .A2(net231323), .ZN(n18344) );
  NAND2_X2 U18777 ( .A1(n10363), .A2(n13163), .ZN(n18350) );
  NAND2_X2 U18778 ( .A1(n18346), .A2(n18345), .ZN(n18349) );
  NAND2_X2 U18779 ( .A1(n18347), .A2(n13159), .ZN(n18348) );
  INV_X4 U18780 ( .A(n18397), .ZN(n18351) );
  NOR2_X4 U18781 ( .A1(n18351), .A2(n13214), .ZN(n18352) );
  NAND4_X2 U18782 ( .A1(n18357), .A2(n18356), .A3(n18355), .A4(n18354), .ZN(
        n7704) );
  OAI211_X2 U18783 ( .C1(n12172), .C2(net231223), .A(n18358), .B(n6751), .ZN(
        n7708) );
  MUX2_X2 U18784 ( .A(DMEM_BUS_OUT[27]), .B(MEM_WB_OUT[64]), .S(net231291), 
        .Z(n7709) );
  NAND2_X2 U18785 ( .A1(n18360), .A2(n18359), .ZN(n18382) );
  NAND2_X2 U18787 ( .A1(n13492), .A2(n18363), .ZN(n18381) );
  INV_X4 U18788 ( .A(n18368), .ZN(n18370) );
  NAND2_X2 U18789 ( .A1(ID_EXEC_OUT[231]), .A2(n13216), .ZN(n18369) );
  OAI21_X4 U18790 ( .B1(n18370), .B2(n13213), .A(n18369), .ZN(n18378) );
  MUX2_X2 U18791 ( .A(n13208), .B(n13490), .S(n18962), .Z(n18375) );
  NAND2_X2 U18792 ( .A1(n10829), .A2(DMEM_BUS_OUT[27]), .ZN(n18371) );
  MUX2_X2 U18793 ( .A(n18375), .B(n18374), .S(n18373), .Z(n18376) );
  NAND4_X2 U18794 ( .A1(n18382), .A2(n18381), .A3(n18380), .A4(n18379), .ZN(
        n7710) );
  MUX2_X2 U18795 ( .A(DMEM_BUS_OUT[25]), .B(MEM_WB_OUT[62]), .S(net231291), 
        .Z(n7715) );
  MUX2_X2 U18796 ( .A(n13209), .B(n13491), .S(n18858), .Z(n18387) );
  MUX2_X2 U18797 ( .A(n18387), .B(n18386), .S(n18967), .Z(n18389) );
  NAND2_X2 U18798 ( .A1(DMEM_BUS_OUT[25]), .A2(net231323), .ZN(n18388) );
  NAND2_X2 U18799 ( .A1(n18389), .A2(n18388), .ZN(n18391) );
  NAND2_X2 U18800 ( .A1(n19118), .A2(n18392), .ZN(n18402) );
  AOI22_X2 U18801 ( .A1(n18394), .A2(n18360), .B1(n17924), .B2(n18393), .ZN(
        n18401) );
  XNOR2_X2 U18802 ( .A(n18396), .B(n18395), .ZN(n18399) );
  NOR2_X4 U18803 ( .A1(n18351), .A2(n13207), .ZN(n18398) );
  NAND4_X2 U18804 ( .A1(n18403), .A2(n18402), .A3(n18401), .A4(n18400), .ZN(
        n7716) );
  NAND2_X2 U18805 ( .A1(n13409), .A2(n13161), .ZN(n18404) );
  OAI211_X2 U18806 ( .C1(n12174), .C2(net231225), .A(n18404), .B(n6749), .ZN(
        n7720) );
  NAND2_X2 U18807 ( .A1(REG_FILE_reg_out_17__29_), .A2(n13434), .ZN(n18410) );
  OAI22_X2 U18808 ( .A1(n13420), .A2(n12822), .B1(n13417), .B2(n11879), .ZN(
        n18413) );
  OAI22_X2 U18809 ( .A1(n13440), .A2(n12598), .B1(n13438), .B2(n12583), .ZN(
        n18412) );
  NOR3_X4 U18810 ( .A1(n18414), .A2(n18413), .A3(n18412), .ZN(n18440) );
  NAND2_X2 U18811 ( .A1(n18493), .A2(REG_FILE_reg_out_6__29_), .ZN(n18418) );
  NAND2_X2 U18812 ( .A1(n13191), .A2(REG_FILE_reg_out_7__29_), .ZN(n18417) );
  NAND2_X2 U18813 ( .A1(n18494), .A2(REG_FILE_reg_out_4__29_), .ZN(n18416) );
  NAND2_X2 U18814 ( .A1(n13189), .A2(REG_FILE_reg_out_5__29_), .ZN(n18415) );
  NAND4_X2 U18815 ( .A1(n18418), .A2(n18417), .A3(n18416), .A4(n18415), .ZN(
        n18421) );
  OAI22_X2 U18816 ( .A1(n11428), .A2(n13445), .B1(n10528), .B2(n13443), .ZN(
        n18420) );
  OAI22_X2 U18817 ( .A1(n12783), .A2(n13451), .B1(n12048), .B2(n13448), .ZN(
        n18419) );
  NAND2_X2 U18818 ( .A1(n13198), .A2(REG_FILE_reg_out_14__29_), .ZN(n18425) );
  NAND2_X2 U18819 ( .A1(n13200), .A2(REG_FILE_reg_out_1__29_), .ZN(n18424) );
  NAND2_X2 U18820 ( .A1(n18502), .A2(REG_FILE_reg_out_11__29_), .ZN(n18423) );
  NAND2_X2 U18821 ( .A1(n13203), .A2(REG_FILE_reg_out_13__29_), .ZN(n18422) );
  NAND4_X2 U18822 ( .A1(n18425), .A2(n18424), .A3(n18423), .A4(n18422), .ZN(
        n18428) );
  OAI22_X2 U18823 ( .A1(n12145), .A2(n13471), .B1(n10299), .B2(n13467), .ZN(
        n18427) );
  OAI22_X2 U18824 ( .A1(n12269), .A2(n13475), .B1(n10925), .B2(n13472), .ZN(
        n18426) );
  NAND2_X2 U18825 ( .A1(n13455), .A2(REG_FILE_reg_out_12__29_), .ZN(n18433) );
  NAND2_X2 U18826 ( .A1(n13194), .A2(REG_FILE_reg_out_19__29_), .ZN(n18432) );
  OAI22_X2 U18827 ( .A1(n13460), .A2(n12916), .B1(n13459), .B2(n12764), .ZN(
        n18435) );
  OAI22_X2 U18828 ( .A1(n13465), .A2(n11894), .B1(n11502), .B2(n13463), .ZN(
        n18434) );
  OAI222_X2 U18829 ( .A1(n10778), .A2(n13476), .B1(n11571), .B2(net231223), 
        .C1(n12039), .C2(n13206), .ZN(n7722) );
  NAND2_X2 U18830 ( .A1(n13411), .A2(ID_EXEC_OUT[189]), .ZN(n18444) );
  NAND2_X2 U18831 ( .A1(DMEM_BUS_OUT[61]), .A2(net231319), .ZN(n18443) );
  NAND2_X2 U18832 ( .A1(n13413), .A2(DMEM_BUS_OUT[29]), .ZN(n18442) );
  NAND2_X2 U18833 ( .A1(n13415), .A2(MEM_WB_OUT[66]), .ZN(n18441) );
  NAND4_X2 U18834 ( .A1(n18444), .A2(n18443), .A3(n18442), .A4(n18441), .ZN(
        n7723) );
  OAI22_X2 U18835 ( .A1(n11535), .A2(net231259), .B1(net230377), .B2(n10778), 
        .ZN(n7724) );
  INV_X4 U18836 ( .A(net137343), .ZN(net223109) );
  XNOR2_X2 U18837 ( .A(n18446), .B(net223109), .ZN(n18448) );
  XNOR2_X2 U18838 ( .A(n18448), .B(n18447), .ZN(n18450) );
  NAND2_X2 U18839 ( .A1(EXEC_MEM_OUT_138), .A2(net231323), .ZN(n18449) );
  OAI221_X2 U18840 ( .B1(n18450), .B2(net231915), .C1(n18455), .C2(net223104), 
        .A(n18449), .ZN(n7729) );
  MUX2_X2 U18841 ( .A(DMEM_BUS_OUT[29]), .B(MEM_WB_OUT[66]), .S(net231291), 
        .Z(n7730) );
  OAI22_X2 U18842 ( .A1(n19114), .A2(n10823), .B1(n18452), .B2(n13213), .ZN(
        n18454) );
  NOR2_X4 U18843 ( .A1(n18454), .A2(n18453), .ZN(n18481) );
  MUX2_X2 U18844 ( .A(n13209), .B(n13491), .S(n18455), .Z(n18459) );
  MUX2_X2 U18846 ( .A(n18459), .B(n18458), .S(n18943), .Z(n18480) );
  NAND2_X2 U18847 ( .A1(n19107), .A2(n13161), .ZN(n18461) );
  NAND2_X2 U18848 ( .A1(n18461), .A2(n18460), .ZN(n18465) );
  INV_X4 U18849 ( .A(net222497), .ZN(net223078) );
  MUX2_X2 U18850 ( .A(n18468), .B(net223077), .S(n18943), .Z(n18471) );
  NOR2_X4 U18851 ( .A1(n18455), .A2(n18469), .ZN(n18470) );
  NOR2_X4 U18852 ( .A1(n18471), .A2(n18470), .ZN(n19099) );
  NAND2_X2 U18853 ( .A1(n13397), .A2(n19096), .ZN(n18474) );
  NAND2_X2 U18854 ( .A1(n13392), .A2(n18472), .ZN(n18473) );
  INV_X4 U18855 ( .A(n18529), .ZN(n18475) );
  NOR2_X4 U18856 ( .A1(n18475), .A2(n13211), .ZN(n18476) );
  AOI21_X4 U18857 ( .B1(n13492), .B2(n18477), .A(n18476), .ZN(n18478) );
  NAND4_X2 U18858 ( .A1(n18481), .A2(n18480), .A3(n18479), .A4(n18478), .ZN(
        n7731) );
  OAI211_X2 U18860 ( .C1(n12175), .C2(net231225), .A(n18482), .B(n6748), .ZN(
        n7735) );
  NAND2_X2 U18861 ( .A1(REG_FILE_reg_out_17__30_), .A2(n13434), .ZN(n18488) );
  NOR2_X4 U18862 ( .A1(n13427), .A2(n12497), .ZN(n18485) );
  OAI22_X2 U18863 ( .A1(n13420), .A2(n12823), .B1(n13418), .B2(n11880), .ZN(
        n18491) );
  OAI22_X2 U18864 ( .A1(n13440), .A2(n12599), .B1(n13438), .B2(n12584), .ZN(
        n18490) );
  NOR3_X4 U18865 ( .A1(n18492), .A2(n18491), .A3(n18490), .ZN(n18521) );
  NAND2_X2 U18866 ( .A1(n18493), .A2(REG_FILE_reg_out_6__30_), .ZN(n18498) );
  NAND2_X2 U18867 ( .A1(n13191), .A2(REG_FILE_reg_out_7__30_), .ZN(n18497) );
  NAND2_X2 U18868 ( .A1(n18494), .A2(REG_FILE_reg_out_4__30_), .ZN(n18496) );
  NAND2_X2 U18869 ( .A1(n13189), .A2(REG_FILE_reg_out_5__30_), .ZN(n18495) );
  NAND4_X2 U18870 ( .A1(n18498), .A2(n18497), .A3(n18496), .A4(n18495), .ZN(
        n18501) );
  OAI22_X2 U18871 ( .A1(n11429), .A2(n13444), .B1(n10529), .B2(n13443), .ZN(
        n18500) );
  OAI22_X2 U18872 ( .A1(n12784), .A2(n13451), .B1(n12049), .B2(n13448), .ZN(
        n18499) );
  NAND2_X2 U18873 ( .A1(n13198), .A2(REG_FILE_reg_out_14__30_), .ZN(n18506) );
  NAND2_X2 U18874 ( .A1(n13200), .A2(REG_FILE_reg_out_1__30_), .ZN(n18505) );
  NAND2_X2 U18875 ( .A1(n18502), .A2(REG_FILE_reg_out_11__30_), .ZN(n18504) );
  NAND2_X2 U18876 ( .A1(n13203), .A2(REG_FILE_reg_out_13__30_), .ZN(n18503) );
  NAND4_X2 U18877 ( .A1(n18506), .A2(n18505), .A3(n18504), .A4(n18503), .ZN(
        n18509) );
  OAI22_X2 U18878 ( .A1(n12146), .A2(n13471), .B1(n10300), .B2(n13467), .ZN(
        n18508) );
  OAI22_X2 U18879 ( .A1(n12270), .A2(n13475), .B1(n10926), .B2(n13472), .ZN(
        n18507) );
  NAND2_X2 U18880 ( .A1(n13455), .A2(REG_FILE_reg_out_12__30_), .ZN(n18514) );
  NAND2_X2 U18881 ( .A1(n13194), .A2(REG_FILE_reg_out_19__30_), .ZN(n18513) );
  OAI22_X2 U18882 ( .A1(n13460), .A2(n12918), .B1(n13459), .B2(n12765), .ZN(
        n18516) );
  OAI22_X2 U18883 ( .A1(n13465), .A2(n11895), .B1(n11503), .B2(n13463), .ZN(
        n18515) );
  OAI222_X2 U18884 ( .A1(n10779), .A2(n13476), .B1(n11562), .B2(net231223), 
        .C1(n12027), .C2(n13206), .ZN(n7737) );
  NAND2_X2 U18885 ( .A1(n13411), .A2(ID_EXEC_OUT[190]), .ZN(n18525) );
  NAND2_X2 U18886 ( .A1(DMEM_BUS_OUT[62]), .A2(net231319), .ZN(n18524) );
  NAND2_X2 U18887 ( .A1(n13413), .A2(DMEM_BUS_OUT[30]), .ZN(n18523) );
  NAND2_X2 U18888 ( .A1(n13415), .A2(MEM_WB_OUT[67]), .ZN(n18522) );
  NAND4_X2 U18889 ( .A1(n18525), .A2(n18524), .A3(n18523), .A4(n18522), .ZN(
        n7738) );
  OAI22_X2 U18890 ( .A1(n11536), .A2(net231259), .B1(net230377), .B2(n10779), 
        .ZN(n7739) );
  OAI22_X2 U18891 ( .A1(n11108), .A2(net231259), .B1(net230377), .B2(net222982), .ZN(n7741) );
  OAI22_X2 U18892 ( .A1(net231251), .A2(net222982), .B1(n11110), .B2(net230383), .ZN(n7742) );
  OAI22_X2 U18893 ( .A1(n11110), .A2(net231259), .B1(n12311), .B2(n13481), 
        .ZN(n7743) );
  NAND2_X2 U18894 ( .A1(net231319), .A2(EXEC_MEM_OUT_139), .ZN(n18527) );
  OAI211_X2 U18896 ( .C1(n18528), .C2(net231915), .A(n18527), .B(n18526), .ZN(
        n7744) );
  MUX2_X2 U18897 ( .A(DMEM_BUS_OUT[30]), .B(MEM_WB_OUT[67]), .S(net231293), 
        .Z(n7745) );
  NAND2_X2 U18898 ( .A1(n19118), .A2(n18529), .ZN(n18557) );
  INV_X4 U18899 ( .A(n19038), .ZN(n18534) );
  INV_X4 U18900 ( .A(n18897), .ZN(n18536) );
  OAI21_X4 U18901 ( .B1(net232817), .B2(n18536), .A(n18535), .ZN(n18537) );
  OAI21_X4 U18902 ( .B1(n18538), .B2(n18537), .A(n18340), .ZN(n18544) );
  AOI22_X2 U18904 ( .A1(n13487), .A2(n18541), .B1(n16061), .B2(n18539), .ZN(
        n18542) );
  NAND4_X2 U18905 ( .A1(n18545), .A2(n18544), .A3(n18543), .A4(n18542), .ZN(
        n19117) );
  NAND2_X2 U18906 ( .A1(DMEM_BUS_OUT[30]), .A2(net231325), .ZN(n18546) );
  NAND4_X2 U18908 ( .A1(n18557), .A2(n18556), .A3(n18555), .A4(n18554), .ZN(
        n7746) );
  NAND2_X2 U18909 ( .A1(n13409), .A2(n18559), .ZN(n18558) );
  OAI211_X2 U18910 ( .C1(n12164), .C2(net231225), .A(n18558), .B(n6762), .ZN(
        n7750) );
  XNOR2_X2 U18911 ( .A(n18901), .B(n18559), .ZN(n18895) );
  INV_X4 U18912 ( .A(n18895), .ZN(n18560) );
  NAND2_X2 U18913 ( .A1(n13490), .A2(n18560), .ZN(n18585) );
  NAND2_X2 U18914 ( .A1(n13492), .A2(n18563), .ZN(n18584) );
  INV_X4 U18915 ( .A(n18564), .ZN(n18565) );
  NAND2_X2 U18916 ( .A1(n18565), .A2(n13208), .ZN(n18568) );
  NAND2_X2 U18917 ( .A1(n18566), .A2(DMEM_BUS_OUT[18]), .ZN(n18567) );
  OAI211_X2 U18918 ( .C1(n18570), .C2(n18569), .A(n18568), .B(n18567), .ZN(
        n18571) );
  NAND2_X2 U18919 ( .A1(n18571), .A2(n18901), .ZN(n18572) );
  NAND2_X2 U18920 ( .A1(DMEM_BUS_OUT[18]), .A2(net231325), .ZN(n18576) );
  INV_X4 U18921 ( .A(n18577), .ZN(n18578) );
  NOR2_X4 U18922 ( .A1(n18578), .A2(n13207), .ZN(n18579) );
  AOI211_X4 U18923 ( .C1(n19118), .C2(n18581), .A(n18580), .B(n18579), .ZN(
        n18582) );
  NAND4_X2 U18924 ( .A1(n18585), .A2(n18584), .A3(n18583), .A4(n18582), .ZN(
        n7752) );
  NAND2_X2 U18926 ( .A1(n18589), .A2(n18870), .ZN(n18591) );
  NAND2_X2 U18927 ( .A1(n18590), .A2(n18591), .ZN(n18593) );
  NAND2_X2 U18928 ( .A1(n18592), .A2(n18591), .ZN(n18596) );
  NAND2_X2 U18929 ( .A1(n18593), .A2(n18596), .ZN(n18606) );
  INV_X4 U18930 ( .A(n18604), .ZN(n18600) );
  INV_X4 U18931 ( .A(n18596), .ZN(n18598) );
  OAI21_X4 U18932 ( .B1(n18598), .B2(n18597), .A(n18606), .ZN(n18603) );
  INV_X4 U18933 ( .A(n18603), .ZN(n18599) );
  NOR3_X4 U18934 ( .A1(n18600), .A2(n18612), .A3(n18599), .ZN(n18609) );
  INV_X4 U18935 ( .A(n18601), .ZN(n18608) );
  INV_X4 U18936 ( .A(n18602), .ZN(n18605) );
  NAND2_X2 U18937 ( .A1(n18604), .A2(n18603), .ZN(n18616) );
  AOI21_X4 U18938 ( .B1(n18609), .B2(n18608), .A(n18607), .ZN(n18617) );
  NAND2_X2 U18939 ( .A1(n18617), .A2(n18610), .ZN(n18619) );
  INV_X4 U18940 ( .A(n18611), .ZN(n18614) );
  INV_X4 U18941 ( .A(n18612), .ZN(n18613) );
  NAND2_X2 U18942 ( .A1(n18614), .A2(n18613), .ZN(n18615) );
  NAND2_X2 U18943 ( .A1(n18617), .A2(n12965), .ZN(n18618) );
  OAI21_X4 U18944 ( .B1(n18620), .B2(n18619), .A(n18618), .ZN(n18621) );
  XNOR2_X2 U18945 ( .A(n18621), .B(n11041), .ZN(n18622) );
  NAND2_X2 U18946 ( .A1(n13399), .A2(n18623), .ZN(n18660) );
  NAND2_X2 U18947 ( .A1(ID_EXEC_OUT[64]), .A2(n13403), .ZN(n18661) );
  NAND2_X2 U18948 ( .A1(n18660), .A2(n18661), .ZN(n18666) );
  INV_X4 U18949 ( .A(n18666), .ZN(n18649) );
  NAND2_X2 U18950 ( .A1(n13484), .A2(DMEM_BUS_OUT[0]), .ZN(n18626) );
  NAND2_X2 U18951 ( .A1(n18649), .A2(n18626), .ZN(n19067) );
  XNOR2_X2 U18952 ( .A(n19067), .B(n19068), .ZN(n19054) );
  INV_X4 U18953 ( .A(n19054), .ZN(n19070) );
  INV_X4 U18954 ( .A(n18629), .ZN(n18632) );
  NOR3_X4 U18955 ( .A1(n18633), .A2(n18632), .A3(n18631), .ZN(n18635) );
  INV_X4 U18956 ( .A(n18636), .ZN(n18638) );
  NAND2_X2 U18957 ( .A1(n18644), .A2(n18643), .ZN(n18646) );
  NAND2_X2 U18958 ( .A1(ID_EXEC_OUT[204]), .A2(n13216), .ZN(n18645) );
  OAI211_X2 U18959 ( .C1(n18647), .C2(n13214), .A(n18646), .B(n18645), .ZN(
        n18682) );
  INV_X4 U18960 ( .A(n6625), .ZN(n18648) );
  NAND2_X2 U18961 ( .A1(n6625), .A2(n13484), .ZN(n18652) );
  NAND2_X2 U18962 ( .A1(n13406), .A2(n18663), .ZN(n18673) );
  NAND2_X2 U18963 ( .A1(n18667), .A2(n18666), .ZN(n18672) );
  INV_X4 U18964 ( .A(n18668), .ZN(n18670) );
  NAND2_X2 U18965 ( .A1(n18670), .A2(n18669), .ZN(n18671) );
  OAI221_X2 U18966 ( .B1(n18680), .B2(n18679), .C1(n18678), .C2(n13211), .A(
        n18676), .ZN(n18681) );
  OAI211_X2 U18968 ( .C1(n12176), .C2(net231227), .A(n18685), .B(n6746), .ZN(
        n7761) );
  NAND2_X2 U18969 ( .A1(n13411), .A2(ID_EXEC_OUT[191]), .ZN(n18689) );
  NAND2_X2 U18970 ( .A1(DMEM_BUS_OUT[63]), .A2(net231319), .ZN(n18688) );
  NAND2_X2 U18971 ( .A1(n13413), .A2(DMEM_BUS_OUT[31]), .ZN(n18687) );
  NAND2_X2 U18972 ( .A1(n13416), .A2(MEM_WB_OUT[68]), .ZN(n18686) );
  NAND4_X2 U18973 ( .A1(n18689), .A2(n18688), .A3(n18687), .A4(n18686), .ZN(
        n7826) );
  OAI22_X2 U18974 ( .A1(n13420), .A2(n12824), .B1(n13418), .B2(n12079), .ZN(
        n18696) );
  OAI22_X2 U18975 ( .A1(n13423), .A2(n12919), .B1(n13422), .B2(n12766), .ZN(
        n18695) );
  NAND2_X2 U18976 ( .A1(REG_FILE_reg_out_24__31_), .A2(n13428), .ZN(n18693) );
  NAND2_X2 U18977 ( .A1(REG_FILE_reg_out_18__31_), .A2(n13433), .ZN(n18692) );
  NAND2_X2 U18978 ( .A1(REG_FILE_reg_out_17__31_), .A2(n13434), .ZN(n18691) );
  AOI22_X2 U18979 ( .A1(REG_FILE_reg_out_25__31_), .A2(n13439), .B1(
        REG_FILE_reg_out_26__31_), .B2(n13441), .ZN(n18710) );
  OAI22_X2 U18980 ( .A1(n11430), .A2(n13444), .B1(n10530), .B2(n13443), .ZN(
        n18704) );
  OAI22_X2 U18981 ( .A1(n10461), .A2(n13190), .B1(n12177), .B2(n18699), .ZN(
        n18703) );
  OAI22_X2 U18982 ( .A1(n11846), .A2(n13192), .B1(n12298), .B2(n13193), .ZN(
        n18702) );
  NAND4_X2 U18983 ( .A1(n18711), .A2(n18710), .A3(n18709), .A4(n18708), .ZN(
        n18744) );
  NAND2_X2 U18984 ( .A1(n13455), .A2(REG_FILE_reg_out_12__31_), .ZN(n18724) );
  AOI22_X2 U18985 ( .A1(n13464), .A2(REG_FILE_reg_out_0__31_), .B1(
        REG_FILE_reg_out_15__31_), .B2(n13466), .ZN(n18722) );
  NAND4_X2 U18986 ( .A1(n18725), .A2(n18724), .A3(n18723), .A4(n18722), .ZN(
        n18743) );
  NAND4_X2 U18987 ( .A1(n18741), .A2(n18740), .A3(n18739), .A4(n18738), .ZN(
        n18742) );
  NOR3_X4 U18988 ( .A1(n18744), .A2(n18743), .A3(n18742), .ZN(n18746) );
  OAI222_X2 U18989 ( .A1(n18746), .A2(n13476), .B1(n12275), .B2(net231223), 
        .C1(n12023), .C2(n13206), .ZN(n7828) );
  OAI22_X2 U18990 ( .A1(n11537), .A2(net231259), .B1(net230377), .B2(n18746), 
        .ZN(n7829) );
  OAI22_X2 U18991 ( .A1(n11109), .A2(net231259), .B1(net230377), .B2(net239557), .ZN(n7831) );
  OAI22_X2 U18992 ( .A1(net231251), .A2(net239557), .B1(n11111), .B2(net230383), .ZN(n7832) );
  OAI22_X2 U18993 ( .A1(n11111), .A2(net231259), .B1(n12312), .B2(n13481), 
        .ZN(n7833) );
  NAND2_X2 U18994 ( .A1(net231317), .A2(EXEC_MEM_OUT_140), .ZN(n18750) );
  MUX2_X2 U18995 ( .A(EXEC_STAGE_imm26_32[31]), .B(EXEC_STAGE_imm16_32[31]), 
        .S(n10140), .Z(n18747) );
  OAI22_X2 U18996 ( .A1(net231251), .A2(n18753), .B1(n10824), .B2(net230383), 
        .ZN(n7839) );
  NAND2_X2 U18997 ( .A1(n18755), .A2(n18754), .ZN(n18758) );
  NAND2_X2 U18998 ( .A1(n18758), .A2(n18757), .ZN(n18761) );
  NOR4_X2 U18999 ( .A1(n18761), .A2(n18760), .A3(n5478), .A4(n18759), .ZN(
        n18763) );
  NAND2_X2 U19000 ( .A1(n13218), .A2(net231325), .ZN(n18762) );
  MUX2_X2 U19001 ( .A(DMEM_BUS_OUT[66]), .B(n13148), .S(net231291), .Z(n7844)
         );
  MUX2_X2 U19002 ( .A(DMEM_BUS_OUT[65]), .B(n13154), .S(net231291), .Z(n7847)
         );
  NAND2_X2 U19003 ( .A1(net231319), .A2(DSize_ex_out_0_), .ZN(n18764) );
  NAND2_X2 U19004 ( .A1(n18765), .A2(n18764), .ZN(n7849) );
  OAI211_X2 U19005 ( .C1(n11102), .C2(net231227), .A(n18846), .B(n12219), .ZN(
        n7852) );
  MUX2_X2 U19006 ( .A(DMEM_BUS_IN[26]), .B(MEM_WB_OUT[95]), .S(net231291), .Z(
        n7853) );
  MUX2_X2 U19007 ( .A(DMEM_BUS_IN[25]), .B(MEM_WB_OUT[94]), .S(net231291), .Z(
        n7854) );
  MUX2_X2 U19008 ( .A(DMEM_BUS_IN[24]), .B(MEM_WB_OUT[93]), .S(net231291), .Z(
        n7855) );
  MUX2_X2 U19009 ( .A(DMEM_BUS_IN[23]), .B(MEM_WB_OUT[92]), .S(net231291), .Z(
        n7856) );
  MUX2_X2 U19010 ( .A(DMEM_BUS_IN[22]), .B(MEM_WB_OUT[91]), .S(net231291), .Z(
        n7857) );
  MUX2_X2 U19011 ( .A(DMEM_BUS_IN[21]), .B(MEM_WB_OUT[90]), .S(net231291), .Z(
        n7858) );
  MUX2_X2 U19012 ( .A(DMEM_BUS_IN[20]), .B(MEM_WB_OUT[89]), .S(net231291), .Z(
        n7859) );
  MUX2_X2 U19013 ( .A(DMEM_BUS_IN[19]), .B(MEM_WB_OUT[88]), .S(net231291), .Z(
        n7860) );
  MUX2_X2 U19014 ( .A(DMEM_BUS_IN[18]), .B(MEM_WB_OUT[87]), .S(net231291), .Z(
        n7861) );
  MUX2_X2 U19015 ( .A(DMEM_BUS_IN[17]), .B(MEM_WB_OUT[86]), .S(net231291), .Z(
        n7862) );
  MUX2_X2 U19016 ( .A(DMEM_BUS_IN[16]), .B(MEM_WB_OUT[85]), .S(net231291), .Z(
        n7863) );
  INV_X4 U19017 ( .A(n10860), .ZN(n18770) );
  MUX2_X2 U19018 ( .A(n18770), .B(RegWrite_wb_out), .S(net231289), .Z(n7870)
         );
  OAI22_X2 U19019 ( .A1(n13477), .A2(n18772), .B1(net231263), .B2(n12017), 
        .ZN(n7873) );
  OAI22_X2 U19020 ( .A1(n12184), .A2(net231259), .B1(net230377), .B2(n18773), 
        .ZN(n7876) );
  MUX2_X2 U19021 ( .A(MEM_WB_REG_MEM_WB_REG_N78), .B(n13878), .S(net231289), 
        .Z(n7879) );
  OAI22_X2 U19022 ( .A1(n12183), .A2(net231261), .B1(net230377), .B2(n18776), 
        .ZN(n7887) );
  OAI22_X2 U19023 ( .A1(n12182), .A2(net231261), .B1(net230377), .B2(n18778), 
        .ZN(n7893) );
  MUX2_X2 U19024 ( .A(MEM_WB_REG_MEM_WB_REG_N76), .B(n13147), .S(net231289), 
        .Z(n7894) );
  OAI22_X2 U19025 ( .A1(net231251), .A2(n18779), .B1(n12064), .B2(net230383), 
        .ZN(n7895) );
  NAND2_X2 U19026 ( .A1(n18782), .A2(n18781), .ZN(n18784) );
  INV_X4 U19027 ( .A(n18785), .ZN(n7896) );
  OAI22_X2 U19028 ( .A1(n12020), .A2(net231261), .B1(n13480), .B2(n18786), 
        .ZN(n7897) );
  OAI22_X2 U19029 ( .A1(net231249), .A2(n12016), .B1(n19170), .B2(n13481), 
        .ZN(n7901) );
  NAND2_X2 U19030 ( .A1(n18787), .A2(net222642), .ZN(n7902) );
  OAI22_X2 U19031 ( .A1(net231249), .A2(n12134), .B1(n19164), .B2(n13481), 
        .ZN(n7906) );
  OAI22_X2 U19032 ( .A1(net231249), .A2(n18790), .B1(n19180), .B2(n13481), 
        .ZN(n7909) );
  NAND2_X2 U19033 ( .A1(ID_STAGE_imm16_aluA[22]), .A2(net230387), .ZN(n18793)
         );
  NAND2_X2 U19034 ( .A1(EXEC_STAGE_imm26_32[22]), .A2(net231325), .ZN(n18791)
         );
  NAND2_X2 U19035 ( .A1(n18793), .A2(n18791), .ZN(n7910) );
  NAND2_X2 U19036 ( .A1(EXEC_STAGE_imm16_32[22]), .A2(net231325), .ZN(n18792)
         );
  NAND2_X2 U19037 ( .A1(n18793), .A2(n18792), .ZN(n7911) );
  OAI22_X2 U19038 ( .A1(net231249), .A2(n18794), .B1(n19179), .B2(n13481), 
        .ZN(n7912) );
  OAI22_X2 U19039 ( .A1(net231249), .A2(n11983), .B1(n19178), .B2(n13481), 
        .ZN(n7915) );
  NAND2_X2 U19040 ( .A1(n2555), .A2(net222629), .ZN(n7919) );
  NAND2_X2 U19041 ( .A1(n2555), .A2(net222628), .ZN(n7920) );
  OAI22_X2 U19042 ( .A1(net231249), .A2(n12021), .B1(n19177), .B2(n13481), 
        .ZN(n7921) );
  NAND2_X2 U19043 ( .A1(EXEC_STAGE_imm16_32[19]), .A2(net231325), .ZN(n18795)
         );
  NAND2_X2 U19044 ( .A1(n2557), .A2(n18795), .ZN(n7925) );
  NAND2_X2 U19045 ( .A1(EXEC_STAGE_imm26_32[19]), .A2(net231325), .ZN(n18796)
         );
  NAND2_X2 U19046 ( .A1(n2557), .A2(n18796), .ZN(n7926) );
  OAI22_X2 U19047 ( .A1(n10806), .A2(net231261), .B1(n19176), .B2(n13481), 
        .ZN(n7927) );
  OAI22_X2 U19048 ( .A1(n11045), .A2(net231261), .B1(n19175), .B2(n13481), 
        .ZN(n7933) );
  NAND2_X2 U19049 ( .A1(EXEC_STAGE_imm16_32[17]), .A2(net231325), .ZN(n18797)
         );
  NAND2_X2 U19050 ( .A1(n2562), .A2(n18797), .ZN(n7937) );
  NAND2_X2 U19051 ( .A1(EXEC_STAGE_imm26_32[17]), .A2(net231325), .ZN(n18798)
         );
  NAND2_X2 U19052 ( .A1(n2562), .A2(n18798), .ZN(n7938) );
  OAI22_X2 U19053 ( .A1(n10807), .A2(net231261), .B1(n19174), .B2(n13481), 
        .ZN(n7939) );
  NAND2_X2 U19054 ( .A1(EXEC_STAGE_imm16_32[16]), .A2(net231325), .ZN(n18799)
         );
  NAND2_X2 U19055 ( .A1(n2564), .A2(n18799), .ZN(n7941) );
  OAI22_X2 U19056 ( .A1(n10816), .A2(net231261), .B1(n19173), .B2(n13481), 
        .ZN(n7945) );
  NAND2_X2 U19057 ( .A1(ID_EXEC_OUT[202]), .A2(net231325), .ZN(n18800) );
  NAND2_X2 U19058 ( .A1(n18801), .A2(n18800), .ZN(n7947) );
  INV_X4 U19059 ( .A(IMEM_BUS_IN[15]), .ZN(n18803) );
  NAND2_X2 U19060 ( .A1(n18805), .A2(n18804), .ZN(n7950) );
  INV_X4 U19061 ( .A(IMEM_BUS_IN[14]), .ZN(n18807) );
  OAI22_X2 U19062 ( .A1(n12214), .A2(net231261), .B1(net230377), .B2(n12953), 
        .ZN(n7952) );
  INV_X4 U19063 ( .A(IMEM_BUS_IN[13]), .ZN(n18809) );
  NAND2_X2 U19064 ( .A1(n13220), .A2(net231325), .ZN(n18808) );
  INV_X4 U19065 ( .A(IMEM_BUS_IN[12]), .ZN(n18812) );
  NAND2_X2 U19066 ( .A1(net231319), .A2(offset_26_id[6]), .ZN(n18811) );
  INV_X4 U19067 ( .A(IMEM_BUS_IN[11]), .ZN(n18815) );
  NAND2_X2 U19068 ( .A1(net231317), .A2(n18813), .ZN(n18814) );
  NAND2_X2 U19069 ( .A1(ID_EXEC_OUT[197]), .A2(net231325), .ZN(n18816) );
  NAND2_X2 U19070 ( .A1(n18817), .A2(n18816), .ZN(n7958) );
  INV_X4 U19071 ( .A(IMEM_BUS_IN[10]), .ZN(n18819) );
  NAND2_X2 U19072 ( .A1(n18821), .A2(n18820), .ZN(n7961) );
  INV_X4 U19073 ( .A(IMEM_BUS_IN[9]), .ZN(n18823) );
  NAND2_X2 U19074 ( .A1(n18825), .A2(n18824), .ZN(n7964) );
  INV_X4 U19075 ( .A(IMEM_BUS_IN[8]), .ZN(n18827) );
  OAI22_X2 U19076 ( .A1(net231249), .A2(n13138), .B1(n10828), .B2(net230373), 
        .ZN(n7967) );
  INV_X4 U19077 ( .A(IMEM_BUS_IN[7]), .ZN(n18828) );
  OAI22_X2 U19078 ( .A1(n10828), .A2(net231261), .B1(n13481), .B2(n18828), 
        .ZN(n7968) );
  OAI22_X2 U19079 ( .A1(net231249), .A2(n18829), .B1(n10360), .B2(net230383), 
        .ZN(n7970) );
  INV_X4 U19080 ( .A(IMEM_BUS_IN[6]), .ZN(n18831) );
  NAND2_X2 U19081 ( .A1(net231317), .A2(offset_26_id[0]), .ZN(n18830) );
  OAI22_X2 U19082 ( .A1(n12029), .A2(net231259), .B1(n19172), .B2(n13481), 
        .ZN(n7972) );
  OAI22_X2 U19083 ( .A1(net231247), .A2(n12027), .B1(n19187), .B2(n13480), 
        .ZN(n7975) );
  OAI22_X2 U19084 ( .A1(net231249), .A2(n12129), .B1(n19171), .B2(n13481), 
        .ZN(n7976) );
  INV_X4 U19085 ( .A(IMEM_BUS_IN[1]), .ZN(n18834) );
  NAND2_X2 U19086 ( .A1(net231317), .A2(n13221), .ZN(n18833) );
  OAI22_X2 U19087 ( .A1(n12039), .A2(net231261), .B1(n19186), .B2(n13481), 
        .ZN(n7980) );
  NAND2_X2 U19088 ( .A1(net230387), .A2(ID_STAGE_imm16_aluA[28]), .ZN(n18837)
         );
  NAND2_X2 U19089 ( .A1(EXEC_STAGE_imm26_32[28]), .A2(net231315), .ZN(n18835)
         );
  NAND2_X2 U19090 ( .A1(n18837), .A2(n18835), .ZN(n7981) );
  NAND2_X2 U19091 ( .A1(n18837), .A2(n18836), .ZN(n7982) );
  OAI22_X2 U19092 ( .A1(n10840), .A2(net231261), .B1(n19185), .B2(n13481), 
        .ZN(n7983) );
  OAI22_X2 U19093 ( .A1(n10838), .A2(net231261), .B1(n19184), .B2(n13481), 
        .ZN(n7986) );
  NAND2_X2 U19094 ( .A1(net230393), .A2(ID_STAGE_imm16_aluA[26]), .ZN(n18840)
         );
  NAND2_X2 U19095 ( .A1(EXEC_STAGE_imm26_32[26]), .A2(net231315), .ZN(n18838)
         );
  NAND2_X2 U19096 ( .A1(n18840), .A2(n18838), .ZN(n7987) );
  NAND2_X2 U19097 ( .A1(EXEC_STAGE_imm16_32[26]), .A2(net231315), .ZN(n18839)
         );
  NAND2_X2 U19098 ( .A1(n18840), .A2(n18839), .ZN(n7988) );
  OAI22_X2 U19099 ( .A1(n10240), .A2(net231261), .B1(n19183), .B2(n13480), 
        .ZN(n7989) );
  OAI22_X2 U19100 ( .A1(n12300), .A2(net231263), .B1(n19182), .B2(n13481), 
        .ZN(n7992) );
  NAND2_X2 U19101 ( .A1(ID_STAGE_imm16_aluA[24]), .A2(net230387), .ZN(n18843)
         );
  NAND2_X2 U19102 ( .A1(EXEC_STAGE_imm26_32[24]), .A2(net231315), .ZN(n18841)
         );
  NAND2_X2 U19103 ( .A1(n18843), .A2(n18841), .ZN(n7993) );
  NAND2_X2 U19104 ( .A1(EXEC_STAGE_imm16_32[24]), .A2(net231315), .ZN(n18842)
         );
  NAND2_X2 U19105 ( .A1(n18843), .A2(n18842), .ZN(n7994) );
  OAI22_X2 U19106 ( .A1(net231249), .A2(n12028), .B1(n19181), .B2(n13480), 
        .ZN(n7995) );
  NAND2_X2 U19107 ( .A1(ID_EXEC_OUT[148]), .A2(net231315), .ZN(n18844) );
  NAND2_X2 U19108 ( .A1(n13476), .A2(n18844), .ZN(n7996) );
  OAI22_X2 U19109 ( .A1(net231247), .A2(n12023), .B1(n19188), .B2(n13481), 
        .ZN(n7999) );
  MUX2_X2 U19110 ( .A(DMEM_BUS_IN[27]), .B(MEM_WB_OUT[96]), .S(net231289), .Z(
        n8012) );
  MUX2_X2 U19111 ( .A(DMEM_BUS_IN[28]), .B(MEM_WB_OUT[97]), .S(net231289), .Z(
        n8013) );
  MUX2_X2 U19112 ( .A(DMEM_BUS_IN[29]), .B(MEM_WB_OUT[98]), .S(net231289), .Z(
        n8014) );
  MUX2_X2 U19113 ( .A(DMEM_BUS_IN[30]), .B(MEM_WB_OUT[99]), .S(net231289), .Z(
        n8015) );
  MUX2_X2 U19114 ( .A(DMEM_BUS_IN[31]), .B(MEM_WB_OUT[100]), .S(net231291), 
        .Z(n8016) );
  NAND2_X2 U19115 ( .A1(net231221), .A2(n18846), .ZN(n8017) );
  NAND2_X2 U19116 ( .A1(n18879), .A2(n18990), .ZN(n18848) );
  NAND2_X2 U19117 ( .A1(n18989), .A2(n18976), .ZN(n18847) );
  NAND2_X2 U19118 ( .A1(n19025), .A2(n19031), .ZN(n18850) );
  NAND2_X2 U19119 ( .A1(n18851), .A2(n19001), .ZN(n18919) );
  INV_X4 U19120 ( .A(n18917), .ZN(n18881) );
  XNOR2_X2 U19121 ( .A(n13151), .B(n19105), .ZN(n19111) );
  NAND4_X2 U19122 ( .A1(n19035), .A2(n19040), .A3(n19044), .A4(n19048), .ZN(
        n18855) );
  NOR3_X4 U19123 ( .A1(n18857), .A2(n18856), .A3(n18855), .ZN(n19058) );
  XNOR2_X2 U19124 ( .A(n18858), .B(n18967), .ZN(n18963) );
  XNOR2_X2 U19125 ( .A(n18925), .B(n18859), .ZN(n18968) );
  XNOR2_X2 U19126 ( .A(n13163), .B(n18860), .ZN(n18951) );
  INV_X4 U19127 ( .A(n18866), .ZN(n18868) );
  NAND2_X2 U19128 ( .A1(n18868), .A2(n18867), .ZN(n19062) );
  INV_X4 U19129 ( .A(n18869), .ZN(n18871) );
  NAND2_X2 U19130 ( .A1(n18871), .A2(n18870), .ZN(n19064) );
  INV_X4 U19131 ( .A(n19064), .ZN(n19073) );
  NAND2_X2 U19132 ( .A1(n19047), .A2(n18872), .ZN(n18876) );
  NAND2_X2 U19133 ( .A1(n18874), .A2(n18873), .ZN(n18875) );
  OAI21_X4 U19134 ( .B1(n18877), .B2(n18876), .A(n18875), .ZN(n19078) );
  INV_X4 U19135 ( .A(n19076), .ZN(n19065) );
  NAND2_X2 U19136 ( .A1(n19064), .A2(n19065), .ZN(n19051) );
  OAI21_X4 U19137 ( .B1(n19073), .B2(n19078), .A(n19051), .ZN(n19049) );
  INV_X4 U19138 ( .A(n18879), .ZN(n18880) );
  NOR2_X4 U19139 ( .A1(n18881), .A2(n18880), .ZN(n18910) );
  OAI21_X4 U19140 ( .B1(n15732), .B2(n18890), .A(n18889), .ZN(n18892) );
  INV_X4 U19141 ( .A(n18896), .ZN(n18898) );
  NAND2_X2 U19142 ( .A1(n18898), .A2(n18897), .ZN(n18913) );
  INV_X4 U19143 ( .A(n18907), .ZN(n18908) );
  NAND2_X2 U19144 ( .A1(n18908), .A2(net222497), .ZN(n18909) );
  INV_X4 U19145 ( .A(n18909), .ZN(n18993) );
  INV_X4 U19146 ( .A(n18911), .ZN(n18915) );
  NAND2_X2 U19147 ( .A1(n18923), .A2(n18922), .ZN(n18975) );
  NAND2_X2 U19148 ( .A1(n13155), .A2(n18926), .ZN(n18937) );
  INV_X4 U19149 ( .A(n13156), .ZN(n18936) );
  INV_X4 U19150 ( .A(n18931), .ZN(n18932) );
  AOI21_X4 U19151 ( .B1(n18934), .B2(n18933), .A(n18932), .ZN(n18935) );
  NOR3_X4 U19152 ( .A1(n18937), .A2(n18936), .A3(n18935), .ZN(n18941) );
  NAND2_X2 U19153 ( .A1(n19100), .A2(n13159), .ZN(n18940) );
  NAND2_X2 U19154 ( .A1(n18943), .A2(n13161), .ZN(n18946) );
  NAND2_X2 U19155 ( .A1(n18946), .A2(n18950), .ZN(n18947) );
  INV_X4 U19156 ( .A(n18950), .ZN(n18952) );
  AOI21_X4 U19157 ( .B1(n18971), .B2(n18970), .A(n18969), .ZN(n18972) );
  INV_X4 U19158 ( .A(n18975), .ZN(n18977) );
  NAND2_X2 U19159 ( .A1(n18981), .A2(n18980), .ZN(n18982) );
  INV_X4 U19160 ( .A(n18990), .ZN(n18997) );
  NOR2_X4 U19161 ( .A1(n18994), .A2(n18993), .ZN(n18996) );
  INV_X4 U19162 ( .A(n18999), .ZN(n19002) );
  NAND3_X2 U19163 ( .A1(n19002), .A2(n19001), .A3(n19000), .ZN(n19007) );
  INV_X4 U19164 ( .A(n19003), .ZN(n19005) );
  NAND2_X2 U19165 ( .A1(n19005), .A2(n19004), .ZN(n19006) );
  NAND2_X2 U19166 ( .A1(n19007), .A2(n19006), .ZN(n19008) );
  AOI21_X4 U19167 ( .B1(n19009), .B2(n19010), .A(n19008), .ZN(n19022) );
  INV_X4 U19168 ( .A(n19011), .ZN(n19021) );
  INV_X4 U19169 ( .A(n19012), .ZN(n19014) );
  NAND2_X2 U19170 ( .A1(n19014), .A2(n19013), .ZN(n19024) );
  INV_X4 U19171 ( .A(n19024), .ZN(n19019) );
  INV_X4 U19172 ( .A(n19015), .ZN(n19017) );
  NOR2_X4 U19173 ( .A1(n19019), .A2(n19018), .ZN(n19020) );
  OAI21_X4 U19174 ( .B1(n19022), .B2(n19021), .A(n19020), .ZN(n19027) );
  INV_X4 U19175 ( .A(n19028), .ZN(n19030) );
  NAND2_X2 U19176 ( .A1(n19030), .A2(n19029), .ZN(n19033) );
  INV_X4 U19177 ( .A(n19031), .ZN(n19032) );
  AOI21_X4 U19178 ( .B1(n19034), .B2(n19033), .A(n19032), .ZN(n19036) );
  NAND2_X2 U19179 ( .A1(n19039), .A2(n19038), .ZN(n19042) );
  INV_X4 U19180 ( .A(n19040), .ZN(n19041) );
  AOI21_X4 U19181 ( .B1(n19043), .B2(n19042), .A(n19041), .ZN(n19045) );
  OAI21_X4 U19182 ( .B1(n19045), .B2(net222353), .A(n19044), .ZN(n19063) );
  NAND3_X4 U19183 ( .A1(n19063), .A2(n19049), .A3(n19062), .ZN(n19046) );
  NAND2_X2 U19184 ( .A1(n19048), .A2(n19047), .ZN(n19061) );
  INV_X4 U19185 ( .A(n19049), .ZN(n19050) );
  AOI21_X4 U19186 ( .B1(n19051), .B2(n19077), .A(n19050), .ZN(n19052) );
  NOR2_X4 U19187 ( .A1(n19053), .A2(n19052), .ZN(n19055) );
  XNOR2_X2 U19188 ( .A(n19055), .B(n19070), .ZN(n19086) );
  INV_X4 U19189 ( .A(n19086), .ZN(n19056) );
  INV_X4 U19190 ( .A(n19061), .ZN(n19077) );
  AOI21_X4 U19191 ( .B1(n19074), .B2(n19077), .A(n19078), .ZN(n19066) );
  OAI21_X4 U19192 ( .B1(n19066), .B2(n19065), .A(n19064), .ZN(n19085) );
  INV_X4 U19193 ( .A(n19067), .ZN(n19069) );
  NAND2_X2 U19194 ( .A1(n19069), .A2(n19068), .ZN(n19071) );
  NAND2_X2 U19195 ( .A1(n19071), .A2(n19070), .ZN(n19075) );
  INV_X4 U19196 ( .A(n19075), .ZN(n19083) );
  INV_X4 U19197 ( .A(n19071), .ZN(n19072) );
  NOR2_X4 U19198 ( .A1(n19073), .A2(n19072), .ZN(n19082) );
  INV_X4 U19199 ( .A(n13074), .ZN(n19081) );
  NAND2_X2 U19200 ( .A1(n12132), .A2(n19077), .ZN(n19080) );
  NAND2_X2 U19201 ( .A1(n12132), .A2(n19078), .ZN(n19079) );
  XNOR2_X2 U19202 ( .A(n19085), .B(n19084), .ZN(n19087) );
  XNOR2_X2 U19203 ( .A(n19087), .B(n19086), .ZN(n19136) );
  INV_X4 U19204 ( .A(n19090), .ZN(n19094) );
  NAND2_X2 U19205 ( .A1(n13487), .A2(n19096), .ZN(n19098) );
  OAI221_X2 U19206 ( .B1(n19102), .B2(n19101), .C1(n19100), .C2(n19099), .A(
        n19098), .ZN(n19103) );
  NAND2_X2 U19207 ( .A1(n13210), .A2(n19103), .ZN(n19122) );
  XNOR2_X2 U19208 ( .A(n19109), .B(n13493), .ZN(n19113) );
  NOR2_X4 U19209 ( .A1(n19111), .A2(n19110), .ZN(n19112) );
  NAND4_X2 U19210 ( .A1(n19122), .A2(n19121), .A3(n19120), .A4(n19119), .ZN(
        n19123) );
  INV_X4 U19211 ( .A(n19123), .ZN(n19139) );
  XNOR2_X2 U19212 ( .A(n13218), .B(ID_EXEC_OUT[157]), .ZN(n19126) );
  NAND2_X2 U19213 ( .A1(n19139), .A2(n19127), .ZN(n19134) );
  AOI21_X4 U19214 ( .B1(n19132), .B2(n19133), .A(n19131), .ZN(n19148) );
  INV_X4 U19215 ( .A(n19134), .ZN(n19135) );
  NAND2_X2 U19216 ( .A1(n19135), .A2(n11915), .ZN(n19144) );
  NAND2_X2 U19217 ( .A1(n19139), .A2(n19138), .ZN(n19143) );
  INV_X4 U19218 ( .A(n19144), .ZN(n19141) );
  INV_X4 U19219 ( .A(IMEM_BUS_IN[2]), .ZN(n19170) );
  INV_X4 U19220 ( .A(IMEM_BUS_IN[3]), .ZN(n19171) );
  INV_X4 U19221 ( .A(IMEM_BUS_IN[4]), .ZN(n19172) );
  INV_X4 U19222 ( .A(IMEM_BUS_IN[16]), .ZN(n19173) );
  INV_X4 U19223 ( .A(IMEM_BUS_IN[17]), .ZN(n19174) );
  INV_X4 U19224 ( .A(IMEM_BUS_IN[18]), .ZN(n19175) );
  INV_X4 U19225 ( .A(IMEM_BUS_IN[19]), .ZN(n19176) );
  INV_X4 U19226 ( .A(IMEM_BUS_IN[20]), .ZN(n19177) );
  INV_X4 U19227 ( .A(IMEM_BUS_IN[21]), .ZN(n19178) );
  INV_X4 U19228 ( .A(IMEM_BUS_IN[22]), .ZN(n19179) );
  INV_X4 U19229 ( .A(IMEM_BUS_IN[23]), .ZN(n19180) );
  INV_X4 U19230 ( .A(IMEM_BUS_IN[24]), .ZN(n19181) );
  INV_X4 U19231 ( .A(IMEM_BUS_IN[25]), .ZN(n19182) );
  INV_X4 U19232 ( .A(IMEM_BUS_IN[26]), .ZN(n19183) );
  INV_X4 U19233 ( .A(IMEM_BUS_IN[27]), .ZN(n19184) );
  INV_X4 U19234 ( .A(IMEM_BUS_IN[28]), .ZN(n19185) );
  INV_X4 U19235 ( .A(IMEM_BUS_IN[29]), .ZN(n19186) );
  INV_X4 U19236 ( .A(IMEM_BUS_IN[30]), .ZN(n19187) );
  INV_X4 U19237 ( .A(IMEM_BUS_IN[31]), .ZN(n19188) );
  INV_X4 U19238 ( .A(n7286), .ZN(n19189) );
  INV_X4 U19239 ( .A(n7288), .ZN(n19190) );
  INV_X4 U19240 ( .A(n7284), .ZN(n19191) );
  INV_X4 U19241 ( .A(n7283), .ZN(n19192) );
  INV_X4 U19242 ( .A(n6815), .ZN(n19193) );
  INV_X4 U19243 ( .A(n6814), .ZN(n19194) );
  INV_X4 U19244 ( .A(n6813), .ZN(n19195) );
  INV_X4 U19245 ( .A(n6812), .ZN(n19196) );
  INV_X4 U19246 ( .A(n6811), .ZN(n19197) );
  INV_X4 U19247 ( .A(n6810), .ZN(n19198) );
  INV_X4 U19248 ( .A(n6809), .ZN(n19199) );
  INV_X4 U19249 ( .A(n6808), .ZN(n19200) );
  INV_X4 U19250 ( .A(n6807), .ZN(n19201) );
  INV_X4 U19251 ( .A(n6806), .ZN(n19202) );
  INV_X4 U19252 ( .A(n6805), .ZN(n19203) );
  INV_X4 U19253 ( .A(n6804), .ZN(n19204) );
  INV_X4 U19254 ( .A(n6803), .ZN(n19205) );
  INV_X4 U19255 ( .A(n6802), .ZN(n19206) );
  INV_X4 U19256 ( .A(n6801), .ZN(n19207) );
  INV_X4 U19257 ( .A(n6800), .ZN(n19208) );
  INV_X4 U19258 ( .A(n6799), .ZN(n19209) );
  INV_X4 U19259 ( .A(n6798), .ZN(n19210) );
  INV_X4 U19260 ( .A(n6797), .ZN(n19211) );
  INV_X4 U19261 ( .A(n6796), .ZN(n19212) );
  INV_X4 U19262 ( .A(n6795), .ZN(n19213) );
  INV_X4 U19263 ( .A(n6794), .ZN(n19214) );
  INV_X4 U19264 ( .A(n6793), .ZN(n19215) );
  INV_X4 U19265 ( .A(n6792), .ZN(n19216) );
  INV_X4 U19266 ( .A(n6791), .ZN(n19217) );
  INV_X4 U19267 ( .A(n6789), .ZN(n19218) );
  INV_X4 U19268 ( .A(n6788), .ZN(n19219) );
  INV_X4 U19269 ( .A(n6787), .ZN(n19220) );
  INV_X4 U19270 ( .A(n6786), .ZN(n19221) );
  INV_X4 U19271 ( .A(n6785), .ZN(n19222) );
  INV_X4 U19272 ( .A(n6784), .ZN(n19223) );
  INV_X4 U19273 ( .A(n6783), .ZN(n19224) );
  INV_X4 U19274 ( .A(n1271), .ZN(n19225) );
  INV_X4 U19275 ( .A(n1290), .ZN(n19226) );
  INV_X4 U19276 ( .A(n1291), .ZN(n19227) );
  INV_X4 U19277 ( .A(n1292), .ZN(n19228) );
  INV_X4 U19278 ( .A(n1293), .ZN(n19229) );
  INV_X4 U19279 ( .A(n1294), .ZN(n19230) );
  INV_X4 U19280 ( .A(n1295), .ZN(n19231) );
  INV_X4 U19281 ( .A(n1298), .ZN(n19232) );
  INV_X4 U19282 ( .A(n1301), .ZN(n19233) );
  INV_X4 U19283 ( .A(n1306), .ZN(n19234) );
  INV_X4 U19284 ( .A(n1307), .ZN(n19235) );
  INV_X4 U19285 ( .A(n1308), .ZN(n19236) );
  INV_X4 U19286 ( .A(n1313), .ZN(n19237) );
  INV_X4 U19287 ( .A(n1316), .ZN(n19238) );
  INV_X4 U19288 ( .A(n1317), .ZN(n19239) );
  INV_X4 U19289 ( .A(n1320), .ZN(n19240) );
  INV_X4 U19290 ( .A(n1338), .ZN(n19241) );
  INV_X4 U19291 ( .A(n1345), .ZN(n19242) );
  INV_X4 U19292 ( .A(n1348), .ZN(n19243) );
  INV_X4 U19293 ( .A(n1351), .ZN(n19244) );
  INV_X4 U19294 ( .A(n1358), .ZN(n19245) );
  INV_X4 U19295 ( .A(n1433), .ZN(n19246) );
  INV_X4 U19296 ( .A(n1434), .ZN(n19247) );
  INV_X4 U19297 ( .A(n1435), .ZN(n19248) );
  INV_X4 U19298 ( .A(n1436), .ZN(n19249) );
  INV_X4 U19299 ( .A(n1437), .ZN(n19250) );
  INV_X4 U19300 ( .A(n1440), .ZN(n19251) );
  INV_X4 U19301 ( .A(n1441), .ZN(n19252) );
  INV_X4 U19302 ( .A(n1442), .ZN(n19253) );
  INV_X4 U19303 ( .A(n1443), .ZN(n19254) );
  INV_X4 U19304 ( .A(n1444), .ZN(n19255) );
  INV_X4 U19305 ( .A(n1445), .ZN(n19256) );
  INV_X4 U19306 ( .A(n1446), .ZN(n19257) );
  INV_X4 U19307 ( .A(n1447), .ZN(n19258) );
  INV_X4 U19308 ( .A(n1448), .ZN(n19259) );
  INV_X4 U19309 ( .A(n1449), .ZN(n19260) );
  INV_X4 U19310 ( .A(n1452), .ZN(n19261) );
  INV_X4 U19311 ( .A(n1453), .ZN(n19262) );
  INV_X4 U19312 ( .A(n1454), .ZN(n19263) );
  INV_X4 U19313 ( .A(n1455), .ZN(n19264) );
  INV_X4 U19314 ( .A(n1456), .ZN(n19265) );
  INV_X4 U19315 ( .A(n1457), .ZN(n19266) );
  INV_X4 U19316 ( .A(n1458), .ZN(n19267) );
  INV_X4 U19317 ( .A(n1459), .ZN(n19268) );
  INV_X4 U19318 ( .A(n1460), .ZN(n19269) );
  INV_X4 U19319 ( .A(n1461), .ZN(n19270) );
  INV_X4 U19320 ( .A(n1464), .ZN(n19271) );
  INV_X4 U19321 ( .A(n1465), .ZN(n19272) );
  INV_X4 U19322 ( .A(n1466), .ZN(n19273) );
  INV_X4 U19323 ( .A(n1467), .ZN(n19274) );
  INV_X4 U19324 ( .A(n1468), .ZN(n19275) );
  INV_X4 U19325 ( .A(n1469), .ZN(n19276) );
  INV_X4 U19326 ( .A(n1470), .ZN(n19277) );
  INV_X4 U19327 ( .A(n1487), .ZN(n19278) );
  INV_X4 U19328 ( .A(n3210), .ZN(n19279) );
  INV_X4 U19329 ( .A(n4674), .ZN(n19280) );
  INV_X4 U19330 ( .A(n5586), .ZN(n19281) );
  INV_X4 U19331 ( .A(n5590), .ZN(n19282) );
  INV_X4 U19332 ( .A(n5595), .ZN(n19283) );
  INV_X4 U19333 ( .A(n5597), .ZN(n19284) );
  INV_X4 U19334 ( .A(n5603), .ZN(n19285) );
  INV_X4 U19335 ( .A(n5608), .ZN(n19286) );
  INV_X4 U19336 ( .A(n5612), .ZN(n19287) );
  INV_X4 U19337 ( .A(n5614), .ZN(n19288) );
  INV_X4 U19338 ( .A(n6744), .ZN(n19289) );
  INV_X4 U19339 ( .A(n6769), .ZN(n19290) );
  INV_X4 U19340 ( .A(n6790), .ZN(n19291) );
  INV_X4 U19341 ( .A(n6816), .ZN(net139967) );
  INV_X4 U19342 ( .A(n5606), .ZN(n19292) );
  INV_X4 U19343 ( .A(n5588), .ZN(n19293) );
  INV_X4 U19344 ( .A(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[26]), .ZN(n19294)
         );
  INV_X4 U19347 ( .A(n5520), .ZN(n19301) );
  INV_X4 U19348 ( .A(n5764), .ZN(n19302) );
  INV_X4 U19349 ( .A(n5724), .ZN(n19303) );
  INV_X4 U19350 ( .A(n5718), .ZN(n19304) );
  INV_X4 U19351 ( .A(n5680), .ZN(n19305) );
  INV_X4 U19352 ( .A(n5676), .ZN(n19306) );
  INV_X4 U19353 ( .A(n5663), .ZN(n19307) );
  INV_X4 U19354 ( .A(n5770), .ZN(n19308) );
  INV_X4 U19355 ( .A(n5669), .ZN(n19309) );
  INV_X4 U19356 ( .A(MEM_WB_REG_MEM_WB_REG_N148), .ZN(n19310) );
  INV_X4 U19357 ( .A(MEM_WB_REG_MEM_WB_REG_N145), .ZN(n19316) );
  INV_X4 U19358 ( .A(EXEC_MEM_IN[105]), .ZN(n19318) );
  INV_X4 U19359 ( .A(nextPC_ex_out[29]), .ZN(net137343) );
  INV_X4 U19361 ( .A(nextPC_ex_out[26]), .ZN(net137303) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_33_ ( .D(n7977), .CK(clk), .RN(reset), 
        .Q(n13221), .QN(n12555) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_44_ ( .D(n7955), .CK(clk), .RN(reset), 
        .Q(offset_26_id[6]), .QN(n11922) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[25]), .QN(n12689) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_56_ ( .D(n7995), .CK(clk), .RN(n13924), 
        .Q(ID_STAGE_imm16_aluA[24]), .QN(n12028) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_54_ ( .D(n7912), .CK(clk), .RN(n13924), 
        .Q(ID_STAGE_imm16_aluA[22]), .QN(n18794) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_0_ ( .D(n7332), .CK(clk), .RN(n13904), 
        .QN(n15638) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_72_ ( .D(n8004), .CK(clk), .RN(n13931), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[19]), .QN(n19297) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_38_ ( .D(n7971), .CK(clk), .RN(n13923), 
        .Q(offset_26_id[0]), .QN(n10360) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_32_ ( .D(n7906), .CK(clk), .RN(n13923), 
        .Q(IF_ID_OUT[32]), .QN(n12134) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_63_ ( .D(n7999), .CK(clk), .RN(n13925), 
        .Q(ID_STAGE_imm16_aluA[31]), .QN(n12023) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_36_ ( .D(n7972), .CK(clk), .RN(n13923), 
        .Q(IF_ID_OUT[36]), .QN(n12029) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_62_ ( .D(n7975), .CK(clk), .RN(n13887), 
        .Q(ID_STAGE_imm16_aluA[30]), .QN(n12027) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_58_ ( .D(n7989), .CK(clk), .RN(n13924), 
        .Q(ID_STAGE_imm16_aluA[26]), .QN(n10240) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_59_ ( .D(n7986), .CK(clk), .RN(n13887), 
        .Q(ID_STAGE_imm16_aluA[27]), .QN(n10838) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_92_ ( .D(n7856), .CK(clk), .RN(n13932), 
        .Q(MEM_WB_OUT[92]), .QN(n11472) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_74_ ( .D(n8006), .CK(clk), .RN(n13931), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[21]), .QN(n19295) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_45_ ( .D(n7954), .CK(clk), .RN(reset), 
        .Q(n13220), .QN(n12953) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_99_ ( .D(n8015), .CK(clk), .RN(n13881), 
        .Q(MEM_WB_OUT[99]), .QN(n11556) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_95_ ( .D(n7853), .CK(clk), .RN(n13881), 
        .Q(MEM_WB_OUT[95]), .QN(n11557) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_70_ ( .D(n8002), .CK(clk), .RN(n13931), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[17]), .QN(n12033) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_71_ ( .D(n8003), .CK(clk), .RN(n13882), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[18]), .QN(n19298) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_69_ ( .D(n8001), .CK(clk), .RN(n13931), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[16]), .QN(n14122) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_34_ ( .D(n7901), .CK(clk), .RN(n13923), 
        .Q(IF_ID_OUT[34]), .QN(n12016) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_158_ ( .D(n7841), .CK(clk), .RN(n13914), 
        .Q(ID_EXEC_OUT[158]), .QN(n11913) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_35_ ( .D(n7976), .CK(clk), .RN(n13888), 
        .Q(IF_ID_OUT[35]), .QN(n12129) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_55_ ( .D(n7909), .CK(clk), .RN(n13887), 
        .Q(ID_STAGE_imm16_aluA[23]), .QN(n18790) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_19_ ( .D(n7573), .CK(clk), .RN(n13916), 
        .Q(nextPC_ex_out[19]), .QN(n10242) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[26]), .QN(n12552) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[27]), .QN(n15478) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[1]), .QN(n12034) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[0]), .QN(n12715) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[29]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_94_ ( .D(n7716), .CK(clk), .RN(
        reset), .Q(DMEM_BUS_OUT[25]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_88_ ( .D(n7634), .CK(clk), .RN(
        reset), .Q(DMEM_BUS_OUT[19]), .QN(n11965) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_35_ ( .D(n7882), .CK(clk), .RN(n13883), 
        .QN(n13128) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_202_ ( .D(n7947), .CK(clk), .RN(n13916), 
        .Q(ID_EXEC_OUT[202]), .QN(n13139) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_91_ ( .D(n7626), .CK(clk), .RN(
        n13912), .Q(DMEM_BUS_OUT[22]), .QN(n11982) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_80_ ( .D(n7403), .CK(clk), .RN(
        n13912), .Q(DMEM_BUS_OUT[11]) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_92_ ( .D(n7645), .CK(clk), .RN(
        n13925), .Q(DMEM_BUS_OUT[23]), .QN(n11969) );
  OAI21_X2 U10189 ( .B1(net225892), .B2(n11921), .A(n10117), .ZN(net225890) );
  NAND2_X1 U10201 ( .A1(n13492), .A2(n17980), .ZN(n18018) );
  AOI221_X4 U10205 ( .B1(net231271), .B2(EXEC_MEM_OUT_121), .C1(n19345), .C2(
        n10361), .A(n19346), .ZN(n19344) );
  INV_X32 U10206 ( .A(n19344), .ZN(n7433) );
  XOR2_X1 U10207 ( .A(net225892), .B(net225821), .Z(n19345) );
  AND2_X2 U10208 ( .A1(net231615), .A2(n19000), .ZN(n19346) );
  NAND2_X4 U10209 ( .A1(n18684), .A2(n18683), .ZN(n7756) );
  XOR2_X2 U10226 ( .A(n13145), .B(n13057), .Z(n15492) );
  INV_X8 U10239 ( .A(n16823), .ZN(n18885) );
  NAND2_X2 U10258 ( .A1(n13359), .A2(n18888), .ZN(n18274) );
  NAND3_X2 U10277 ( .A1(n14106), .A2(n14107), .A3(n14108), .ZN(n19347) );
  NAND3_X2 U10290 ( .A1(n14106), .A2(n14107), .A3(n14108), .ZN(n16810) );
  INV_X1 U10297 ( .A(n13113), .ZN(n19348) );
  INV_X8 U10299 ( .A(n15562), .ZN(n10113) );
  INV_X4 U10302 ( .A(net224850), .ZN(n19349) );
  INV_X2 U10315 ( .A(net224850), .ZN(net225162) );
  INV_X2 U10323 ( .A(net225207), .ZN(n10112) );
  NAND2_X1 U10324 ( .A1(net223666), .A2(net239761), .ZN(n19350) );
  BUF_X32 U10328 ( .A(net225453), .Z(n10109) );
  AOI21_X4 U10331 ( .B1(net227019), .B2(n11994), .A(net227020), .ZN(net227008)
         );
  NOR2_X4 U10351 ( .A1(n10131), .A2(net225162), .ZN(net227019) );
  OAI21_X4 U10352 ( .B1(net225201), .B2(net224713), .A(net225202), .ZN(n7494)
         );
  BUF_X32 U10413 ( .A(n12987), .Z(n19351) );
  NOR3_X4 U10478 ( .A1(n12315), .A2(n11097), .A3(n15412), .ZN(n19352) );
  INV_X4 U10495 ( .A(n19352), .ZN(n15437) );
  INV_X4 U10516 ( .A(n15412), .ZN(n15435) );
  NAND3_X2 U10641 ( .A1(n17993), .A2(n18629), .A3(n16794), .ZN(n19353) );
  AOI21_X4 U10671 ( .B1(n18654), .B2(DMEM_BUS_OUT[0]), .A(n18653), .ZN(n19354)
         );
  OAI221_X1 U10839 ( .B1(n19354), .B2(n18586), .C1(n12178), .C2(net231221), 
        .A(n6782), .ZN(n7754) );
  NAND3_X1 U11169 ( .A1(n5464), .A2(RegWrite_wb_out), .A3(n5463), .ZN(n15582)
         );
  NAND2_X1 U11226 ( .A1(n2536), .A2(RegWrite_wb_out), .ZN(n14977) );
  NOR2_X2 U11421 ( .A1(n14046), .A2(n14045), .ZN(n14047) );
  NAND2_X1 U12696 ( .A1(n17911), .A2(n16061), .ZN(n17912) );
  NAND2_X1 U12780 ( .A1(n13389), .A2(n19353), .ZN(n16801) );
  NAND2_X1 U12781 ( .A1(n13488), .A2(n17911), .ZN(n17521) );
  NAND2_X1 U12851 ( .A1(n13393), .A2(n19353), .ZN(n17850) );
  NAND3_X2 U13096 ( .A1(n17993), .A2(n18629), .A3(n16794), .ZN(n17911) );
  CLKBUF_X3 U13539 ( .A(net225452), .Z(n10141) );
  BUF_X8 U13630 ( .A(net227143), .Z(n10136) );
  NAND3_X4 U13739 ( .A1(n12987), .A2(IMEM_BUS_OUT[12]), .A3(IMEM_BUS_OUT[11]), 
        .ZN(n15412) );
  NOR3_X4 U13768 ( .A1(n15422), .A2(n12989), .A3(n12988), .ZN(n12987) );
  BUF_X16 U13771 ( .A(n17502), .Z(n10121) );
  INV_X16 U13823 ( .A(n13118), .ZN(n13879) );
  INV_X32 U13956 ( .A(n13879), .ZN(n13877) );
  NOR2_X2 U13983 ( .A1(n13878), .A2(n13073), .ZN(n14176) );
  CLKBUF_X3 U14037 ( .A(net225528), .Z(net239597) );
  AOI22_X2 U14058 ( .A1(n13987), .A2(n14081), .B1(n13985), .B2(n13986), .ZN(
        n13993) );
  INV_X8 U14061 ( .A(n18939), .ZN(n13158) );
  INV_X2 U14075 ( .A(n15700), .ZN(n18510) );
  INV_X16 U14080 ( .A(n13879), .ZN(n13878) );
  AOI21_X2 U14095 ( .B1(n13990), .B2(n14079), .A(n13989), .ZN(n13991) );
  AOI22_X1 U14102 ( .A1(n13490), .A2(n18457), .B1(n10829), .B2(
        DMEM_BUS_OUT[29]), .ZN(n18458) );
  INV_X8 U14103 ( .A(n18942), .ZN(n13160) );
  XNOR2_X1 U14116 ( .A(n18362), .B(n18361), .ZN(n18363) );
  XNOR2_X2 U14174 ( .A(n13122), .B(n13113), .ZN(n13144) );
  INV_X2 U14202 ( .A(n13122), .ZN(n13123) );
  AND3_X4 U14204 ( .A1(n13142), .A2(n13143), .A3(n13144), .ZN(n19355) );
  INV_X16 U14209 ( .A(n13158), .ZN(n13159) );
  NAND2_X4 U14215 ( .A1(n15830), .A2(n13159), .ZN(n15831) );
  NAND2_X2 U14247 ( .A1(net232816), .A2(n13159), .ZN(n16048) );
  NAND2_X1 U14266 ( .A1(n13409), .A2(n13159), .ZN(n18482) );
  NAND2_X1 U14270 ( .A1(n19107), .A2(n13159), .ZN(n18543) );
  NAND2_X1 U14311 ( .A1(net231615), .A2(n13159), .ZN(n18526) );
  NAND2_X1 U14323 ( .A1(n18360), .A2(n13159), .ZN(n18266) );
  XNOR2_X2 U14348 ( .A(n13150), .B(n19356), .ZN(n15828) );
  INV_X32 U14382 ( .A(n13494), .ZN(n19356) );
  INV_X4 U14385 ( .A(n13150), .ZN(n13151) );
  INV_X4 U14388 ( .A(n18548), .ZN(n15832) );
  XNOR2_X1 U14424 ( .A(n18549), .B(n18548), .ZN(n18551) );
  NAND2_X2 U14443 ( .A1(n13492), .A2(n16789), .ZN(n16828) );
  NAND4_X4 U14457 ( .A1(n16161), .A2(n16160), .A3(n16159), .A4(n16158), .ZN(
        n7374) );
  NAND2_X4 U14464 ( .A1(n16143), .A2(n13492), .ZN(n16161) );
  CLKBUF_X2 U14563 ( .A(net225684), .Z(net239718) );
  AOI21_X2 U14626 ( .B1(n16085), .B2(n13492), .A(n16084), .ZN(n16086) );
  BUF_X32 U14629 ( .A(n15775), .Z(n19358) );
  BUF_X32 U14634 ( .A(n15669), .Z(n19359) );
  NAND2_X1 U14677 ( .A1(DMEM_BUS_OUT[25]), .A2(n18927), .ZN(n15787) );
  NAND2_X4 U14706 ( .A1(n18628), .A2(n13095), .ZN(n13096) );
  NAND2_X2 U15190 ( .A1(n16078), .A2(n16077), .ZN(n16079) );
  NAND3_X1 U15339 ( .A1(ID_EXEC_OUT[87]), .A2(n13092), .A3(n15836), .ZN(n15764) );
  NAND2_X2 U15520 ( .A1(n13092), .A2(n15836), .ZN(n15677) );
  INV_X2 U15584 ( .A(net225163), .ZN(n10131) );
  XNOR2_X2 U15590 ( .A(n13053), .B(n13128), .ZN(n15500) );
  INV_X8 U16830 ( .A(n14000), .ZN(n14125) );
  NOR2_X4 U16923 ( .A1(n13154), .A2(n13148), .ZN(n14081) );
  INV_X2 U16980 ( .A(n18959), .ZN(n18961) );
  NAND2_X2 U17034 ( .A1(n18953), .A2(n18959), .ZN(n18954) );
  INV_X16 U17037 ( .A(n14068), .ZN(n14104) );
  INV_X8 U17038 ( .A(n14103), .ZN(n14105) );
  AOI22_X4 U17235 ( .A1(MEM_WB_OUT[29]), .A2(n13877), .B1(MEM_WB_OUT[98]), 
        .B2(n14102), .ZN(n14057) );
  AOI21_X4 U17280 ( .B1(n18949), .B2(n18948), .A(n18947), .ZN(n18957) );
  XNOR2_X1 U17313 ( .A(n18884), .B(n18885), .ZN(n19360) );
  INV_X1 U17344 ( .A(n18885), .ZN(n13051) );
  INV_X4 U17565 ( .A(net227045), .ZN(net225075) );
  NAND3_X4 U17566 ( .A1(n15816), .A2(n15817), .A3(n15818), .ZN(n18882) );
  XNOR2_X2 U17745 ( .A(n13054), .B(n13105), .ZN(n15499) );
  INV_X2 U17746 ( .A(n13105), .ZN(n13152) );
  NAND2_X4 U18213 ( .A1(n19362), .A2(n19363), .ZN(n19361) );
  XNOR2_X2 U18432 ( .A(n13129), .B(n13130), .ZN(n19362) );
  XNOR2_X2 U18464 ( .A(n13139), .B(n13140), .ZN(n19363) );
  NAND2_X4 U18508 ( .A1(ID_EXEC_OUT[93]), .A2(n18625), .ZN(n15689) );
  XNOR2_X2 U18722 ( .A(n18882), .B(n19091), .ZN(n19364) );
  AOI21_X4 U18786 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[17]), .B2(
        n14019), .A(n14104), .ZN(n14020) );
  NAND2_X4 U18845 ( .A1(n18664), .A2(n17094), .ZN(n14023) );
  INV_X8 U18859 ( .A(n18888), .ZN(n15732) );
  BUF_X32 U18895 ( .A(n18887), .Z(n13050) );
  NAND3_X2 U18903 ( .A1(n12936), .A2(n15651), .A3(n15648), .ZN(n15657) );
  AND2_X4 EXEC_STAGE_mul_ex_add_88_U2 ( .A1(ID_EXEC_OUT[235]), .A2(
        ID_EXEC_OUT[219]), .ZN(EXEC_STAGE_mul_ex_add_88_n2) );
  XOR2_X2 EXEC_STAGE_mul_ex_add_88_U1 ( .A(ID_EXEC_OUT[235]), .B(
        ID_EXEC_OUT[219]), .Z(EXEC_STAGE_mul_ex_N120) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_U1_1 ( .A(ID_EXEC_OUT[218]), .B(
        ID_EXEC_OUT[234]), .CI(EXEC_STAGE_mul_ex_add_88_n2), .CO(
        EXEC_STAGE_mul_ex_add_88_carry[2]), .S(EXEC_STAGE_mul_ex_N121) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_U1_2 ( .A(ID_EXEC_OUT[217]), .B(
        ID_EXEC_OUT[233]), .CI(EXEC_STAGE_mul_ex_add_88_carry[2]), .CO(
        EXEC_STAGE_mul_ex_add_88_carry[3]), .S(EXEC_STAGE_mul_ex_N122) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_U1_3 ( .A(ID_EXEC_OUT[216]), .B(
        ID_EXEC_OUT[232]), .CI(EXEC_STAGE_mul_ex_add_88_carry[3]), .CO(
        EXEC_STAGE_mul_ex_add_88_carry[4]), .S(EXEC_STAGE_mul_ex_N123) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_U1_4 ( .A(ID_EXEC_OUT[215]), .B(
        ID_EXEC_OUT[231]), .CI(EXEC_STAGE_mul_ex_add_88_carry[4]), .CO(
        EXEC_STAGE_mul_ex_add_88_carry[5]), .S(EXEC_STAGE_mul_ex_N124) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_U1_5 ( .A(ID_EXEC_OUT[214]), .B(
        ID_EXEC_OUT[230]), .CI(EXEC_STAGE_mul_ex_add_88_carry[5]), .CO(
        EXEC_STAGE_mul_ex_add_88_carry[6]), .S(EXEC_STAGE_mul_ex_N125) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_U1_6 ( .A(ID_EXEC_OUT[213]), .B(
        ID_EXEC_OUT[229]), .CI(EXEC_STAGE_mul_ex_add_88_carry[6]), .CO(
        EXEC_STAGE_mul_ex_add_88_carry[7]), .S(EXEC_STAGE_mul_ex_N126) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_U1_7 ( .A(ID_EXEC_OUT[212]), .B(
        ID_EXEC_OUT[228]), .CI(EXEC_STAGE_mul_ex_add_88_carry[7]), .CO(
        EXEC_STAGE_mul_ex_add_88_carry[8]), .S(EXEC_STAGE_mul_ex_N127) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_U1_8 ( .A(ID_EXEC_OUT[211]), .B(
        ID_EXEC_OUT[227]), .CI(EXEC_STAGE_mul_ex_add_88_carry[8]), .CO(
        EXEC_STAGE_mul_ex_add_88_carry[9]), .S(EXEC_STAGE_mul_ex_N128) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_U1_9 ( .A(ID_EXEC_OUT[210]), .B(
        ID_EXEC_OUT[226]), .CI(EXEC_STAGE_mul_ex_add_88_carry[9]), .CO(
        EXEC_STAGE_mul_ex_add_88_carry[10]), .S(EXEC_STAGE_mul_ex_N129) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_U1_10 ( .A(ID_EXEC_OUT[209]), .B(
        ID_EXEC_OUT[225]), .CI(EXEC_STAGE_mul_ex_add_88_carry[10]), .CO(
        EXEC_STAGE_mul_ex_add_88_carry[11]), .S(EXEC_STAGE_mul_ex_N130) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_U1_11 ( .A(ID_EXEC_OUT[208]), .B(
        ID_EXEC_OUT[224]), .CI(EXEC_STAGE_mul_ex_add_88_carry[11]), .CO(
        EXEC_STAGE_mul_ex_add_88_carry[12]), .S(EXEC_STAGE_mul_ex_N131) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_U1_12 ( .A(ID_EXEC_OUT[207]), .B(
        ID_EXEC_OUT[223]), .CI(EXEC_STAGE_mul_ex_add_88_carry[12]), .CO(
        EXEC_STAGE_mul_ex_add_88_carry[13]), .S(EXEC_STAGE_mul_ex_N132) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_U1_13 ( .A(ID_EXEC_OUT[206]), .B(
        ID_EXEC_OUT[222]), .CI(EXEC_STAGE_mul_ex_add_88_carry[13]), .CO(
        EXEC_STAGE_mul_ex_add_88_carry[14]), .S(EXEC_STAGE_mul_ex_N133) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_U1_14 ( .A(ID_EXEC_OUT[205]), .B(
        ID_EXEC_OUT[221]), .CI(EXEC_STAGE_mul_ex_add_88_carry[14]), .CO(
        EXEC_STAGE_mul_ex_add_88_carry[15]), .S(EXEC_STAGE_mul_ex_N134) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_U1_15 ( .A(ID_EXEC_OUT[204]), .B(
        ID_EXEC_OUT[220]), .CI(EXEC_STAGE_mul_ex_add_88_carry[15]), .CO(
        EXEC_STAGE_mul_ex_N136), .S(EXEC_STAGE_mul_ex_N135) );
  AND2_X4 EXEC_STAGE_mul_ex_add_88_2_U2 ( .A1(ID_EXEC_OUT[267]), .A2(
        ID_EXEC_OUT[251]), .ZN(EXEC_STAGE_mul_ex_add_88_2_n2) );
  XOR2_X2 EXEC_STAGE_mul_ex_add_88_2_U1 ( .A(ID_EXEC_OUT[267]), .B(
        ID_EXEC_OUT[251]), .Z(EXEC_STAGE_mul_ex_N137) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_2_U1_1 ( .A(ID_EXEC_OUT[250]), .B(
        ID_EXEC_OUT[266]), .CI(EXEC_STAGE_mul_ex_add_88_2_n2), .CO(
        EXEC_STAGE_mul_ex_add_88_2_carry[2]), .S(EXEC_STAGE_mul_ex_N138) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_2_U1_2 ( .A(ID_EXEC_OUT[249]), .B(
        ID_EXEC_OUT[265]), .CI(EXEC_STAGE_mul_ex_add_88_2_carry[2]), .CO(
        EXEC_STAGE_mul_ex_add_88_2_carry[3]), .S(EXEC_STAGE_mul_ex_N139) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_2_U1_3 ( .A(ID_EXEC_OUT[248]), .B(
        ID_EXEC_OUT[264]), .CI(EXEC_STAGE_mul_ex_add_88_2_carry[3]), .CO(
        EXEC_STAGE_mul_ex_add_88_2_carry[4]), .S(EXEC_STAGE_mul_ex_N140) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_2_U1_4 ( .A(ID_EXEC_OUT[247]), .B(
        ID_EXEC_OUT[263]), .CI(EXEC_STAGE_mul_ex_add_88_2_carry[4]), .CO(
        EXEC_STAGE_mul_ex_add_88_2_carry[5]), .S(EXEC_STAGE_mul_ex_N141) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_2_U1_5 ( .A(ID_EXEC_OUT[246]), .B(
        ID_EXEC_OUT[262]), .CI(EXEC_STAGE_mul_ex_add_88_2_carry[5]), .CO(
        EXEC_STAGE_mul_ex_add_88_2_carry[6]), .S(EXEC_STAGE_mul_ex_N142) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_2_U1_6 ( .A(ID_EXEC_OUT[245]), .B(
        ID_EXEC_OUT[261]), .CI(EXEC_STAGE_mul_ex_add_88_2_carry[6]), .CO(
        EXEC_STAGE_mul_ex_add_88_2_carry[7]), .S(EXEC_STAGE_mul_ex_N143) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_2_U1_7 ( .A(ID_EXEC_OUT[244]), .B(
        ID_EXEC_OUT[260]), .CI(EXEC_STAGE_mul_ex_add_88_2_carry[7]), .CO(
        EXEC_STAGE_mul_ex_add_88_2_carry[8]), .S(EXEC_STAGE_mul_ex_N144) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_2_U1_8 ( .A(ID_EXEC_OUT[243]), .B(
        ID_EXEC_OUT[259]), .CI(EXEC_STAGE_mul_ex_add_88_2_carry[8]), .CO(
        EXEC_STAGE_mul_ex_add_88_2_carry[9]), .S(EXEC_STAGE_mul_ex_N145) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_2_U1_9 ( .A(ID_EXEC_OUT[242]), .B(
        ID_EXEC_OUT[258]), .CI(EXEC_STAGE_mul_ex_add_88_2_carry[9]), .CO(
        EXEC_STAGE_mul_ex_add_88_2_carry[10]), .S(EXEC_STAGE_mul_ex_N146) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_2_U1_10 ( .A(ID_EXEC_OUT[241]), .B(
        ID_EXEC_OUT[257]), .CI(EXEC_STAGE_mul_ex_add_88_2_carry[10]), .CO(
        EXEC_STAGE_mul_ex_add_88_2_carry[11]), .S(EXEC_STAGE_mul_ex_N147) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_2_U1_11 ( .A(ID_EXEC_OUT[240]), .B(
        ID_EXEC_OUT[256]), .CI(EXEC_STAGE_mul_ex_add_88_2_carry[11]), .CO(
        EXEC_STAGE_mul_ex_add_88_2_carry[12]), .S(EXEC_STAGE_mul_ex_N148) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_2_U1_12 ( .A(ID_EXEC_OUT[239]), .B(
        ID_EXEC_OUT[255]), .CI(EXEC_STAGE_mul_ex_add_88_2_carry[12]), .CO(
        EXEC_STAGE_mul_ex_add_88_2_carry[13]), .S(EXEC_STAGE_mul_ex_N149) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_2_U1_13 ( .A(ID_EXEC_OUT[238]), .B(
        ID_EXEC_OUT[254]), .CI(EXEC_STAGE_mul_ex_add_88_2_carry[13]), .CO(
        EXEC_STAGE_mul_ex_add_88_2_carry[14]), .S(EXEC_STAGE_mul_ex_N150) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_2_U1_14 ( .A(ID_EXEC_OUT[237]), .B(
        ID_EXEC_OUT[253]), .CI(EXEC_STAGE_mul_ex_add_88_2_carry[14]), .CO(
        EXEC_STAGE_mul_ex_add_88_2_carry[15]), .S(EXEC_STAGE_mul_ex_N151) );
  FA_X1 EXEC_STAGE_mul_ex_add_88_2_U1_15 ( .A(ID_EXEC_OUT[236]), .B(
        ID_EXEC_OUT[252]), .CI(EXEC_STAGE_mul_ex_add_88_2_carry[15]), .CO(
        EXEC_STAGE_mul_ex_N153), .S(EXEC_STAGE_mul_ex_N152) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U389 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(EXEC_STAGE_mul_ex_N154) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U388 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U387 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U386 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U385 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U384 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U383 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U382 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U381 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U380 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U379 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U378 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U377 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U376 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U375 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U374 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U373 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_0__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U372 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U371 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U370 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U369 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U368 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U367 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U366 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U365 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U364 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U363 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U362 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U361 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U360 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U359 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U358 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U357 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U356 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_10__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U355 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U354 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U353 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U352 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U351 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U350 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U349 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U348 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U347 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U346 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U345 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U344 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U343 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U342 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U341 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U340 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U339 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_11__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U338 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U337 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U336 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U335 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U334 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U333 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U332 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U331 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U330 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U329 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U328 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U327 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U326 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U325 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U324 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U323 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U322 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_12__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U321 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U320 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U319 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U318 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U317 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U316 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U315 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U314 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U313 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U312 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U311 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U310 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U309 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U308 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U307 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U306 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U305 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_13__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U304 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U303 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U302 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U301 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U300 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U299 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U298 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U297 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U296 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U295 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U294 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U293 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U292 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U291 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U290 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U289 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U288 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_14__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U287 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U286 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U285 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U284 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U283 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U282 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U281 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U280 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U279 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U278 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U277 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U276 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U275 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U274 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U273 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U272 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U271 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_15__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U270 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U269 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U268 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U267 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U266 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U265 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U264 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U263 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U262 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U261 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U260 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U259 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U258 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U257 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U256 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U255 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U254 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_16__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U253 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U252 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U251 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U250 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U249 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U248 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U247 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U246 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U245 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U244 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U243 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U242 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U241 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U240 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U239 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U238 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U237 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_1__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U236 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U235 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U234 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U233 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U232 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U231 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U230 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U229 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U228 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U227 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U226 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U225 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U224 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U223 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U222 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U221 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U220 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_2__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U219 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U218 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U217 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U216 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U215 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U214 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U213 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U212 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U211 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U210 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U209 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U208 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U207 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U206 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U205 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U204 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U203 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_3__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U202 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U201 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U200 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U199 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U198 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U197 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U196 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U195 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U194 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U193 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U192 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U191 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U190 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U189 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U188 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U187 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U186 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_4__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U185 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U184 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U183 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U182 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U181 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U180 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U179 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U178 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U177 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U176 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U175 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U174 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U173 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U172 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U171 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U170 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U169 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_5__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U168 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U167 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U166 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U165 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U164 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U163 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U162 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U161 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U160 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U159 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U158 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U157 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U156 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U155 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U154 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U153 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U152 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_6__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U151 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U150 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U149 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U148 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U147 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U146 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U145 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U144 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U143 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U142 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U141 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U140 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U139 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U138 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U137 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U136 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U135 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_7__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U134 ( .A1(EXEC_STAGE_mul_ex_mult_88_n100), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U133 ( .A1(EXEC_STAGE_mul_ex_mult_88_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U132 ( .A1(EXEC_STAGE_mul_ex_mult_88_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U131 ( .A1(EXEC_STAGE_mul_ex_mult_88_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U130 ( .A1(EXEC_STAGE_mul_ex_mult_88_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U129 ( .A1(EXEC_STAGE_mul_ex_mult_88_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U128 ( .A1(EXEC_STAGE_mul_ex_mult_88_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U127 ( .A1(EXEC_STAGE_mul_ex_mult_88_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U126 ( .A1(EXEC_STAGE_mul_ex_mult_88_n99), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U125 ( .A1(EXEC_STAGE_mul_ex_mult_88_n98), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U124 ( .A1(EXEC_STAGE_mul_ex_mult_88_n97), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U123 ( .A1(EXEC_STAGE_mul_ex_mult_88_n96), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U122 ( .A1(EXEC_STAGE_mul_ex_mult_88_n95), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U121 ( .A1(EXEC_STAGE_mul_ex_mult_88_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U120 ( .A1(EXEC_STAGE_mul_ex_mult_88_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U119 ( .A1(EXEC_STAGE_mul_ex_mult_88_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U118 ( .A1(EXEC_STAGE_mul_ex_mult_88_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_8__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U117 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n100), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U116 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U115 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U114 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U113 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U112 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U111 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U110 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U109 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n99), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U108 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n98), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U107 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n97), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U106 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n96), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U105 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n95), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U104 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n94), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U103 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U102 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_U101 ( .A1(EXEC_STAGE_mul_ex_mult_88_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_88_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_88_ab_9__9_) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U99 ( .A(EXEC_STAGE_mul_ex_N137), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n100) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U98 ( .A(EXEC_STAGE_mul_ex_N138), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n99) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U97 ( .A(EXEC_STAGE_mul_ex_N139), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n98) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U96 ( .A(EXEC_STAGE_mul_ex_N140), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n97) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U95 ( .A(EXEC_STAGE_mul_ex_N141), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n96) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U94 ( .A(EXEC_STAGE_mul_ex_N142), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n95) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U93 ( .A(EXEC_STAGE_mul_ex_N143), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n94) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U92 ( .A(EXEC_STAGE_mul_ex_N144), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n93) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U91 ( .A(EXEC_STAGE_mul_ex_N145), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n92) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U90 ( .A(EXEC_STAGE_mul_ex_N146), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n91) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U89 ( .A(EXEC_STAGE_mul_ex_N147), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n90) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U88 ( .A(EXEC_STAGE_mul_ex_N148), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n89) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U87 ( .A(EXEC_STAGE_mul_ex_N149), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n88) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U86 ( .A(EXEC_STAGE_mul_ex_N150), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n87) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U85 ( .A(EXEC_STAGE_mul_ex_N151), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n86) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U84 ( .A(EXEC_STAGE_mul_ex_N152), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n85) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U83 ( .A(EXEC_STAGE_mul_ex_N120), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n83) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U82 ( .A(EXEC_STAGE_mul_ex_N121), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n82) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U81 ( .A(EXEC_STAGE_mul_ex_N122), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n81) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U80 ( .A(EXEC_STAGE_mul_ex_N123), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n80) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U79 ( .A(EXEC_STAGE_mul_ex_N124), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n79) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U78 ( .A(EXEC_STAGE_mul_ex_N125), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n78) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U77 ( .A(EXEC_STAGE_mul_ex_N126), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n77) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U76 ( .A(EXEC_STAGE_mul_ex_N127), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n76) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U75 ( .A(EXEC_STAGE_mul_ex_N128), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n75) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U74 ( .A(EXEC_STAGE_mul_ex_N129), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n74) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U73 ( .A(EXEC_STAGE_mul_ex_N130), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n73) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U72 ( .A(EXEC_STAGE_mul_ex_N131), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n72) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U71 ( .A(EXEC_STAGE_mul_ex_N132), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n71) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U70 ( .A(EXEC_STAGE_mul_ex_N133), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n70) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U69 ( .A(EXEC_STAGE_mul_ex_N134), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n69) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U68 ( .A(EXEC_STAGE_mul_ex_N135), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n68) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U67 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__1_), .Z(
        EXEC_STAGE_mul_ex_mult_88_n66) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U66 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__13_), .A2(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__14_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n65) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U65 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__1_), .Z(EXEC_STAGE_mul_ex_N155) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U64 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__0_), .A2(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n63) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U63 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__2_), .A2(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n62) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U62 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__4_), .A2(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n61) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U61 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__6_), .A2(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n60) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U60 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__8_), .A2(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n59) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U59 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__10_), .A2(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__11_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n58) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U58 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__12_), .A2(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__13_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n57) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U57 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__1_), .A2(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n56) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U56 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__3_), .A2(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n55) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U55 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__5_), .A2(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n54) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U54 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__7_), .A2(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n53) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U53 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__9_), .A2(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n52) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U52 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__11_), .A2(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__12_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n51) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U51 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__2_), .Z(EXEC_STAGE_mul_ex_mult_88_n50)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U50 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__3_), .Z(EXEC_STAGE_mul_ex_mult_88_n49)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U49 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__4_), .Z(EXEC_STAGE_mul_ex_mult_88_n48)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U48 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__5_), .Z(EXEC_STAGE_mul_ex_mult_88_n47)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U47 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__6_), .Z(EXEC_STAGE_mul_ex_mult_88_n46)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U46 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__7_), .Z(EXEC_STAGE_mul_ex_mult_88_n45)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U45 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__8_), .Z(EXEC_STAGE_mul_ex_mult_88_n44)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U44 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__9_), .Z(EXEC_STAGE_mul_ex_mult_88_n43)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U43 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__10_), .Z(EXEC_STAGE_mul_ex_mult_88_n42) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U42 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__11_), .Z(EXEC_STAGE_mul_ex_mult_88_n41) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U41 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__12_), .Z(EXEC_STAGE_mul_ex_mult_88_n40) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U40 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__13_), .Z(EXEC_STAGE_mul_ex_mult_88_n39) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U39 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__14_), .Z(EXEC_STAGE_mul_ex_mult_88_n38) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U38 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__15_), .Z(EXEC_STAGE_mul_ex_mult_88_n37) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U37 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_1__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_0__16_), .Z(EXEC_STAGE_mul_ex_mult_88_n36) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U36 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__16_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__15_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n35) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U35 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__15_), .Z(
        EXEC_STAGE_mul_ex_mult_88_n34) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U34 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__4_), .Z(
        EXEC_STAGE_mul_ex_mult_88_n33) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U33 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__6_), .Z(
        EXEC_STAGE_mul_ex_mult_88_n32) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U32 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__8_), .Z(
        EXEC_STAGE_mul_ex_mult_88_n31) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U31 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__10_), .Z(
        EXEC_STAGE_mul_ex_mult_88_n30) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U30 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__12_), .Z(
        EXEC_STAGE_mul_ex_mult_88_n29) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U29 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__14_), .Z(
        EXEC_STAGE_mul_ex_mult_88_n28) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U28 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__2_), .Z(
        EXEC_STAGE_mul_ex_mult_88_n27) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U27 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__3_), .Z(
        EXEC_STAGE_mul_ex_mult_88_n26) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U26 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__5_), .Z(
        EXEC_STAGE_mul_ex_mult_88_n25) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U25 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__7_), .Z(
        EXEC_STAGE_mul_ex_mult_88_n24) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U24 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__9_), .Z(
        EXEC_STAGE_mul_ex_mult_88_n23) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U23 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__11_), .Z(
        EXEC_STAGE_mul_ex_mult_88_n22) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U22 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__13_), .Z(
        EXEC_STAGE_mul_ex_mult_88_n21) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U21 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__1_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__0_), .ZN(EXEC_STAGE_mul_ex_mult_88_n20) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U20 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__2_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__1_), .ZN(EXEC_STAGE_mul_ex_mult_88_n19) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U19 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__3_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__2_), .ZN(EXEC_STAGE_mul_ex_mult_88_n18) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U18 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__4_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__3_), .ZN(EXEC_STAGE_mul_ex_mult_88_n17) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U17 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__5_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__4_), .ZN(EXEC_STAGE_mul_ex_mult_88_n16) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U16 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__6_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__5_), .ZN(EXEC_STAGE_mul_ex_mult_88_n15) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U15 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__7_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__6_), .ZN(EXEC_STAGE_mul_ex_mult_88_n14) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U14 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__8_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__7_), .ZN(EXEC_STAGE_mul_ex_mult_88_n13) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U13 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__9_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__8_), .ZN(EXEC_STAGE_mul_ex_mult_88_n12) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U12 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__10_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__9_), .ZN(EXEC_STAGE_mul_ex_mult_88_n11) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U11 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__11_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n10) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U10 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__12_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__11_), .ZN(EXEC_STAGE_mul_ex_mult_88_n9) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U9 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__13_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__12_), .ZN(EXEC_STAGE_mul_ex_mult_88_n8) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U8 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__14_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__13_), .ZN(EXEC_STAGE_mul_ex_mult_88_n7) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U7 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_ab_0__15_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_1__14_), .ZN(EXEC_STAGE_mul_ex_mult_88_n6) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_88_U6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_ab_16__16_), .Z(EXEC_STAGE_mul_ex_mult_88_n5) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U5 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__15_), .A2(
        EXEC_STAGE_mul_ex_mult_88_ab_16__16_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n4) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_U4 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__14_), .A2(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__15_), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n3) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U3 ( .A(EXEC_STAGE_mul_ex_N136), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n67) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_U2 ( .A(EXEC_STAGE_mul_ex_N153), .ZN(
        EXEC_STAGE_mul_ex_mult_88_n84) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S3_2_15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__15_), .B(EXEC_STAGE_mul_ex_mult_88_n35), .CI(EXEC_STAGE_mul_ex_mult_88_ab_1__16_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__15_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_2_14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__14_), .B(EXEC_STAGE_mul_ex_mult_88_n6), 
        .CI(EXEC_STAGE_mul_ex_mult_88_n36), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__14_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_2_13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__13_), .B(EXEC_STAGE_mul_ex_mult_88_n7), 
        .CI(EXEC_STAGE_mul_ex_mult_88_n37), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__13_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_2_12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__12_), .B(EXEC_STAGE_mul_ex_mult_88_n8), 
        .CI(EXEC_STAGE_mul_ex_mult_88_n38), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__12_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_2_11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__11_), .B(EXEC_STAGE_mul_ex_mult_88_n9), 
        .CI(EXEC_STAGE_mul_ex_mult_88_n39), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__11_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_2_10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__10_), .B(EXEC_STAGE_mul_ex_mult_88_n10), .CI(EXEC_STAGE_mul_ex_mult_88_n40), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__10_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_2_9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__9_), .B(EXEC_STAGE_mul_ex_mult_88_n11), 
        .CI(EXEC_STAGE_mul_ex_mult_88_n41), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__9_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_2_8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__8_), .B(EXEC_STAGE_mul_ex_mult_88_n12), 
        .CI(EXEC_STAGE_mul_ex_mult_88_n42), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__8_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_2_7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__7_), .B(EXEC_STAGE_mul_ex_mult_88_n13), 
        .CI(EXEC_STAGE_mul_ex_mult_88_n43), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__7_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_2_6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__6_), .B(EXEC_STAGE_mul_ex_mult_88_n14), 
        .CI(EXEC_STAGE_mul_ex_mult_88_n44), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__6_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_2_5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__5_), .B(EXEC_STAGE_mul_ex_mult_88_n15), 
        .CI(EXEC_STAGE_mul_ex_mult_88_n45), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__5_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_2_4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__4_), .B(EXEC_STAGE_mul_ex_mult_88_n16), 
        .CI(EXEC_STAGE_mul_ex_mult_88_n46), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__4_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_2_3 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__3_), .B(EXEC_STAGE_mul_ex_mult_88_n17), 
        .CI(EXEC_STAGE_mul_ex_mult_88_n47), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__3_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_2_2 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__2_), .B(EXEC_STAGE_mul_ex_mult_88_n18), 
        .CI(EXEC_STAGE_mul_ex_mult_88_n48), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__2_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_2_1 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__1_), .B(EXEC_STAGE_mul_ex_mult_88_n19), 
        .CI(EXEC_STAGE_mul_ex_mult_88_n49), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__1_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S1_2_0 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_2__0_), .B(EXEC_STAGE_mul_ex_mult_88_n20), 
        .CI(EXEC_STAGE_mul_ex_mult_88_n50), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__0_), .S(
        EXEC_STAGE_mul_ex_mult_88_A1_0_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S3_3_15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__15_), .CI(
        EXEC_STAGE_mul_ex_mult_88_ab_2__16_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__15_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_3_14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__14_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__15_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__14_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_3_13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__13_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__14_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__13_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_3_12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__12_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__13_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__12_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_3_11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__11_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__12_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__11_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_3_10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__10_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__11_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__10_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_3_9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__9_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__10_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__9_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_3_8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__8_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__9_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__8_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_3_7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__7_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__8_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__7_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_3_6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__6_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__7_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__6_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_3_5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__5_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__6_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__5_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_3_4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__4_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__5_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__4_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_3_3 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__3_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__4_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__3_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_3_2 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__2_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__3_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__2_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_3_1 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__1_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__2_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__1_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S1_3_0 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_3__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_2__0_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_2__1_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__0_), .S(
        EXEC_STAGE_mul_ex_mult_88_A1_1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S3_4_15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__15_), .CI(
        EXEC_STAGE_mul_ex_mult_88_ab_3__16_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__15_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_4_14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__14_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__15_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__14_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_4_13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__13_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__14_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__13_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_4_12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__12_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__13_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__12_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_4_11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__11_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__12_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__11_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_4_10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__10_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__11_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__10_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_4_9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__9_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__10_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__9_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_4_8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__8_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__9_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__8_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_4_7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__7_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__8_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__7_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_4_6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__6_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__7_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__6_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_4_5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__5_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__6_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__5_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_4_4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__4_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__5_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__4_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_4_3 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__3_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__4_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__3_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_4_2 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__2_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__3_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__2_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_4_1 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__1_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__2_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__1_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S1_4_0 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_4__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_3__0_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_3__1_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__0_), .S(
        EXEC_STAGE_mul_ex_mult_88_A1_2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S3_5_15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__15_), .CI(
        EXEC_STAGE_mul_ex_mult_88_ab_4__16_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__15_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_5_14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__14_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__15_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__14_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_5_13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__13_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__14_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__13_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_5_12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__12_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__13_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__12_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_5_11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__11_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__12_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__11_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_5_10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__10_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__11_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__10_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_5_9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__9_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__10_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__9_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_5_8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__8_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__9_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__8_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_5_7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__7_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__8_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__7_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_5_6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__6_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__7_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__6_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_5_5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__5_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__6_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__5_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_5_4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__4_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__5_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__4_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_5_3 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__3_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__4_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__3_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_5_2 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__2_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__3_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__2_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_5_1 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__1_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__2_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__1_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S1_5_0 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_5__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_4__0_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_4__1_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__0_), .S(
        EXEC_STAGE_mul_ex_mult_88_A1_3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S3_6_15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__15_), .CI(
        EXEC_STAGE_mul_ex_mult_88_ab_5__16_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__15_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_6_14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__14_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__15_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__14_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_6_13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__13_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__14_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__13_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_6_12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__12_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__13_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__12_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_6_11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__11_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__12_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__11_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_6_10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__10_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__11_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__10_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_6_9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__9_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__10_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__9_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_6_8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__8_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__9_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__8_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_6_7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__7_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__8_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__7_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_6_6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__6_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__7_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__6_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_6_5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__5_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__6_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__5_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_6_4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__4_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__5_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__4_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_6_3 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__3_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__4_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__3_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_6_2 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__2_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__3_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__2_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_6_1 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__1_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__2_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__1_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S1_6_0 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_6__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_5__0_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_5__1_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__0_), .S(
        EXEC_STAGE_mul_ex_mult_88_A1_4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S3_7_15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__15_), .CI(
        EXEC_STAGE_mul_ex_mult_88_ab_6__16_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__15_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_7_14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__14_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__15_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__14_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_7_13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__13_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__14_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__13_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_7_12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__12_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__13_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__12_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_7_11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__11_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__12_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__11_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_7_10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__10_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__11_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__10_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_7_9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__9_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__10_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__9_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_7_8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__8_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__9_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__8_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_7_7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__7_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__8_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__7_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_7_6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__6_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__7_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__6_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_7_5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__5_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__6_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__5_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_7_4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__4_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__5_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__4_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_7_3 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__3_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__4_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__3_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_7_2 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__2_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__3_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__2_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_7_1 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__1_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__2_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__1_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S1_7_0 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_7__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_6__0_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_6__1_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__0_), .S(
        EXEC_STAGE_mul_ex_mult_88_A1_5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S3_8_15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__15_), .CI(
        EXEC_STAGE_mul_ex_mult_88_ab_7__16_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__15_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_8_14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__14_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__15_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__14_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_8_13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__13_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__14_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__13_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_8_12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__12_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__13_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__12_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_8_11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__11_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__12_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__11_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_8_10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__10_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__11_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__10_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_8_9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__9_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__10_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__9_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_8_8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__8_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__9_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__8_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_8_7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__7_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__8_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__7_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_8_6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__6_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__7_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__6_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_8_5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__5_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__6_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__5_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_8_4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__4_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__5_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__4_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_8_3 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__3_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__4_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__3_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_8_2 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__2_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__3_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__2_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_8_1 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__1_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__2_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__1_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S1_8_0 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_8__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_7__0_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_7__1_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__0_), .S(
        EXEC_STAGE_mul_ex_mult_88_A1_6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S3_9_15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__15_), .CI(
        EXEC_STAGE_mul_ex_mult_88_ab_8__16_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__15_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_9_14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__14_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__15_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__14_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_9_13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__13_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__14_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__13_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_9_12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__12_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__13_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__12_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_9_11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__11_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__12_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__11_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_9_10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__10_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__11_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__10_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_9_9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__9_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__10_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__9_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_9_8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__8_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__9_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__8_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_9_7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__7_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__8_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__7_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_9_6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__6_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__7_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__6_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_9_5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__5_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__6_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__5_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_9_4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__4_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__5_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__4_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_9_3 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__3_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__4_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__3_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_9_2 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__2_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__3_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__2_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_9_1 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__1_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__2_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__1_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S1_9_0 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_9__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_8__0_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_8__1_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__0_), .S(
        EXEC_STAGE_mul_ex_mult_88_A1_7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S3_10_15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__15_), .CI(
        EXEC_STAGE_mul_ex_mult_88_ab_9__16_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__15_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_10_14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__14_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__15_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__14_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_10_13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__13_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__14_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__13_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_10_12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__12_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__13_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__12_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_10_11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__11_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__12_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__11_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_10_10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__10_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__11_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__10_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_10_9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__9_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__10_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__9_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_10_8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__8_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__9_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__8_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_10_7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__7_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__8_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__7_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_10_6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__6_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__7_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__6_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_10_5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__5_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__6_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__5_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_10_4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__4_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__5_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__4_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_10_3 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__3_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__4_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__3_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_10_2 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__2_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__3_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__2_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_10_1 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__1_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__2_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__1_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S1_10_0 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_10__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_9__0_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_9__1_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__0_), .S(
        EXEC_STAGE_mul_ex_mult_88_A1_8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S3_11_15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__15_), .CI(
        EXEC_STAGE_mul_ex_mult_88_ab_10__16_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__15_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_11_14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__14_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__15_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__14_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_11_13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__13_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__14_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__13_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_11_12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__12_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__13_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__12_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_11_11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__11_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__12_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__11_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_11_10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__10_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__11_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__10_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_11_9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__9_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__10_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__9_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_11_8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__8_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__9_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__8_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_11_7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__7_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__8_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__7_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_11_6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__6_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__7_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__6_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_11_5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__5_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__6_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__5_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_11_4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__4_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__5_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__4_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_11_3 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__3_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__4_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__3_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_11_2 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__2_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__3_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__2_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_11_1 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__1_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__2_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__1_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S1_11_0 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_11__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_10__0_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_10__1_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__0_), .S(
        EXEC_STAGE_mul_ex_mult_88_A1_9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S3_12_15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__15_), .CI(
        EXEC_STAGE_mul_ex_mult_88_ab_11__16_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__15_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_12_14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__14_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__15_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__14_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_12_13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__13_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__14_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__13_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_12_12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__12_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__13_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__12_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_12_11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__11_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__12_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__11_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_12_10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__10_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__11_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__10_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_12_9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__9_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__10_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__9_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_12_8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__8_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__9_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__8_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_12_7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__7_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__8_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__7_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_12_6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__6_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__7_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__6_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_12_5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__5_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__6_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__5_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_12_4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__4_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__5_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__4_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_12_3 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__3_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__4_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__3_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_12_2 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__2_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__3_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__2_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_12_1 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__1_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__2_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__1_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S1_12_0 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_12__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_11__0_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_11__1_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__0_), .S(
        EXEC_STAGE_mul_ex_mult_88_A1_10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S3_13_15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__15_), .CI(
        EXEC_STAGE_mul_ex_mult_88_ab_12__16_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__15_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_13_14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__14_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__15_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__14_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_13_13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__13_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__14_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__13_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_13_12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__12_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__13_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__12_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_13_11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__11_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__12_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__11_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_13_10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__10_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__11_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__10_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_13_9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__9_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__10_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__9_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_13_8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__8_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__9_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__8_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_13_7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__7_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__8_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__7_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_13_6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__6_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__7_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__6_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_13_5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__5_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__6_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__5_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_13_4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__4_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__5_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__4_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_13_3 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__3_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__4_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__3_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_13_2 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__2_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__3_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__2_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_13_1 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__1_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__2_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__1_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S1_13_0 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_13__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_12__0_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_12__1_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__0_), .S(
        EXEC_STAGE_mul_ex_mult_88_A1_11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S3_14_15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__15_), .CI(
        EXEC_STAGE_mul_ex_mult_88_ab_13__16_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__15_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_14_14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__14_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__15_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__14_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_14_13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__13_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__14_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__13_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_14_12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__12_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__13_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__12_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_14_11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__11_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__12_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__11_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_14_10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__10_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__11_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__10_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_14_9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__9_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__10_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__9_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_14_8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__8_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__9_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__8_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_14_7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__7_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__8_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__7_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_14_6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__6_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__7_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__6_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_14_5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__5_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__6_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__5_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_14_4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__4_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__5_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__4_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_14_3 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__3_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__4_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__3_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_14_2 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__2_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__3_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__2_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_14_1 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__1_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__2_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__1_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S1_14_0 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_14__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_13__0_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_13__1_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__0_), .S(
        EXEC_STAGE_mul_ex_mult_88_A1_12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S3_15_15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__15_), .CI(
        EXEC_STAGE_mul_ex_mult_88_ab_14__16_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__15_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_15_14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__14_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__15_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__14_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_15_13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__13_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__14_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__13_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_15_12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__12_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__13_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__12_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_15_11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__11_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__12_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__11_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_15_10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__10_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__11_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__10_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_15_9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__9_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__10_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__9_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_15_8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__8_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__9_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__8_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_15_7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__7_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__8_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__7_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_15_6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__6_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__7_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__6_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_15_5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__5_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__6_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__5_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_15_4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__4_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__5_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__4_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_15_3 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__3_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__4_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__3_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_15_2 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__2_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__3_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__2_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S2_15_1 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__1_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__2_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__1_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S1_15_0 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_15__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_14__0_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_14__1_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__0_), .S(
        EXEC_STAGE_mul_ex_mult_88_A1_13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S5_15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__15_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__15_), .CI(
        EXEC_STAGE_mul_ex_mult_88_ab_15__16_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__15_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S4_14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__14_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__14_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__15_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__14_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S4_13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__13_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__13_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__14_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__13_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S4_12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__12_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__12_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__13_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__12_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S4_11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__11_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__11_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__12_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__11_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S4_10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__10_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__10_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__11_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__10_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S4_9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__9_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__9_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__10_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__9_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S4_8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__8_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__8_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__9_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__8_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S4_7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__7_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__7_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__8_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__7_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S4_6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__6_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__6_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__7_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__6_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S4_5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__5_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__5_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__6_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__5_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S4_4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__4_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__4_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__5_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__4_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S4_3 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__3_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__3_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__4_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__3_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S4_2 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__2_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__2_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__3_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__2_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S4_1 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__1_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__1_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__2_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__1_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_88_S4_0 ( .A(
        EXEC_STAGE_mul_ex_mult_88_ab_16__0_), .B(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_15__0_), .CI(
        EXEC_STAGE_mul_ex_mult_88_SUMB_15__1_), .CO(
        EXEC_STAGE_mul_ex_mult_88_CARRYB_16__0_), .S(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__0_) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U95 ( .A(
        EXEC_STAGE_mul_ex_mult_88_n66), .Z(EXEC_STAGE_mul_ex_N171) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U94 ( .A(
        EXEC_STAGE_mul_ex_mult_88_SUMB_16__0_), .Z(EXEC_STAGE_mul_ex_N170) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U93 ( .A(
        EXEC_STAGE_mul_ex_mult_88_A1_13_), .Z(EXEC_STAGE_mul_ex_N169) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U92 ( .A(
        EXEC_STAGE_mul_ex_mult_88_A1_12_), .Z(EXEC_STAGE_mul_ex_N168) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U91 ( .A(
        EXEC_STAGE_mul_ex_mult_88_A1_11_), .Z(EXEC_STAGE_mul_ex_N167) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U90 ( .A(
        EXEC_STAGE_mul_ex_mult_88_A1_10_), .Z(EXEC_STAGE_mul_ex_N166) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U89 ( .A(
        EXEC_STAGE_mul_ex_mult_88_A1_9_), .Z(EXEC_STAGE_mul_ex_N165) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U88 ( .A(
        EXEC_STAGE_mul_ex_mult_88_A1_8_), .Z(EXEC_STAGE_mul_ex_N164) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U87 ( .A(
        EXEC_STAGE_mul_ex_mult_88_A1_7_), .Z(EXEC_STAGE_mul_ex_N163) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U86 ( .A(
        EXEC_STAGE_mul_ex_mult_88_A1_6_), .Z(EXEC_STAGE_mul_ex_N162) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U85 ( .A(
        EXEC_STAGE_mul_ex_mult_88_A1_5_), .Z(EXEC_STAGE_mul_ex_N161) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U84 ( .A(
        EXEC_STAGE_mul_ex_mult_88_A1_4_), .Z(EXEC_STAGE_mul_ex_N160) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U83 ( .A(
        EXEC_STAGE_mul_ex_mult_88_A1_3_), .Z(EXEC_STAGE_mul_ex_N159) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U82 ( .A(
        EXEC_STAGE_mul_ex_mult_88_A1_2_), .Z(EXEC_STAGE_mul_ex_N158) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U81 ( .A(
        EXEC_STAGE_mul_ex_mult_88_A1_1_), .Z(EXEC_STAGE_mul_ex_N157) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_88_FS_1_U80 ( .A(
        EXEC_STAGE_mul_ex_mult_88_A1_0_), .Z(EXEC_STAGE_mul_ex_N156) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U79 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n63), .A2(EXEC_STAGE_mul_ex_mult_88_n27), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n65) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U78 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n56), .A2(EXEC_STAGE_mul_ex_mult_88_n26), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n62) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U77 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n56), .A2(EXEC_STAGE_mul_ex_mult_88_n26), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n63) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U76 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n62), .A2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n64) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U75 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n3), .B(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n64), .Z(EXEC_STAGE_mul_ex_N173) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U74 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n62), .A2(EXEC_STAGE_mul_ex_mult_88_n33), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n58) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U73 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n62), .A2(EXEC_STAGE_mul_ex_mult_88_n33), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n60) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U72 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n10), .A2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n60), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n61) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U71 ( .B1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n9), .B2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n3), .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n59) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U70 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n61), .B(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n59), .Z(EXEC_STAGE_mul_ex_N174) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U69 ( .B1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n58), .B2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n59), .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n60), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n54) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U68 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n55), .A2(EXEC_STAGE_mul_ex_mult_88_n25), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n55) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U67 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n55), .A2(EXEC_STAGE_mul_ex_mult_88_n25), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n56) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U66 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n55), .A2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n56), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n57) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U65 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n54), .B(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n57), .Z(EXEC_STAGE_mul_ex_N175) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U64 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n61), .A2(EXEC_STAGE_mul_ex_mult_88_n32), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n50) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U63 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n61), .A2(EXEC_STAGE_mul_ex_mult_88_n32), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n52) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U62 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n12), .A2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n53) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U61 ( .B1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n11), .B2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n54), .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n55), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n51) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U60 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n53), .B(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n51), .Z(EXEC_STAGE_mul_ex_N176) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U59 ( .B1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n50), .B2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n51), .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n46) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U58 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n54), .A2(EXEC_STAGE_mul_ex_mult_88_n24), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n47) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U57 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n54), .A2(EXEC_STAGE_mul_ex_mult_88_n24), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n48) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U56 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n47), .A2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n48), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n49) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U55 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n46), .B(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n49), .Z(EXEC_STAGE_mul_ex_N177) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U54 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n60), .A2(EXEC_STAGE_mul_ex_mult_88_n31), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n42) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U53 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n60), .A2(EXEC_STAGE_mul_ex_mult_88_n31), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n44) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U52 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n14), .A2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n44), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n45) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U51 ( .B1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n13), .B2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n46), .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n47), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n43) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U50 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n45), .B(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n43), .Z(EXEC_STAGE_mul_ex_N178) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U49 ( .B1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n42), .B2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n43), .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n44), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n38) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U48 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n53), .A2(EXEC_STAGE_mul_ex_mult_88_n23), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n39) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U47 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n53), .A2(EXEC_STAGE_mul_ex_mult_88_n23), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n40) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U46 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n39), .A2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n40), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n41) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U45 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n38), .B(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n41), .Z(EXEC_STAGE_mul_ex_N179) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U44 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n59), .A2(EXEC_STAGE_mul_ex_mult_88_n30), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n34) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U43 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n59), .A2(EXEC_STAGE_mul_ex_mult_88_n30), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n36) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U42 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n6), .A2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n36), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n37) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U41 ( .B1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n15), .B2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n38), .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n39), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n35) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U40 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n37), .B(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n35), .Z(EXEC_STAGE_mul_ex_N180) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U39 ( .B1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n34), .B2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n35), .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n36), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n30) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U38 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n52), .A2(EXEC_STAGE_mul_ex_mult_88_n22), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n31) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U37 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n52), .A2(EXEC_STAGE_mul_ex_mult_88_n22), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n32) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U36 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n31), .A2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n32), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n33) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U35 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n30), .B(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n33), .Z(EXEC_STAGE_mul_ex_N181) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U34 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n58), .A2(EXEC_STAGE_mul_ex_mult_88_n29), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n26) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U33 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n58), .A2(EXEC_STAGE_mul_ex_mult_88_n29), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n28) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U32 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n4), .A2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n28), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n29) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U31 ( .B1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n5), .B2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n30), .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n31), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n27) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U30 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n29), .B(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n27), .Z(EXEC_STAGE_mul_ex_N182) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U29 ( .B1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n26), .B2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n27), .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n28), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n22) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U28 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n51), .A2(EXEC_STAGE_mul_ex_mult_88_n21), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n23) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U27 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n51), .A2(EXEC_STAGE_mul_ex_mult_88_n21), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n24) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U26 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n23), .A2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n24), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n25) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U25 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n22), .B(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n25), .Z(EXEC_STAGE_mul_ex_N183) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U24 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n57), .A2(EXEC_STAGE_mul_ex_mult_88_n28), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n18) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U23 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_n57), .A2(EXEC_STAGE_mul_ex_mult_88_n28), 
        .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n20) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U22 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n8), .A2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n20), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n21) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U21 ( .B1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n7), .B2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n22), .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n23), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n19) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U20 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n21), .B(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n19), .Z(EXEC_STAGE_mul_ex_N184) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U19 ( .B1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n18), .B2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n19), .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n20), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n16) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U18 ( .A(
        EXEC_STAGE_mul_ex_mult_88_n65), .B(EXEC_STAGE_mul_ex_mult_88_n34), .Z(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n17) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_88_FS_1_U17 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n16), .B(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n17), .Z(EXEC_STAGE_mul_ex_N185) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_FS_1_U16 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n40), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n15) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_FS_1_U15 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n42), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n14) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_FS_1_U14 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n48), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n13) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_FS_1_U13 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n50), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n12) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_FS_1_U12 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n56), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n11) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_FS_1_U11 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n58), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n10) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_FS_1_U10 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n9) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_FS_1_U9 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n18), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n8) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_FS_1_U8 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n24), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n7) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_FS_1_U7 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n34), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n6) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_FS_1_U6 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n32), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n5) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_FS_1_U5 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n26), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n4) );
  INV_X4 EXEC_STAGE_mul_ex_mult_88_FS_1_U4 ( .A(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n3) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_88_FS_1_U3 ( .A1(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n1), .A2(
        EXEC_STAGE_mul_ex_mult_88_FS_1_n65), .ZN(EXEC_STAGE_mul_ex_N172) );
  OR2_X4 EXEC_STAGE_mul_ex_mult_88_FS_1_U2 ( .A1(EXEC_STAGE_mul_ex_mult_88_n63), .A2(EXEC_STAGE_mul_ex_mult_88_n27), .ZN(EXEC_STAGE_mul_ex_mult_88_FS_1_n1)
         );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U35 ( .A(
        EXEC_STAGE_mul_ex_L_31_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n33) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U34 ( .A(
        EXEC_STAGE_mul_ex_L_30_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n32) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U33 ( .A(
        EXEC_STAGE_mul_ex_L_29_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n31) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U32 ( .A(
        EXEC_STAGE_mul_ex_L_28_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n30) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U31 ( .A(
        EXEC_STAGE_mul_ex_L_27_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n29) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U30 ( .A(
        EXEC_STAGE_mul_ex_L_26_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n28) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U29 ( .A(
        EXEC_STAGE_mul_ex_L_25_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n27) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U28 ( .A(
        EXEC_STAGE_mul_ex_L_24_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n26) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U27 ( .A(
        EXEC_STAGE_mul_ex_L_23_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n25) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U26 ( .A(
        EXEC_STAGE_mul_ex_L_22_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n24) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U25 ( .A(
        EXEC_STAGE_mul_ex_L_21_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n23) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U24 ( .A(
        EXEC_STAGE_mul_ex_L_20_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n22) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U23 ( .A(
        EXEC_STAGE_mul_ex_L_19_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n21) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U22 ( .A(
        EXEC_STAGE_mul_ex_L_18_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n20) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U21 ( .A(
        EXEC_STAGE_mul_ex_L_17_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n19) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U20 ( .A(
        EXEC_STAGE_mul_ex_L_16_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n18) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U19 ( .A(
        EXEC_STAGE_mul_ex_L_15_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n17) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U18 ( .A(
        EXEC_STAGE_mul_ex_L_14_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n16) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U17 ( .A(
        EXEC_STAGE_mul_ex_L_13_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n15) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U16 ( .A(
        EXEC_STAGE_mul_ex_L_12_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n14) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U15 ( .A(
        EXEC_STAGE_mul_ex_L_11_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n13) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U14 ( .A(
        EXEC_STAGE_mul_ex_L_10_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n12) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U13 ( .A(
        EXEC_STAGE_mul_ex_L_9_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n11) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U12 ( .A(
        EXEC_STAGE_mul_ex_L_8_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n10) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U11 ( .A(
        EXEC_STAGE_mul_ex_L_7_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n9) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U10 ( .A(
        EXEC_STAGE_mul_ex_L_6_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n8) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U9 ( .A(
        EXEC_STAGE_mul_ex_L_5_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n7) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U8 ( .A(
        EXEC_STAGE_mul_ex_L_4_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n6) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U7 ( .A(
        EXEC_STAGE_mul_ex_L_3_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n5) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U6 ( .A(
        EXEC_STAGE_mul_ex_L_2_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n4) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U5 ( .A(
        EXEC_STAGE_mul_ex_L_1_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n3) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U4 ( .A(
        EXEC_STAGE_mul_ex_L_0_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n2) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U3 ( .A(
        EXEC_STAGE_mul_ex_P[31]), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n1) );
  XNOR2_X2 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2 ( .A(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n33), .B(
        EXEC_STAGE_mul_ex_P[31]), .ZN(EXEC_STAGE_mul_ex_N186) );
  NAND2_X2 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U1 ( .A1(
        EXEC_STAGE_mul_ex_L_31_), .A2(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n1), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[1]) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_1 ( .A(
        EXEC_STAGE_mul_ex_P[30]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n32), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[1]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[2]), .S(
        EXEC_STAGE_mul_ex_N187) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_2 ( .A(
        EXEC_STAGE_mul_ex_P[29]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n31), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[2]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[3]), .S(
        EXEC_STAGE_mul_ex_N188) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_3 ( .A(
        EXEC_STAGE_mul_ex_P[28]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n30), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[3]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[4]), .S(
        EXEC_STAGE_mul_ex_N189) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_4 ( .A(
        EXEC_STAGE_mul_ex_P[27]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n29), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[4]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[5]), .S(
        EXEC_STAGE_mul_ex_N190) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_5 ( .A(
        EXEC_STAGE_mul_ex_P[26]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n28), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[5]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[6]), .S(
        EXEC_STAGE_mul_ex_N191) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_6 ( .A(
        EXEC_STAGE_mul_ex_P[25]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n27), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[6]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[7]), .S(
        EXEC_STAGE_mul_ex_N192) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_7 ( .A(
        EXEC_STAGE_mul_ex_P[24]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n26), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[7]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[8]), .S(
        EXEC_STAGE_mul_ex_N193) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_8 ( .A(
        EXEC_STAGE_mul_ex_P[23]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n25), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[8]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[9]), .S(
        EXEC_STAGE_mul_ex_N194) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_9 ( .A(
        EXEC_STAGE_mul_ex_P[22]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n24), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[9]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[10]), .S(
        EXEC_STAGE_mul_ex_N195) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_10 ( .A(
        EXEC_STAGE_mul_ex_P[21]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n23), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[10]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[11]), .S(
        EXEC_STAGE_mul_ex_N196) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_11 ( .A(
        EXEC_STAGE_mul_ex_P[20]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n22), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[11]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[12]), .S(
        EXEC_STAGE_mul_ex_N197) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_12 ( .A(
        EXEC_STAGE_mul_ex_P[19]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n21), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[12]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[13]), .S(
        EXEC_STAGE_mul_ex_N198) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_13 ( .A(
        EXEC_STAGE_mul_ex_P[18]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n20), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[13]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[14]), .S(
        EXEC_STAGE_mul_ex_N199) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_14 ( .A(
        EXEC_STAGE_mul_ex_P[17]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n19), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[14]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[15]), .S(
        EXEC_STAGE_mul_ex_N200) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_15 ( .A(
        EXEC_STAGE_mul_ex_P[16]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n18), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[15]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[16]), .S(
        EXEC_STAGE_mul_ex_N201) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_16 ( .A(
        EXEC_STAGE_mul_ex_P[15]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n17), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[16]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[17]), .S(
        EXEC_STAGE_mul_ex_N202) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_17 ( .A(
        EXEC_STAGE_mul_ex_P[14]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n16), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[17]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[18]), .S(
        EXEC_STAGE_mul_ex_N203) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_18 ( .A(
        EXEC_STAGE_mul_ex_P[13]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n15), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[18]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[19]), .S(
        EXEC_STAGE_mul_ex_N204) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_19 ( .A(
        EXEC_STAGE_mul_ex_P[12]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n14), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[19]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[20]), .S(
        EXEC_STAGE_mul_ex_N205) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_20 ( .A(
        EXEC_STAGE_mul_ex_P[11]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n13), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[20]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[21]), .S(
        EXEC_STAGE_mul_ex_N206) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_21 ( .A(
        EXEC_STAGE_mul_ex_P[10]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n12), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[21]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[22]), .S(
        EXEC_STAGE_mul_ex_N207) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_22 ( .A(
        EXEC_STAGE_mul_ex_P[9]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n11), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[22]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[23]), .S(
        EXEC_STAGE_mul_ex_N208) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_23 ( .A(
        EXEC_STAGE_mul_ex_P[8]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n10), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[23]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[24]), .S(
        EXEC_STAGE_mul_ex_N209) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_24 ( .A(
        EXEC_STAGE_mul_ex_P[7]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n9), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[24]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[25]), .S(
        EXEC_STAGE_mul_ex_N210) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_25 ( .A(
        EXEC_STAGE_mul_ex_P[6]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n8), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[25]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[26]), .S(
        EXEC_STAGE_mul_ex_N211) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_26 ( .A(
        EXEC_STAGE_mul_ex_P[5]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n7), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[26]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[27]), .S(
        EXEC_STAGE_mul_ex_N212) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_27 ( .A(
        EXEC_STAGE_mul_ex_P[4]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n6), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[27]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[28]), .S(
        EXEC_STAGE_mul_ex_N213) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_28 ( .A(
        EXEC_STAGE_mul_ex_P[3]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n5), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[28]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[29]), .S(
        EXEC_STAGE_mul_ex_N214) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_29 ( .A(
        EXEC_STAGE_mul_ex_P[2]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n4), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[29]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[30]), .S(
        EXEC_STAGE_mul_ex_N215) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_30 ( .A(
        EXEC_STAGE_mul_ex_P[1]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n3), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[30]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[31]), .S(
        EXEC_STAGE_mul_ex_N216) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_31 ( .A(
        EXEC_STAGE_mul_ex_P[0]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n2), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[31]), .S(
        EXEC_STAGE_mul_ex_N217) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U35 ( .A(
        EXEC_STAGE_mul_ex_H[0]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n33) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U34 ( .A(
        EXEC_STAGE_mul_ex_H[1]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n32) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U33 ( .A(
        EXEC_STAGE_mul_ex_H[2]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n31) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U32 ( .A(
        EXEC_STAGE_mul_ex_H[3]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n30) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U31 ( .A(
        EXEC_STAGE_mul_ex_H[4]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n29) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U30 ( .A(
        EXEC_STAGE_mul_ex_H[5]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n28) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U29 ( .A(
        EXEC_STAGE_mul_ex_H[6]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n27) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U28 ( .A(
        EXEC_STAGE_mul_ex_H[7]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n26) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U27 ( .A(
        EXEC_STAGE_mul_ex_H[8]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n25) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U26 ( .A(
        EXEC_STAGE_mul_ex_H[9]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n24) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U25 ( .A(
        EXEC_STAGE_mul_ex_H[10]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n23) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U24 ( .A(
        EXEC_STAGE_mul_ex_H[11]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n22) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U23 ( .A(
        EXEC_STAGE_mul_ex_H[12]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n21) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U22 ( .A(
        EXEC_STAGE_mul_ex_H[13]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n20) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U21 ( .A(
        EXEC_STAGE_mul_ex_H[14]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n19) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U20 ( .A(
        EXEC_STAGE_mul_ex_H[15]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n18) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U19 ( .A(
        EXEC_STAGE_mul_ex_H[16]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n17) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U18 ( .A(
        EXEC_STAGE_mul_ex_H[17]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n16) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U17 ( .A(
        EXEC_STAGE_mul_ex_H[18]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n15) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U16 ( .A(
        EXEC_STAGE_mul_ex_H[19]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n14) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U15 ( .A(
        EXEC_STAGE_mul_ex_H[20]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n13) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U14 ( .A(
        EXEC_STAGE_mul_ex_H[21]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n12) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U13 ( .A(
        EXEC_STAGE_mul_ex_H[22]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n11) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U12 ( .A(
        EXEC_STAGE_mul_ex_H[23]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n10) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U11 ( .A(
        EXEC_STAGE_mul_ex_H[24]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n9) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U10 ( .A(
        EXEC_STAGE_mul_ex_H[25]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n8) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U9 ( .A(
        EXEC_STAGE_mul_ex_H[26]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n7) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U8 ( .A(
        EXEC_STAGE_mul_ex_H[27]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n6) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U7 ( .A(
        EXEC_STAGE_mul_ex_H[28]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n5) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U6 ( .A(
        EXEC_STAGE_mul_ex_H[29]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n4) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U5 ( .A(
        EXEC_STAGE_mul_ex_H[30]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n3) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U4 ( .A(
        EXEC_STAGE_mul_ex_H[31]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n2) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U3 ( .A(
        EXEC_STAGE_mul_ex_N186), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n1) );
  XNOR2_X2 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2 ( .A(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n2), .B(
        EXEC_STAGE_mul_ex_N186), .ZN(EXEC_STAGE_mul_ex_N218) );
  NAND2_X2 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U1 ( .A1(
        EXEC_STAGE_mul_ex_H[31]), .A2(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n1), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[1]) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_1 ( .A(
        EXEC_STAGE_mul_ex_N187), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n3), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[1]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[2]), .S(
        EXEC_STAGE_mul_ex_N219) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_2 ( .A(
        EXEC_STAGE_mul_ex_N188), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n4), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[2]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[3]), .S(
        EXEC_STAGE_mul_ex_N220) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_3 ( .A(
        EXEC_STAGE_mul_ex_N189), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n5), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[3]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[4]), .S(
        EXEC_STAGE_mul_ex_N221) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_4 ( .A(
        EXEC_STAGE_mul_ex_N190), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n6), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[4]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[5]), .S(
        EXEC_STAGE_mul_ex_N222) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_5 ( .A(
        EXEC_STAGE_mul_ex_N191), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n7), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[5]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[6]), .S(
        EXEC_STAGE_mul_ex_N223) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_6 ( .A(
        EXEC_STAGE_mul_ex_N192), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n8), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[6]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[7]), .S(
        EXEC_STAGE_mul_ex_N224) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_7 ( .A(
        EXEC_STAGE_mul_ex_N193), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n9), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[7]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[8]), .S(
        EXEC_STAGE_mul_ex_N225) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_8 ( .A(
        EXEC_STAGE_mul_ex_N194), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n10), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[8]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[9]), .S(
        EXEC_STAGE_mul_ex_N226) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_9 ( .A(
        EXEC_STAGE_mul_ex_N195), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n11), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[9]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[10]), .S(
        EXEC_STAGE_mul_ex_N227) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_10 ( .A(
        EXEC_STAGE_mul_ex_N196), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n12), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[10]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[11]), .S(
        EXEC_STAGE_mul_ex_N228) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_11 ( .A(
        EXEC_STAGE_mul_ex_N197), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n13), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[11]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[12]), .S(
        EXEC_STAGE_mul_ex_N229) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_12 ( .A(
        EXEC_STAGE_mul_ex_N198), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n14), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[12]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[13]), .S(
        EXEC_STAGE_mul_ex_N230) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_13 ( .A(
        EXEC_STAGE_mul_ex_N199), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n15), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[13]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[14]), .S(
        EXEC_STAGE_mul_ex_N231) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_14 ( .A(
        EXEC_STAGE_mul_ex_N200), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n16), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[14]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[15]), .S(
        EXEC_STAGE_mul_ex_N232) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_15 ( .A(
        EXEC_STAGE_mul_ex_N201), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n17), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[15]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[16]), .S(
        EXEC_STAGE_mul_ex_N233) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_16 ( .A(
        EXEC_STAGE_mul_ex_N202), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n18), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[16]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[17]), .S(
        EXEC_STAGE_mul_ex_N234) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_17 ( .A(
        EXEC_STAGE_mul_ex_N203), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n19), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[17]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[18]), .S(
        EXEC_STAGE_mul_ex_N235) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_18 ( .A(
        EXEC_STAGE_mul_ex_N204), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n20), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[18]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[19]), .S(
        EXEC_STAGE_mul_ex_N236) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_19 ( .A(
        EXEC_STAGE_mul_ex_N205), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n21), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[19]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[20]), .S(
        EXEC_STAGE_mul_ex_N237) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_20 ( .A(
        EXEC_STAGE_mul_ex_N206), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n22), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[20]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[21]), .S(
        EXEC_STAGE_mul_ex_N238) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_21 ( .A(
        EXEC_STAGE_mul_ex_N207), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n23), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[21]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[22]), .S(
        EXEC_STAGE_mul_ex_N239) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_22 ( .A(
        EXEC_STAGE_mul_ex_N208), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n24), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[22]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[23]), .S(
        EXEC_STAGE_mul_ex_N240) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_23 ( .A(
        EXEC_STAGE_mul_ex_N209), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n25), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[23]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[24]), .S(
        EXEC_STAGE_mul_ex_N241) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_24 ( .A(
        EXEC_STAGE_mul_ex_N210), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n26), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[24]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[25]), .S(
        EXEC_STAGE_mul_ex_N242) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_25 ( .A(
        EXEC_STAGE_mul_ex_N211), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n27), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[25]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[26]), .S(
        EXEC_STAGE_mul_ex_N243) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_26 ( .A(
        EXEC_STAGE_mul_ex_N212), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n28), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[26]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[27]), .S(
        EXEC_STAGE_mul_ex_N244) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_27 ( .A(
        EXEC_STAGE_mul_ex_N213), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n29), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[27]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[28]), .S(
        EXEC_STAGE_mul_ex_N245) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_28 ( .A(
        EXEC_STAGE_mul_ex_N214), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n30), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[28]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[29]), .S(
        EXEC_STAGE_mul_ex_N246) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_29 ( .A(
        EXEC_STAGE_mul_ex_N215), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n31), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[29]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[30]), .S(
        EXEC_STAGE_mul_ex_N247) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_30 ( .A(
        EXEC_STAGE_mul_ex_N216), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n32), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[30]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[31]), .S(
        EXEC_STAGE_mul_ex_N248) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_U2_31 ( .A(
        EXEC_STAGE_mul_ex_N217), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_n33), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_92_2_carry[31]), .S(
        EXEC_STAGE_mul_ex_N249) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U50 ( .A(
        EXEC_STAGE_mul_ex_L_31_), .Z(EXEC_STAGE_mul_ex_N250) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U49 ( .A(
        EXEC_STAGE_mul_ex_L_30_), .Z(EXEC_STAGE_mul_ex_N251) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U48 ( .A(
        EXEC_STAGE_mul_ex_L_29_), .Z(EXEC_STAGE_mul_ex_N252) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U47 ( .A(
        EXEC_STAGE_mul_ex_L_28_), .Z(EXEC_STAGE_mul_ex_N253) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U46 ( .A(
        EXEC_STAGE_mul_ex_L_27_), .Z(EXEC_STAGE_mul_ex_N254) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U45 ( .A(
        EXEC_STAGE_mul_ex_L_26_), .Z(EXEC_STAGE_mul_ex_N255) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U44 ( .A(
        EXEC_STAGE_mul_ex_L_25_), .Z(EXEC_STAGE_mul_ex_N256) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U43 ( .A(
        EXEC_STAGE_mul_ex_L_24_), .Z(EXEC_STAGE_mul_ex_N257) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U42 ( .A(
        EXEC_STAGE_mul_ex_L_23_), .Z(EXEC_STAGE_mul_ex_N258) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U41 ( .A(
        EXEC_STAGE_mul_ex_L_22_), .Z(EXEC_STAGE_mul_ex_N259) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U40 ( .A(
        EXEC_STAGE_mul_ex_L_21_), .Z(EXEC_STAGE_mul_ex_N260) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U39 ( .A(
        EXEC_STAGE_mul_ex_L_20_), .Z(EXEC_STAGE_mul_ex_N261) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U38 ( .A(
        EXEC_STAGE_mul_ex_L_19_), .Z(EXEC_STAGE_mul_ex_N262) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U37 ( .A(
        EXEC_STAGE_mul_ex_L_18_), .Z(EXEC_STAGE_mul_ex_N263) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U36 ( .A(
        EXEC_STAGE_mul_ex_L_17_), .Z(EXEC_STAGE_mul_ex_N264) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U35 ( .A(
        EXEC_STAGE_mul_ex_L_16_), .Z(EXEC_STAGE_mul_ex_N265) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U34 ( .A(
        EXEC_STAGE_mul_ex_Z_31_), .B(EXEC_STAGE_mul_ex_L_15_), .Z(
        EXEC_STAGE_mul_ex_N266) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U33 ( .A1(
        EXEC_STAGE_mul_ex_Z_31_), .A2(EXEC_STAGE_mul_ex_L_15_), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n33) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U32 ( .A1(
        EXEC_STAGE_mul_ex_Z_0_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n10), .ZN(
        EXEC_STAGE_mul_ex_N298) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U31 ( .A(
        EXEC_STAGE_mul_ex_Z_0_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n10), .Z(
        EXEC_STAGE_mul_ex_N297) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U30 ( .A(
        EXEC_STAGE_mul_ex_Z_1_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n3), .Z(
        EXEC_STAGE_mul_ex_N296) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U29 ( .A(
        EXEC_STAGE_mul_ex_Z_2_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n11), .Z(
        EXEC_STAGE_mul_ex_N295) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U28 ( .A(
        EXEC_STAGE_mul_ex_Z_3_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n4), .Z(
        EXEC_STAGE_mul_ex_N294) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U27 ( .A(
        EXEC_STAGE_mul_ex_Z_4_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n12), .Z(
        EXEC_STAGE_mul_ex_N293) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U26 ( .A(
        EXEC_STAGE_mul_ex_Z_5_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n5), .Z(
        EXEC_STAGE_mul_ex_N292) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U25 ( .A(
        EXEC_STAGE_mul_ex_Z_6_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n13), .Z(
        EXEC_STAGE_mul_ex_N291) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U24 ( .A(
        EXEC_STAGE_mul_ex_Z_7_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n6), .Z(
        EXEC_STAGE_mul_ex_N290) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U23 ( .A(
        EXEC_STAGE_mul_ex_Z_8_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n14), .Z(
        EXEC_STAGE_mul_ex_N289) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U22 ( .A(
        EXEC_STAGE_mul_ex_Z_9_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n7), .Z(
        EXEC_STAGE_mul_ex_N288) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U21 ( .A(
        EXEC_STAGE_mul_ex_Z_10_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n15), .Z(
        EXEC_STAGE_mul_ex_N287) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U20 ( .A(
        EXEC_STAGE_mul_ex_Z_11_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n2), .Z(
        EXEC_STAGE_mul_ex_N286) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U19 ( .A(
        EXEC_STAGE_mul_ex_Z_12_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n16), .Z(
        EXEC_STAGE_mul_ex_N285) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U18 ( .A(
        EXEC_STAGE_mul_ex_Z_13_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n8), .Z(
        EXEC_STAGE_mul_ex_N284) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U17 ( .A1(
        EXEC_STAGE_mul_ex_Z_15_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_32_), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n17) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U16 ( .A1(
        EXEC_STAGE_mul_ex_Z_13_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n8), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n16) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U15 ( .A1(
        EXEC_STAGE_mul_ex_Z_11_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n2), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n15) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U14 ( .A1(
        EXEC_STAGE_mul_ex_Z_9_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n7), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n14) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U13 ( .A1(
        EXEC_STAGE_mul_ex_Z_7_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n6), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n13) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U12 ( .A1(
        EXEC_STAGE_mul_ex_Z_5_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n5), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n12) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U11 ( .A1(
        EXEC_STAGE_mul_ex_Z_3_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n4), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n11) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U10 ( .A1(
        EXEC_STAGE_mul_ex_Z_1_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n3), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n10) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U9 ( .A(
        EXEC_STAGE_mul_ex_Z_15_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_32_), .Z(
        EXEC_STAGE_mul_ex_N282) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U8 ( .A1(
        EXEC_STAGE_mul_ex_Z_14_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n17), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n8) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U7 ( .A1(
        EXEC_STAGE_mul_ex_Z_10_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n15), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n7) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U6 ( .A1(
        EXEC_STAGE_mul_ex_Z_8_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n14), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n6) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U5 ( .A1(
        EXEC_STAGE_mul_ex_Z_6_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n13), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n5) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U4 ( .A1(
        EXEC_STAGE_mul_ex_Z_4_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n12), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n4) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U3 ( .A1(
        EXEC_STAGE_mul_ex_Z_2_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n11), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n3) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U2 ( .A1(
        EXEC_STAGE_mul_ex_Z_12_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n16), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n2) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1 ( .A(
        EXEC_STAGE_mul_ex_Z_14_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n17), .Z(
        EXEC_STAGE_mul_ex_N283) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_17 ( .A(
        EXEC_STAGE_mul_ex_L_14_), .B(EXEC_STAGE_mul_ex_Z_30_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n33), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_18_), .S(
        EXEC_STAGE_mul_ex_N267) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_18 ( .A(
        EXEC_STAGE_mul_ex_L_13_), .B(EXEC_STAGE_mul_ex_Z_29_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_18_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_19_), .S(
        EXEC_STAGE_mul_ex_N268) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_19 ( .A(
        EXEC_STAGE_mul_ex_L_12_), .B(EXEC_STAGE_mul_ex_Z_28_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_19_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_20_), .S(
        EXEC_STAGE_mul_ex_N269) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_20 ( .A(
        EXEC_STAGE_mul_ex_L_11_), .B(EXEC_STAGE_mul_ex_Z_27_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_20_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_21_), .S(
        EXEC_STAGE_mul_ex_N270) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_21 ( .A(
        EXEC_STAGE_mul_ex_L_10_), .B(EXEC_STAGE_mul_ex_Z_26_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_21_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_22_), .S(
        EXEC_STAGE_mul_ex_N271) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_22 ( .A(
        EXEC_STAGE_mul_ex_L_9_), .B(EXEC_STAGE_mul_ex_Z_25_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_22_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_23_), .S(
        EXEC_STAGE_mul_ex_N272) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_23 ( .A(
        EXEC_STAGE_mul_ex_L_8_), .B(EXEC_STAGE_mul_ex_Z_24_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_23_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_24_), .S(
        EXEC_STAGE_mul_ex_N273) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_24 ( .A(
        EXEC_STAGE_mul_ex_L_7_), .B(EXEC_STAGE_mul_ex_Z_23_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_24_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_25_), .S(
        EXEC_STAGE_mul_ex_N274) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_25 ( .A(
        EXEC_STAGE_mul_ex_L_6_), .B(EXEC_STAGE_mul_ex_Z_22_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_25_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_26_), .S(
        EXEC_STAGE_mul_ex_N275) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_26 ( .A(
        EXEC_STAGE_mul_ex_L_5_), .B(EXEC_STAGE_mul_ex_Z_21_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_26_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_27_), .S(
        EXEC_STAGE_mul_ex_N276) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_27 ( .A(
        EXEC_STAGE_mul_ex_L_4_), .B(EXEC_STAGE_mul_ex_Z_20_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_27_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_28_), .S(
        EXEC_STAGE_mul_ex_N277) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_28 ( .A(
        EXEC_STAGE_mul_ex_L_3_), .B(EXEC_STAGE_mul_ex_Z_19_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_28_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_29_), .S(
        EXEC_STAGE_mul_ex_N278) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_29 ( .A(
        EXEC_STAGE_mul_ex_L_2_), .B(EXEC_STAGE_mul_ex_Z_18_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_29_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_30_), .S(
        EXEC_STAGE_mul_ex_N279) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_30 ( .A(
        EXEC_STAGE_mul_ex_L_1_), .B(EXEC_STAGE_mul_ex_Z_17_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_30_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_31_), .S(
        EXEC_STAGE_mul_ex_N280) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_31 ( .A(
        EXEC_STAGE_mul_ex_L_0_), .B(EXEC_STAGE_mul_ex_Z_16_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_31_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_32_), .S(
        EXEC_STAGE_mul_ex_N281) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U63 ( .A(
        EXEC_STAGE_mul_ex_N274), .Z(EXEC_STAGE_mul_ex_N338) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U62 ( .A(
        EXEC_STAGE_mul_ex_N273), .Z(EXEC_STAGE_mul_ex_N337) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U61 ( .A(
        EXEC_STAGE_mul_ex_N272), .Z(EXEC_STAGE_mul_ex_N336) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U60 ( .A(
        EXEC_STAGE_mul_ex_N271), .Z(EXEC_STAGE_mul_ex_N335) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U59 ( .A(
        EXEC_STAGE_mul_ex_N270), .Z(EXEC_STAGE_mul_ex_N334) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U58 ( .A(
        EXEC_STAGE_mul_ex_N269), .Z(EXEC_STAGE_mul_ex_N333) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U57 ( .A(
        EXEC_STAGE_mul_ex_N268), .Z(EXEC_STAGE_mul_ex_N332) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U56 ( .A(
        EXEC_STAGE_mul_ex_N267), .Z(EXEC_STAGE_mul_ex_N331) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U55 ( .A(
        EXEC_STAGE_mul_ex_N266), .Z(EXEC_STAGE_mul_ex_N330) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U54 ( .A(
        EXEC_STAGE_mul_ex_N265), .Z(EXEC_STAGE_mul_ex_N329) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U53 ( .A(
        EXEC_STAGE_mul_ex_N264), .Z(EXEC_STAGE_mul_ex_N328) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U52 ( .A(
        EXEC_STAGE_mul_ex_N263), .Z(EXEC_STAGE_mul_ex_N327) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U51 ( .A(
        EXEC_STAGE_mul_ex_N262), .Z(EXEC_STAGE_mul_ex_N326) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U50 ( .A(
        EXEC_STAGE_mul_ex_N261), .Z(EXEC_STAGE_mul_ex_N325) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U49 ( .A(
        EXEC_STAGE_mul_ex_N260), .Z(EXEC_STAGE_mul_ex_N324) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U48 ( .A(
        EXEC_STAGE_mul_ex_N259), .Z(EXEC_STAGE_mul_ex_N323) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U47 ( .A(
        EXEC_STAGE_mul_ex_N258), .Z(EXEC_STAGE_mul_ex_N322) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U46 ( .A(
        EXEC_STAGE_mul_ex_N257), .Z(EXEC_STAGE_mul_ex_N321) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U45 ( .A(
        EXEC_STAGE_mul_ex_N256), .Z(EXEC_STAGE_mul_ex_N320) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U44 ( .A(
        EXEC_STAGE_mul_ex_N255), .Z(EXEC_STAGE_mul_ex_N319) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U43 ( .A(
        EXEC_STAGE_mul_ex_N254), .Z(EXEC_STAGE_mul_ex_N318) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U42 ( .A(
        EXEC_STAGE_mul_ex_N253), .Z(EXEC_STAGE_mul_ex_N317) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U41 ( .A(
        EXEC_STAGE_mul_ex_N252), .Z(EXEC_STAGE_mul_ex_N316) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U40 ( .A(
        EXEC_STAGE_mul_ex_N251), .Z(EXEC_STAGE_mul_ex_N315) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U39 ( .A(
        EXEC_STAGE_mul_ex_N250), .Z(EXEC_STAGE_mul_ex_N314) );
  BUF_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U38 ( .A(
        EXEC_STAGE_mul_ex_N275), .Z(EXEC_STAGE_mul_ex_N339) );
  BUF_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U37 ( .A(
        EXEC_STAGE_mul_ex_N276), .Z(EXEC_STAGE_mul_ex_N340) );
  BUF_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U36 ( .A(
        EXEC_STAGE_mul_ex_N277), .Z(EXEC_STAGE_mul_ex_N341) );
  BUF_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U35 ( .A(
        EXEC_STAGE_mul_ex_N278), .Z(EXEC_STAGE_mul_ex_N342) );
  BUF_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U34 ( .A(
        EXEC_STAGE_mul_ex_N279), .Z(EXEC_STAGE_mul_ex_N343) );
  BUF_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U33 ( .A(
        EXEC_STAGE_mul_ex_N280), .Z(EXEC_STAGE_mul_ex_N344) );
  BUF_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U32 ( .A(
        EXEC_STAGE_mul_ex_N281), .Z(EXEC_STAGE_mul_ex_N345) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U31 ( .A(
        EXEC_STAGE_mul_ex_Z_0_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n25), .Z(
        EXEC_STAGE_mul_ex_N377) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U30 ( .A(
        EXEC_STAGE_mul_ex_Z_11_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n22), .Z(
        EXEC_STAGE_mul_ex_N366) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U29 ( .A(
        EXEC_STAGE_mul_ex_Z_12_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n1), .Z(
        EXEC_STAGE_mul_ex_N365) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U28 ( .A(
        EXEC_STAGE_mul_ex_Z_13_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n23), .Z(
        EXEC_STAGE_mul_ex_N364) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U27 ( .A(
        EXEC_STAGE_mul_ex_N282), .B(EXEC_STAGE_mul_ex_Z_31_), .Z(
        EXEC_STAGE_mul_ex_N346) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U26 ( .A(
        EXEC_STAGE_mul_ex_Z_14_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_49_), .Z(
        EXEC_STAGE_mul_ex_N363) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U25 ( .A1(
        EXEC_STAGE_mul_ex_Z_1_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n17), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n25) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U24 ( .A1(
        EXEC_STAGE_mul_ex_N282), .A2(EXEC_STAGE_mul_ex_Z_31_), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n24) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U23 ( .A1(
        EXEC_STAGE_mul_ex_Z_14_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_49_), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n23) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U22 ( .A1(
        EXEC_STAGE_mul_ex_Z_12_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n1), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n22) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U21 ( .A1(
        EXEC_STAGE_mul_ex_Z_10_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n2), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n21) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U20 ( .A1(
        EXEC_STAGE_mul_ex_Z_8_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n6), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n20) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U19 ( .A1(
        EXEC_STAGE_mul_ex_Z_6_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n5), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n19) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U18 ( .A1(
        EXEC_STAGE_mul_ex_Z_4_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n4), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n18) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U17 ( .A1(
        EXEC_STAGE_mul_ex_Z_2_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n3), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n17) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U16 ( .A(
        EXEC_STAGE_mul_ex_Z_1_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n17), .Z(
        EXEC_STAGE_mul_ex_N376) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U15 ( .A(
        EXEC_STAGE_mul_ex_Z_2_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n3), .Z(
        EXEC_STAGE_mul_ex_N375) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U14 ( .A(
        EXEC_STAGE_mul_ex_Z_3_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n18), .Z(
        EXEC_STAGE_mul_ex_N374) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U13 ( .A(
        EXEC_STAGE_mul_ex_Z_4_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n4), .Z(
        EXEC_STAGE_mul_ex_N373) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U12 ( .A(
        EXEC_STAGE_mul_ex_Z_5_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n19), .Z(
        EXEC_STAGE_mul_ex_N372) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U11 ( .A(
        EXEC_STAGE_mul_ex_Z_6_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n5), .Z(
        EXEC_STAGE_mul_ex_N371) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U10 ( .A(
        EXEC_STAGE_mul_ex_Z_7_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n20), .Z(
        EXEC_STAGE_mul_ex_N370) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U9 ( .A(
        EXEC_STAGE_mul_ex_Z_8_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n6), .Z(
        EXEC_STAGE_mul_ex_N369) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U8 ( .A(
        EXEC_STAGE_mul_ex_Z_9_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n21), .Z(
        EXEC_STAGE_mul_ex_N368) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U7 ( .A(
        EXEC_STAGE_mul_ex_Z_10_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n2), .Z(
        EXEC_STAGE_mul_ex_N367) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U6 ( .A1(
        EXEC_STAGE_mul_ex_Z_9_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n21), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n6) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U5 ( .A1(
        EXEC_STAGE_mul_ex_Z_7_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n20), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n5) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U4 ( .A1(
        EXEC_STAGE_mul_ex_Z_5_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n19), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n4) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U3 ( .A1(
        EXEC_STAGE_mul_ex_Z_3_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n18), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n3) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U2 ( .A1(
        EXEC_STAGE_mul_ex_Z_11_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n22), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n2) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1 ( .A1(
        EXEC_STAGE_mul_ex_Z_13_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n23), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n1) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_33 ( .A(
        EXEC_STAGE_mul_ex_Z_30_), .B(EXEC_STAGE_mul_ex_N283), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_n24), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_34_), .S(
        EXEC_STAGE_mul_ex_N347) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_34 ( .A(
        EXEC_STAGE_mul_ex_Z_29_), .B(EXEC_STAGE_mul_ex_N284), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_34_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_35_), .S(
        EXEC_STAGE_mul_ex_N348) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_35 ( .A(
        EXEC_STAGE_mul_ex_Z_28_), .B(EXEC_STAGE_mul_ex_N285), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_35_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_36_), .S(
        EXEC_STAGE_mul_ex_N349) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_36 ( .A(
        EXEC_STAGE_mul_ex_Z_27_), .B(EXEC_STAGE_mul_ex_N286), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_36_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_37_), .S(
        EXEC_STAGE_mul_ex_N350) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_37 ( .A(
        EXEC_STAGE_mul_ex_Z_26_), .B(EXEC_STAGE_mul_ex_N287), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_37_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_38_), .S(
        EXEC_STAGE_mul_ex_N351) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_38 ( .A(
        EXEC_STAGE_mul_ex_Z_25_), .B(EXEC_STAGE_mul_ex_N288), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_38_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_39_), .S(
        EXEC_STAGE_mul_ex_N352) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_39 ( .A(
        EXEC_STAGE_mul_ex_Z_24_), .B(EXEC_STAGE_mul_ex_N289), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_39_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_40_), .S(
        EXEC_STAGE_mul_ex_N353) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_40 ( .A(
        EXEC_STAGE_mul_ex_Z_23_), .B(EXEC_STAGE_mul_ex_N290), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_40_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_41_), .S(
        EXEC_STAGE_mul_ex_N354) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_41 ( .A(
        EXEC_STAGE_mul_ex_Z_22_), .B(EXEC_STAGE_mul_ex_N291), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_41_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_42_), .S(
        EXEC_STAGE_mul_ex_N355) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_42 ( .A(
        EXEC_STAGE_mul_ex_Z_21_), .B(EXEC_STAGE_mul_ex_N292), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_42_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_43_), .S(
        EXEC_STAGE_mul_ex_N356) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_43 ( .A(
        EXEC_STAGE_mul_ex_Z_20_), .B(EXEC_STAGE_mul_ex_N293), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_43_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_44_), .S(
        EXEC_STAGE_mul_ex_N357) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_44 ( .A(
        EXEC_STAGE_mul_ex_Z_19_), .B(EXEC_STAGE_mul_ex_N294), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_44_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_45_), .S(
        EXEC_STAGE_mul_ex_N358) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_45 ( .A(
        EXEC_STAGE_mul_ex_Z_18_), .B(EXEC_STAGE_mul_ex_N295), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_45_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_46_), .S(
        EXEC_STAGE_mul_ex_N359) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_46 ( .A(
        EXEC_STAGE_mul_ex_Z_17_), .B(EXEC_STAGE_mul_ex_N296), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_46_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_47_), .S(
        EXEC_STAGE_mul_ex_N360) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_47 ( .A(
        EXEC_STAGE_mul_ex_Z_16_), .B(EXEC_STAGE_mul_ex_N297), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_47_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_48_), .S(
        EXEC_STAGE_mul_ex_N361) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_U1_48 ( .A(
        EXEC_STAGE_mul_ex_Z_15_), .B(EXEC_STAGE_mul_ex_N298), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_48_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_96_2_carry_49_), .S(
        EXEC_STAGE_mul_ex_N362) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U350 ( .A1(EXEC_STAGE_mul_ex_mult_84_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(EXEC_STAGE_mul_ex_N88) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U349 ( .A1(EXEC_STAGE_mul_ex_mult_84_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_0__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U348 ( .A1(EXEC_STAGE_mul_ex_mult_84_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_0__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U347 ( .A1(EXEC_STAGE_mul_ex_mult_84_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_0__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U346 ( .A1(EXEC_STAGE_mul_ex_mult_84_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_0__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U345 ( .A1(EXEC_STAGE_mul_ex_mult_84_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_0__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U344 ( .A1(EXEC_STAGE_mul_ex_mult_84_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_0__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U343 ( .A1(EXEC_STAGE_mul_ex_mult_84_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_0__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U342 ( .A1(EXEC_STAGE_mul_ex_mult_84_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_0__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U341 ( .A1(EXEC_STAGE_mul_ex_mult_84_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_0__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U340 ( .A1(EXEC_STAGE_mul_ex_mult_84_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_0__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U339 ( .A1(EXEC_STAGE_mul_ex_mult_84_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_0__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U338 ( .A1(EXEC_STAGE_mul_ex_mult_84_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_0__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U337 ( .A1(EXEC_STAGE_mul_ex_mult_84_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_0__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U336 ( .A1(EXEC_STAGE_mul_ex_mult_84_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_0__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U335 ( .A1(EXEC_STAGE_mul_ex_mult_84_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_0__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U334 ( .A1(EXEC_STAGE_mul_ex_mult_84_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U333 ( .A1(EXEC_STAGE_mul_ex_mult_84_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U332 ( .A1(EXEC_STAGE_mul_ex_mult_84_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U331 ( .A1(EXEC_STAGE_mul_ex_mult_84_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U330 ( .A1(EXEC_STAGE_mul_ex_mult_84_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U329 ( .A1(EXEC_STAGE_mul_ex_mult_84_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U328 ( .A1(EXEC_STAGE_mul_ex_mult_84_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U327 ( .A1(EXEC_STAGE_mul_ex_mult_84_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U326 ( .A1(EXEC_STAGE_mul_ex_mult_84_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U325 ( .A1(EXEC_STAGE_mul_ex_mult_84_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U324 ( .A1(EXEC_STAGE_mul_ex_mult_84_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U323 ( .A1(EXEC_STAGE_mul_ex_mult_84_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U322 ( .A1(EXEC_STAGE_mul_ex_mult_84_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U321 ( .A1(EXEC_STAGE_mul_ex_mult_84_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U320 ( .A1(EXEC_STAGE_mul_ex_mult_84_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U319 ( .A1(EXEC_STAGE_mul_ex_mult_84_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_10__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U318 ( .A1(EXEC_STAGE_mul_ex_mult_84_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U317 ( .A1(EXEC_STAGE_mul_ex_mult_84_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U316 ( .A1(EXEC_STAGE_mul_ex_mult_84_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U315 ( .A1(EXEC_STAGE_mul_ex_mult_84_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U314 ( .A1(EXEC_STAGE_mul_ex_mult_84_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U313 ( .A1(EXEC_STAGE_mul_ex_mult_84_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U312 ( .A1(EXEC_STAGE_mul_ex_mult_84_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U311 ( .A1(EXEC_STAGE_mul_ex_mult_84_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U310 ( .A1(EXEC_STAGE_mul_ex_mult_84_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U309 ( .A1(EXEC_STAGE_mul_ex_mult_84_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U308 ( .A1(EXEC_STAGE_mul_ex_mult_84_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U307 ( .A1(EXEC_STAGE_mul_ex_mult_84_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U306 ( .A1(EXEC_STAGE_mul_ex_mult_84_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U305 ( .A1(EXEC_STAGE_mul_ex_mult_84_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U304 ( .A1(EXEC_STAGE_mul_ex_mult_84_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U303 ( .A1(EXEC_STAGE_mul_ex_mult_84_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_11__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U302 ( .A1(EXEC_STAGE_mul_ex_mult_84_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U301 ( .A1(EXEC_STAGE_mul_ex_mult_84_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U300 ( .A1(EXEC_STAGE_mul_ex_mult_84_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U299 ( .A1(EXEC_STAGE_mul_ex_mult_84_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U298 ( .A1(EXEC_STAGE_mul_ex_mult_84_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U297 ( .A1(EXEC_STAGE_mul_ex_mult_84_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U296 ( .A1(EXEC_STAGE_mul_ex_mult_84_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U295 ( .A1(EXEC_STAGE_mul_ex_mult_84_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U294 ( .A1(EXEC_STAGE_mul_ex_mult_84_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U293 ( .A1(EXEC_STAGE_mul_ex_mult_84_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U292 ( .A1(EXEC_STAGE_mul_ex_mult_84_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U291 ( .A1(EXEC_STAGE_mul_ex_mult_84_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U290 ( .A1(EXEC_STAGE_mul_ex_mult_84_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U289 ( .A1(EXEC_STAGE_mul_ex_mult_84_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U288 ( .A1(EXEC_STAGE_mul_ex_mult_84_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U287 ( .A1(EXEC_STAGE_mul_ex_mult_84_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_12__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U286 ( .A1(EXEC_STAGE_mul_ex_mult_84_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U285 ( .A1(EXEC_STAGE_mul_ex_mult_84_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U284 ( .A1(EXEC_STAGE_mul_ex_mult_84_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U283 ( .A1(EXEC_STAGE_mul_ex_mult_84_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U282 ( .A1(EXEC_STAGE_mul_ex_mult_84_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U281 ( .A1(EXEC_STAGE_mul_ex_mult_84_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U280 ( .A1(EXEC_STAGE_mul_ex_mult_84_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U279 ( .A1(EXEC_STAGE_mul_ex_mult_84_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U278 ( .A1(EXEC_STAGE_mul_ex_mult_84_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U277 ( .A1(EXEC_STAGE_mul_ex_mult_84_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U276 ( .A1(EXEC_STAGE_mul_ex_mult_84_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U275 ( .A1(EXEC_STAGE_mul_ex_mult_84_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U274 ( .A1(EXEC_STAGE_mul_ex_mult_84_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U273 ( .A1(EXEC_STAGE_mul_ex_mult_84_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U272 ( .A1(EXEC_STAGE_mul_ex_mult_84_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U271 ( .A1(EXEC_STAGE_mul_ex_mult_84_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_13__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U270 ( .A1(EXEC_STAGE_mul_ex_mult_84_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U269 ( .A1(EXEC_STAGE_mul_ex_mult_84_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U268 ( .A1(EXEC_STAGE_mul_ex_mult_84_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U267 ( .A1(EXEC_STAGE_mul_ex_mult_84_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U266 ( .A1(EXEC_STAGE_mul_ex_mult_84_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U265 ( .A1(EXEC_STAGE_mul_ex_mult_84_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U264 ( .A1(EXEC_STAGE_mul_ex_mult_84_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U263 ( .A1(EXEC_STAGE_mul_ex_mult_84_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U262 ( .A1(EXEC_STAGE_mul_ex_mult_84_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U261 ( .A1(EXEC_STAGE_mul_ex_mult_84_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U260 ( .A1(EXEC_STAGE_mul_ex_mult_84_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U259 ( .A1(EXEC_STAGE_mul_ex_mult_84_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U258 ( .A1(EXEC_STAGE_mul_ex_mult_84_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U257 ( .A1(EXEC_STAGE_mul_ex_mult_84_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U256 ( .A1(EXEC_STAGE_mul_ex_mult_84_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U255 ( .A1(EXEC_STAGE_mul_ex_mult_84_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_14__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U254 ( .A1(EXEC_STAGE_mul_ex_mult_84_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U253 ( .A1(EXEC_STAGE_mul_ex_mult_84_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U252 ( .A1(EXEC_STAGE_mul_ex_mult_84_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U251 ( .A1(EXEC_STAGE_mul_ex_mult_84_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U250 ( .A1(EXEC_STAGE_mul_ex_mult_84_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U249 ( .A1(EXEC_STAGE_mul_ex_mult_84_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U248 ( .A1(EXEC_STAGE_mul_ex_mult_84_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U247 ( .A1(EXEC_STAGE_mul_ex_mult_84_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U246 ( .A1(EXEC_STAGE_mul_ex_mult_84_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U245 ( .A1(EXEC_STAGE_mul_ex_mult_84_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U244 ( .A1(EXEC_STAGE_mul_ex_mult_84_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U243 ( .A1(EXEC_STAGE_mul_ex_mult_84_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U242 ( .A1(EXEC_STAGE_mul_ex_mult_84_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U241 ( .A1(EXEC_STAGE_mul_ex_mult_84_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U240 ( .A1(EXEC_STAGE_mul_ex_mult_84_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U239 ( .A1(EXEC_STAGE_mul_ex_mult_84_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_15__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U238 ( .A1(EXEC_STAGE_mul_ex_mult_84_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U237 ( .A1(EXEC_STAGE_mul_ex_mult_84_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U236 ( .A1(EXEC_STAGE_mul_ex_mult_84_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U235 ( .A1(EXEC_STAGE_mul_ex_mult_84_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U234 ( .A1(EXEC_STAGE_mul_ex_mult_84_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U233 ( .A1(EXEC_STAGE_mul_ex_mult_84_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U232 ( .A1(EXEC_STAGE_mul_ex_mult_84_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U231 ( .A1(EXEC_STAGE_mul_ex_mult_84_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U230 ( .A1(EXEC_STAGE_mul_ex_mult_84_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U229 ( .A1(EXEC_STAGE_mul_ex_mult_84_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U228 ( .A1(EXEC_STAGE_mul_ex_mult_84_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U227 ( .A1(EXEC_STAGE_mul_ex_mult_84_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U226 ( .A1(EXEC_STAGE_mul_ex_mult_84_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U225 ( .A1(EXEC_STAGE_mul_ex_mult_84_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U224 ( .A1(EXEC_STAGE_mul_ex_mult_84_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U223 ( .A1(EXEC_STAGE_mul_ex_mult_84_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_1__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U222 ( .A1(EXEC_STAGE_mul_ex_mult_84_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U221 ( .A1(EXEC_STAGE_mul_ex_mult_84_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U220 ( .A1(EXEC_STAGE_mul_ex_mult_84_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U219 ( .A1(EXEC_STAGE_mul_ex_mult_84_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U218 ( .A1(EXEC_STAGE_mul_ex_mult_84_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U217 ( .A1(EXEC_STAGE_mul_ex_mult_84_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U216 ( .A1(EXEC_STAGE_mul_ex_mult_84_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U215 ( .A1(EXEC_STAGE_mul_ex_mult_84_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U214 ( .A1(EXEC_STAGE_mul_ex_mult_84_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U213 ( .A1(EXEC_STAGE_mul_ex_mult_84_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U212 ( .A1(EXEC_STAGE_mul_ex_mult_84_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U211 ( .A1(EXEC_STAGE_mul_ex_mult_84_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U210 ( .A1(EXEC_STAGE_mul_ex_mult_84_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U209 ( .A1(EXEC_STAGE_mul_ex_mult_84_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U208 ( .A1(EXEC_STAGE_mul_ex_mult_84_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U207 ( .A1(EXEC_STAGE_mul_ex_mult_84_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_2__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U206 ( .A1(EXEC_STAGE_mul_ex_mult_84_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U205 ( .A1(EXEC_STAGE_mul_ex_mult_84_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U204 ( .A1(EXEC_STAGE_mul_ex_mult_84_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U203 ( .A1(EXEC_STAGE_mul_ex_mult_84_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U202 ( .A1(EXEC_STAGE_mul_ex_mult_84_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U201 ( .A1(EXEC_STAGE_mul_ex_mult_84_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U200 ( .A1(EXEC_STAGE_mul_ex_mult_84_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U199 ( .A1(EXEC_STAGE_mul_ex_mult_84_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U198 ( .A1(EXEC_STAGE_mul_ex_mult_84_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U197 ( .A1(EXEC_STAGE_mul_ex_mult_84_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U196 ( .A1(EXEC_STAGE_mul_ex_mult_84_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U195 ( .A1(EXEC_STAGE_mul_ex_mult_84_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U194 ( .A1(EXEC_STAGE_mul_ex_mult_84_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U193 ( .A1(EXEC_STAGE_mul_ex_mult_84_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U192 ( .A1(EXEC_STAGE_mul_ex_mult_84_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U191 ( .A1(EXEC_STAGE_mul_ex_mult_84_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_3__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U190 ( .A1(EXEC_STAGE_mul_ex_mult_84_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U189 ( .A1(EXEC_STAGE_mul_ex_mult_84_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U188 ( .A1(EXEC_STAGE_mul_ex_mult_84_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U187 ( .A1(EXEC_STAGE_mul_ex_mult_84_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U186 ( .A1(EXEC_STAGE_mul_ex_mult_84_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U185 ( .A1(EXEC_STAGE_mul_ex_mult_84_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U184 ( .A1(EXEC_STAGE_mul_ex_mult_84_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U183 ( .A1(EXEC_STAGE_mul_ex_mult_84_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U182 ( .A1(EXEC_STAGE_mul_ex_mult_84_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U181 ( .A1(EXEC_STAGE_mul_ex_mult_84_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U180 ( .A1(EXEC_STAGE_mul_ex_mult_84_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U179 ( .A1(EXEC_STAGE_mul_ex_mult_84_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U178 ( .A1(EXEC_STAGE_mul_ex_mult_84_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U177 ( .A1(EXEC_STAGE_mul_ex_mult_84_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U176 ( .A1(EXEC_STAGE_mul_ex_mult_84_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U175 ( .A1(EXEC_STAGE_mul_ex_mult_84_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_4__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U174 ( .A1(EXEC_STAGE_mul_ex_mult_84_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U173 ( .A1(EXEC_STAGE_mul_ex_mult_84_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U172 ( .A1(EXEC_STAGE_mul_ex_mult_84_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U171 ( .A1(EXEC_STAGE_mul_ex_mult_84_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U170 ( .A1(EXEC_STAGE_mul_ex_mult_84_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U169 ( .A1(EXEC_STAGE_mul_ex_mult_84_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U168 ( .A1(EXEC_STAGE_mul_ex_mult_84_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U167 ( .A1(EXEC_STAGE_mul_ex_mult_84_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U166 ( .A1(EXEC_STAGE_mul_ex_mult_84_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U165 ( .A1(EXEC_STAGE_mul_ex_mult_84_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U164 ( .A1(EXEC_STAGE_mul_ex_mult_84_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U163 ( .A1(EXEC_STAGE_mul_ex_mult_84_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U162 ( .A1(EXEC_STAGE_mul_ex_mult_84_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U161 ( .A1(EXEC_STAGE_mul_ex_mult_84_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U160 ( .A1(EXEC_STAGE_mul_ex_mult_84_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U159 ( .A1(EXEC_STAGE_mul_ex_mult_84_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_5__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U158 ( .A1(EXEC_STAGE_mul_ex_mult_84_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U157 ( .A1(EXEC_STAGE_mul_ex_mult_84_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U156 ( .A1(EXEC_STAGE_mul_ex_mult_84_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U155 ( .A1(EXEC_STAGE_mul_ex_mult_84_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U154 ( .A1(EXEC_STAGE_mul_ex_mult_84_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U153 ( .A1(EXEC_STAGE_mul_ex_mult_84_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U152 ( .A1(EXEC_STAGE_mul_ex_mult_84_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U151 ( .A1(EXEC_STAGE_mul_ex_mult_84_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U150 ( .A1(EXEC_STAGE_mul_ex_mult_84_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U149 ( .A1(EXEC_STAGE_mul_ex_mult_84_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U148 ( .A1(EXEC_STAGE_mul_ex_mult_84_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U147 ( .A1(EXEC_STAGE_mul_ex_mult_84_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U146 ( .A1(EXEC_STAGE_mul_ex_mult_84_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U145 ( .A1(EXEC_STAGE_mul_ex_mult_84_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U144 ( .A1(EXEC_STAGE_mul_ex_mult_84_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U143 ( .A1(EXEC_STAGE_mul_ex_mult_84_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_6__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U142 ( .A1(EXEC_STAGE_mul_ex_mult_84_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U141 ( .A1(EXEC_STAGE_mul_ex_mult_84_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U140 ( .A1(EXEC_STAGE_mul_ex_mult_84_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U139 ( .A1(EXEC_STAGE_mul_ex_mult_84_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U138 ( .A1(EXEC_STAGE_mul_ex_mult_84_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U137 ( .A1(EXEC_STAGE_mul_ex_mult_84_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U136 ( .A1(EXEC_STAGE_mul_ex_mult_84_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U135 ( .A1(EXEC_STAGE_mul_ex_mult_84_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U134 ( .A1(EXEC_STAGE_mul_ex_mult_84_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U133 ( .A1(EXEC_STAGE_mul_ex_mult_84_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U132 ( .A1(EXEC_STAGE_mul_ex_mult_84_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U131 ( .A1(EXEC_STAGE_mul_ex_mult_84_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U130 ( .A1(EXEC_STAGE_mul_ex_mult_84_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U129 ( .A1(EXEC_STAGE_mul_ex_mult_84_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U128 ( .A1(EXEC_STAGE_mul_ex_mult_84_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U127 ( .A1(EXEC_STAGE_mul_ex_mult_84_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_7__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U126 ( .A1(EXEC_STAGE_mul_ex_mult_84_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U125 ( .A1(EXEC_STAGE_mul_ex_mult_84_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U124 ( .A1(EXEC_STAGE_mul_ex_mult_84_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U123 ( .A1(EXEC_STAGE_mul_ex_mult_84_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U122 ( .A1(EXEC_STAGE_mul_ex_mult_84_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U121 ( .A1(EXEC_STAGE_mul_ex_mult_84_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U120 ( .A1(EXEC_STAGE_mul_ex_mult_84_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U119 ( .A1(EXEC_STAGE_mul_ex_mult_84_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U118 ( .A1(EXEC_STAGE_mul_ex_mult_84_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U117 ( .A1(EXEC_STAGE_mul_ex_mult_84_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U116 ( .A1(EXEC_STAGE_mul_ex_mult_84_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U115 ( .A1(EXEC_STAGE_mul_ex_mult_84_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U114 ( .A1(EXEC_STAGE_mul_ex_mult_84_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U113 ( .A1(EXEC_STAGE_mul_ex_mult_84_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U112 ( .A1(EXEC_STAGE_mul_ex_mult_84_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U111 ( .A1(EXEC_STAGE_mul_ex_mult_84_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_8__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U110 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n94), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U109 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U108 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U107 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U106 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U105 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U104 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U103 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U102 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U101 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U100 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U99 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U98 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U97 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U96 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_U95 ( .A1(EXEC_STAGE_mul_ex_mult_84_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_84_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_84_ab_9__9_) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U93 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__14_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_15__15_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n62) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U92 ( .A(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__0_), .B(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__1_), .Z(
        EXEC_STAGE_mul_ex_mult_84_n61) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U91 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_1__0_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_0__1_), .Z(EXEC_STAGE_mul_ex_N89) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U90 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__0_), .A2(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n59) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U89 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__2_), .A2(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n58) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U88 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__4_), .A2(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n57) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U87 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__6_), .A2(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n56) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U86 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__8_), .A2(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n55) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U85 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__10_), .A2(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__11_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n54) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U84 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__12_), .A2(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__13_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n53) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U83 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__1_), .A2(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n52) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U82 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__3_), .A2(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n51) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U81 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__5_), .A2(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n50) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U80 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__7_), .A2(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n49) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U79 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__9_), .A2(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n48) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U78 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__11_), .A2(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__12_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n47) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U77 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__13_), .A2(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__14_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n46) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U76 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_1__1_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_0__2_), .Z(EXEC_STAGE_mul_ex_mult_84_n45)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U75 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_1__2_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_0__3_), .Z(EXEC_STAGE_mul_ex_mult_84_n44)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U74 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_1__3_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_0__4_), .Z(EXEC_STAGE_mul_ex_mult_84_n43)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U73 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_1__4_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_0__5_), .Z(EXEC_STAGE_mul_ex_mult_84_n42)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U72 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_1__5_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_0__6_), .Z(EXEC_STAGE_mul_ex_mult_84_n41)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U71 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_1__6_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_0__7_), .Z(EXEC_STAGE_mul_ex_mult_84_n40)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U70 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_1__7_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_0__8_), .Z(EXEC_STAGE_mul_ex_mult_84_n39)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U69 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_1__8_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_0__9_), .Z(EXEC_STAGE_mul_ex_mult_84_n38)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U68 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_1__9_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_0__10_), .Z(EXEC_STAGE_mul_ex_mult_84_n37) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U67 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_1__10_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_0__11_), .Z(EXEC_STAGE_mul_ex_mult_84_n36) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U66 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_1__11_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_0__12_), .Z(EXEC_STAGE_mul_ex_mult_84_n35) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U65 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_1__12_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_0__13_), .Z(EXEC_STAGE_mul_ex_mult_84_n34) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U64 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_1__13_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_0__14_), .Z(EXEC_STAGE_mul_ex_mult_84_n33) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U63 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_1__14_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_0__15_), .Z(EXEC_STAGE_mul_ex_mult_84_n32) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U62 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_ab_0__15_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_1__14_), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n31) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U61 ( .A(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__3_), .B(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__4_), .Z(
        EXEC_STAGE_mul_ex_mult_84_n30) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U60 ( .A(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__5_), .B(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__6_), .Z(
        EXEC_STAGE_mul_ex_mult_84_n29) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U59 ( .A(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__7_), .B(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__8_), .Z(
        EXEC_STAGE_mul_ex_mult_84_n28) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U58 ( .A(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__9_), .B(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__10_), .Z(
        EXEC_STAGE_mul_ex_mult_84_n27) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U57 ( .A(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__11_), .B(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__12_), .Z(
        EXEC_STAGE_mul_ex_mult_84_n26) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U56 ( .A(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__13_), .B(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__14_), .Z(
        EXEC_STAGE_mul_ex_mult_84_n25) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U55 ( .A(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__1_), .B(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__2_), .Z(
        EXEC_STAGE_mul_ex_mult_84_n24) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U54 ( .A(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__2_), .B(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__3_), .Z(
        EXEC_STAGE_mul_ex_mult_84_n23) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U53 ( .A(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__4_), .B(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__5_), .Z(
        EXEC_STAGE_mul_ex_mult_84_n22) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U52 ( .A(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__6_), .B(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__7_), .Z(
        EXEC_STAGE_mul_ex_mult_84_n21) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U51 ( .A(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__8_), .B(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__9_), .Z(
        EXEC_STAGE_mul_ex_mult_84_n20) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U50 ( .A(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__10_), .B(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__11_), .Z(
        EXEC_STAGE_mul_ex_mult_84_n19) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U49 ( .A(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__12_), .B(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__13_), .Z(
        EXEC_STAGE_mul_ex_mult_84_n18) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_84_U48 ( .A(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__14_), .B(
        EXEC_STAGE_mul_ex_mult_84_ab_15__15_), .Z(
        EXEC_STAGE_mul_ex_mult_84_n17) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U47 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_ab_0__1_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_1__0_), .ZN(EXEC_STAGE_mul_ex_mult_84_n16) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U46 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_ab_0__2_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_1__1_), .ZN(EXEC_STAGE_mul_ex_mult_84_n15) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U45 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_ab_0__3_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_1__2_), .ZN(EXEC_STAGE_mul_ex_mult_84_n14) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U44 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_ab_0__4_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_1__3_), .ZN(EXEC_STAGE_mul_ex_mult_84_n13) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U43 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_ab_0__5_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_1__4_), .ZN(EXEC_STAGE_mul_ex_mult_84_n12) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U42 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_ab_0__6_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_1__5_), .ZN(EXEC_STAGE_mul_ex_mult_84_n11) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U41 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_ab_0__7_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_1__6_), .ZN(EXEC_STAGE_mul_ex_mult_84_n10) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U40 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_ab_0__8_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_1__7_), .ZN(EXEC_STAGE_mul_ex_mult_84_n9)
         );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U39 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_ab_0__9_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_1__8_), .ZN(EXEC_STAGE_mul_ex_mult_84_n8)
         );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U38 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_ab_0__10_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_1__9_), .ZN(EXEC_STAGE_mul_ex_mult_84_n7)
         );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U37 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_ab_0__11_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_1__10_), .ZN(EXEC_STAGE_mul_ex_mult_84_n6) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U36 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_ab_0__12_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_1__11_), .ZN(EXEC_STAGE_mul_ex_mult_84_n5) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U35 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_ab_0__13_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_1__12_), .ZN(EXEC_STAGE_mul_ex_mult_84_n4) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_U34 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_ab_0__14_), .A2(
        EXEC_STAGE_mul_ex_mult_84_ab_1__13_), .ZN(EXEC_STAGE_mul_ex_mult_84_n3) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U33 ( .A(ID_EXEC_OUT[267]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n94) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U32 ( .A(ID_EXEC_OUT[235]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n63) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U31 ( .A(ID_EXEC_OUT[220]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n78) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U30 ( .A(ID_EXEC_OUT[266]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n67) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U29 ( .A(ID_EXEC_OUT[221]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n80) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U28 ( .A(ID_EXEC_OUT[222]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n64) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U27 ( .A(ID_EXEC_OUT[223]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n88) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U26 ( .A(ID_EXEC_OUT[224]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n82) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U25 ( .A(ID_EXEC_OUT[225]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n84) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U24 ( .A(ID_EXEC_OUT[226]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n86) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U23 ( .A(ID_EXEC_OUT[227]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n90) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U22 ( .A(ID_EXEC_OUT[228]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n92) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U21 ( .A(ID_EXEC_OUT[229]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n70) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U20 ( .A(ID_EXEC_OUT[230]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n74) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U19 ( .A(ID_EXEC_OUT[231]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n72) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U18 ( .A(ID_EXEC_OUT[232]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n76) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U17 ( .A(ID_EXEC_OUT[233]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n68) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U16 ( .A(ID_EXEC_OUT[234]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n66) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U15 ( .A(ID_EXEC_OUT[252]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n79) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U14 ( .A(ID_EXEC_OUT[253]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n81) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U13 ( .A(ID_EXEC_OUT[265]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n69) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U12 ( .A(ID_EXEC_OUT[254]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n65) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U11 ( .A(ID_EXEC_OUT[255]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n89) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U10 ( .A(ID_EXEC_OUT[256]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n83) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U9 ( .A(ID_EXEC_OUT[257]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n85) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U8 ( .A(ID_EXEC_OUT[258]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n87) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U7 ( .A(ID_EXEC_OUT[259]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n91) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U6 ( .A(ID_EXEC_OUT[260]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n93) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U5 ( .A(ID_EXEC_OUT[261]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n71) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U4 ( .A(ID_EXEC_OUT[262]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n75) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U3 ( .A(ID_EXEC_OUT[263]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n73) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_U2 ( .A(ID_EXEC_OUT[264]), .ZN(
        EXEC_STAGE_mul_ex_mult_84_n77) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S3_2_14 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_2__14_), .B(EXEC_STAGE_mul_ex_mult_84_n31), .CI(EXEC_STAGE_mul_ex_mult_84_ab_1__15_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__14_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_2_13 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_2__13_), .B(EXEC_STAGE_mul_ex_mult_84_n3), 
        .CI(EXEC_STAGE_mul_ex_mult_84_n32), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__13_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_2_12 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_2__12_), .B(EXEC_STAGE_mul_ex_mult_84_n4), 
        .CI(EXEC_STAGE_mul_ex_mult_84_n33), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__12_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_2_11 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_2__11_), .B(EXEC_STAGE_mul_ex_mult_84_n5), 
        .CI(EXEC_STAGE_mul_ex_mult_84_n34), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__11_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_2_10 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_2__10_), .B(EXEC_STAGE_mul_ex_mult_84_n6), 
        .CI(EXEC_STAGE_mul_ex_mult_84_n35), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__10_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_2_9 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_2__9_), .B(EXEC_STAGE_mul_ex_mult_84_n7), 
        .CI(EXEC_STAGE_mul_ex_mult_84_n36), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__9_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_2_8 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_2__8_), .B(EXEC_STAGE_mul_ex_mult_84_n8), 
        .CI(EXEC_STAGE_mul_ex_mult_84_n37), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__8_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_2_7 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_2__7_), .B(EXEC_STAGE_mul_ex_mult_84_n9), 
        .CI(EXEC_STAGE_mul_ex_mult_84_n38), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__7_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_2_6 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_2__6_), .B(EXEC_STAGE_mul_ex_mult_84_n10), 
        .CI(EXEC_STAGE_mul_ex_mult_84_n39), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__6_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_2_5 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_2__5_), .B(EXEC_STAGE_mul_ex_mult_84_n11), 
        .CI(EXEC_STAGE_mul_ex_mult_84_n40), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__5_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_2_4 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_2__4_), .B(EXEC_STAGE_mul_ex_mult_84_n12), 
        .CI(EXEC_STAGE_mul_ex_mult_84_n41), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__4_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_2_3 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_2__3_), .B(EXEC_STAGE_mul_ex_mult_84_n13), 
        .CI(EXEC_STAGE_mul_ex_mult_84_n42), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__3_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_2_2 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_2__2_), .B(EXEC_STAGE_mul_ex_mult_84_n14), 
        .CI(EXEC_STAGE_mul_ex_mult_84_n43), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__2_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_2_1 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_2__1_), .B(EXEC_STAGE_mul_ex_mult_84_n15), 
        .CI(EXEC_STAGE_mul_ex_mult_84_n44), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__1_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S1_2_0 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_2__0_), .B(EXEC_STAGE_mul_ex_mult_84_n16), 
        .CI(EXEC_STAGE_mul_ex_mult_84_n45), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__0_), .S(
        EXEC_STAGE_mul_ex_mult_84_A1_0_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S3_3_14 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_3__14_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__14_), .CI(
        EXEC_STAGE_mul_ex_mult_84_ab_2__15_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__14_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_3_13 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_3__13_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__13_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__14_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__13_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_3_12 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_3__12_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__12_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__13_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__12_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_3_11 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_3__11_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__11_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__12_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__11_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_3_10 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_3__10_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__10_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__11_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__10_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_3_9 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_3__9_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__9_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__10_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__9_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_3_8 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_3__8_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__8_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__9_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__8_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_3_7 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_3__7_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__7_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__8_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__7_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_3_6 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_3__6_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__6_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__7_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__6_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_3_5 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_3__5_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__5_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__6_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__5_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_3_4 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_3__4_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__4_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__5_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__4_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_3_3 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_3__3_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__3_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__4_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__3_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_3_2 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_3__2_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__2_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__3_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__2_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_3_1 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_3__1_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__1_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__2_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__1_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S1_3_0 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_3__0_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_2__0_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_2__1_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__0_), .S(
        EXEC_STAGE_mul_ex_mult_84_A1_1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S3_4_14 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_4__14_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__14_), .CI(
        EXEC_STAGE_mul_ex_mult_84_ab_3__15_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__14_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_4_13 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_4__13_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__13_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__14_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__13_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_4_12 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_4__12_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__12_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__13_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__12_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_4_11 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_4__11_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__11_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__12_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__11_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_4_10 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_4__10_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__10_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__11_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__10_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_4_9 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_4__9_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__9_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__10_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__9_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_4_8 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_4__8_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__8_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__9_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__8_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_4_7 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_4__7_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__7_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__8_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__7_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_4_6 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_4__6_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__6_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__7_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__6_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_4_5 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_4__5_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__5_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__6_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__5_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_4_4 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_4__4_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__4_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__5_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__4_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_4_3 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_4__3_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__3_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__4_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__3_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_4_2 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_4__2_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__2_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__3_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__2_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_4_1 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_4__1_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__1_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__2_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__1_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S1_4_0 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_4__0_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_3__0_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_3__1_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__0_), .S(
        EXEC_STAGE_mul_ex_mult_84_A1_2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S3_5_14 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_5__14_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__14_), .CI(
        EXEC_STAGE_mul_ex_mult_84_ab_4__15_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__14_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_5_13 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_5__13_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__13_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__14_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__13_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_5_12 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_5__12_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__12_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__13_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__12_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_5_11 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_5__11_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__11_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__12_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__11_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_5_10 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_5__10_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__10_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__11_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__10_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_5_9 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_5__9_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__9_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__10_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__9_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_5_8 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_5__8_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__8_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__9_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__8_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_5_7 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_5__7_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__7_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__8_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__7_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_5_6 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_5__6_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__6_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__7_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__6_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_5_5 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_5__5_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__5_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__6_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__5_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_5_4 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_5__4_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__4_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__5_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__4_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_5_3 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_5__3_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__3_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__4_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__3_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_5_2 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_5__2_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__2_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__3_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__2_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_5_1 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_5__1_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__1_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__2_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__1_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S1_5_0 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_5__0_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_4__0_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_4__1_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__0_), .S(
        EXEC_STAGE_mul_ex_mult_84_A1_3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S3_6_14 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_6__14_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__14_), .CI(
        EXEC_STAGE_mul_ex_mult_84_ab_5__15_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__14_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_6_13 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_6__13_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__13_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__14_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__13_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_6_12 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_6__12_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__12_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__13_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__12_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_6_11 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_6__11_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__11_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__12_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__11_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_6_10 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_6__10_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__10_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__11_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__10_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_6_9 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_6__9_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__9_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__10_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__9_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_6_8 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_6__8_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__8_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__9_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__8_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_6_7 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_6__7_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__7_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__8_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__7_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_6_6 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_6__6_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__6_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__7_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__6_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_6_5 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_6__5_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__5_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__6_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__5_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_6_4 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_6__4_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__4_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__5_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__4_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_6_3 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_6__3_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__3_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__4_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__3_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_6_2 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_6__2_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__2_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__3_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__2_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_6_1 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_6__1_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__1_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__2_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__1_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S1_6_0 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_6__0_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_5__0_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_5__1_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__0_), .S(
        EXEC_STAGE_mul_ex_mult_84_A1_4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S3_7_14 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_7__14_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__14_), .CI(
        EXEC_STAGE_mul_ex_mult_84_ab_6__15_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__14_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_7_13 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_7__13_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__13_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__14_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__13_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_7_12 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_7__12_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__12_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__13_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__12_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_7_11 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_7__11_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__11_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__12_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__11_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_7_10 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_7__10_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__10_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__11_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__10_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_7_9 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_7__9_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__9_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__10_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__9_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_7_8 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_7__8_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__8_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__9_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__8_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_7_7 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_7__7_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__7_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__8_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__7_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_7_6 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_7__6_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__6_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__7_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__6_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_7_5 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_7__5_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__5_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__6_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__5_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_7_4 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_7__4_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__4_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__5_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__4_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_7_3 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_7__3_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__3_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__4_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__3_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_7_2 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_7__2_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__2_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__3_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__2_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_7_1 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_7__1_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__1_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__2_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__1_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S1_7_0 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_7__0_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_6__0_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_6__1_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__0_), .S(
        EXEC_STAGE_mul_ex_mult_84_A1_5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S3_8_14 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_8__14_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__14_), .CI(
        EXEC_STAGE_mul_ex_mult_84_ab_7__15_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__14_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_8_13 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_8__13_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__13_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__14_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__13_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_8_12 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_8__12_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__12_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__13_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__12_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_8_11 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_8__11_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__11_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__12_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__11_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_8_10 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_8__10_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__10_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__11_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__10_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_8_9 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_8__9_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__9_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__10_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__9_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_8_8 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_8__8_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__8_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__9_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__8_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_8_7 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_8__7_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__7_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__8_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__7_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_8_6 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_8__6_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__6_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__7_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__6_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_8_5 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_8__5_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__5_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__6_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__5_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_8_4 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_8__4_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__4_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__5_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__4_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_8_3 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_8__3_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__3_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__4_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__3_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_8_2 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_8__2_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__2_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__3_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__2_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_8_1 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_8__1_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__1_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__2_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__1_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S1_8_0 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_8__0_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_7__0_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_7__1_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__0_), .S(
        EXEC_STAGE_mul_ex_mult_84_A1_6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S3_9_14 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_9__14_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__14_), .CI(
        EXEC_STAGE_mul_ex_mult_84_ab_8__15_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__14_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_9_13 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_9__13_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__13_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__14_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__13_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_9_12 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_9__12_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__12_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__13_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__12_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_9_11 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_9__11_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__11_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__12_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__11_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_9_10 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_9__10_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__10_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__11_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__10_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_9_9 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_9__9_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__9_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__10_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__9_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_9_8 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_9__8_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__8_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__9_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__8_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_9_7 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_9__7_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__7_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__8_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__7_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_9_6 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_9__6_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__6_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__7_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__6_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_9_5 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_9__5_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__5_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__6_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__5_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_9_4 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_9__4_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__4_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__5_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__4_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_9_3 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_9__3_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__3_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__4_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__3_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_9_2 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_9__2_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__2_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__3_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__2_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_9_1 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_9__1_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__1_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__2_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__1_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S1_9_0 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_9__0_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_8__0_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_8__1_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__0_), .S(
        EXEC_STAGE_mul_ex_mult_84_A1_7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S3_10_14 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_10__14_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__14_), .CI(
        EXEC_STAGE_mul_ex_mult_84_ab_9__15_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__14_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_10_13 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_10__13_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__13_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__14_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__13_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_10_12 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_10__12_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__12_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__13_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__12_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_10_11 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_10__11_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__11_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__12_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__11_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_10_10 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_10__10_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__10_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__11_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__10_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_10_9 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_10__9_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__9_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__10_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__9_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_10_8 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_10__8_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__8_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__9_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__8_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_10_7 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_10__7_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__7_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__8_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__7_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_10_6 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_10__6_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__6_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__7_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__6_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_10_5 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_10__5_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__5_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__6_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__5_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_10_4 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_10__4_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__4_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__5_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__4_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_10_3 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_10__3_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__3_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__4_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__3_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_10_2 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_10__2_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__2_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__3_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__2_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_10_1 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_10__1_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__1_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__2_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__1_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S1_10_0 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_10__0_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_9__0_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_9__1_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__0_), .S(
        EXEC_STAGE_mul_ex_mult_84_A1_8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S3_11_14 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_11__14_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__14_), .CI(
        EXEC_STAGE_mul_ex_mult_84_ab_10__15_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__14_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_11_13 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_11__13_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__13_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__14_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__13_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_11_12 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_11__12_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__12_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__13_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__12_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_11_11 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_11__11_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__11_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__12_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__11_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_11_10 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_11__10_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__10_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__11_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__10_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_11_9 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_11__9_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__9_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__10_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__9_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_11_8 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_11__8_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__8_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__9_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__8_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_11_7 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_11__7_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__7_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__8_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__7_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_11_6 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_11__6_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__6_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__7_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__6_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_11_5 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_11__5_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__5_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__6_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__5_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_11_4 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_11__4_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__4_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__5_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__4_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_11_3 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_11__3_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__3_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__4_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__3_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_11_2 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_11__2_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__2_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__3_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__2_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_11_1 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_11__1_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__1_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__2_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__1_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S1_11_0 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_11__0_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_10__0_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_10__1_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__0_), .S(
        EXEC_STAGE_mul_ex_mult_84_A1_9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S3_12_14 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_12__14_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__14_), .CI(
        EXEC_STAGE_mul_ex_mult_84_ab_11__15_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__14_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_12_13 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_12__13_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__13_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__14_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__13_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_12_12 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_12__12_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__12_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__13_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__12_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_12_11 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_12__11_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__11_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__12_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__11_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_12_10 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_12__10_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__10_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__11_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__10_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_12_9 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_12__9_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__9_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__10_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__9_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_12_8 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_12__8_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__8_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__9_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__8_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_12_7 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_12__7_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__7_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__8_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__7_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_12_6 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_12__6_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__6_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__7_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__6_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_12_5 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_12__5_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__5_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__6_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__5_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_12_4 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_12__4_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__4_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__5_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__4_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_12_3 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_12__3_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__3_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__4_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__3_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_12_2 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_12__2_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__2_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__3_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__2_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_12_1 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_12__1_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__1_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__2_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__1_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S1_12_0 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_12__0_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_11__0_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_11__1_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__0_), .S(
        EXEC_STAGE_mul_ex_mult_84_A1_10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S3_13_14 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_13__14_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__14_), .CI(
        EXEC_STAGE_mul_ex_mult_84_ab_12__15_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__14_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_13_13 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_13__13_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__13_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__14_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__13_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_13_12 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_13__12_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__12_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__13_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__12_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_13_11 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_13__11_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__11_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__12_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__11_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_13_10 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_13__10_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__10_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__11_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__10_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_13_9 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_13__9_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__9_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__10_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__9_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_13_8 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_13__8_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__8_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__9_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__8_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_13_7 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_13__7_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__7_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__8_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__7_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_13_6 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_13__6_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__6_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__7_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__6_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_13_5 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_13__5_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__5_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__6_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__5_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_13_4 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_13__4_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__4_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__5_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__4_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_13_3 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_13__3_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__3_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__4_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__3_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_13_2 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_13__2_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__2_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__3_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__2_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_13_1 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_13__1_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__1_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__2_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__1_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S1_13_0 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_13__0_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_12__0_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_12__1_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__0_), .S(
        EXEC_STAGE_mul_ex_mult_84_A1_11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S3_14_14 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_14__14_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__14_), .CI(
        EXEC_STAGE_mul_ex_mult_84_ab_13__15_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__14_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_14_13 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_14__13_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__13_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__14_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__13_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_14_12 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_14__12_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__12_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__13_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__12_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_14_11 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_14__11_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__11_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__12_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__11_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_14_10 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_14__10_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__10_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__11_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__10_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_14_9 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_14__9_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__9_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__10_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__9_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_14_8 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_14__8_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__8_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__9_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__8_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_14_7 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_14__7_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__7_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__8_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__7_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_14_6 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_14__6_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__6_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__7_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__6_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_14_5 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_14__5_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__5_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__6_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__5_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_14_4 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_14__4_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__4_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__5_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__4_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_14_3 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_14__3_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__3_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__4_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__3_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_14_2 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_14__2_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__2_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__3_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__2_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S2_14_1 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_14__1_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__1_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__2_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__1_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S1_14_0 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_14__0_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_13__0_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_13__1_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__0_), .S(
        EXEC_STAGE_mul_ex_mult_84_A1_12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S5_14 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_15__14_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__14_), .CI(
        EXEC_STAGE_mul_ex_mult_84_ab_14__15_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__14_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S4_13 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_15__13_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__13_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__14_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__13_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S4_12 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_15__12_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__12_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__13_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__12_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S4_11 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_15__11_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__11_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__12_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__11_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S4_10 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_15__10_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__10_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__11_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__10_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S4_9 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_15__9_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__9_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__10_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__9_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S4_8 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_15__8_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__8_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__9_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__8_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S4_7 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_15__7_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__7_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__8_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__7_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S4_6 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_15__6_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__6_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__7_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__6_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S4_5 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_15__5_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__5_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__6_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__5_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S4_4 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_15__4_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__4_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__5_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__4_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S4_3 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_15__3_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__3_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__4_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__3_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S4_2 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_15__2_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__2_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__3_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__2_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S4_1 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_15__1_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__1_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__2_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__1_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_84_S4_0 ( .A(
        EXEC_STAGE_mul_ex_mult_84_ab_15__0_), .B(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_14__0_), .CI(
        EXEC_STAGE_mul_ex_mult_84_SUMB_14__1_), .CO(
        EXEC_STAGE_mul_ex_mult_84_CARRYB_15__0_), .S(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__0_) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_84_FS_1_U100 ( .A(
        EXEC_STAGE_mul_ex_mult_84_n61), .Z(EXEC_STAGE_mul_ex_N104) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_84_FS_1_U99 ( .A(
        EXEC_STAGE_mul_ex_mult_84_SUMB_15__0_), .Z(EXEC_STAGE_mul_ex_N103) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_84_FS_1_U98 ( .A(
        EXEC_STAGE_mul_ex_mult_84_A1_12_), .Z(EXEC_STAGE_mul_ex_N102) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_84_FS_1_U97 ( .A(
        EXEC_STAGE_mul_ex_mult_84_A1_11_), .Z(EXEC_STAGE_mul_ex_N101) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_84_FS_1_U96 ( .A(
        EXEC_STAGE_mul_ex_mult_84_A1_10_), .Z(EXEC_STAGE_mul_ex_N100) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_84_FS_1_U95 ( .A(
        EXEC_STAGE_mul_ex_mult_84_A1_9_), .Z(EXEC_STAGE_mul_ex_N99) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_84_FS_1_U94 ( .A(
        EXEC_STAGE_mul_ex_mult_84_A1_8_), .Z(EXEC_STAGE_mul_ex_N98) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_84_FS_1_U93 ( .A(
        EXEC_STAGE_mul_ex_mult_84_A1_7_), .Z(EXEC_STAGE_mul_ex_N97) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_84_FS_1_U92 ( .A(
        EXEC_STAGE_mul_ex_mult_84_A1_6_), .Z(EXEC_STAGE_mul_ex_N96) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_84_FS_1_U91 ( .A(
        EXEC_STAGE_mul_ex_mult_84_A1_5_), .Z(EXEC_STAGE_mul_ex_N95) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_84_FS_1_U90 ( .A(
        EXEC_STAGE_mul_ex_mult_84_A1_4_), .Z(EXEC_STAGE_mul_ex_N94) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_84_FS_1_U89 ( .A(
        EXEC_STAGE_mul_ex_mult_84_A1_3_), .Z(EXEC_STAGE_mul_ex_N93) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_84_FS_1_U88 ( .A(
        EXEC_STAGE_mul_ex_mult_84_A1_2_), .Z(EXEC_STAGE_mul_ex_N92) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_84_FS_1_U87 ( .A(
        EXEC_STAGE_mul_ex_mult_84_A1_1_), .Z(EXEC_STAGE_mul_ex_N91) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_84_FS_1_U86 ( .A(
        EXEC_STAGE_mul_ex_mult_84_A1_0_), .Z(EXEC_STAGE_mul_ex_N90) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U85 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n59), .A2(EXEC_STAGE_mul_ex_mult_84_n24), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n70) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U84 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n52), .A2(EXEC_STAGE_mul_ex_mult_84_n23), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n67) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U83 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n52), .A2(EXEC_STAGE_mul_ex_mult_84_n23), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n68) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U82 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n67), .A2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n69) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U81 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n17), .B(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n69), .Z(EXEC_STAGE_mul_ex_N106) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U80 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n58), .A2(EXEC_STAGE_mul_ex_mult_84_n30), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n63) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U79 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n58), .A2(EXEC_STAGE_mul_ex_mult_84_n30), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n65) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U78 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n15), .A2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n66) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U77 ( .B1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n16), .B2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n17), .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n64) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U76 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n66), .B(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n64), .Z(EXEC_STAGE_mul_ex_N107) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U75 ( .B1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n63), .B2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n64), .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n59) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U74 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n51), .A2(EXEC_STAGE_mul_ex_mult_84_n22), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n60) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U73 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n51), .A2(EXEC_STAGE_mul_ex_mult_84_n22), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n61) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U72 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n60), .A2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n61), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n62) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U71 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n59), .B(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n62), .Z(EXEC_STAGE_mul_ex_N108) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U70 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n57), .A2(EXEC_STAGE_mul_ex_mult_84_n29), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n55) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U69 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n57), .A2(EXEC_STAGE_mul_ex_mult_84_n29), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n57) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U68 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n13), .A2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n57), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n58) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U67 ( .B1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n14), .B2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n59), .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n60), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n56) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U66 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n58), .B(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n56), .Z(EXEC_STAGE_mul_ex_N109) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U65 ( .B1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n55), .B2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n56), .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n57), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n51) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U64 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n50), .A2(EXEC_STAGE_mul_ex_mult_84_n21), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n52) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U63 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n50), .A2(EXEC_STAGE_mul_ex_mult_84_n21), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n53) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U62 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n52), .A2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n54) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U61 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n51), .B(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n54), .Z(EXEC_STAGE_mul_ex_N110) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U60 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n56), .A2(EXEC_STAGE_mul_ex_mult_84_n28), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n47) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U59 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n56), .A2(EXEC_STAGE_mul_ex_mult_84_n28), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n49) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U58 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n11), .A2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n49), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n50) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U57 ( .B1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n12), .B2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n51), .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n48) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U56 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n50), .B(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n48), .Z(EXEC_STAGE_mul_ex_N111) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U55 ( .B1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n47), .B2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n48), .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n49), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n43) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U54 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n49), .A2(EXEC_STAGE_mul_ex_mult_84_n20), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n44) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U53 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n49), .A2(EXEC_STAGE_mul_ex_mult_84_n20), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n45) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U52 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n44), .A2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n45), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n46) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U51 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n43), .B(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n46), .Z(EXEC_STAGE_mul_ex_N112) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U50 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n55), .A2(EXEC_STAGE_mul_ex_mult_84_n27), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n39) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U49 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n55), .A2(EXEC_STAGE_mul_ex_mult_84_n27), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n41) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U48 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n9), .A2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n41), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n42) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U47 ( .B1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n10), .B2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n43), .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n44), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n40) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U46 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n42), .B(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n40), .Z(EXEC_STAGE_mul_ex_N113) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U45 ( .B1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n39), .B2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n40), .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n41), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n35) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U44 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n48), .A2(EXEC_STAGE_mul_ex_mult_84_n19), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n36) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U43 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n48), .A2(EXEC_STAGE_mul_ex_mult_84_n19), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n37) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U42 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n36), .A2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n37), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n38) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U41 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n35), .B(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n38), .Z(EXEC_STAGE_mul_ex_N114) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U40 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n54), .A2(EXEC_STAGE_mul_ex_mult_84_n26), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n31) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U39 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n54), .A2(EXEC_STAGE_mul_ex_mult_84_n26), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n33) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U38 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n7), .A2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n33), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n34) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U37 ( .B1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n8), .B2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n35), .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n36), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n32) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U36 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n34), .B(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n32), .Z(EXEC_STAGE_mul_ex_N115) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U35 ( .B1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n31), .B2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n32), .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n33), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n27) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U34 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n47), .A2(EXEC_STAGE_mul_ex_mult_84_n18), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n28) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U33 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n47), .A2(EXEC_STAGE_mul_ex_mult_84_n18), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n29) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U32 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n28), .A2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n29), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n30) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U31 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n27), .B(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n30), .Z(EXEC_STAGE_mul_ex_N116) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U30 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n53), .A2(EXEC_STAGE_mul_ex_mult_84_n25), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n23) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U29 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n53), .A2(EXEC_STAGE_mul_ex_mult_84_n25), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n25) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U28 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n5), .A2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n25), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n26) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U27 ( .B1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n6), .B2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n27), .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n28), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n24) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U26 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n26), .B(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n24), .Z(EXEC_STAGE_mul_ex_N117) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U25 ( .B1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n23), .B2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n24), .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n25), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n19) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U24 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n46), .A2(EXEC_STAGE_mul_ex_mult_84_n17), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n20) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U23 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_n46), .A2(EXEC_STAGE_mul_ex_mult_84_n17), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n21) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U22 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n20), .A2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n21), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n22) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U21 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n19), .B(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n22), .Z(EXEC_STAGE_mul_ex_N118) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U20 ( .B1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n19), .B2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n4), .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n20), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n18) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_84_FS_1_U19 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n3), .B(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n18), .Z(EXEC_STAGE_mul_ex_N119) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U18 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n17) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U17 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n16) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U16 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n15) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U15 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n61), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n14) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U14 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n55), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n13) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U13 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n12) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U12 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n47), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n11) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U11 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n45), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n10) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U10 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n39), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n9) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U9 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n37), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n8) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U8 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n31), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n7) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U7 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n29), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n6) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U6 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n23), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n5) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U5 ( .A(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n21), .ZN(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n4) );
  INV_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U4 ( .A(EXEC_STAGE_mul_ex_mult_84_n62), 
        .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n3) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U3 ( .A1(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n1), .A2(
        EXEC_STAGE_mul_ex_mult_84_FS_1_n70), .ZN(EXEC_STAGE_mul_ex_N105) );
  OR2_X4 EXEC_STAGE_mul_ex_mult_84_FS_1_U2 ( .A1(EXEC_STAGE_mul_ex_mult_84_n59), .A2(EXEC_STAGE_mul_ex_mult_84_n24), .ZN(EXEC_STAGE_mul_ex_mult_84_FS_1_n1)
         );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U350 ( .A1(EXEC_STAGE_mul_ex_mult_76_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(EXEC_STAGE_mul_ex_N56) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U349 ( .A1(EXEC_STAGE_mul_ex_mult_76_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U348 ( .A1(EXEC_STAGE_mul_ex_mult_76_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U347 ( .A1(EXEC_STAGE_mul_ex_mult_76_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U346 ( .A1(EXEC_STAGE_mul_ex_mult_76_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U345 ( .A1(EXEC_STAGE_mul_ex_mult_76_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U344 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U343 ( .A1(EXEC_STAGE_mul_ex_mult_76_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U342 ( .A1(EXEC_STAGE_mul_ex_mult_76_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U341 ( .A1(EXEC_STAGE_mul_ex_mult_76_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U340 ( .A1(EXEC_STAGE_mul_ex_mult_76_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U339 ( .A1(EXEC_STAGE_mul_ex_mult_76_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U338 ( .A1(EXEC_STAGE_mul_ex_mult_76_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U337 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U336 ( .A1(EXEC_STAGE_mul_ex_mult_76_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U335 ( .A1(EXEC_STAGE_mul_ex_mult_76_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U334 ( .A1(EXEC_STAGE_mul_ex_mult_76_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U333 ( .A1(EXEC_STAGE_mul_ex_mult_76_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U332 ( .A1(EXEC_STAGE_mul_ex_mult_76_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U331 ( .A1(EXEC_STAGE_mul_ex_mult_76_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U330 ( .A1(EXEC_STAGE_mul_ex_mult_76_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U329 ( .A1(EXEC_STAGE_mul_ex_mult_76_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U328 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U327 ( .A1(EXEC_STAGE_mul_ex_mult_76_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U326 ( .A1(EXEC_STAGE_mul_ex_mult_76_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U325 ( .A1(EXEC_STAGE_mul_ex_mult_76_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U324 ( .A1(EXEC_STAGE_mul_ex_mult_76_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U323 ( .A1(EXEC_STAGE_mul_ex_mult_76_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U322 ( .A1(EXEC_STAGE_mul_ex_mult_76_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U321 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U320 ( .A1(EXEC_STAGE_mul_ex_mult_76_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U319 ( .A1(EXEC_STAGE_mul_ex_mult_76_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U318 ( .A1(EXEC_STAGE_mul_ex_mult_76_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U317 ( .A1(EXEC_STAGE_mul_ex_mult_76_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U316 ( .A1(EXEC_STAGE_mul_ex_mult_76_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U315 ( .A1(EXEC_STAGE_mul_ex_mult_76_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U314 ( .A1(EXEC_STAGE_mul_ex_mult_76_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U313 ( .A1(EXEC_STAGE_mul_ex_mult_76_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U312 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U311 ( .A1(EXEC_STAGE_mul_ex_mult_76_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U310 ( .A1(EXEC_STAGE_mul_ex_mult_76_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U309 ( .A1(EXEC_STAGE_mul_ex_mult_76_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U308 ( .A1(EXEC_STAGE_mul_ex_mult_76_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U307 ( .A1(EXEC_STAGE_mul_ex_mult_76_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U306 ( .A1(EXEC_STAGE_mul_ex_mult_76_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U305 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U304 ( .A1(EXEC_STAGE_mul_ex_mult_76_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U303 ( .A1(EXEC_STAGE_mul_ex_mult_76_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U302 ( .A1(EXEC_STAGE_mul_ex_mult_76_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U301 ( .A1(EXEC_STAGE_mul_ex_mult_76_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U300 ( .A1(EXEC_STAGE_mul_ex_mult_76_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U299 ( .A1(EXEC_STAGE_mul_ex_mult_76_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U298 ( .A1(EXEC_STAGE_mul_ex_mult_76_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U297 ( .A1(EXEC_STAGE_mul_ex_mult_76_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U296 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U295 ( .A1(EXEC_STAGE_mul_ex_mult_76_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U294 ( .A1(EXEC_STAGE_mul_ex_mult_76_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U293 ( .A1(EXEC_STAGE_mul_ex_mult_76_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U292 ( .A1(EXEC_STAGE_mul_ex_mult_76_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U291 ( .A1(EXEC_STAGE_mul_ex_mult_76_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U290 ( .A1(EXEC_STAGE_mul_ex_mult_76_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U289 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U288 ( .A1(EXEC_STAGE_mul_ex_mult_76_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U287 ( .A1(EXEC_STAGE_mul_ex_mult_76_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U286 ( .A1(EXEC_STAGE_mul_ex_mult_76_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U285 ( .A1(EXEC_STAGE_mul_ex_mult_76_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U284 ( .A1(EXEC_STAGE_mul_ex_mult_76_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U283 ( .A1(EXEC_STAGE_mul_ex_mult_76_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U282 ( .A1(EXEC_STAGE_mul_ex_mult_76_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U281 ( .A1(EXEC_STAGE_mul_ex_mult_76_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U280 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U279 ( .A1(EXEC_STAGE_mul_ex_mult_76_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U278 ( .A1(EXEC_STAGE_mul_ex_mult_76_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U277 ( .A1(EXEC_STAGE_mul_ex_mult_76_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U276 ( .A1(EXEC_STAGE_mul_ex_mult_76_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U275 ( .A1(EXEC_STAGE_mul_ex_mult_76_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U274 ( .A1(EXEC_STAGE_mul_ex_mult_76_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U273 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U272 ( .A1(EXEC_STAGE_mul_ex_mult_76_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U271 ( .A1(EXEC_STAGE_mul_ex_mult_76_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U270 ( .A1(EXEC_STAGE_mul_ex_mult_76_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U269 ( .A1(EXEC_STAGE_mul_ex_mult_76_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U268 ( .A1(EXEC_STAGE_mul_ex_mult_76_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U267 ( .A1(EXEC_STAGE_mul_ex_mult_76_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U266 ( .A1(EXEC_STAGE_mul_ex_mult_76_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U265 ( .A1(EXEC_STAGE_mul_ex_mult_76_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U264 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U263 ( .A1(EXEC_STAGE_mul_ex_mult_76_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U262 ( .A1(EXEC_STAGE_mul_ex_mult_76_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U261 ( .A1(EXEC_STAGE_mul_ex_mult_76_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U260 ( .A1(EXEC_STAGE_mul_ex_mult_76_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U259 ( .A1(EXEC_STAGE_mul_ex_mult_76_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U258 ( .A1(EXEC_STAGE_mul_ex_mult_76_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U257 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U256 ( .A1(EXEC_STAGE_mul_ex_mult_76_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U255 ( .A1(EXEC_STAGE_mul_ex_mult_76_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U254 ( .A1(EXEC_STAGE_mul_ex_mult_76_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U253 ( .A1(EXEC_STAGE_mul_ex_mult_76_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U252 ( .A1(EXEC_STAGE_mul_ex_mult_76_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U251 ( .A1(EXEC_STAGE_mul_ex_mult_76_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U250 ( .A1(EXEC_STAGE_mul_ex_mult_76_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U249 ( .A1(EXEC_STAGE_mul_ex_mult_76_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U248 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U247 ( .A1(EXEC_STAGE_mul_ex_mult_76_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U246 ( .A1(EXEC_STAGE_mul_ex_mult_76_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U245 ( .A1(EXEC_STAGE_mul_ex_mult_76_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U244 ( .A1(EXEC_STAGE_mul_ex_mult_76_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U243 ( .A1(EXEC_STAGE_mul_ex_mult_76_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U242 ( .A1(EXEC_STAGE_mul_ex_mult_76_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U241 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U240 ( .A1(EXEC_STAGE_mul_ex_mult_76_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U239 ( .A1(EXEC_STAGE_mul_ex_mult_76_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U238 ( .A1(EXEC_STAGE_mul_ex_mult_76_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U237 ( .A1(EXEC_STAGE_mul_ex_mult_76_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U236 ( .A1(EXEC_STAGE_mul_ex_mult_76_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U235 ( .A1(EXEC_STAGE_mul_ex_mult_76_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U234 ( .A1(EXEC_STAGE_mul_ex_mult_76_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U233 ( .A1(EXEC_STAGE_mul_ex_mult_76_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U232 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U231 ( .A1(EXEC_STAGE_mul_ex_mult_76_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U230 ( .A1(EXEC_STAGE_mul_ex_mult_76_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U229 ( .A1(EXEC_STAGE_mul_ex_mult_76_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U228 ( .A1(EXEC_STAGE_mul_ex_mult_76_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U227 ( .A1(EXEC_STAGE_mul_ex_mult_76_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U226 ( .A1(EXEC_STAGE_mul_ex_mult_76_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U225 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U224 ( .A1(EXEC_STAGE_mul_ex_mult_76_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U223 ( .A1(EXEC_STAGE_mul_ex_mult_76_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U222 ( .A1(EXEC_STAGE_mul_ex_mult_76_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U221 ( .A1(EXEC_STAGE_mul_ex_mult_76_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U220 ( .A1(EXEC_STAGE_mul_ex_mult_76_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U219 ( .A1(EXEC_STAGE_mul_ex_mult_76_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U218 ( .A1(EXEC_STAGE_mul_ex_mult_76_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U217 ( .A1(EXEC_STAGE_mul_ex_mult_76_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U216 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U215 ( .A1(EXEC_STAGE_mul_ex_mult_76_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U214 ( .A1(EXEC_STAGE_mul_ex_mult_76_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U213 ( .A1(EXEC_STAGE_mul_ex_mult_76_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U212 ( .A1(EXEC_STAGE_mul_ex_mult_76_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U211 ( .A1(EXEC_STAGE_mul_ex_mult_76_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U210 ( .A1(EXEC_STAGE_mul_ex_mult_76_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U209 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U208 ( .A1(EXEC_STAGE_mul_ex_mult_76_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U207 ( .A1(EXEC_STAGE_mul_ex_mult_76_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U206 ( .A1(EXEC_STAGE_mul_ex_mult_76_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U205 ( .A1(EXEC_STAGE_mul_ex_mult_76_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U204 ( .A1(EXEC_STAGE_mul_ex_mult_76_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U203 ( .A1(EXEC_STAGE_mul_ex_mult_76_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U202 ( .A1(EXEC_STAGE_mul_ex_mult_76_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U201 ( .A1(EXEC_STAGE_mul_ex_mult_76_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U200 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U199 ( .A1(EXEC_STAGE_mul_ex_mult_76_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U198 ( .A1(EXEC_STAGE_mul_ex_mult_76_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U197 ( .A1(EXEC_STAGE_mul_ex_mult_76_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U196 ( .A1(EXEC_STAGE_mul_ex_mult_76_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U195 ( .A1(EXEC_STAGE_mul_ex_mult_76_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U194 ( .A1(EXEC_STAGE_mul_ex_mult_76_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U193 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U192 ( .A1(EXEC_STAGE_mul_ex_mult_76_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U191 ( .A1(EXEC_STAGE_mul_ex_mult_76_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U190 ( .A1(EXEC_STAGE_mul_ex_mult_76_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U189 ( .A1(EXEC_STAGE_mul_ex_mult_76_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U188 ( .A1(EXEC_STAGE_mul_ex_mult_76_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U187 ( .A1(EXEC_STAGE_mul_ex_mult_76_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U186 ( .A1(EXEC_STAGE_mul_ex_mult_76_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U185 ( .A1(EXEC_STAGE_mul_ex_mult_76_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U184 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U183 ( .A1(EXEC_STAGE_mul_ex_mult_76_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U182 ( .A1(EXEC_STAGE_mul_ex_mult_76_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U181 ( .A1(EXEC_STAGE_mul_ex_mult_76_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U180 ( .A1(EXEC_STAGE_mul_ex_mult_76_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U179 ( .A1(EXEC_STAGE_mul_ex_mult_76_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U178 ( .A1(EXEC_STAGE_mul_ex_mult_76_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U177 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U176 ( .A1(EXEC_STAGE_mul_ex_mult_76_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U175 ( .A1(EXEC_STAGE_mul_ex_mult_76_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U174 ( .A1(EXEC_STAGE_mul_ex_mult_76_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U173 ( .A1(EXEC_STAGE_mul_ex_mult_76_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U172 ( .A1(EXEC_STAGE_mul_ex_mult_76_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U171 ( .A1(EXEC_STAGE_mul_ex_mult_76_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U170 ( .A1(EXEC_STAGE_mul_ex_mult_76_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U169 ( .A1(EXEC_STAGE_mul_ex_mult_76_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U168 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U167 ( .A1(EXEC_STAGE_mul_ex_mult_76_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U166 ( .A1(EXEC_STAGE_mul_ex_mult_76_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U165 ( .A1(EXEC_STAGE_mul_ex_mult_76_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U164 ( .A1(EXEC_STAGE_mul_ex_mult_76_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U163 ( .A1(EXEC_STAGE_mul_ex_mult_76_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U162 ( .A1(EXEC_STAGE_mul_ex_mult_76_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U161 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U160 ( .A1(EXEC_STAGE_mul_ex_mult_76_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U159 ( .A1(EXEC_STAGE_mul_ex_mult_76_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U158 ( .A1(EXEC_STAGE_mul_ex_mult_76_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U157 ( .A1(EXEC_STAGE_mul_ex_mult_76_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U156 ( .A1(EXEC_STAGE_mul_ex_mult_76_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U155 ( .A1(EXEC_STAGE_mul_ex_mult_76_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U154 ( .A1(EXEC_STAGE_mul_ex_mult_76_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U153 ( .A1(EXEC_STAGE_mul_ex_mult_76_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U152 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U151 ( .A1(EXEC_STAGE_mul_ex_mult_76_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U150 ( .A1(EXEC_STAGE_mul_ex_mult_76_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U149 ( .A1(EXEC_STAGE_mul_ex_mult_76_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U148 ( .A1(EXEC_STAGE_mul_ex_mult_76_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U147 ( .A1(EXEC_STAGE_mul_ex_mult_76_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U146 ( .A1(EXEC_STAGE_mul_ex_mult_76_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U145 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U144 ( .A1(EXEC_STAGE_mul_ex_mult_76_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U143 ( .A1(EXEC_STAGE_mul_ex_mult_76_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U142 ( .A1(EXEC_STAGE_mul_ex_mult_76_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U141 ( .A1(EXEC_STAGE_mul_ex_mult_76_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U140 ( .A1(EXEC_STAGE_mul_ex_mult_76_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U139 ( .A1(EXEC_STAGE_mul_ex_mult_76_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U138 ( .A1(EXEC_STAGE_mul_ex_mult_76_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U137 ( .A1(EXEC_STAGE_mul_ex_mult_76_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U136 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U135 ( .A1(EXEC_STAGE_mul_ex_mult_76_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U134 ( .A1(EXEC_STAGE_mul_ex_mult_76_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U133 ( .A1(EXEC_STAGE_mul_ex_mult_76_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U132 ( .A1(EXEC_STAGE_mul_ex_mult_76_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U131 ( .A1(EXEC_STAGE_mul_ex_mult_76_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U130 ( .A1(EXEC_STAGE_mul_ex_mult_76_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U129 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U128 ( .A1(EXEC_STAGE_mul_ex_mult_76_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U127 ( .A1(EXEC_STAGE_mul_ex_mult_76_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U126 ( .A1(EXEC_STAGE_mul_ex_mult_76_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U125 ( .A1(EXEC_STAGE_mul_ex_mult_76_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U124 ( .A1(EXEC_STAGE_mul_ex_mult_76_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U123 ( .A1(EXEC_STAGE_mul_ex_mult_76_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U122 ( .A1(EXEC_STAGE_mul_ex_mult_76_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U121 ( .A1(EXEC_STAGE_mul_ex_mult_76_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U120 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U119 ( .A1(EXEC_STAGE_mul_ex_mult_76_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U118 ( .A1(EXEC_STAGE_mul_ex_mult_76_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U117 ( .A1(EXEC_STAGE_mul_ex_mult_76_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U116 ( .A1(EXEC_STAGE_mul_ex_mult_76_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U115 ( .A1(EXEC_STAGE_mul_ex_mult_76_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U114 ( .A1(EXEC_STAGE_mul_ex_mult_76_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U113 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U112 ( .A1(EXEC_STAGE_mul_ex_mult_76_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U111 ( .A1(EXEC_STAGE_mul_ex_mult_76_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U110 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U109 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U108 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U107 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U106 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U105 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U104 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n94), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U103 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U102 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U101 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U100 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U99 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U98 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U97 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U96 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U95 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__9_) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U93 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__14_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_15__15_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n62) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U92 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__1_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n61) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U91 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__0_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n60) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U90 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__2_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n59) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U89 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__4_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n58) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U88 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__6_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n57) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U87 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__8_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n56) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U86 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__10_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__11_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n55) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U85 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__12_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__13_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n54) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U84 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__1_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n53) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U83 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__3_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n52) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U82 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__5_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n51) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U81 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__7_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n50) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U80 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__9_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n49) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U79 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__11_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__12_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n48) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U78 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__13_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__14_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n47) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U77 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__1_), .Z(EXEC_STAGE_mul_ex_N57) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U76 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__2_), .Z(EXEC_STAGE_mul_ex_mult_76_n45)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U75 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__3_), .Z(EXEC_STAGE_mul_ex_mult_76_n44)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U74 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__4_), .Z(EXEC_STAGE_mul_ex_mult_76_n43)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U73 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__5_), .Z(EXEC_STAGE_mul_ex_mult_76_n42)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U72 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__6_), .Z(EXEC_STAGE_mul_ex_mult_76_n41)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U71 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__7_), .Z(EXEC_STAGE_mul_ex_mult_76_n40)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U70 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__8_), .Z(EXEC_STAGE_mul_ex_mult_76_n39)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U69 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__9_), .Z(EXEC_STAGE_mul_ex_mult_76_n38)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U68 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__10_), .Z(EXEC_STAGE_mul_ex_mult_76_n37) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U67 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__11_), .Z(EXEC_STAGE_mul_ex_mult_76_n36) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U66 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__12_), .Z(EXEC_STAGE_mul_ex_mult_76_n35) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U65 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__13_), .Z(EXEC_STAGE_mul_ex_mult_76_n34) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U64 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__14_), .Z(EXEC_STAGE_mul_ex_mult_76_n33) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U63 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__15_), .Z(EXEC_STAGE_mul_ex_mult_76_n32) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U62 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__15_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__14_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n31) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U61 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__4_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n30) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U60 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__6_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n29) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U59 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__8_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n28) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U58 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__10_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n27) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U57 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__12_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n26) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U56 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__14_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n25) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U55 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__2_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n24) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U54 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__3_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n23) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U53 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__5_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n22) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U52 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__7_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n21) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U51 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__9_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n20) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U50 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__11_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n19) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U49 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__13_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n18) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U48 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_15__15_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n17) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U47 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__1_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__0_), .ZN(EXEC_STAGE_mul_ex_mult_76_n16) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U46 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__2_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__1_), .ZN(EXEC_STAGE_mul_ex_mult_76_n15) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U45 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__3_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__2_), .ZN(EXEC_STAGE_mul_ex_mult_76_n14) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U44 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__4_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__3_), .ZN(EXEC_STAGE_mul_ex_mult_76_n13) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U43 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__5_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__4_), .ZN(EXEC_STAGE_mul_ex_mult_76_n12) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U42 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__6_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__5_), .ZN(EXEC_STAGE_mul_ex_mult_76_n11) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U41 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__7_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__6_), .ZN(EXEC_STAGE_mul_ex_mult_76_n10) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U40 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__8_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__7_), .ZN(EXEC_STAGE_mul_ex_mult_76_n9)
         );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U39 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__9_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__8_), .ZN(EXEC_STAGE_mul_ex_mult_76_n8)
         );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U38 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__10_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__9_), .ZN(EXEC_STAGE_mul_ex_mult_76_n7)
         );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U37 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__11_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__10_), .ZN(EXEC_STAGE_mul_ex_mult_76_n6) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U36 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__12_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__11_), .ZN(EXEC_STAGE_mul_ex_mult_76_n5) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U35 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__13_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__12_), .ZN(EXEC_STAGE_mul_ex_mult_76_n4) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U34 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__14_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__13_), .ZN(EXEC_STAGE_mul_ex_mult_76_n3) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U33 ( .A(ID_EXEC_OUT[251]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n65) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U32 ( .A(ID_EXEC_OUT[219]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n64) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U31 ( .A(ID_EXEC_OUT[217]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n68) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U30 ( .A(ID_EXEC_OUT[216]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n88) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U29 ( .A(ID_EXEC_OUT[215]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n78) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U28 ( .A(ID_EXEC_OUT[214]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n80) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U27 ( .A(ID_EXEC_OUT[213]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n90) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U26 ( .A(ID_EXEC_OUT[212]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n82) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U25 ( .A(ID_EXEC_OUT[211]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n76) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U24 ( .A(ID_EXEC_OUT[210]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n86) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U23 ( .A(ID_EXEC_OUT[209]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n84) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U22 ( .A(ID_EXEC_OUT[208]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n92) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U21 ( .A(ID_EXEC_OUT[207]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n70) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U20 ( .A(ID_EXEC_OUT[206]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n74) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U19 ( .A(ID_EXEC_OUT[205]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n72) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U18 ( .A(ID_EXEC_OUT[204]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n63) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U17 ( .A(ID_EXEC_OUT[218]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n66) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U16 ( .A(ID_EXEC_OUT[250]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n67) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U15 ( .A(ID_EXEC_OUT[249]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n69) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U14 ( .A(ID_EXEC_OUT[236]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n94) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U13 ( .A(ID_EXEC_OUT[237]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n73) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U12 ( .A(ID_EXEC_OUT[248]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n89) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U11 ( .A(ID_EXEC_OUT[247]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n79) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U10 ( .A(ID_EXEC_OUT[246]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n81) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U9 ( .A(ID_EXEC_OUT[245]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n91) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U8 ( .A(ID_EXEC_OUT[244]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n83) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U7 ( .A(ID_EXEC_OUT[243]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n77) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U6 ( .A(ID_EXEC_OUT[242]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n87) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U5 ( .A(ID_EXEC_OUT[241]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n85) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U4 ( .A(ID_EXEC_OUT[240]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n93) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U3 ( .A(ID_EXEC_OUT[239]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n71) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U2 ( .A(ID_EXEC_OUT[238]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n75) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_2_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__14_), .B(EXEC_STAGE_mul_ex_mult_76_n31), .CI(EXEC_STAGE_mul_ex_mult_76_ab_1__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__13_), .B(EXEC_STAGE_mul_ex_mult_76_n3), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n32), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__12_), .B(EXEC_STAGE_mul_ex_mult_76_n4), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n33), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__11_), .B(EXEC_STAGE_mul_ex_mult_76_n5), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n34), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__10_), .B(EXEC_STAGE_mul_ex_mult_76_n6), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n35), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__9_), .B(EXEC_STAGE_mul_ex_mult_76_n7), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n36), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__8_), .B(EXEC_STAGE_mul_ex_mult_76_n8), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n37), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__7_), .B(EXEC_STAGE_mul_ex_mult_76_n9), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n38), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__6_), .B(EXEC_STAGE_mul_ex_mult_76_n10), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n39), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__5_), .B(EXEC_STAGE_mul_ex_mult_76_n11), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n40), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__4_), .B(EXEC_STAGE_mul_ex_mult_76_n12), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n41), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__3_), .B(EXEC_STAGE_mul_ex_mult_76_n13), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n42), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__2_), .B(EXEC_STAGE_mul_ex_mult_76_n14), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n43), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__1_), .B(EXEC_STAGE_mul_ex_mult_76_n15), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n44), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_2_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__0_), .B(EXEC_STAGE_mul_ex_mult_76_n16), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n45), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_0_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_3_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_2__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_3_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_4_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_3__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_4_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_5_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_4__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_5_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_6_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_5__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_6_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_7_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_6__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_7_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_8_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_7__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_8_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_9_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_8__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_9_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_10_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_9__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_10_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_11_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_10__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_11_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_12_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_11__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_12_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_13_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_12__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_13_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_14_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_13__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_14_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S5_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_14__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__0_) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U100 ( .A(
        EXEC_STAGE_mul_ex_mult_76_n61), .Z(EXEC_STAGE_mul_ex_N72) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U99 ( .A(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__0_), .Z(EXEC_STAGE_mul_ex_N71) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U98 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_12_), .Z(EXEC_STAGE_mul_ex_N70) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U97 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_11_), .Z(EXEC_STAGE_mul_ex_N69) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U96 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_10_), .Z(EXEC_STAGE_mul_ex_N68) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U95 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_9_), .Z(EXEC_STAGE_mul_ex_N67) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U94 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_8_), .Z(EXEC_STAGE_mul_ex_N66) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U93 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_7_), .Z(EXEC_STAGE_mul_ex_N65) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U92 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_6_), .Z(EXEC_STAGE_mul_ex_N64) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U91 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_5_), .Z(EXEC_STAGE_mul_ex_N63) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U90 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_4_), .Z(EXEC_STAGE_mul_ex_N62) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U89 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_3_), .Z(EXEC_STAGE_mul_ex_N61) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U88 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_2_), .Z(EXEC_STAGE_mul_ex_N60) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U87 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_1_), .Z(EXEC_STAGE_mul_ex_N59) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U86 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_0_), .Z(EXEC_STAGE_mul_ex_N58) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U85 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n60), .A2(EXEC_STAGE_mul_ex_mult_76_n24), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n70) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U84 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n53), .A2(EXEC_STAGE_mul_ex_mult_76_n23), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n67) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U83 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n53), .A2(EXEC_STAGE_mul_ex_mult_76_n23), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n68) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U82 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n67), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n69) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U81 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n17), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n69), .Z(EXEC_STAGE_mul_ex_N74) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U80 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n59), .A2(EXEC_STAGE_mul_ex_mult_76_n30), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n63) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U79 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n59), .A2(EXEC_STAGE_mul_ex_mult_76_n30), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n65) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U78 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n15), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n66) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U77 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n16), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n17), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n64) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U76 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n66), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n64), .Z(EXEC_STAGE_mul_ex_N75) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U75 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n63), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n64), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n59) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U74 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n52), .A2(EXEC_STAGE_mul_ex_mult_76_n22), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n60) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U73 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n52), .A2(EXEC_STAGE_mul_ex_mult_76_n22), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n61) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U72 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n60), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n61), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n62) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U71 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n59), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n62), .Z(EXEC_STAGE_mul_ex_N76) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U70 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n58), .A2(EXEC_STAGE_mul_ex_mult_76_n29), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n55) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U69 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n58), .A2(EXEC_STAGE_mul_ex_mult_76_n29), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n57) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U68 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n13), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n57), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n58) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U67 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n14), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n59), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n60), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n56) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U66 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n58), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n56), .Z(EXEC_STAGE_mul_ex_N77) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U65 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n55), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n56), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n57), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n51) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U64 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n51), .A2(EXEC_STAGE_mul_ex_mult_76_n21), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n52) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U63 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n51), .A2(EXEC_STAGE_mul_ex_mult_76_n21), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n53) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U62 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n52), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n54) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U61 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n51), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n54), .Z(EXEC_STAGE_mul_ex_N78) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U60 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n57), .A2(EXEC_STAGE_mul_ex_mult_76_n28), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n47) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U59 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n57), .A2(EXEC_STAGE_mul_ex_mult_76_n28), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n49) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U58 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n11), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n49), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n50) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U57 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n12), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n51), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n48) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U56 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n50), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n48), .Z(EXEC_STAGE_mul_ex_N79) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U55 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n47), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n48), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n49), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n43) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U54 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n50), .A2(EXEC_STAGE_mul_ex_mult_76_n20), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n44) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U53 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n50), .A2(EXEC_STAGE_mul_ex_mult_76_n20), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n45) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U52 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n44), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n45), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n46) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U51 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n43), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n46), .Z(EXEC_STAGE_mul_ex_N80) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U50 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n56), .A2(EXEC_STAGE_mul_ex_mult_76_n27), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n39) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U49 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n56), .A2(EXEC_STAGE_mul_ex_mult_76_n27), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n41) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U48 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n9), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n41), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n42) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U47 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n10), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n43), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n44), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n40) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U46 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n42), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n40), .Z(EXEC_STAGE_mul_ex_N81) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U45 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n39), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n40), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n41), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n35) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U44 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n49), .A2(EXEC_STAGE_mul_ex_mult_76_n19), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n36) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U43 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n49), .A2(EXEC_STAGE_mul_ex_mult_76_n19), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n37) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U42 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n36), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n37), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n38) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U41 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n35), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n38), .Z(EXEC_STAGE_mul_ex_N82) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U40 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n55), .A2(EXEC_STAGE_mul_ex_mult_76_n26), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n31) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U39 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n55), .A2(EXEC_STAGE_mul_ex_mult_76_n26), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n33) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U38 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n7), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n33), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n34) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U37 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n8), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n35), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n36), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n32) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U36 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n34), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n32), .Z(EXEC_STAGE_mul_ex_N83) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U35 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n31), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n32), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n33), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n27) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U34 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n48), .A2(EXEC_STAGE_mul_ex_mult_76_n18), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n28) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U33 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n48), .A2(EXEC_STAGE_mul_ex_mult_76_n18), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n29) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U32 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n28), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n29), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n30) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U31 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n27), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n30), .Z(EXEC_STAGE_mul_ex_N84) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U30 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n54), .A2(EXEC_STAGE_mul_ex_mult_76_n25), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n23) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U29 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n54), .A2(EXEC_STAGE_mul_ex_mult_76_n25), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n25) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U28 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n5), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n25), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n26) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U27 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n6), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n27), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n28), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n24) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U26 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n26), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n24), .Z(EXEC_STAGE_mul_ex_N85) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U25 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n23), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n24), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n25), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n19) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U24 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n47), .A2(EXEC_STAGE_mul_ex_mult_76_n17), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n20) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U23 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n47), .A2(EXEC_STAGE_mul_ex_mult_76_n17), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n21) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U22 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n20), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n21), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n22) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U21 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n19), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n22), .Z(EXEC_STAGE_mul_ex_N86) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U20 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n19), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n4), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n20), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n18) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U19 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n3), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n18), .Z(EXEC_STAGE_mul_ex_N87) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U18 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n17) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U17 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n16) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U16 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n15) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U15 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n61), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n14) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n55), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n13) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n12) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n47), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n11) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n45), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n10) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n39), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n9) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n37), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n8) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n31), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n7) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n29), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n6) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n23), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n5) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n21), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n4) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U4 ( .A(EXEC_STAGE_mul_ex_mult_76_n62), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n3) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U3 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n1), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n70), .ZN(EXEC_STAGE_mul_ex_N73) );
  OR2_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U2 ( .A1(EXEC_STAGE_mul_ex_mult_76_n60), .A2(EXEC_STAGE_mul_ex_mult_76_n24), .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n1)
         );
endmodule

