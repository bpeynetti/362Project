module execute (
    //inputs
    nextPC_in,opA_in,opB_in,offset26_in,offset16_in,destReg_in,PCtoReg_in,
    RegToPC_in,jump_in,branch_in,branchZero_in,RType_in,RegWrite_in,MemToReg_in,
    MemWrite_in,loadSign_in,mul_in,DSize_in,ALUCtrl_in,
    //basic clk, reset input
    clk,reset,
    //outputs
    aluResult_out, leapAddr_out, destReg_out, leap_out,
    PCtoReg_out, RegToPC_out, 
    // jump_out, branch_out, branchZero_out,
    RegWrite_out, MemToReg_out, MemWrite_out, loadSign_out, DSize_out
    );
    
    input [0:31] nextPC_in;
    input [0:31] opA_in;
    input [0:31] opB_in;
    input [0:25] offset_26_in;
    input [0:15] offset_16_in;
    input [0:4] destReg_in;
    input PCtoReg_in;
    input RegToPC_in;
    input jump_in;
    input branch_in;
    input branchZero_in;
    input RType_in;
    input RegWrite_in;
    input MemToReg_in;
    input MemWrite_in;
    input loadSign_in;
    input mul_in;
    input [0:1] DSize_in;
    input [0:3] ALUCtrl_in;
    input clk,reset;
    
    output [0:31] nextPC_out;
    output [0:31] aluResult_out;
    output [0:31] leapAddr_out;
    output [0:4] destReg_out;
    output leap_out;
    output PCtoReg_out;
    output RegToPC_out;
    output RegWrite_out;
    output MemToReg_out;
    output MemWrite_out;
    output loadSign_out;
    output [0:1] DSize_out;
    
    wire [0:31] imm16_32, imm26_32, imm_final;
    wire sum_cout, sum_of;
    wire zero, of;
    wire not_mul_result, mul_result;
    
    assign PCtoReg_out = PCtoReg_in;
    assign RegToPC_out = RegToPC_in;
    assign RegWrite_out = RegWrite_in;
    assign MemToReg_out = MemToReg_in;
    assign MemWrite_out = MemWrite_in;
    assign loadSign_out = loadSign_in;
    assign DSize_out = DSize_in;
    
    alu alu_ex(
       .A(opA),
       .B(opB),
       .ctrl(ALUCtrl),
       .ALUout(not_mul_result),
       .zero(zero),
       .of(of)
    );
    
    multiplier mul_ex(
        .X(opA),
        .Y(opB),
        .Z(mul_result)
    );
    
    mux2to1_32bit choose_result(
        .X(not_mul_result),
        .Y(mul_result),
        .sel(mul),
        .Z(aluResult)
    );
    
    check_branch decide_if_leap(
        .busA(not_mul_result),
        .branchZero(branchZero),
        .branch(branch),
        .jump(jump),
        .leap(leap)
    );
    
    //SHOULDN'T THESE BY SIGN EXTEND? RIGHT NOW THEY ARE BOTH ZERO EXTEND (taken from PC LOGIC)
    extend_16to32 EXTEND_IMM16(offset16, 1'b0, imm16_32);
    extend_26to32 EXTEND_IMM26(offset26, 1'b0, imm26_32);
    mux2to1_32bit CHOOSE_IMMEDIATE(imm26_32, imm16_32, branch, imm_final);
    
    fa_nbit ADD_IMM(imm_final, nextPC, 1'b0, pc_nonreg, sum_cout, sum_of);
    mux2to1_32bit IMM_OR_REG(pc_nonreg, opA, regToPC, leapAddr);
        
endmodule