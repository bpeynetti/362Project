
module execute ( nextPC_in, opA_in, opB_in, offset26_in, offset16_in, 
        destReg_in, PCtoReg_in, RegToPC_in, jump_in, branch_in, branchZero_in, 
        RType_in, RegWrite_in, MemToReg_in, MemWrite_in, loadSign_in, mul_in, 
        DSize_in, ALUCtrl_in, memVal_in, f1_in, f2_in, fDestReg_in, FPRType_in, 
        FPRegWrite_in, movfp2i_in, movi2fp_in, clk, reset, nextPC_out, 
        aluResult_out, leapAddr_out, destReg_out, leap_out, PCtoReg_out, 
        RegToPC_out, RegWrite_out, MemToReg_out, MemWrite_out, loadSign_out, 
        DSize_out, memVal_out, stall_out, fDestReg_out, fbusW, FPRegWrite_out, 
        mul_out );
  input [0:31] nextPC_in;
  input [0:31] opA_in;
  input [0:31] opB_in;
  input [0:25] offset26_in;
  input [0:15] offset16_in;
  input [0:4] destReg_in;
  input [0:1] DSize_in;
  input [0:3] ALUCtrl_in;
  input [0:31] memVal_in;
  input [0:31] f1_in;
  input [0:31] f2_in;
  input [0:4] fDestReg_in;
  output [0:31] nextPC_out;
  output [0:31] aluResult_out;
  output [0:31] leapAddr_out;
  output [0:4] destReg_out;
  output [0:1] DSize_out;
  output [0:31] memVal_out;
  output [0:4] fDestReg_out;
  output [0:63] fbusW;
  input PCtoReg_in, RegToPC_in, jump_in, branch_in, branchZero_in, RType_in,
         RegWrite_in, MemToReg_in, MemWrite_in, loadSign_in, mul_in,
         FPRType_in, FPRegWrite_in, movfp2i_in, movi2fp_in, clk, reset;
  output leap_out, PCtoReg_out, RegToPC_out, RegWrite_out, MemToReg_out,
         MemWrite_out, loadSign_out, stall_out, FPRegWrite_out, mul_out;
  wire   mul_done, n2, alu_ex_n4, alu_ex_n1, alu_ex_sgt_out_31_,
         alu_ex_sge_out_31_, alu_ex_slt_out_31_, alu_ex_sle_out_31_,
         alu_ex_sne_out_31_, alu_ex_seq_out_31_, alu_ex_sgt_1bit,
         alu_ex_sge_1bit, alu_ex_slt_1bit, alu_ex_sle_1bit, alu_ex_sne_1bit,
         alu_ex_shift_out_31_, alu_ex_shift_out_30_, alu_ex_shift_out_29_,
         alu_ex_shift_out_28_, alu_ex_shift_out_27_, alu_ex_shift_out_26_,
         alu_ex_shift_out_25_, alu_ex_shift_out_24_, alu_ex_shift_out_23_,
         alu_ex_shift_out_22_, alu_ex_shift_out_21_, alu_ex_shift_out_20_,
         alu_ex_shift_out_19_, alu_ex_shift_out_18_, alu_ex_shift_out_17_,
         alu_ex_shift_out_16_, alu_ex_shift_out_15_, alu_ex_shift_out_14_,
         alu_ex_shift_out_13_, alu_ex_shift_out_12_, alu_ex_shift_out_11_,
         alu_ex_shift_out_10_, alu_ex_shift_out_9_, alu_ex_shift_out_8_,
         alu_ex_shift_out_7_, alu_ex_shift_out_6_, alu_ex_shift_out_5_,
         alu_ex_shift_out_4_, alu_ex_shift_out_3_, alu_ex_shift_out_2_,
         alu_ex_shift_out_1_, alu_ex_shift_out_0_, alu_ex_add_sub_out_31_,
         alu_ex_add_sub_out_30_, alu_ex_add_sub_out_29_,
         alu_ex_add_sub_out_28_, alu_ex_add_sub_out_27_,
         alu_ex_add_sub_out_26_, alu_ex_add_sub_out_25_,
         alu_ex_add_sub_out_24_, alu_ex_add_sub_out_23_,
         alu_ex_add_sub_out_22_, alu_ex_add_sub_out_21_,
         alu_ex_add_sub_out_20_, alu_ex_add_sub_out_19_,
         alu_ex_add_sub_out_18_, alu_ex_add_sub_out_17_,
         alu_ex_add_sub_out_16_, alu_ex_add_sub_out_15_,
         alu_ex_add_sub_out_14_, alu_ex_add_sub_out_13_,
         alu_ex_add_sub_out_12_, alu_ex_add_sub_out_11_,
         alu_ex_add_sub_out_10_, alu_ex_add_sub_out_9_, alu_ex_add_sub_out_8_,
         alu_ex_add_sub_out_7_, alu_ex_add_sub_out_6_, alu_ex_add_sub_out_5_,
         alu_ex_add_sub_out_4_, alu_ex_add_sub_out_3_, alu_ex_add_sub_out_2_,
         alu_ex_add_sub_out_1_, alu_ex_add_sub_out_0_, alu_ex_and_out_31_,
         alu_ex_and_out_30_, alu_ex_and_out_29_, alu_ex_and_out_28_,
         alu_ex_and_out_27_, alu_ex_and_out_26_, alu_ex_and_out_25_,
         alu_ex_and_out_24_, alu_ex_and_out_23_, alu_ex_and_out_22_,
         alu_ex_and_out_21_, alu_ex_and_out_20_, alu_ex_and_out_19_,
         alu_ex_and_out_18_, alu_ex_and_out_17_, alu_ex_and_out_16_,
         alu_ex_and_out_15_, alu_ex_and_out_14_, alu_ex_and_out_13_,
         alu_ex_and_out_12_, alu_ex_and_out_11_, alu_ex_and_out_10_,
         alu_ex_and_out_9_, alu_ex_and_out_8_, alu_ex_and_out_7_,
         alu_ex_and_out_6_, alu_ex_and_out_5_, alu_ex_and_out_4_,
         alu_ex_and_out_3_, alu_ex_and_out_2_, alu_ex_and_out_1_,
         alu_ex_and_out_0_, alu_ex_n3, alu_ex_ADD_OR_SUB_n4,
         alu_ex_ADD_OR_SUB_n3, alu_ex_ADD_OR_SUB_n2, alu_ex_ADD_OR_SUB_n1,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_30__MUX_n3,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_30__MUX_n2,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_31__MUX_n3,
         alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_31__MUX_n2,
         alu_ex_FULL_ADDER_FA_NBIT_0__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_1__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_1__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_1__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_1__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_2__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_2__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_2__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_2__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_3__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_3__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_3__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_3__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_4__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_4__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_4__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_4__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_5__FA_n6,
         alu_ex_FULL_ADDER_FA_NBIT_5__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_5__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_5__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_6__FA_n6,
         alu_ex_FULL_ADDER_FA_NBIT_6__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_6__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_6__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_6__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_6__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_7__FA_n8,
         alu_ex_FULL_ADDER_FA_NBIT_7__FA_n6,
         alu_ex_FULL_ADDER_FA_NBIT_7__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_7__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_7__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_7__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_7__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_8__FA_n8,
         alu_ex_FULL_ADDER_FA_NBIT_8__FA_n6,
         alu_ex_FULL_ADDER_FA_NBIT_8__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_8__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_8__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_8__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_8__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_9__FA_n6,
         alu_ex_FULL_ADDER_FA_NBIT_9__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_9__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_9__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_9__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_9__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_10__FA_n8,
         alu_ex_FULL_ADDER_FA_NBIT_10__FA_n6,
         alu_ex_FULL_ADDER_FA_NBIT_10__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_10__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_10__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_10__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_10__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_11__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_11__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_11__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_11__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_11__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_12__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_12__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_12__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_12__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_12__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_13__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_13__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_13__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_13__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_13__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_14__FA_n8,
         alu_ex_FULL_ADDER_FA_NBIT_14__FA_n6,
         alu_ex_FULL_ADDER_FA_NBIT_14__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_14__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_14__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_14__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_14__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_15__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_15__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_15__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_15__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_15__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_16__FA_n8,
         alu_ex_FULL_ADDER_FA_NBIT_16__FA_n6,
         alu_ex_FULL_ADDER_FA_NBIT_16__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_16__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_16__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_16__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_16__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_17__FA_n8,
         alu_ex_FULL_ADDER_FA_NBIT_17__FA_n6,
         alu_ex_FULL_ADDER_FA_NBIT_17__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_17__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_17__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_17__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_17__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_18__FA_n8,
         alu_ex_FULL_ADDER_FA_NBIT_18__FA_n6,
         alu_ex_FULL_ADDER_FA_NBIT_18__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_18__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_18__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_18__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_18__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_19__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_19__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_19__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_19__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_19__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_20__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_20__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_20__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_20__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_20__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_21__FA_n7,
         alu_ex_FULL_ADDER_FA_NBIT_21__FA_n6,
         alu_ex_FULL_ADDER_FA_NBIT_21__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_21__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_21__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_21__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_21__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_22__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_22__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_22__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_22__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_22__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_23__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_23__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_23__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_23__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_23__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_24__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_24__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_24__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_24__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_24__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_25__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_25__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_25__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_25__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_25__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_26__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_26__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_26__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_26__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_26__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_27__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_27__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_27__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_27__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_27__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_28__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_28__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_28__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_28__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_28__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_29__FA_n6,
         alu_ex_FULL_ADDER_FA_NBIT_29__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_29__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_29__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_29__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_29__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_30__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_30__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_30__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_30__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_30__FA_n1,
         alu_ex_FULL_ADDER_FA_NBIT_31__FA_n5,
         alu_ex_FULL_ADDER_FA_NBIT_31__FA_n4,
         alu_ex_FULL_ADDER_FA_NBIT_31__FA_n3,
         alu_ex_FULL_ADDER_FA_NBIT_31__FA_n2,
         alu_ex_FULL_ADDER_FA_NBIT_31__FA_n1, alu_ex_SHIFTER_n12,
         alu_ex_SHIFTER_n11, alu_ex_SHIFTER_n10, alu_ex_SHIFTER_n9,
         alu_ex_SHIFTER_n8, alu_ex_SHIFTER_n7, alu_ex_SHIFTER_n6,
         alu_ex_SHIFTER_n5, alu_ex_SHIFTER_n4, alu_ex_SHIFTER_n3,
         alu_ex_SHIFTER_n2, alu_ex_SHIFTER_n1, alu_ex_SHIFTER_rtemp3_31_,
         alu_ex_SHIFTER_rtemp3_30_, alu_ex_SHIFTER_rtemp3_29_,
         alu_ex_SHIFTER_rtemp3_28_, alu_ex_SHIFTER_rtemp3_27_,
         alu_ex_SHIFTER_rtemp3_26_, alu_ex_SHIFTER_rtemp3_25_,
         alu_ex_SHIFTER_rtemp3_24_, alu_ex_SHIFTER_rtemp3_23_,
         alu_ex_SHIFTER_rtemp3_22_, alu_ex_SHIFTER_rtemp3_21_,
         alu_ex_SHIFTER_rtemp3_20_, alu_ex_SHIFTER_rtemp3_19_,
         alu_ex_SHIFTER_rtemp3_18_, alu_ex_SHIFTER_rtemp3_17_,
         alu_ex_SHIFTER_rtemp3_16_, alu_ex_SHIFTER_rtemp3_15_,
         alu_ex_SHIFTER_rtemp3_14_, alu_ex_SHIFTER_rtemp3_13_,
         alu_ex_SHIFTER_rtemp3_12_, alu_ex_SHIFTER_rtemp3_11_,
         alu_ex_SHIFTER_rtemp3_10_, alu_ex_SHIFTER_rtemp3_9_,
         alu_ex_SHIFTER_rtemp3_8_, alu_ex_SHIFTER_rtemp3_7_,
         alu_ex_SHIFTER_rtemp3_6_, alu_ex_SHIFTER_rtemp3_5_,
         alu_ex_SHIFTER_rtemp3_4_, alu_ex_SHIFTER_rtemp3_3_,
         alu_ex_SHIFTER_rtemp3_2_, alu_ex_SHIFTER_rtemp3_1_,
         alu_ex_SHIFTER_rtemp3_0_, alu_ex_SHIFTER_rtemp2_31_,
         alu_ex_SHIFTER_rtemp2_30_, alu_ex_SHIFTER_rtemp2_29_,
         alu_ex_SHIFTER_rtemp2_28_, alu_ex_SHIFTER_rtemp2_27_,
         alu_ex_SHIFTER_rtemp2_26_, alu_ex_SHIFTER_rtemp2_25_,
         alu_ex_SHIFTER_rtemp2_24_, alu_ex_SHIFTER_rtemp2_23_,
         alu_ex_SHIFTER_rtemp2_22_, alu_ex_SHIFTER_rtemp2_21_,
         alu_ex_SHIFTER_rtemp2_20_, alu_ex_SHIFTER_rtemp2_19_,
         alu_ex_SHIFTER_rtemp2_18_, alu_ex_SHIFTER_rtemp2_17_,
         alu_ex_SHIFTER_rtemp2_16_, alu_ex_SHIFTER_rtemp2_15_,
         alu_ex_SHIFTER_rtemp2_14_, alu_ex_SHIFTER_rtemp2_13_,
         alu_ex_SHIFTER_rtemp2_12_, alu_ex_SHIFTER_rtemp2_11_,
         alu_ex_SHIFTER_rtemp2_10_, alu_ex_SHIFTER_rtemp2_9_,
         alu_ex_SHIFTER_rtemp2_8_, alu_ex_SHIFTER_rtemp2_7_,
         alu_ex_SHIFTER_rtemp2_6_, alu_ex_SHIFTER_rtemp2_5_,
         alu_ex_SHIFTER_rtemp2_4_, alu_ex_SHIFTER_rtemp2_3_,
         alu_ex_SHIFTER_rtemp2_2_, alu_ex_SHIFTER_rtemp2_1_,
         alu_ex_SHIFTER_rtemp2_0_, alu_ex_SHIFTER_rtemp1_31_,
         alu_ex_SHIFTER_rtemp1_30_, alu_ex_SHIFTER_rtemp1_29_,
         alu_ex_SHIFTER_rtemp1_28_, alu_ex_SHIFTER_rtemp1_27_,
         alu_ex_SHIFTER_rtemp1_26_, alu_ex_SHIFTER_rtemp1_25_,
         alu_ex_SHIFTER_rtemp1_24_, alu_ex_SHIFTER_rtemp1_23_,
         alu_ex_SHIFTER_rtemp1_22_, alu_ex_SHIFTER_rtemp1_21_,
         alu_ex_SHIFTER_rtemp1_20_, alu_ex_SHIFTER_rtemp1_19_,
         alu_ex_SHIFTER_rtemp1_18_, alu_ex_SHIFTER_rtemp1_17_,
         alu_ex_SHIFTER_rtemp1_16_, alu_ex_SHIFTER_rtemp1_15_,
         alu_ex_SHIFTER_rtemp1_14_, alu_ex_SHIFTER_rtemp1_13_,
         alu_ex_SHIFTER_rtemp1_12_, alu_ex_SHIFTER_rtemp1_11_,
         alu_ex_SHIFTER_rtemp1_10_, alu_ex_SHIFTER_rtemp1_9_,
         alu_ex_SHIFTER_rtemp1_8_, alu_ex_SHIFTER_rtemp1_7_,
         alu_ex_SHIFTER_rtemp1_6_, alu_ex_SHIFTER_rtemp1_5_,
         alu_ex_SHIFTER_rtemp1_4_, alu_ex_SHIFTER_rtemp1_3_,
         alu_ex_SHIFTER_rtemp1_2_, alu_ex_SHIFTER_rtemp1_1_,
         alu_ex_SHIFTER_rtemp1_0_, alu_ex_SHIFTER_rtemp0_31_,
         alu_ex_SHIFTER_rtemp0_30_, alu_ex_SHIFTER_rtemp0_29_,
         alu_ex_SHIFTER_rtemp0_28_, alu_ex_SHIFTER_rtemp0_27_,
         alu_ex_SHIFTER_rtemp0_26_, alu_ex_SHIFTER_rtemp0_25_,
         alu_ex_SHIFTER_rtemp0_24_, alu_ex_SHIFTER_rtemp0_23_,
         alu_ex_SHIFTER_rtemp0_22_, alu_ex_SHIFTER_rtemp0_21_,
         alu_ex_SHIFTER_rtemp0_20_, alu_ex_SHIFTER_rtemp0_19_,
         alu_ex_SHIFTER_rtemp0_18_, alu_ex_SHIFTER_rtemp0_17_,
         alu_ex_SHIFTER_rtemp0_16_, alu_ex_SHIFTER_rtemp0_15_,
         alu_ex_SHIFTER_rtemp0_14_, alu_ex_SHIFTER_rtemp0_13_,
         alu_ex_SHIFTER_rtemp0_12_, alu_ex_SHIFTER_rtemp0_11_,
         alu_ex_SHIFTER_rtemp0_10_, alu_ex_SHIFTER_rtemp0_9_,
         alu_ex_SHIFTER_rtemp0_8_, alu_ex_SHIFTER_rtemp0_7_,
         alu_ex_SHIFTER_rtemp0_6_, alu_ex_SHIFTER_rtemp0_5_,
         alu_ex_SHIFTER_rtemp0_4_, alu_ex_SHIFTER_rtemp0_3_,
         alu_ex_SHIFTER_rtemp0_2_, alu_ex_SHIFTER_rtemp0_1_,
         alu_ex_SHIFTER_rtemp0_0_, alu_ex_SHIFTER_ltemp3_31_,
         alu_ex_SHIFTER_ltemp3_30_, alu_ex_SHIFTER_ltemp3_29_,
         alu_ex_SHIFTER_ltemp3_28_, alu_ex_SHIFTER_ltemp3_27_,
         alu_ex_SHIFTER_ltemp3_26_, alu_ex_SHIFTER_ltemp3_25_,
         alu_ex_SHIFTER_ltemp3_24_, alu_ex_SHIFTER_ltemp3_23_,
         alu_ex_SHIFTER_ltemp3_22_, alu_ex_SHIFTER_ltemp3_21_,
         alu_ex_SHIFTER_ltemp3_20_, alu_ex_SHIFTER_ltemp3_19_,
         alu_ex_SHIFTER_ltemp3_18_, alu_ex_SHIFTER_ltemp3_17_,
         alu_ex_SHIFTER_ltemp3_16_, alu_ex_SHIFTER_ltemp3_15_,
         alu_ex_SHIFTER_ltemp3_14_, alu_ex_SHIFTER_ltemp3_13_,
         alu_ex_SHIFTER_ltemp3_12_, alu_ex_SHIFTER_ltemp3_11_,
         alu_ex_SHIFTER_ltemp3_10_, alu_ex_SHIFTER_ltemp3_9_,
         alu_ex_SHIFTER_ltemp3_8_, alu_ex_SHIFTER_ltemp3_7_,
         alu_ex_SHIFTER_ltemp3_6_, alu_ex_SHIFTER_ltemp3_5_,
         alu_ex_SHIFTER_ltemp3_4_, alu_ex_SHIFTER_ltemp3_3_,
         alu_ex_SHIFTER_ltemp3_2_, alu_ex_SHIFTER_ltemp3_1_,
         alu_ex_SHIFTER_ltemp3_0_, alu_ex_SHIFTER_ltemp2_31_,
         alu_ex_SHIFTER_ltemp2_30_, alu_ex_SHIFTER_ltemp2_29_,
         alu_ex_SHIFTER_ltemp2_28_, alu_ex_SHIFTER_ltemp2_27_,
         alu_ex_SHIFTER_ltemp2_26_, alu_ex_SHIFTER_ltemp2_25_,
         alu_ex_SHIFTER_ltemp2_24_, alu_ex_SHIFTER_ltemp2_23_,
         alu_ex_SHIFTER_ltemp2_22_, alu_ex_SHIFTER_ltemp2_21_,
         alu_ex_SHIFTER_ltemp2_20_, alu_ex_SHIFTER_ltemp2_19_,
         alu_ex_SHIFTER_ltemp2_18_, alu_ex_SHIFTER_ltemp2_17_,
         alu_ex_SHIFTER_ltemp2_16_, alu_ex_SHIFTER_ltemp2_15_,
         alu_ex_SHIFTER_ltemp2_14_, alu_ex_SHIFTER_ltemp2_13_,
         alu_ex_SHIFTER_ltemp2_12_, alu_ex_SHIFTER_ltemp2_11_,
         alu_ex_SHIFTER_ltemp2_10_, alu_ex_SHIFTER_ltemp2_9_,
         alu_ex_SHIFTER_ltemp2_8_, alu_ex_SHIFTER_ltemp2_7_,
         alu_ex_SHIFTER_ltemp2_6_, alu_ex_SHIFTER_ltemp2_5_,
         alu_ex_SHIFTER_ltemp2_4_, alu_ex_SHIFTER_ltemp2_3_,
         alu_ex_SHIFTER_ltemp2_2_, alu_ex_SHIFTER_ltemp2_1_,
         alu_ex_SHIFTER_ltemp2_0_, alu_ex_SHIFTER_ltemp1_31_,
         alu_ex_SHIFTER_ltemp1_30_, alu_ex_SHIFTER_ltemp1_29_,
         alu_ex_SHIFTER_ltemp1_28_, alu_ex_SHIFTER_ltemp1_27_,
         alu_ex_SHIFTER_ltemp1_26_, alu_ex_SHIFTER_ltemp1_25_,
         alu_ex_SHIFTER_ltemp1_24_, alu_ex_SHIFTER_ltemp1_23_,
         alu_ex_SHIFTER_ltemp1_22_, alu_ex_SHIFTER_ltemp1_21_,
         alu_ex_SHIFTER_ltemp1_20_, alu_ex_SHIFTER_ltemp1_19_,
         alu_ex_SHIFTER_ltemp1_18_, alu_ex_SHIFTER_ltemp1_17_,
         alu_ex_SHIFTER_ltemp1_16_, alu_ex_SHIFTER_ltemp1_15_,
         alu_ex_SHIFTER_ltemp1_14_, alu_ex_SHIFTER_ltemp1_13_,
         alu_ex_SHIFTER_ltemp1_12_, alu_ex_SHIFTER_ltemp1_11_,
         alu_ex_SHIFTER_ltemp1_10_, alu_ex_SHIFTER_ltemp1_9_,
         alu_ex_SHIFTER_ltemp1_8_, alu_ex_SHIFTER_ltemp1_7_,
         alu_ex_SHIFTER_ltemp1_6_, alu_ex_SHIFTER_ltemp1_5_,
         alu_ex_SHIFTER_ltemp1_4_, alu_ex_SHIFTER_ltemp1_3_,
         alu_ex_SHIFTER_ltemp1_2_, alu_ex_SHIFTER_ltemp1_1_,
         alu_ex_SHIFTER_ltemp1_0_, alu_ex_SHIFTER_ltemp0_31_,
         alu_ex_SHIFTER_ltemp0_30_, alu_ex_SHIFTER_ltemp0_29_,
         alu_ex_SHIFTER_ltemp0_28_, alu_ex_SHIFTER_ltemp0_27_,
         alu_ex_SHIFTER_ltemp0_26_, alu_ex_SHIFTER_ltemp0_25_,
         alu_ex_SHIFTER_ltemp0_24_, alu_ex_SHIFTER_ltemp0_23_,
         alu_ex_SHIFTER_ltemp0_22_, alu_ex_SHIFTER_ltemp0_21_,
         alu_ex_SHIFTER_ltemp0_20_, alu_ex_SHIFTER_ltemp0_19_,
         alu_ex_SHIFTER_ltemp0_18_, alu_ex_SHIFTER_ltemp0_17_,
         alu_ex_SHIFTER_ltemp0_16_, alu_ex_SHIFTER_ltemp0_15_,
         alu_ex_SHIFTER_ltemp0_14_, alu_ex_SHIFTER_ltemp0_13_,
         alu_ex_SHIFTER_ltemp0_12_, alu_ex_SHIFTER_ltemp0_11_,
         alu_ex_SHIFTER_ltemp0_10_, alu_ex_SHIFTER_ltemp0_9_,
         alu_ex_SHIFTER_ltemp0_8_, alu_ex_SHIFTER_ltemp0_7_,
         alu_ex_SHIFTER_ltemp0_6_, alu_ex_SHIFTER_ltemp0_5_,
         alu_ex_SHIFTER_ltemp0_4_, alu_ex_SHIFTER_ltemp0_3_,
         alu_ex_SHIFTER_ltemp0_2_, alu_ex_SHIFTER_ltemp0_1_,
         alu_ex_SHIFTER_ltemp0_0_, alu_ex_SHIFTER_SHIFTLEFT16_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_n3, alu_ex_SHIFTER_SHIFTLEFT16_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_16__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_17__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_18__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_19__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_20__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_21__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_22__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_23__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_24__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_25__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_26__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_27__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_28__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_29__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_30__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_31__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT8_n3, alu_ex_SHIFTER_SHIFTLEFT8_n2,
         alu_ex_SHIFTER_SHIFTLEFT8_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_24__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_25__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_26__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_27__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_28__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_29__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_30__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_31__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT4_n3, alu_ex_SHIFTER_SHIFTLEFT4_n2,
         alu_ex_SHIFTER_SHIFTLEFT4_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_28__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_29__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_30__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_31__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT2_n4, alu_ex_SHIFTER_SHIFTLEFT2_n3,
         alu_ex_SHIFTER_SHIFTLEFT2_n2, alu_ex_SHIFTER_SHIFTLEFT2_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_30__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_31__MUX_n2,
         alu_ex_SHIFTER_SHIFTLEFT1_n3, alu_ex_SHIFTER_SHIFTLEFT1_n2,
         alu_ex_SHIFTER_SHIFTLEFT1_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_31__MUX_n2,
         alu_ex_SHIFTER_SHIFTRIGHT16_n3, alu_ex_SHIFTER_SHIFTRIGHT16_n2,
         alu_ex_SHIFTER_SHIFTRIGHT16_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_31__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_n4, alu_ex_SHIFTER_SHIFTRIGHT8_n3,
         alu_ex_SHIFTER_SHIFTRIGHT8_n2, alu_ex_SHIFTER_SHIFTRIGHT8_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_31__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_n4, alu_ex_SHIFTER_SHIFTRIGHT4_n3,
         alu_ex_SHIFTER_SHIFTRIGHT4_n2, alu_ex_SHIFTER_SHIFTRIGHT4_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_31__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_n4, alu_ex_SHIFTER_SHIFTRIGHT2_n3,
         alu_ex_SHIFTER_SHIFTRIGHT2_n2, alu_ex_SHIFTER_SHIFTRIGHT2_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_31__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_n4, alu_ex_SHIFTER_SHIFTRIGHT1_n3,
         alu_ex_SHIFTER_SHIFTRIGHT1_n2, alu_ex_SHIFTER_SHIFTRIGHT1_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_31__MUX_n4,
         alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_n4, alu_ex_SHIFTER_LEFTORRIGHT_n3,
         alu_ex_SHIFTER_LEFTORRIGHT_n2, alu_ex_SHIFTER_LEFTORRIGHT_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_31__MUX_n4,
         alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_SET_FLAGS_n6, alu_ex_SET_FLAGS_n5, alu_ex_SET_FLAGS_n4,
         alu_ex_SET_FLAGS_n3, alu_ex_SET_FLAGS_n2, alu_ex_SET_FLAGS_n1,
         alu_ex_SET_FLAGS_n12, alu_ex_SET_FLAGS_sub_of,
         alu_ex_SET_FLAGS_difference_31_, alu_ex_SET_FLAGS_difference_30_,
         alu_ex_SET_FLAGS_difference_29_, alu_ex_SET_FLAGS_difference_28_,
         alu_ex_SET_FLAGS_difference_27_, alu_ex_SET_FLAGS_difference_26_,
         alu_ex_SET_FLAGS_difference_25_, alu_ex_SET_FLAGS_difference_24_,
         alu_ex_SET_FLAGS_difference_23_, alu_ex_SET_FLAGS_difference_22_,
         alu_ex_SET_FLAGS_difference_21_, alu_ex_SET_FLAGS_difference_20_,
         alu_ex_SET_FLAGS_difference_19_, alu_ex_SET_FLAGS_difference_18_,
         alu_ex_SET_FLAGS_difference_17_, alu_ex_SET_FLAGS_difference_16_,
         alu_ex_SET_FLAGS_difference_15_, alu_ex_SET_FLAGS_difference_14_,
         alu_ex_SET_FLAGS_difference_13_, alu_ex_SET_FLAGS_difference_12_,
         alu_ex_SET_FLAGS_difference_11_, alu_ex_SET_FLAGS_difference_10_,
         alu_ex_SET_FLAGS_difference_9_, alu_ex_SET_FLAGS_difference_8_,
         alu_ex_SET_FLAGS_difference_7_, alu_ex_SET_FLAGS_difference_6_,
         alu_ex_SET_FLAGS_difference_5_, alu_ex_SET_FLAGS_difference_4_,
         alu_ex_SET_FLAGS_difference_3_, alu_ex_SET_FLAGS_difference_2_,
         alu_ex_SET_FLAGS_difference_1_, alu_ex_SET_FLAGS_difference_0_,
         alu_ex_SET_FLAGS_FULL_ADDER_n7, alu_ex_SET_FLAGS_FULL_ADDER_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_n5, alu_ex_SET_FLAGS_FULL_ADDER_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_n1, alu_ex_SET_FLAGS_FULL_ADDER_carry_31_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_30_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_29_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_28_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_27_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_26_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_25_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_24_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_23_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_22_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_21_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_20_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_19_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_18_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_17_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_16_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_15_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_14_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_13_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_12_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_11_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_10_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_9_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_8_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_7_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_6_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_5_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_4_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_3_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_2_,
         alu_ex_SET_FLAGS_FULL_ADDER_carry_1_, alu_ex_SET_FLAGS_FULL_ADDER_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n15,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n14,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n13,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n12,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n10,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n8,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n7,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n8,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n7,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n9,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n8,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n7,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n10,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n9,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n8,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n9,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n8,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n7,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n10,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n9,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n8,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n7,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n4,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n1,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n14,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n13,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n12,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n10,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n9,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n8,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n7,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n6,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n3,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_31__FA_n5,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_31__FA_n2,
         alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_31__FA_n1,
         alu_ex_SET_FLAGS_CHECK_EQ_n19, alu_ex_SET_FLAGS_CHECK_EQ_n18,
         alu_ex_SET_FLAGS_CHECK_EQ_n17, alu_ex_SET_FLAGS_CHECK_EQ_n16,
         alu_ex_SET_FLAGS_CHECK_EQ_n15, alu_ex_SET_FLAGS_CHECK_EQ_n14,
         alu_ex_SET_FLAGS_CHECK_EQ_n13, alu_ex_SET_FLAGS_CHECK_EQ_n12,
         alu_ex_SET_FLAGS_CHECK_EQ_n11, alu_ex_SET_FLAGS_CHECK_EQ_n10,
         alu_ex_SET_FLAGS_CHECK_EQ_n9, alu_ex_SET_FLAGS_CHECK_EQ_n8,
         alu_ex_SET_FLAGS_CHECK_EQ_n7, alu_ex_SET_FLAGS_CHECK_EQ_n6,
         alu_ex_SET_FLAGS_CHECK_EQ_n5, alu_ex_SET_FLAGS_CHECK_EQ_n4,
         alu_ex_SET_FLAGS_CHECK_EQ_n3, alu_ex_SET_FLAGS_CHECK_EQ_n2,
         alu_ex_SET_FLAGS_CHECK_EQ_n1, alu_ex_EXTEND_SEQ_n1,
         alu_ex_EXTEND_SNE_n1, alu_ex_EXTEND_SLE_n1, alu_ex_EXTEND_SLT_n1,
         alu_ex_EXTEND_SGE_n1, alu_ex_EXTEND_SGT_n1, alu_ex_FINAL_MUX_n2,
         alu_ex_FINAL_MUX_n1, alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus2_31_,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_n3,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_n3,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n3,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n6,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n5,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n3,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n3,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus1_31_,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n3,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n3,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n3,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n3,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n3,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_0__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_1__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_2__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_3__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_4__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_5__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_6__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_7__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_8__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_9__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_10__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_11__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_12__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_13__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_14__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_15__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_16__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_17__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_18__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_19__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_20__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_21__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_22__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_23__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_24__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_25__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_26__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_27__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_28__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_29__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_30__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n3,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n3,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n3,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n6,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n5,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n3,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n3,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n2,
         alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n1,
         alu_ex_FINAL_MUX_MUX_OUT_n4, alu_ex_FINAL_MUX_MUX_OUT_n3,
         alu_ex_FINAL_MUX_MUX_OUT_n2, alu_ex_FINAL_MUX_MUX_OUT_n1,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_0__MUX_n2,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_0__MUX_n1,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_1__MUX_n3,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_1__MUX_n2,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_19__MUX_n4,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_19__MUX_n1,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_20__MUX_n4,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_20__MUX_n1,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_21__MUX_n4,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_21__MUX_n1,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_22__MUX_n4,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_22__MUX_n1,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_23__MUX_n4,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_23__MUX_n1,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_24__MUX_n4,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_24__MUX_n1,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_25__MUX_n4,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_25__MUX_n1,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_26__MUX_n4,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_26__MUX_n1,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_27__MUX_n4,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_27__MUX_n1,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_28__MUX_n4,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_28__MUX_n1,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_29__MUX_n4,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_29__MUX_n1,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_30__MUX_n4,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_30__MUX_n1,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_31__MUX_n3,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_31__MUX_n2,
         alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_31__MUX_n1,
         CHOOSE_FP_OR_NOTMUL_n3, CHOOSE_FP_OR_NOTMUL_n2,
         CHOOSE_FP_OR_NOTMUL_n1, CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_0__MUX_n3,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_0__MUX_n2,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_0__MUX_n1,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_19__MUX_n4,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_19__MUX_n1,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_20__MUX_n4,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_20__MUX_n1,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_21__MUX_n4,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_21__MUX_n1,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_22__MUX_n4,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_22__MUX_n1,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_23__MUX_n4,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_23__MUX_n1,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_24__MUX_n4,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_24__MUX_n1,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_25__MUX_n4,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_25__MUX_n1,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_26__MUX_n4,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_26__MUX_n1,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_27__MUX_n4,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_27__MUX_n1,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_28__MUX_n4,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_28__MUX_n1,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_29__MUX_n4,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_29__MUX_n1,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_30__MUX_n4,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_30__MUX_n1,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_31__MUX_n3,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_31__MUX_n2,
         CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_31__MUX_n1, mul_ex_n40, mul_ex_n39,
         mul_ex_n37, mul_ex_n32, mul_ex_n31, mul_ex_n30, mul_ex_n29,
         mul_ex_n28, mul_ex_n27, mul_ex_n26, mul_ex_n25, mul_ex_n24,
         mul_ex_n23, mul_ex_n22, mul_ex_n21, mul_ex_n20, mul_ex_n19,
         mul_ex_n18, mul_ex_n17, mul_ex_n16, mul_ex_n15, mul_ex_n14,
         mul_ex_n13, mul_ex_n12, mul_ex_n11, mul_ex_n10, mul_ex_n9, mul_ex_n8,
         mul_ex_n7, mul_ex_n6, mul_ex_n5, mul_ex_n4, mul_ex_n3, mul_ex_N186,
         mul_ex_N187, mul_ex_N188, mul_ex_N189, mul_ex_N190, mul_ex_N191,
         mul_ex_N192, mul_ex_N193, mul_ex_N194, mul_ex_N195, mul_ex_N196,
         mul_ex_N197, mul_ex_N198, mul_ex_N199, mul_ex_N200, mul_ex_N201,
         mul_ex_N202, mul_ex_N203, mul_ex_N204, mul_ex_N205, mul_ex_N206,
         mul_ex_N207, mul_ex_N208, mul_ex_N209, mul_ex_N210, mul_ex_N211,
         mul_ex_N212, mul_ex_N213, mul_ex_N214, mul_ex_N215, mul_ex_N216,
         mul_ex_N217, mul_ex_N250, mul_ex_N251, mul_ex_N252, mul_ex_N253,
         mul_ex_N254, mul_ex_N255, mul_ex_N256, mul_ex_N257, mul_ex_N258,
         mul_ex_N259, mul_ex_N260, mul_ex_N261, mul_ex_N262, mul_ex_N263,
         mul_ex_N264, mul_ex_N265, mul_ex_N266, mul_ex_N267, mul_ex_N268,
         mul_ex_N269, mul_ex_N270, mul_ex_N271, mul_ex_N272, mul_ex_N273,
         mul_ex_N274, mul_ex_N275, mul_ex_N276, mul_ex_N277, mul_ex_N278,
         mul_ex_N279, mul_ex_N280, mul_ex_N281, mul_ex_N282, mul_ex_N283,
         mul_ex_N284, mul_ex_N285, mul_ex_N286, mul_ex_N287, mul_ex_N288,
         mul_ex_N289, mul_ex_N290, mul_ex_N291, mul_ex_N292, mul_ex_N293,
         mul_ex_N294, mul_ex_N295, mul_ex_N296, mul_ex_N297, mul_ex_N298,
         mul_ex_n36, mul_ex_n35, mul_ex_n34, mul_ex_n33, mul_ex_N476,
         mul_ex_N475, mul_ex_N474, mul_ex_N473, mul_ex_N472, mul_ex_N471,
         mul_ex_N470, mul_ex_N469, mul_ex_N468, mul_ex_N467, mul_ex_N466,
         mul_ex_N465, mul_ex_N464, mul_ex_N463, mul_ex_N462, mul_ex_N461,
         mul_ex_N460, mul_ex_N459, mul_ex_N458, mul_ex_N457, mul_ex_N456,
         mul_ex_N455, mul_ex_N454, mul_ex_N453, mul_ex_N452, mul_ex_N451,
         mul_ex_N450, mul_ex_N449, mul_ex_N448, mul_ex_N447, mul_ex_N446,
         mul_ex_N445, mul_ex_N443, mul_ex_N442, mul_ex_N441, mul_ex_N440,
         mul_ex_N439, mul_ex_N438, mul_ex_N437, mul_ex_N436, mul_ex_N435,
         mul_ex_N434, mul_ex_N433, mul_ex_N432, mul_ex_N431, mul_ex_N430,
         mul_ex_N429, mul_ex_N428, mul_ex_N427, mul_ex_N426, mul_ex_N425,
         mul_ex_N424, mul_ex_N423, mul_ex_N422, mul_ex_N421, mul_ex_N420,
         mul_ex_N419, mul_ex_N418, mul_ex_N417, mul_ex_N416, mul_ex_N415,
         mul_ex_N414, mul_ex_N413, mul_ex_N412, mul_ex_N410, mul_ex_N409,
         mul_ex_N408, mul_ex_N407, mul_ex_N406, mul_ex_N405, mul_ex_N404,
         mul_ex_N403, mul_ex_N402, mul_ex_N401, mul_ex_N400, mul_ex_N399,
         mul_ex_N398, mul_ex_N397, mul_ex_N396, mul_ex_N395, mul_ex_N394,
         mul_ex_N393, mul_ex_N392, mul_ex_N391, mul_ex_N390, mul_ex_N389,
         mul_ex_N388, mul_ex_N387, mul_ex_N386, mul_ex_N385, mul_ex_N384,
         mul_ex_N383, mul_ex_N382, mul_ex_N381, mul_ex_N380, mul_ex_N379,
         mul_ex_N377, mul_ex_N376, mul_ex_N375, mul_ex_N374, mul_ex_N373,
         mul_ex_N372, mul_ex_N371, mul_ex_N370, mul_ex_N369, mul_ex_N368,
         mul_ex_N367, mul_ex_N366, mul_ex_N365, mul_ex_N364, mul_ex_N363,
         mul_ex_N362, mul_ex_N361, mul_ex_N360, mul_ex_N359, mul_ex_N358,
         mul_ex_N357, mul_ex_N356, mul_ex_N355, mul_ex_N354, mul_ex_N353,
         mul_ex_N352, mul_ex_N351, mul_ex_N350, mul_ex_N349, mul_ex_N348,
         mul_ex_N347, mul_ex_N346, mul_ex_N345, mul_ex_N344, mul_ex_N343,
         mul_ex_N342, mul_ex_N341, mul_ex_N340, mul_ex_N339, mul_ex_N338,
         mul_ex_N337, mul_ex_N336, mul_ex_N335, mul_ex_N334, mul_ex_N333,
         mul_ex_N332, mul_ex_N331, mul_ex_N330, mul_ex_N329, mul_ex_N328,
         mul_ex_N327, mul_ex_N326, mul_ex_N325, mul_ex_N324, mul_ex_N323,
         mul_ex_N322, mul_ex_N321, mul_ex_N320, mul_ex_N319, mul_ex_N318,
         mul_ex_N317, mul_ex_N316, mul_ex_N315, mul_ex_N314, mul_ex_N249,
         mul_ex_N248, mul_ex_N247, mul_ex_N246, mul_ex_N245, mul_ex_N244,
         mul_ex_N243, mul_ex_N242, mul_ex_N241, mul_ex_N240, mul_ex_N239,
         mul_ex_N238, mul_ex_N237, mul_ex_N236, mul_ex_N235, mul_ex_N234,
         mul_ex_N233, mul_ex_N232, mul_ex_N231, mul_ex_N230, mul_ex_N229,
         mul_ex_N228, mul_ex_N227, mul_ex_N226, mul_ex_N225, mul_ex_N224,
         mul_ex_N223, mul_ex_N222, mul_ex_N221, mul_ex_N220, mul_ex_N219,
         mul_ex_N218, mul_ex_N185, mul_ex_N184, mul_ex_N183, mul_ex_N182,
         mul_ex_N181, mul_ex_N180, mul_ex_N179, mul_ex_N178, mul_ex_N177,
         mul_ex_N176, mul_ex_N175, mul_ex_N174, mul_ex_N173, mul_ex_N172,
         mul_ex_N171, mul_ex_N170, mul_ex_N169, mul_ex_N168, mul_ex_N167,
         mul_ex_N166, mul_ex_N165, mul_ex_N164, mul_ex_N163, mul_ex_N162,
         mul_ex_N161, mul_ex_N160, mul_ex_N159, mul_ex_N158, mul_ex_N157,
         mul_ex_N156, mul_ex_N155, mul_ex_N154, mul_ex_N153, mul_ex_N152,
         mul_ex_N151, mul_ex_N150, mul_ex_N149, mul_ex_N148, mul_ex_N147,
         mul_ex_N146, mul_ex_N145, mul_ex_N144, mul_ex_N143, mul_ex_N142,
         mul_ex_N141, mul_ex_N140, mul_ex_N139, mul_ex_N138, mul_ex_N137,
         mul_ex_N136, mul_ex_N135, mul_ex_N134, mul_ex_N133, mul_ex_N132,
         mul_ex_N131, mul_ex_N130, mul_ex_N129, mul_ex_N128, mul_ex_N127,
         mul_ex_N126, mul_ex_N125, mul_ex_N124, mul_ex_N123, mul_ex_N122,
         mul_ex_N121, mul_ex_N120, mul_ex_N119, mul_ex_N118, mul_ex_N117,
         mul_ex_N116, mul_ex_N115, mul_ex_N114, mul_ex_N113, mul_ex_N112,
         mul_ex_N111, mul_ex_N110, mul_ex_N109, mul_ex_N108, mul_ex_N107,
         mul_ex_N106, mul_ex_N105, mul_ex_N104, mul_ex_N103, mul_ex_N102,
         mul_ex_N101, mul_ex_N100, mul_ex_N99, mul_ex_N98, mul_ex_N97,
         mul_ex_N96, mul_ex_N95, mul_ex_N94, mul_ex_N93, mul_ex_N92,
         mul_ex_N91, mul_ex_N90, mul_ex_N89, mul_ex_N88, mul_ex_N87,
         mul_ex_N86, mul_ex_N85, mul_ex_N84, mul_ex_N83, mul_ex_N82,
         mul_ex_N81, mul_ex_N80, mul_ex_N79, mul_ex_N78, mul_ex_N77,
         mul_ex_N76, mul_ex_N75, mul_ex_N74, mul_ex_N73, mul_ex_N72,
         mul_ex_N71, mul_ex_N70, mul_ex_N69, mul_ex_N68, mul_ex_N67,
         mul_ex_N66, mul_ex_N65, mul_ex_N64, mul_ex_N63, mul_ex_N62,
         mul_ex_N61, mul_ex_N60, mul_ex_N59, mul_ex_N58, mul_ex_N57,
         mul_ex_N56, mul_ex_N43, mul_ex_Z_31_, mul_ex_Z_30_, mul_ex_Z_29_,
         mul_ex_Z_28_, mul_ex_Z_27_, mul_ex_Z_26_, mul_ex_Z_25_, mul_ex_Z_24_,
         mul_ex_Z_23_, mul_ex_Z_22_, mul_ex_Z_21_, mul_ex_Z_20_, mul_ex_Z_19_,
         mul_ex_Z_18_, mul_ex_Z_17_, mul_ex_Z_16_, mul_ex_Z_15_, mul_ex_Z_14_,
         mul_ex_Z_13_, mul_ex_Z_12_, mul_ex_Z_11_, mul_ex_Z_10_, mul_ex_Z_9_,
         mul_ex_Z_8_, mul_ex_Z_7_, mul_ex_Z_6_, mul_ex_Z_5_, mul_ex_Z_4_,
         mul_ex_Z_3_, mul_ex_Z_2_, mul_ex_Z_1_, mul_ex_Z_0_, mul_ex_L_31_,
         mul_ex_L_30_, mul_ex_L_29_, mul_ex_L_28_, mul_ex_L_27_, mul_ex_L_26_,
         mul_ex_L_25_, mul_ex_L_24_, mul_ex_L_23_, mul_ex_L_22_, mul_ex_L_21_,
         mul_ex_L_20_, mul_ex_L_19_, mul_ex_L_18_, mul_ex_L_17_, mul_ex_L_16_,
         mul_ex_L_15_, mul_ex_L_14_, mul_ex_L_13_, mul_ex_L_12_, mul_ex_L_11_,
         mul_ex_L_10_, mul_ex_L_9_, mul_ex_L_8_, mul_ex_L_7_, mul_ex_L_6_,
         mul_ex_L_5_, mul_ex_L_4_, mul_ex_L_3_, mul_ex_L_2_, mul_ex_L_1_,
         mul_ex_L_0_, mul_ex_N16, mul_ex_N15, mul_ex_N14,
         mul_ex_CurrentState_2_, mul_ex_CurrentState_1_,
         mul_ex_CurrentState_0_, mul_ex_add_85_n2, mul_ex_add_77_n2,
         mul_ex_add_1_root_add_0_root_add_98_2_n33,
         mul_ex_add_1_root_add_0_root_add_98_2_n17,
         mul_ex_add_1_root_add_0_root_add_98_2_n16,
         mul_ex_add_1_root_add_0_root_add_98_2_n15,
         mul_ex_add_1_root_add_0_root_add_98_2_n14,
         mul_ex_add_1_root_add_0_root_add_98_2_n13,
         mul_ex_add_1_root_add_0_root_add_98_2_n12,
         mul_ex_add_1_root_add_0_root_add_98_2_n11,
         mul_ex_add_1_root_add_0_root_add_98_2_n10,
         mul_ex_add_1_root_add_0_root_add_98_2_n8,
         mul_ex_add_1_root_add_0_root_add_98_2_n7,
         mul_ex_add_1_root_add_0_root_add_98_2_n6,
         mul_ex_add_1_root_add_0_root_add_98_2_n5,
         mul_ex_add_1_root_add_0_root_add_98_2_n4,
         mul_ex_add_1_root_add_0_root_add_98_2_n3,
         mul_ex_add_1_root_add_0_root_add_98_2_n2,
         mul_ex_add_1_root_add_0_root_add_98_2_carry_18_,
         mul_ex_add_1_root_add_0_root_add_98_2_carry_19_,
         mul_ex_add_1_root_add_0_root_add_98_2_carry_20_,
         mul_ex_add_1_root_add_0_root_add_98_2_carry_21_,
         mul_ex_add_1_root_add_0_root_add_98_2_carry_22_,
         mul_ex_add_1_root_add_0_root_add_98_2_carry_23_,
         mul_ex_add_1_root_add_0_root_add_98_2_carry_24_,
         mul_ex_add_1_root_add_0_root_add_98_2_carry_25_,
         mul_ex_add_1_root_add_0_root_add_98_2_carry_26_,
         mul_ex_add_1_root_add_0_root_add_98_2_carry_27_,
         mul_ex_add_1_root_add_0_root_add_98_2_carry_28_,
         mul_ex_add_1_root_add_0_root_add_98_2_carry_29_,
         mul_ex_add_1_root_add_0_root_add_98_2_carry_30_,
         mul_ex_add_1_root_add_0_root_add_98_2_carry_31_,
         mul_ex_add_1_root_add_0_root_add_98_2_carry_32_,
         mul_ex_add_0_root_add_0_root_add_98_2_n15,
         mul_ex_add_0_root_add_0_root_add_98_2_n14,
         mul_ex_add_0_root_add_0_root_add_98_2_n13,
         mul_ex_add_0_root_add_0_root_add_98_2_n12,
         mul_ex_add_0_root_add_0_root_add_98_2_n11,
         mul_ex_add_0_root_add_0_root_add_98_2_n10,
         mul_ex_add_0_root_add_0_root_add_98_2_n9,
         mul_ex_add_0_root_add_0_root_add_98_2_n8,
         mul_ex_add_0_root_add_0_root_add_98_2_n7,
         mul_ex_add_0_root_add_0_root_add_98_2_n6,
         mul_ex_add_0_root_add_0_root_add_98_2_n5,
         mul_ex_add_0_root_add_0_root_add_98_2_n4,
         mul_ex_add_0_root_add_0_root_add_98_2_n3,
         mul_ex_add_0_root_add_0_root_add_98_2_n2,
         mul_ex_add_0_root_add_0_root_add_98_2_n1,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_34_,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_35_,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_36_,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_37_,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_38_,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_39_,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_40_,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_41_,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_42_,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_43_,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_44_,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_45_,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_46_,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_47_,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_48_,
         mul_ex_add_0_root_add_0_root_add_98_2_carry_49_,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n33,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n32,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n31,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n30,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n29,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n28,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n27,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n26,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n25,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n24,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n23,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n22,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n21,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n20,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n19,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n18,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n17,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n16,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n15,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n14,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n13,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n12,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n11,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n10,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n9,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n8,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n7,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n6,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n5,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n4,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n3,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n2,
         mul_ex_sub_1_root_sub_0_root_sub_94_2_n1,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n33,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n32,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n31,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n30,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n29,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n28,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n27,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n26,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n25,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n24,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n23,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n22,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n21,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n20,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n19,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n18,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n17,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n16,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n15,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n14,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n13,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n12,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n11,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n10,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n9,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n8,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n7,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n6,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n5,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n4,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n3,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n2,
         mul_ex_sub_0_root_sub_0_root_sub_94_2_n1, mul_ex_mult_90_n299,
         mul_ex_mult_90_n298, mul_ex_mult_90_n297, mul_ex_mult_90_n296,
         mul_ex_mult_90_n295, mul_ex_mult_90_n294, mul_ex_mult_90_n293,
         mul_ex_mult_90_n292, mul_ex_mult_90_n291, mul_ex_mult_90_n290,
         mul_ex_mult_90_n289, mul_ex_mult_90_n288, mul_ex_mult_90_n287,
         mul_ex_mult_90_n286, mul_ex_mult_90_n285, mul_ex_mult_90_n284,
         mul_ex_mult_90_n283, mul_ex_mult_90_n282, mul_ex_mult_90_n281,
         mul_ex_mult_90_n280, mul_ex_mult_90_n279, mul_ex_mult_90_n278,
         mul_ex_mult_90_n277, mul_ex_mult_90_n276, mul_ex_mult_90_n275,
         mul_ex_mult_90_n274, mul_ex_mult_90_n273, mul_ex_mult_90_n272,
         mul_ex_mult_90_n271, mul_ex_mult_90_n270, mul_ex_mult_90_n269,
         mul_ex_mult_90_n268, mul_ex_mult_90_n267, mul_ex_mult_90_n266,
         mul_ex_mult_90_n265, mul_ex_mult_90_n264, mul_ex_mult_90_n263,
         mul_ex_mult_90_n262, mul_ex_mult_90_n261, mul_ex_mult_90_n260,
         mul_ex_mult_90_n259, mul_ex_mult_90_n258, mul_ex_mult_90_n257,
         mul_ex_mult_90_n256, mul_ex_mult_90_n255, mul_ex_mult_90_n254,
         mul_ex_mult_90_n253, mul_ex_mult_90_n252, mul_ex_mult_90_n251,
         mul_ex_mult_90_n250, mul_ex_mult_90_n249, mul_ex_mult_90_n248,
         mul_ex_mult_90_n247, mul_ex_mult_90_n246, mul_ex_mult_90_n245,
         mul_ex_mult_90_n244, mul_ex_mult_90_n243, mul_ex_mult_90_n242,
         mul_ex_mult_90_n241, mul_ex_mult_90_n240, mul_ex_mult_90_n239,
         mul_ex_mult_90_n238, mul_ex_mult_90_n237, mul_ex_mult_90_n236,
         mul_ex_mult_90_n235, mul_ex_mult_90_n234, mul_ex_mult_90_n233,
         mul_ex_mult_90_n232, mul_ex_mult_90_n231, mul_ex_mult_90_n230,
         mul_ex_mult_90_n229, mul_ex_mult_90_n228, mul_ex_mult_90_n227,
         mul_ex_mult_90_n226, mul_ex_mult_90_n225, mul_ex_mult_90_n224,
         mul_ex_mult_90_n223, mul_ex_mult_90_n222, mul_ex_mult_90_n221,
         mul_ex_mult_90_n220, mul_ex_mult_90_n219, mul_ex_mult_90_n218,
         mul_ex_mult_90_n217, mul_ex_mult_90_n216, mul_ex_mult_90_n215,
         mul_ex_mult_90_n214, mul_ex_mult_90_n213, mul_ex_mult_90_n212,
         mul_ex_mult_90_n211, mul_ex_mult_90_n210, mul_ex_mult_90_n209,
         mul_ex_mult_90_n208, mul_ex_mult_90_n207, mul_ex_mult_90_n206,
         mul_ex_mult_90_n205, mul_ex_mult_90_n204, mul_ex_mult_90_n203,
         mul_ex_mult_90_n202, mul_ex_mult_90_n201, mul_ex_mult_90_n200,
         mul_ex_mult_90_n199, mul_ex_mult_90_n198, mul_ex_mult_90_n197,
         mul_ex_mult_90_n196, mul_ex_mult_90_n195, mul_ex_mult_90_n194,
         mul_ex_mult_90_n193, mul_ex_mult_90_n192, mul_ex_mult_90_n191,
         mul_ex_mult_90_n190, mul_ex_mult_90_n189, mul_ex_mult_90_n188,
         mul_ex_mult_90_n187, mul_ex_mult_90_n186, mul_ex_mult_90_n185,
         mul_ex_mult_90_n184, mul_ex_mult_90_n183, mul_ex_mult_90_n182,
         mul_ex_mult_90_n181, mul_ex_mult_90_n180, mul_ex_mult_90_n179,
         mul_ex_mult_90_n178, mul_ex_mult_90_n177, mul_ex_mult_90_n176,
         mul_ex_mult_90_n175, mul_ex_mult_90_n174, mul_ex_mult_90_n173,
         mul_ex_mult_90_n172, mul_ex_mult_90_n171, mul_ex_mult_90_n170,
         mul_ex_mult_90_n169, mul_ex_mult_90_n168, mul_ex_mult_90_n167,
         mul_ex_mult_90_n166, mul_ex_mult_90_n165, mul_ex_mult_90_n164,
         mul_ex_mult_90_n163, mul_ex_mult_90_n162, mul_ex_mult_90_n161,
         mul_ex_mult_90_n160, mul_ex_mult_90_n159, mul_ex_mult_90_n158,
         mul_ex_mult_90_n157, mul_ex_mult_90_n156, mul_ex_mult_90_n155,
         mul_ex_mult_90_n154, mul_ex_mult_90_n153, mul_ex_mult_90_n152,
         mul_ex_mult_90_n151, mul_ex_mult_90_n150, mul_ex_mult_90_n149,
         mul_ex_mult_90_n148, mul_ex_mult_90_n147, mul_ex_mult_90_n146,
         mul_ex_mult_90_n145, mul_ex_mult_90_n144, mul_ex_mult_90_n143,
         mul_ex_mult_90_n142, mul_ex_mult_90_n141, mul_ex_mult_90_n140,
         mul_ex_mult_90_n139, mul_ex_mult_90_n138, mul_ex_mult_90_n137,
         mul_ex_mult_90_n136, mul_ex_mult_90_n135, mul_ex_mult_90_n134,
         mul_ex_mult_90_n133, mul_ex_mult_90_n132, mul_ex_mult_90_n131,
         mul_ex_mult_90_n130, mul_ex_mult_90_n129, mul_ex_mult_90_n128,
         mul_ex_mult_90_n127, mul_ex_mult_90_n126, mul_ex_mult_90_n125,
         mul_ex_mult_90_n124, mul_ex_mult_90_n123, mul_ex_mult_90_n122,
         mul_ex_mult_90_n121, mul_ex_mult_90_n120, mul_ex_mult_90_n119,
         mul_ex_mult_90_n118, mul_ex_mult_90_n117, mul_ex_mult_90_n116,
         mul_ex_mult_90_n115, mul_ex_mult_90_n114, mul_ex_mult_90_n113,
         mul_ex_mult_90_n112, mul_ex_mult_90_n111, mul_ex_mult_90_n110,
         mul_ex_mult_90_n109, mul_ex_mult_90_n108, mul_ex_mult_90_n107,
         mul_ex_mult_90_n106, mul_ex_mult_90_n105, mul_ex_mult_90_n104,
         mul_ex_mult_90_n103, mul_ex_mult_90_n102, mul_ex_mult_90_n101,
         mul_ex_mult_90_n100, mul_ex_mult_90_n99, mul_ex_mult_90_n98,
         mul_ex_mult_90_n97, mul_ex_mult_90_n96, mul_ex_mult_90_n95,
         mul_ex_mult_90_n94, mul_ex_mult_90_n93, mul_ex_mult_90_n92,
         mul_ex_mult_90_n91, mul_ex_mult_90_n90, mul_ex_mult_90_n89,
         mul_ex_mult_90_n88, mul_ex_mult_90_n87, mul_ex_mult_90_n86,
         mul_ex_mult_90_n85, mul_ex_mult_90_n84, mul_ex_mult_90_n83,
         mul_ex_mult_90_n82, mul_ex_mult_90_n81, mul_ex_mult_90_n80,
         mul_ex_mult_90_n79, mul_ex_mult_90_n78, mul_ex_mult_90_n77,
         mul_ex_mult_90_n76, mul_ex_mult_90_n75, mul_ex_mult_90_n74,
         mul_ex_mult_90_n73, mul_ex_mult_90_n72, mul_ex_mult_90_n71,
         mul_ex_mult_90_n70, mul_ex_mult_90_n69, mul_ex_mult_90_n68,
         mul_ex_mult_90_n67, mul_ex_mult_90_n66, mul_ex_mult_90_n65,
         mul_ex_mult_90_n64, mul_ex_mult_90_n63, mul_ex_mult_90_n62,
         mul_ex_mult_90_n61, mul_ex_mult_90_n60, mul_ex_mult_90_n59,
         mul_ex_mult_90_n58, mul_ex_mult_90_n57, mul_ex_mult_90_n56,
         mul_ex_mult_90_n55, mul_ex_mult_90_n54, mul_ex_mult_90_n53,
         mul_ex_mult_90_n52, mul_ex_mult_90_n51, mul_ex_mult_90_n50,
         mul_ex_mult_90_n48, mul_ex_mult_90_n47, mul_ex_mult_90_n46,
         mul_ex_mult_90_n45, mul_ex_mult_90_n44, mul_ex_mult_90_n43,
         mul_ex_mult_90_n42, mul_ex_mult_90_n41, mul_ex_mult_90_n40,
         mul_ex_mult_90_n39, mul_ex_mult_90_n38, mul_ex_mult_90_n37,
         mul_ex_mult_90_n36, mul_ex_mult_90_n35, mul_ex_mult_90_n34,
         mul_ex_mult_90_n33, mul_ex_mult_90_n32, mul_ex_mult_90_n31,
         mul_ex_mult_90_n30, mul_ex_mult_90_n29, mul_ex_mult_90_n28,
         mul_ex_mult_90_n27, mul_ex_mult_90_n26, mul_ex_mult_90_n25,
         mul_ex_mult_90_n24, mul_ex_mult_90_n23, mul_ex_mult_90_n22,
         mul_ex_mult_90_n21, mul_ex_mult_90_n20, mul_ex_mult_90_n19,
         mul_ex_mult_90_n18, mul_ex_mult_90_n17, mul_ex_mult_90_n16,
         mul_ex_mult_90_n15, mul_ex_mult_90_n14, mul_ex_mult_90_n13,
         mul_ex_mult_90_n12, mul_ex_mult_90_n11, mul_ex_mult_90_n10,
         mul_ex_mult_90_n9, mul_ex_mult_90_n8, mul_ex_mult_90_n7,
         mul_ex_mult_90_n6, mul_ex_mult_90_n5, mul_ex_mult_90_n4,
         mul_ex_mult_90_n3, mul_ex_mult_90_SUMB_16__1_,
         mul_ex_mult_90_SUMB_16__2_, mul_ex_mult_90_SUMB_16__3_,
         mul_ex_mult_90_SUMB_16__4_, mul_ex_mult_90_SUMB_16__5_,
         mul_ex_mult_90_SUMB_16__6_, mul_ex_mult_90_SUMB_16__7_,
         mul_ex_mult_90_SUMB_16__8_, mul_ex_mult_90_SUMB_16__9_,
         mul_ex_mult_90_SUMB_16__10_, mul_ex_mult_90_SUMB_16__11_,
         mul_ex_mult_90_SUMB_16__12_, mul_ex_mult_90_SUMB_16__13_,
         mul_ex_mult_90_SUMB_16__14_, mul_ex_mult_90_SUMB_16__15_,
         mul_ex_mult_90_SUMB_17__1_, mul_ex_mult_90_SUMB_17__2_,
         mul_ex_mult_90_SUMB_17__3_, mul_ex_mult_90_SUMB_17__4_,
         mul_ex_mult_90_SUMB_17__5_, mul_ex_mult_90_SUMB_17__6_,
         mul_ex_mult_90_SUMB_17__7_, mul_ex_mult_90_SUMB_17__8_,
         mul_ex_mult_90_SUMB_17__9_, mul_ex_mult_90_SUMB_17__10_,
         mul_ex_mult_90_SUMB_17__11_, mul_ex_mult_90_SUMB_17__12_,
         mul_ex_mult_90_SUMB_17__13_, mul_ex_mult_90_SUMB_17__14_,
         mul_ex_mult_90_SUMB_18__1_, mul_ex_mult_90_SUMB_18__2_,
         mul_ex_mult_90_SUMB_18__3_, mul_ex_mult_90_SUMB_18__4_,
         mul_ex_mult_90_SUMB_18__5_, mul_ex_mult_90_SUMB_18__6_,
         mul_ex_mult_90_SUMB_18__7_, mul_ex_mult_90_SUMB_18__8_,
         mul_ex_mult_90_SUMB_18__9_, mul_ex_mult_90_SUMB_18__10_,
         mul_ex_mult_90_SUMB_18__11_, mul_ex_mult_90_SUMB_18__12_,
         mul_ex_mult_90_SUMB_18__13_, mul_ex_mult_90_SUMB_19__1_,
         mul_ex_mult_90_SUMB_19__2_, mul_ex_mult_90_SUMB_19__3_,
         mul_ex_mult_90_SUMB_19__4_, mul_ex_mult_90_SUMB_19__5_,
         mul_ex_mult_90_SUMB_19__6_, mul_ex_mult_90_SUMB_19__7_,
         mul_ex_mult_90_SUMB_19__8_, mul_ex_mult_90_SUMB_19__9_,
         mul_ex_mult_90_SUMB_19__10_, mul_ex_mult_90_SUMB_19__11_,
         mul_ex_mult_90_SUMB_19__12_, mul_ex_mult_90_SUMB_20__1_,
         mul_ex_mult_90_SUMB_20__2_, mul_ex_mult_90_SUMB_20__3_,
         mul_ex_mult_90_SUMB_20__4_, mul_ex_mult_90_SUMB_20__5_,
         mul_ex_mult_90_SUMB_20__6_, mul_ex_mult_90_SUMB_20__7_,
         mul_ex_mult_90_SUMB_20__8_, mul_ex_mult_90_SUMB_20__9_,
         mul_ex_mult_90_SUMB_20__10_, mul_ex_mult_90_SUMB_20__11_,
         mul_ex_mult_90_SUMB_21__1_, mul_ex_mult_90_SUMB_21__2_,
         mul_ex_mult_90_SUMB_21__3_, mul_ex_mult_90_SUMB_21__4_,
         mul_ex_mult_90_SUMB_21__5_, mul_ex_mult_90_SUMB_21__6_,
         mul_ex_mult_90_SUMB_21__7_, mul_ex_mult_90_SUMB_21__8_,
         mul_ex_mult_90_SUMB_21__9_, mul_ex_mult_90_SUMB_21__10_,
         mul_ex_mult_90_SUMB_22__1_, mul_ex_mult_90_SUMB_22__2_,
         mul_ex_mult_90_SUMB_22__3_, mul_ex_mult_90_SUMB_22__4_,
         mul_ex_mult_90_SUMB_22__5_, mul_ex_mult_90_SUMB_22__6_,
         mul_ex_mult_90_SUMB_22__7_, mul_ex_mult_90_SUMB_22__8_,
         mul_ex_mult_90_SUMB_22__9_, mul_ex_mult_90_SUMB_23__1_,
         mul_ex_mult_90_SUMB_23__2_, mul_ex_mult_90_SUMB_23__3_,
         mul_ex_mult_90_SUMB_23__4_, mul_ex_mult_90_SUMB_23__5_,
         mul_ex_mult_90_SUMB_23__6_, mul_ex_mult_90_SUMB_23__7_,
         mul_ex_mult_90_SUMB_23__8_, mul_ex_mult_90_SUMB_24__1_,
         mul_ex_mult_90_SUMB_24__2_, mul_ex_mult_90_SUMB_24__3_,
         mul_ex_mult_90_SUMB_24__4_, mul_ex_mult_90_SUMB_24__5_,
         mul_ex_mult_90_SUMB_24__6_, mul_ex_mult_90_SUMB_24__7_,
         mul_ex_mult_90_SUMB_25__1_, mul_ex_mult_90_SUMB_25__2_,
         mul_ex_mult_90_SUMB_25__3_, mul_ex_mult_90_SUMB_25__4_,
         mul_ex_mult_90_SUMB_25__5_, mul_ex_mult_90_SUMB_25__6_,
         mul_ex_mult_90_SUMB_26__1_, mul_ex_mult_90_SUMB_26__2_,
         mul_ex_mult_90_SUMB_26__3_, mul_ex_mult_90_SUMB_26__4_,
         mul_ex_mult_90_SUMB_26__5_, mul_ex_mult_90_SUMB_27__1_,
         mul_ex_mult_90_SUMB_27__2_, mul_ex_mult_90_SUMB_27__3_,
         mul_ex_mult_90_SUMB_27__4_, mul_ex_mult_90_SUMB_28__1_,
         mul_ex_mult_90_SUMB_28__2_, mul_ex_mult_90_SUMB_28__3_,
         mul_ex_mult_90_SUMB_29__1_, mul_ex_mult_90_SUMB_29__2_,
         mul_ex_mult_90_SUMB_30__1_, mul_ex_mult_90_CARRYB_16__0_,
         mul_ex_mult_90_CARRYB_16__1_, mul_ex_mult_90_CARRYB_16__2_,
         mul_ex_mult_90_CARRYB_16__3_, mul_ex_mult_90_CARRYB_16__4_,
         mul_ex_mult_90_CARRYB_16__5_, mul_ex_mult_90_CARRYB_16__6_,
         mul_ex_mult_90_CARRYB_16__7_, mul_ex_mult_90_CARRYB_16__8_,
         mul_ex_mult_90_CARRYB_16__9_, mul_ex_mult_90_CARRYB_16__10_,
         mul_ex_mult_90_CARRYB_16__11_, mul_ex_mult_90_CARRYB_16__12_,
         mul_ex_mult_90_CARRYB_16__13_, mul_ex_mult_90_CARRYB_16__14_,
         mul_ex_mult_90_CARRYB_17__0_, mul_ex_mult_90_CARRYB_17__1_,
         mul_ex_mult_90_CARRYB_17__2_, mul_ex_mult_90_CARRYB_17__3_,
         mul_ex_mult_90_CARRYB_17__4_, mul_ex_mult_90_CARRYB_17__5_,
         mul_ex_mult_90_CARRYB_17__6_, mul_ex_mult_90_CARRYB_17__7_,
         mul_ex_mult_90_CARRYB_17__8_, mul_ex_mult_90_CARRYB_17__9_,
         mul_ex_mult_90_CARRYB_17__10_, mul_ex_mult_90_CARRYB_17__11_,
         mul_ex_mult_90_CARRYB_17__12_, mul_ex_mult_90_CARRYB_17__13_,
         mul_ex_mult_90_CARRYB_18__0_, mul_ex_mult_90_CARRYB_18__1_,
         mul_ex_mult_90_CARRYB_18__2_, mul_ex_mult_90_CARRYB_18__3_,
         mul_ex_mult_90_CARRYB_18__4_, mul_ex_mult_90_CARRYB_18__5_,
         mul_ex_mult_90_CARRYB_18__6_, mul_ex_mult_90_CARRYB_18__7_,
         mul_ex_mult_90_CARRYB_18__8_, mul_ex_mult_90_CARRYB_18__9_,
         mul_ex_mult_90_CARRYB_18__10_, mul_ex_mult_90_CARRYB_18__11_,
         mul_ex_mult_90_CARRYB_18__12_, mul_ex_mult_90_CARRYB_19__0_,
         mul_ex_mult_90_CARRYB_19__1_, mul_ex_mult_90_CARRYB_19__2_,
         mul_ex_mult_90_CARRYB_19__3_, mul_ex_mult_90_CARRYB_19__4_,
         mul_ex_mult_90_CARRYB_19__5_, mul_ex_mult_90_CARRYB_19__6_,
         mul_ex_mult_90_CARRYB_19__7_, mul_ex_mult_90_CARRYB_19__8_,
         mul_ex_mult_90_CARRYB_19__9_, mul_ex_mult_90_CARRYB_19__10_,
         mul_ex_mult_90_CARRYB_19__11_, mul_ex_mult_90_CARRYB_20__0_,
         mul_ex_mult_90_CARRYB_20__1_, mul_ex_mult_90_CARRYB_20__2_,
         mul_ex_mult_90_CARRYB_20__3_, mul_ex_mult_90_CARRYB_20__4_,
         mul_ex_mult_90_CARRYB_20__5_, mul_ex_mult_90_CARRYB_20__6_,
         mul_ex_mult_90_CARRYB_20__7_, mul_ex_mult_90_CARRYB_20__8_,
         mul_ex_mult_90_CARRYB_20__9_, mul_ex_mult_90_CARRYB_20__10_,
         mul_ex_mult_90_CARRYB_21__0_, mul_ex_mult_90_CARRYB_21__1_,
         mul_ex_mult_90_CARRYB_21__2_, mul_ex_mult_90_CARRYB_21__3_,
         mul_ex_mult_90_CARRYB_21__4_, mul_ex_mult_90_CARRYB_21__5_,
         mul_ex_mult_90_CARRYB_21__6_, mul_ex_mult_90_CARRYB_21__7_,
         mul_ex_mult_90_CARRYB_21__8_, mul_ex_mult_90_CARRYB_21__9_,
         mul_ex_mult_90_CARRYB_22__0_, mul_ex_mult_90_CARRYB_22__1_,
         mul_ex_mult_90_CARRYB_22__2_, mul_ex_mult_90_CARRYB_22__3_,
         mul_ex_mult_90_CARRYB_22__4_, mul_ex_mult_90_CARRYB_22__5_,
         mul_ex_mult_90_CARRYB_22__6_, mul_ex_mult_90_CARRYB_22__7_,
         mul_ex_mult_90_CARRYB_22__8_, mul_ex_mult_90_CARRYB_23__0_,
         mul_ex_mult_90_CARRYB_23__1_, mul_ex_mult_90_CARRYB_23__2_,
         mul_ex_mult_90_CARRYB_23__3_, mul_ex_mult_90_CARRYB_23__4_,
         mul_ex_mult_90_CARRYB_23__5_, mul_ex_mult_90_CARRYB_23__6_,
         mul_ex_mult_90_CARRYB_23__7_, mul_ex_mult_90_CARRYB_24__0_,
         mul_ex_mult_90_CARRYB_24__1_, mul_ex_mult_90_CARRYB_24__2_,
         mul_ex_mult_90_CARRYB_24__3_, mul_ex_mult_90_CARRYB_24__4_,
         mul_ex_mult_90_CARRYB_24__5_, mul_ex_mult_90_CARRYB_24__6_,
         mul_ex_mult_90_CARRYB_25__0_, mul_ex_mult_90_CARRYB_25__1_,
         mul_ex_mult_90_CARRYB_25__2_, mul_ex_mult_90_CARRYB_25__3_,
         mul_ex_mult_90_CARRYB_25__4_, mul_ex_mult_90_CARRYB_25__5_,
         mul_ex_mult_90_CARRYB_26__0_, mul_ex_mult_90_CARRYB_26__1_,
         mul_ex_mult_90_CARRYB_26__2_, mul_ex_mult_90_CARRYB_26__3_,
         mul_ex_mult_90_CARRYB_26__4_, mul_ex_mult_90_CARRYB_27__0_,
         mul_ex_mult_90_CARRYB_27__1_, mul_ex_mult_90_CARRYB_27__2_,
         mul_ex_mult_90_CARRYB_27__3_, mul_ex_mult_90_CARRYB_28__0_,
         mul_ex_mult_90_CARRYB_28__1_, mul_ex_mult_90_CARRYB_28__2_,
         mul_ex_mult_90_CARRYB_29__0_, mul_ex_mult_90_CARRYB_29__1_,
         mul_ex_mult_90_CARRYB_30__0_, mul_ex_mult_90_SUMB_2__1_,
         mul_ex_mult_90_SUMB_2__2_, mul_ex_mult_90_SUMB_2__3_,
         mul_ex_mult_90_SUMB_2__4_, mul_ex_mult_90_SUMB_2__5_,
         mul_ex_mult_90_SUMB_2__6_, mul_ex_mult_90_SUMB_2__7_,
         mul_ex_mult_90_SUMB_2__8_, mul_ex_mult_90_SUMB_2__9_,
         mul_ex_mult_90_SUMB_2__10_, mul_ex_mult_90_SUMB_2__11_,
         mul_ex_mult_90_SUMB_2__12_, mul_ex_mult_90_SUMB_2__13_,
         mul_ex_mult_90_SUMB_2__14_, mul_ex_mult_90_SUMB_2__15_,
         mul_ex_mult_90_SUMB_2__16_, mul_ex_mult_90_SUMB_3__1_,
         mul_ex_mult_90_SUMB_3__2_, mul_ex_mult_90_SUMB_3__3_,
         mul_ex_mult_90_SUMB_3__4_, mul_ex_mult_90_SUMB_3__5_,
         mul_ex_mult_90_SUMB_3__6_, mul_ex_mult_90_SUMB_3__7_,
         mul_ex_mult_90_SUMB_3__8_, mul_ex_mult_90_SUMB_3__9_,
         mul_ex_mult_90_SUMB_3__10_, mul_ex_mult_90_SUMB_3__11_,
         mul_ex_mult_90_SUMB_3__12_, mul_ex_mult_90_SUMB_3__13_,
         mul_ex_mult_90_SUMB_3__14_, mul_ex_mult_90_SUMB_3__15_,
         mul_ex_mult_90_SUMB_3__16_, mul_ex_mult_90_SUMB_4__1_,
         mul_ex_mult_90_SUMB_4__2_, mul_ex_mult_90_SUMB_4__3_,
         mul_ex_mult_90_SUMB_4__4_, mul_ex_mult_90_SUMB_4__5_,
         mul_ex_mult_90_SUMB_4__6_, mul_ex_mult_90_SUMB_4__7_,
         mul_ex_mult_90_SUMB_4__8_, mul_ex_mult_90_SUMB_4__9_,
         mul_ex_mult_90_SUMB_4__10_, mul_ex_mult_90_SUMB_4__11_,
         mul_ex_mult_90_SUMB_4__12_, mul_ex_mult_90_SUMB_4__13_,
         mul_ex_mult_90_SUMB_4__14_, mul_ex_mult_90_SUMB_4__15_,
         mul_ex_mult_90_SUMB_4__16_, mul_ex_mult_90_SUMB_5__1_,
         mul_ex_mult_90_SUMB_5__2_, mul_ex_mult_90_SUMB_5__3_,
         mul_ex_mult_90_SUMB_5__4_, mul_ex_mult_90_SUMB_5__5_,
         mul_ex_mult_90_SUMB_5__6_, mul_ex_mult_90_SUMB_5__7_,
         mul_ex_mult_90_SUMB_5__8_, mul_ex_mult_90_SUMB_5__9_,
         mul_ex_mult_90_SUMB_5__10_, mul_ex_mult_90_SUMB_5__11_,
         mul_ex_mult_90_SUMB_5__12_, mul_ex_mult_90_SUMB_5__13_,
         mul_ex_mult_90_SUMB_5__14_, mul_ex_mult_90_SUMB_5__15_,
         mul_ex_mult_90_SUMB_5__16_, mul_ex_mult_90_SUMB_6__1_,
         mul_ex_mult_90_SUMB_6__2_, mul_ex_mult_90_SUMB_6__3_,
         mul_ex_mult_90_SUMB_6__4_, mul_ex_mult_90_SUMB_6__5_,
         mul_ex_mult_90_SUMB_6__6_, mul_ex_mult_90_SUMB_6__7_,
         mul_ex_mult_90_SUMB_6__8_, mul_ex_mult_90_SUMB_6__9_,
         mul_ex_mult_90_SUMB_6__10_, mul_ex_mult_90_SUMB_6__11_,
         mul_ex_mult_90_SUMB_6__12_, mul_ex_mult_90_SUMB_6__13_,
         mul_ex_mult_90_SUMB_6__14_, mul_ex_mult_90_SUMB_6__15_,
         mul_ex_mult_90_SUMB_6__16_, mul_ex_mult_90_SUMB_7__1_,
         mul_ex_mult_90_SUMB_7__2_, mul_ex_mult_90_SUMB_7__3_,
         mul_ex_mult_90_SUMB_7__4_, mul_ex_mult_90_SUMB_7__5_,
         mul_ex_mult_90_SUMB_7__6_, mul_ex_mult_90_SUMB_7__7_,
         mul_ex_mult_90_SUMB_7__8_, mul_ex_mult_90_SUMB_7__9_,
         mul_ex_mult_90_SUMB_7__10_, mul_ex_mult_90_SUMB_7__11_,
         mul_ex_mult_90_SUMB_7__12_, mul_ex_mult_90_SUMB_7__13_,
         mul_ex_mult_90_SUMB_7__14_, mul_ex_mult_90_SUMB_7__15_,
         mul_ex_mult_90_SUMB_7__16_, mul_ex_mult_90_SUMB_8__1_,
         mul_ex_mult_90_SUMB_8__2_, mul_ex_mult_90_SUMB_8__3_,
         mul_ex_mult_90_SUMB_8__4_, mul_ex_mult_90_SUMB_8__5_,
         mul_ex_mult_90_SUMB_8__6_, mul_ex_mult_90_SUMB_8__7_,
         mul_ex_mult_90_SUMB_8__8_, mul_ex_mult_90_SUMB_8__9_,
         mul_ex_mult_90_SUMB_8__10_, mul_ex_mult_90_SUMB_8__11_,
         mul_ex_mult_90_SUMB_8__12_, mul_ex_mult_90_SUMB_8__13_,
         mul_ex_mult_90_SUMB_8__14_, mul_ex_mult_90_SUMB_8__15_,
         mul_ex_mult_90_SUMB_8__16_, mul_ex_mult_90_SUMB_9__1_,
         mul_ex_mult_90_SUMB_9__2_, mul_ex_mult_90_SUMB_9__3_,
         mul_ex_mult_90_SUMB_9__4_, mul_ex_mult_90_SUMB_9__5_,
         mul_ex_mult_90_SUMB_9__6_, mul_ex_mult_90_SUMB_9__7_,
         mul_ex_mult_90_SUMB_9__8_, mul_ex_mult_90_SUMB_9__9_,
         mul_ex_mult_90_SUMB_9__10_, mul_ex_mult_90_SUMB_9__11_,
         mul_ex_mult_90_SUMB_9__12_, mul_ex_mult_90_SUMB_9__13_,
         mul_ex_mult_90_SUMB_9__14_, mul_ex_mult_90_SUMB_9__15_,
         mul_ex_mult_90_SUMB_9__16_, mul_ex_mult_90_SUMB_10__1_,
         mul_ex_mult_90_SUMB_10__2_, mul_ex_mult_90_SUMB_10__3_,
         mul_ex_mult_90_SUMB_10__4_, mul_ex_mult_90_SUMB_10__5_,
         mul_ex_mult_90_SUMB_10__6_, mul_ex_mult_90_SUMB_10__7_,
         mul_ex_mult_90_SUMB_10__8_, mul_ex_mult_90_SUMB_10__9_,
         mul_ex_mult_90_SUMB_10__10_, mul_ex_mult_90_SUMB_10__11_,
         mul_ex_mult_90_SUMB_10__12_, mul_ex_mult_90_SUMB_10__13_,
         mul_ex_mult_90_SUMB_10__14_, mul_ex_mult_90_SUMB_10__15_,
         mul_ex_mult_90_SUMB_10__16_, mul_ex_mult_90_SUMB_11__1_,
         mul_ex_mult_90_SUMB_11__2_, mul_ex_mult_90_SUMB_11__3_,
         mul_ex_mult_90_SUMB_11__4_, mul_ex_mult_90_SUMB_11__5_,
         mul_ex_mult_90_SUMB_11__6_, mul_ex_mult_90_SUMB_11__7_,
         mul_ex_mult_90_SUMB_11__8_, mul_ex_mult_90_SUMB_11__9_,
         mul_ex_mult_90_SUMB_11__10_, mul_ex_mult_90_SUMB_11__11_,
         mul_ex_mult_90_SUMB_11__12_, mul_ex_mult_90_SUMB_11__13_,
         mul_ex_mult_90_SUMB_11__14_, mul_ex_mult_90_SUMB_11__15_,
         mul_ex_mult_90_SUMB_11__16_, mul_ex_mult_90_SUMB_12__1_,
         mul_ex_mult_90_SUMB_12__2_, mul_ex_mult_90_SUMB_12__3_,
         mul_ex_mult_90_SUMB_12__4_, mul_ex_mult_90_SUMB_12__5_,
         mul_ex_mult_90_SUMB_12__6_, mul_ex_mult_90_SUMB_12__7_,
         mul_ex_mult_90_SUMB_12__8_, mul_ex_mult_90_SUMB_12__9_,
         mul_ex_mult_90_SUMB_12__10_, mul_ex_mult_90_SUMB_12__11_,
         mul_ex_mult_90_SUMB_12__12_, mul_ex_mult_90_SUMB_12__13_,
         mul_ex_mult_90_SUMB_12__14_, mul_ex_mult_90_SUMB_12__15_,
         mul_ex_mult_90_SUMB_12__16_, mul_ex_mult_90_SUMB_13__1_,
         mul_ex_mult_90_SUMB_13__2_, mul_ex_mult_90_SUMB_13__3_,
         mul_ex_mult_90_SUMB_13__4_, mul_ex_mult_90_SUMB_13__5_,
         mul_ex_mult_90_SUMB_13__6_, mul_ex_mult_90_SUMB_13__7_,
         mul_ex_mult_90_SUMB_13__8_, mul_ex_mult_90_SUMB_13__9_,
         mul_ex_mult_90_SUMB_13__10_, mul_ex_mult_90_SUMB_13__11_,
         mul_ex_mult_90_SUMB_13__12_, mul_ex_mult_90_SUMB_13__13_,
         mul_ex_mult_90_SUMB_13__14_, mul_ex_mult_90_SUMB_13__15_,
         mul_ex_mult_90_SUMB_13__16_, mul_ex_mult_90_SUMB_14__1_,
         mul_ex_mult_90_SUMB_14__2_, mul_ex_mult_90_SUMB_14__3_,
         mul_ex_mult_90_SUMB_14__4_, mul_ex_mult_90_SUMB_14__5_,
         mul_ex_mult_90_SUMB_14__6_, mul_ex_mult_90_SUMB_14__7_,
         mul_ex_mult_90_SUMB_14__8_, mul_ex_mult_90_SUMB_14__9_,
         mul_ex_mult_90_SUMB_14__10_, mul_ex_mult_90_SUMB_14__11_,
         mul_ex_mult_90_SUMB_14__12_, mul_ex_mult_90_SUMB_14__13_,
         mul_ex_mult_90_SUMB_14__14_, mul_ex_mult_90_SUMB_14__15_,
         mul_ex_mult_90_SUMB_14__16_, mul_ex_mult_90_SUMB_15__1_,
         mul_ex_mult_90_SUMB_15__2_, mul_ex_mult_90_SUMB_15__3_,
         mul_ex_mult_90_SUMB_15__4_, mul_ex_mult_90_SUMB_15__5_,
         mul_ex_mult_90_SUMB_15__6_, mul_ex_mult_90_SUMB_15__7_,
         mul_ex_mult_90_SUMB_15__8_, mul_ex_mult_90_SUMB_15__9_,
         mul_ex_mult_90_SUMB_15__10_, mul_ex_mult_90_SUMB_15__11_,
         mul_ex_mult_90_SUMB_15__12_, mul_ex_mult_90_SUMB_15__13_,
         mul_ex_mult_90_SUMB_15__14_, mul_ex_mult_90_SUMB_15__15_,
         mul_ex_mult_90_SUMB_15__16_, mul_ex_mult_90_CARRYB_2__0_,
         mul_ex_mult_90_CARRYB_2__1_, mul_ex_mult_90_CARRYB_2__2_,
         mul_ex_mult_90_CARRYB_2__3_, mul_ex_mult_90_CARRYB_2__4_,
         mul_ex_mult_90_CARRYB_2__5_, mul_ex_mult_90_CARRYB_2__6_,
         mul_ex_mult_90_CARRYB_2__7_, mul_ex_mult_90_CARRYB_2__8_,
         mul_ex_mult_90_CARRYB_2__9_, mul_ex_mult_90_CARRYB_2__10_,
         mul_ex_mult_90_CARRYB_2__11_, mul_ex_mult_90_CARRYB_2__12_,
         mul_ex_mult_90_CARRYB_2__13_, mul_ex_mult_90_CARRYB_2__14_,
         mul_ex_mult_90_CARRYB_2__15_, mul_ex_mult_90_CARRYB_3__0_,
         mul_ex_mult_90_CARRYB_3__1_, mul_ex_mult_90_CARRYB_3__2_,
         mul_ex_mult_90_CARRYB_3__3_, mul_ex_mult_90_CARRYB_3__4_,
         mul_ex_mult_90_CARRYB_3__5_, mul_ex_mult_90_CARRYB_3__6_,
         mul_ex_mult_90_CARRYB_3__7_, mul_ex_mult_90_CARRYB_3__8_,
         mul_ex_mult_90_CARRYB_3__9_, mul_ex_mult_90_CARRYB_3__10_,
         mul_ex_mult_90_CARRYB_3__11_, mul_ex_mult_90_CARRYB_3__12_,
         mul_ex_mult_90_CARRYB_3__13_, mul_ex_mult_90_CARRYB_3__14_,
         mul_ex_mult_90_CARRYB_3__15_, mul_ex_mult_90_CARRYB_4__0_,
         mul_ex_mult_90_CARRYB_4__1_, mul_ex_mult_90_CARRYB_4__2_,
         mul_ex_mult_90_CARRYB_4__3_, mul_ex_mult_90_CARRYB_4__4_,
         mul_ex_mult_90_CARRYB_4__5_, mul_ex_mult_90_CARRYB_4__6_,
         mul_ex_mult_90_CARRYB_4__7_, mul_ex_mult_90_CARRYB_4__8_,
         mul_ex_mult_90_CARRYB_4__9_, mul_ex_mult_90_CARRYB_4__10_,
         mul_ex_mult_90_CARRYB_4__11_, mul_ex_mult_90_CARRYB_4__12_,
         mul_ex_mult_90_CARRYB_4__13_, mul_ex_mult_90_CARRYB_4__14_,
         mul_ex_mult_90_CARRYB_4__15_, mul_ex_mult_90_CARRYB_5__0_,
         mul_ex_mult_90_CARRYB_5__1_, mul_ex_mult_90_CARRYB_5__2_,
         mul_ex_mult_90_CARRYB_5__3_, mul_ex_mult_90_CARRYB_5__4_,
         mul_ex_mult_90_CARRYB_5__5_, mul_ex_mult_90_CARRYB_5__6_,
         mul_ex_mult_90_CARRYB_5__7_, mul_ex_mult_90_CARRYB_5__8_,
         mul_ex_mult_90_CARRYB_5__9_, mul_ex_mult_90_CARRYB_5__10_,
         mul_ex_mult_90_CARRYB_5__11_, mul_ex_mult_90_CARRYB_5__12_,
         mul_ex_mult_90_CARRYB_5__13_, mul_ex_mult_90_CARRYB_5__14_,
         mul_ex_mult_90_CARRYB_5__15_, mul_ex_mult_90_CARRYB_6__0_,
         mul_ex_mult_90_CARRYB_6__1_, mul_ex_mult_90_CARRYB_6__2_,
         mul_ex_mult_90_CARRYB_6__3_, mul_ex_mult_90_CARRYB_6__4_,
         mul_ex_mult_90_CARRYB_6__5_, mul_ex_mult_90_CARRYB_6__6_,
         mul_ex_mult_90_CARRYB_6__7_, mul_ex_mult_90_CARRYB_6__8_,
         mul_ex_mult_90_CARRYB_6__9_, mul_ex_mult_90_CARRYB_6__10_,
         mul_ex_mult_90_CARRYB_6__11_, mul_ex_mult_90_CARRYB_6__12_,
         mul_ex_mult_90_CARRYB_6__13_, mul_ex_mult_90_CARRYB_6__14_,
         mul_ex_mult_90_CARRYB_6__15_, mul_ex_mult_90_CARRYB_7__0_,
         mul_ex_mult_90_CARRYB_7__1_, mul_ex_mult_90_CARRYB_7__2_,
         mul_ex_mult_90_CARRYB_7__3_, mul_ex_mult_90_CARRYB_7__4_,
         mul_ex_mult_90_CARRYB_7__5_, mul_ex_mult_90_CARRYB_7__6_,
         mul_ex_mult_90_CARRYB_7__7_, mul_ex_mult_90_CARRYB_7__8_,
         mul_ex_mult_90_CARRYB_7__9_, mul_ex_mult_90_CARRYB_7__10_,
         mul_ex_mult_90_CARRYB_7__11_, mul_ex_mult_90_CARRYB_7__12_,
         mul_ex_mult_90_CARRYB_7__13_, mul_ex_mult_90_CARRYB_7__14_,
         mul_ex_mult_90_CARRYB_7__15_, mul_ex_mult_90_CARRYB_8__0_,
         mul_ex_mult_90_CARRYB_8__1_, mul_ex_mult_90_CARRYB_8__2_,
         mul_ex_mult_90_CARRYB_8__3_, mul_ex_mult_90_CARRYB_8__4_,
         mul_ex_mult_90_CARRYB_8__5_, mul_ex_mult_90_CARRYB_8__6_,
         mul_ex_mult_90_CARRYB_8__7_, mul_ex_mult_90_CARRYB_8__8_,
         mul_ex_mult_90_CARRYB_8__9_, mul_ex_mult_90_CARRYB_8__10_,
         mul_ex_mult_90_CARRYB_8__11_, mul_ex_mult_90_CARRYB_8__12_,
         mul_ex_mult_90_CARRYB_8__13_, mul_ex_mult_90_CARRYB_8__14_,
         mul_ex_mult_90_CARRYB_8__15_, mul_ex_mult_90_CARRYB_9__0_,
         mul_ex_mult_90_CARRYB_9__1_, mul_ex_mult_90_CARRYB_9__2_,
         mul_ex_mult_90_CARRYB_9__3_, mul_ex_mult_90_CARRYB_9__4_,
         mul_ex_mult_90_CARRYB_9__5_, mul_ex_mult_90_CARRYB_9__6_,
         mul_ex_mult_90_CARRYB_9__7_, mul_ex_mult_90_CARRYB_9__8_,
         mul_ex_mult_90_CARRYB_9__9_, mul_ex_mult_90_CARRYB_9__10_,
         mul_ex_mult_90_CARRYB_9__11_, mul_ex_mult_90_CARRYB_9__12_,
         mul_ex_mult_90_CARRYB_9__13_, mul_ex_mult_90_CARRYB_9__14_,
         mul_ex_mult_90_CARRYB_9__15_, mul_ex_mult_90_CARRYB_10__0_,
         mul_ex_mult_90_CARRYB_10__1_, mul_ex_mult_90_CARRYB_10__2_,
         mul_ex_mult_90_CARRYB_10__3_, mul_ex_mult_90_CARRYB_10__4_,
         mul_ex_mult_90_CARRYB_10__5_, mul_ex_mult_90_CARRYB_10__6_,
         mul_ex_mult_90_CARRYB_10__7_, mul_ex_mult_90_CARRYB_10__8_,
         mul_ex_mult_90_CARRYB_10__9_, mul_ex_mult_90_CARRYB_10__10_,
         mul_ex_mult_90_CARRYB_10__11_, mul_ex_mult_90_CARRYB_10__12_,
         mul_ex_mult_90_CARRYB_10__13_, mul_ex_mult_90_CARRYB_10__14_,
         mul_ex_mult_90_CARRYB_10__15_, mul_ex_mult_90_CARRYB_11__0_,
         mul_ex_mult_90_CARRYB_11__1_, mul_ex_mult_90_CARRYB_11__2_,
         mul_ex_mult_90_CARRYB_11__3_, mul_ex_mult_90_CARRYB_11__4_,
         mul_ex_mult_90_CARRYB_11__5_, mul_ex_mult_90_CARRYB_11__6_,
         mul_ex_mult_90_CARRYB_11__7_, mul_ex_mult_90_CARRYB_11__8_,
         mul_ex_mult_90_CARRYB_11__9_, mul_ex_mult_90_CARRYB_11__10_,
         mul_ex_mult_90_CARRYB_11__11_, mul_ex_mult_90_CARRYB_11__12_,
         mul_ex_mult_90_CARRYB_11__13_, mul_ex_mult_90_CARRYB_11__14_,
         mul_ex_mult_90_CARRYB_11__15_, mul_ex_mult_90_CARRYB_12__0_,
         mul_ex_mult_90_CARRYB_12__1_, mul_ex_mult_90_CARRYB_12__2_,
         mul_ex_mult_90_CARRYB_12__3_, mul_ex_mult_90_CARRYB_12__4_,
         mul_ex_mult_90_CARRYB_12__5_, mul_ex_mult_90_CARRYB_12__6_,
         mul_ex_mult_90_CARRYB_12__7_, mul_ex_mult_90_CARRYB_12__8_,
         mul_ex_mult_90_CARRYB_12__9_, mul_ex_mult_90_CARRYB_12__10_,
         mul_ex_mult_90_CARRYB_12__11_, mul_ex_mult_90_CARRYB_12__12_,
         mul_ex_mult_90_CARRYB_12__13_, mul_ex_mult_90_CARRYB_12__14_,
         mul_ex_mult_90_CARRYB_12__15_, mul_ex_mult_90_CARRYB_13__0_,
         mul_ex_mult_90_CARRYB_13__1_, mul_ex_mult_90_CARRYB_13__2_,
         mul_ex_mult_90_CARRYB_13__3_, mul_ex_mult_90_CARRYB_13__4_,
         mul_ex_mult_90_CARRYB_13__5_, mul_ex_mult_90_CARRYB_13__6_,
         mul_ex_mult_90_CARRYB_13__7_, mul_ex_mult_90_CARRYB_13__8_,
         mul_ex_mult_90_CARRYB_13__9_, mul_ex_mult_90_CARRYB_13__10_,
         mul_ex_mult_90_CARRYB_13__11_, mul_ex_mult_90_CARRYB_13__12_,
         mul_ex_mult_90_CARRYB_13__13_, mul_ex_mult_90_CARRYB_13__14_,
         mul_ex_mult_90_CARRYB_13__15_, mul_ex_mult_90_CARRYB_14__0_,
         mul_ex_mult_90_CARRYB_14__1_, mul_ex_mult_90_CARRYB_14__2_,
         mul_ex_mult_90_CARRYB_14__3_, mul_ex_mult_90_CARRYB_14__4_,
         mul_ex_mult_90_CARRYB_14__5_, mul_ex_mult_90_CARRYB_14__6_,
         mul_ex_mult_90_CARRYB_14__7_, mul_ex_mult_90_CARRYB_14__8_,
         mul_ex_mult_90_CARRYB_14__9_, mul_ex_mult_90_CARRYB_14__10_,
         mul_ex_mult_90_CARRYB_14__11_, mul_ex_mult_90_CARRYB_14__12_,
         mul_ex_mult_90_CARRYB_14__13_, mul_ex_mult_90_CARRYB_14__14_,
         mul_ex_mult_90_CARRYB_14__15_, mul_ex_mult_90_CARRYB_15__0_,
         mul_ex_mult_90_CARRYB_15__1_, mul_ex_mult_90_CARRYB_15__2_,
         mul_ex_mult_90_CARRYB_15__3_, mul_ex_mult_90_CARRYB_15__4_,
         mul_ex_mult_90_CARRYB_15__5_, mul_ex_mult_90_CARRYB_15__6_,
         mul_ex_mult_90_CARRYB_15__7_, mul_ex_mult_90_CARRYB_15__8_,
         mul_ex_mult_90_CARRYB_15__9_, mul_ex_mult_90_CARRYB_15__10_,
         mul_ex_mult_90_CARRYB_15__11_, mul_ex_mult_90_CARRYB_15__12_,
         mul_ex_mult_90_CARRYB_15__13_, mul_ex_mult_90_CARRYB_15__14_,
         mul_ex_mult_90_CARRYB_15__15_, mul_ex_mult_90_ab_0__1_,
         mul_ex_mult_90_ab_0__2_, mul_ex_mult_90_ab_0__3_,
         mul_ex_mult_90_ab_0__4_, mul_ex_mult_90_ab_0__5_,
         mul_ex_mult_90_ab_0__6_, mul_ex_mult_90_ab_0__7_,
         mul_ex_mult_90_ab_0__8_, mul_ex_mult_90_ab_0__9_,
         mul_ex_mult_90_ab_0__10_, mul_ex_mult_90_ab_0__11_,
         mul_ex_mult_90_ab_0__12_, mul_ex_mult_90_ab_0__13_,
         mul_ex_mult_90_ab_0__14_, mul_ex_mult_90_ab_0__15_,
         mul_ex_mult_90_ab_0__16_, mul_ex_mult_90_ab_1__0_,
         mul_ex_mult_90_ab_1__1_, mul_ex_mult_90_ab_1__2_,
         mul_ex_mult_90_ab_1__3_, mul_ex_mult_90_ab_1__4_,
         mul_ex_mult_90_ab_1__5_, mul_ex_mult_90_ab_1__6_,
         mul_ex_mult_90_ab_1__7_, mul_ex_mult_90_ab_1__8_,
         mul_ex_mult_90_ab_1__9_, mul_ex_mult_90_ab_1__10_,
         mul_ex_mult_90_ab_1__11_, mul_ex_mult_90_ab_1__12_,
         mul_ex_mult_90_ab_1__13_, mul_ex_mult_90_ab_1__14_,
         mul_ex_mult_90_ab_1__15_, mul_ex_mult_90_ab_1__16_,
         mul_ex_mult_90_ab_2__0_, mul_ex_mult_90_ab_2__1_,
         mul_ex_mult_90_ab_2__2_, mul_ex_mult_90_ab_2__3_,
         mul_ex_mult_90_ab_2__4_, mul_ex_mult_90_ab_2__5_,
         mul_ex_mult_90_ab_2__6_, mul_ex_mult_90_ab_2__7_,
         mul_ex_mult_90_ab_2__8_, mul_ex_mult_90_ab_2__9_,
         mul_ex_mult_90_ab_2__10_, mul_ex_mult_90_ab_2__11_,
         mul_ex_mult_90_ab_2__12_, mul_ex_mult_90_ab_2__13_,
         mul_ex_mult_90_ab_2__14_, mul_ex_mult_90_ab_2__15_,
         mul_ex_mult_90_ab_3__0_, mul_ex_mult_90_ab_3__1_,
         mul_ex_mult_90_ab_3__2_, mul_ex_mult_90_ab_3__3_,
         mul_ex_mult_90_ab_3__4_, mul_ex_mult_90_ab_3__5_,
         mul_ex_mult_90_ab_3__6_, mul_ex_mult_90_ab_3__7_,
         mul_ex_mult_90_ab_3__8_, mul_ex_mult_90_ab_3__9_,
         mul_ex_mult_90_ab_3__10_, mul_ex_mult_90_ab_3__11_,
         mul_ex_mult_90_ab_3__12_, mul_ex_mult_90_ab_3__13_,
         mul_ex_mult_90_ab_3__14_, mul_ex_mult_90_ab_3__15_,
         mul_ex_mult_90_ab_4__0_, mul_ex_mult_90_ab_4__1_,
         mul_ex_mult_90_ab_4__2_, mul_ex_mult_90_ab_4__3_,
         mul_ex_mult_90_ab_4__4_, mul_ex_mult_90_ab_4__5_,
         mul_ex_mult_90_ab_4__6_, mul_ex_mult_90_ab_4__7_,
         mul_ex_mult_90_ab_4__8_, mul_ex_mult_90_ab_4__9_,
         mul_ex_mult_90_ab_4__10_, mul_ex_mult_90_ab_4__11_,
         mul_ex_mult_90_ab_4__12_, mul_ex_mult_90_ab_4__13_,
         mul_ex_mult_90_ab_4__14_, mul_ex_mult_90_ab_4__15_,
         mul_ex_mult_90_ab_5__0_, mul_ex_mult_90_ab_5__1_,
         mul_ex_mult_90_ab_5__2_, mul_ex_mult_90_ab_5__3_,
         mul_ex_mult_90_ab_5__4_, mul_ex_mult_90_ab_5__5_,
         mul_ex_mult_90_ab_5__6_, mul_ex_mult_90_ab_5__7_,
         mul_ex_mult_90_ab_5__8_, mul_ex_mult_90_ab_5__9_,
         mul_ex_mult_90_ab_5__10_, mul_ex_mult_90_ab_5__11_,
         mul_ex_mult_90_ab_5__12_, mul_ex_mult_90_ab_5__13_,
         mul_ex_mult_90_ab_5__14_, mul_ex_mult_90_ab_5__15_,
         mul_ex_mult_90_ab_6__0_, mul_ex_mult_90_ab_6__1_,
         mul_ex_mult_90_ab_6__2_, mul_ex_mult_90_ab_6__3_,
         mul_ex_mult_90_ab_6__4_, mul_ex_mult_90_ab_6__5_,
         mul_ex_mult_90_ab_6__6_, mul_ex_mult_90_ab_6__7_,
         mul_ex_mult_90_ab_6__8_, mul_ex_mult_90_ab_6__9_,
         mul_ex_mult_90_ab_6__10_, mul_ex_mult_90_ab_6__11_,
         mul_ex_mult_90_ab_6__12_, mul_ex_mult_90_ab_6__13_,
         mul_ex_mult_90_ab_6__14_, mul_ex_mult_90_ab_6__15_,
         mul_ex_mult_90_ab_7__0_, mul_ex_mult_90_ab_7__1_,
         mul_ex_mult_90_ab_7__2_, mul_ex_mult_90_ab_7__3_,
         mul_ex_mult_90_ab_7__4_, mul_ex_mult_90_ab_7__5_,
         mul_ex_mult_90_ab_7__6_, mul_ex_mult_90_ab_7__7_,
         mul_ex_mult_90_ab_7__8_, mul_ex_mult_90_ab_7__9_,
         mul_ex_mult_90_ab_7__10_, mul_ex_mult_90_ab_7__11_,
         mul_ex_mult_90_ab_7__12_, mul_ex_mult_90_ab_7__13_,
         mul_ex_mult_90_ab_7__14_, mul_ex_mult_90_ab_7__15_,
         mul_ex_mult_90_ab_8__0_, mul_ex_mult_90_ab_8__1_,
         mul_ex_mult_90_ab_8__2_, mul_ex_mult_90_ab_8__3_,
         mul_ex_mult_90_ab_8__4_, mul_ex_mult_90_ab_8__5_,
         mul_ex_mult_90_ab_8__6_, mul_ex_mult_90_ab_8__7_,
         mul_ex_mult_90_ab_8__8_, mul_ex_mult_90_ab_8__9_,
         mul_ex_mult_90_ab_8__10_, mul_ex_mult_90_ab_8__11_,
         mul_ex_mult_90_ab_8__12_, mul_ex_mult_90_ab_8__13_,
         mul_ex_mult_90_ab_8__14_, mul_ex_mult_90_ab_8__15_,
         mul_ex_mult_90_ab_9__0_, mul_ex_mult_90_ab_9__1_,
         mul_ex_mult_90_ab_9__2_, mul_ex_mult_90_ab_9__3_,
         mul_ex_mult_90_ab_9__4_, mul_ex_mult_90_ab_9__5_,
         mul_ex_mult_90_ab_9__6_, mul_ex_mult_90_ab_9__7_,
         mul_ex_mult_90_ab_9__8_, mul_ex_mult_90_ab_9__9_,
         mul_ex_mult_90_ab_9__10_, mul_ex_mult_90_ab_9__11_,
         mul_ex_mult_90_ab_9__12_, mul_ex_mult_90_ab_9__13_,
         mul_ex_mult_90_ab_9__14_, mul_ex_mult_90_ab_9__15_,
         mul_ex_mult_90_ab_10__0_, mul_ex_mult_90_ab_10__1_,
         mul_ex_mult_90_ab_10__2_, mul_ex_mult_90_ab_10__3_,
         mul_ex_mult_90_ab_10__4_, mul_ex_mult_90_ab_10__5_,
         mul_ex_mult_90_ab_10__6_, mul_ex_mult_90_ab_10__7_,
         mul_ex_mult_90_ab_10__8_, mul_ex_mult_90_ab_10__9_,
         mul_ex_mult_90_ab_10__10_, mul_ex_mult_90_ab_10__11_,
         mul_ex_mult_90_ab_10__12_, mul_ex_mult_90_ab_10__13_,
         mul_ex_mult_90_ab_10__14_, mul_ex_mult_90_ab_10__15_,
         mul_ex_mult_90_ab_11__0_, mul_ex_mult_90_ab_11__1_,
         mul_ex_mult_90_ab_11__2_, mul_ex_mult_90_ab_11__3_,
         mul_ex_mult_90_ab_11__4_, mul_ex_mult_90_ab_11__5_,
         mul_ex_mult_90_ab_11__6_, mul_ex_mult_90_ab_11__7_,
         mul_ex_mult_90_ab_11__8_, mul_ex_mult_90_ab_11__9_,
         mul_ex_mult_90_ab_11__10_, mul_ex_mult_90_ab_11__11_,
         mul_ex_mult_90_ab_11__12_, mul_ex_mult_90_ab_11__13_,
         mul_ex_mult_90_ab_11__14_, mul_ex_mult_90_ab_11__15_,
         mul_ex_mult_90_ab_12__0_, mul_ex_mult_90_ab_12__1_,
         mul_ex_mult_90_ab_12__2_, mul_ex_mult_90_ab_12__3_,
         mul_ex_mult_90_ab_12__4_, mul_ex_mult_90_ab_12__5_,
         mul_ex_mult_90_ab_12__6_, mul_ex_mult_90_ab_12__7_,
         mul_ex_mult_90_ab_12__8_, mul_ex_mult_90_ab_12__9_,
         mul_ex_mult_90_ab_12__10_, mul_ex_mult_90_ab_12__11_,
         mul_ex_mult_90_ab_12__12_, mul_ex_mult_90_ab_12__13_,
         mul_ex_mult_90_ab_12__14_, mul_ex_mult_90_ab_12__15_,
         mul_ex_mult_90_ab_13__0_, mul_ex_mult_90_ab_13__1_,
         mul_ex_mult_90_ab_13__2_, mul_ex_mult_90_ab_13__3_,
         mul_ex_mult_90_ab_13__4_, mul_ex_mult_90_ab_13__5_,
         mul_ex_mult_90_ab_13__6_, mul_ex_mult_90_ab_13__7_,
         mul_ex_mult_90_ab_13__8_, mul_ex_mult_90_ab_13__9_,
         mul_ex_mult_90_ab_13__10_, mul_ex_mult_90_ab_13__11_,
         mul_ex_mult_90_ab_13__12_, mul_ex_mult_90_ab_13__13_,
         mul_ex_mult_90_ab_13__14_, mul_ex_mult_90_ab_13__15_,
         mul_ex_mult_90_ab_14__0_, mul_ex_mult_90_ab_14__1_,
         mul_ex_mult_90_ab_14__2_, mul_ex_mult_90_ab_14__3_,
         mul_ex_mult_90_ab_14__4_, mul_ex_mult_90_ab_14__5_,
         mul_ex_mult_90_ab_14__6_, mul_ex_mult_90_ab_14__7_,
         mul_ex_mult_90_ab_14__8_, mul_ex_mult_90_ab_14__9_,
         mul_ex_mult_90_ab_14__10_, mul_ex_mult_90_ab_14__11_,
         mul_ex_mult_90_ab_14__12_, mul_ex_mult_90_ab_14__13_,
         mul_ex_mult_90_ab_14__14_, mul_ex_mult_90_ab_14__15_,
         mul_ex_mult_90_ab_15__0_, mul_ex_mult_90_ab_15__1_,
         mul_ex_mult_90_ab_15__2_, mul_ex_mult_90_ab_15__3_,
         mul_ex_mult_90_ab_15__4_, mul_ex_mult_90_ab_15__5_,
         mul_ex_mult_90_ab_15__6_, mul_ex_mult_90_ab_15__7_,
         mul_ex_mult_90_ab_15__8_, mul_ex_mult_90_ab_15__9_,
         mul_ex_mult_90_ab_15__10_, mul_ex_mult_90_ab_15__11_,
         mul_ex_mult_90_ab_15__12_, mul_ex_mult_90_ab_15__13_,
         mul_ex_mult_90_ab_15__14_, mul_ex_mult_90_ab_15__15_,
         mul_ex_mult_90_ab_16__0_, mul_ex_mult_90_ab_16__1_,
         mul_ex_mult_90_ab_16__2_, mul_ex_mult_90_ab_16__3_,
         mul_ex_mult_90_ab_16__4_, mul_ex_mult_90_ab_16__5_,
         mul_ex_mult_90_ab_16__6_, mul_ex_mult_90_ab_16__7_,
         mul_ex_mult_90_ab_16__8_, mul_ex_mult_90_ab_16__9_,
         mul_ex_mult_90_ab_16__10_, mul_ex_mult_90_ab_16__11_,
         mul_ex_mult_90_ab_16__12_, mul_ex_mult_90_ab_16__13_,
         mul_ex_mult_90_ab_16__14_, mul_ex_mult_90_ab_16__15_,
         mul_ex_mult_76_n94, mul_ex_mult_76_n93, mul_ex_mult_76_n92,
         mul_ex_mult_76_n91, mul_ex_mult_76_n90, mul_ex_mult_76_n89,
         mul_ex_mult_76_n88, mul_ex_mult_76_n87, mul_ex_mult_76_n86,
         mul_ex_mult_76_n85, mul_ex_mult_76_n84, mul_ex_mult_76_n83,
         mul_ex_mult_76_n82, mul_ex_mult_76_n81, mul_ex_mult_76_n80,
         mul_ex_mult_76_n79, mul_ex_mult_76_n78, mul_ex_mult_76_n77,
         mul_ex_mult_76_n76, mul_ex_mult_76_n75, mul_ex_mult_76_n74,
         mul_ex_mult_76_n73, mul_ex_mult_76_n72, mul_ex_mult_76_n71,
         mul_ex_mult_76_n70, mul_ex_mult_76_n69, mul_ex_mult_76_n68,
         mul_ex_mult_76_n67, mul_ex_mult_76_n66, mul_ex_mult_76_n65,
         mul_ex_mult_76_n64, mul_ex_mult_76_n63, mul_ex_mult_76_n62,
         mul_ex_mult_76_n61, mul_ex_mult_76_n60, mul_ex_mult_76_n59,
         mul_ex_mult_76_n58, mul_ex_mult_76_n57, mul_ex_mult_76_n56,
         mul_ex_mult_76_n55, mul_ex_mult_76_n54, mul_ex_mult_76_n53,
         mul_ex_mult_76_n52, mul_ex_mult_76_n51, mul_ex_mult_76_n50,
         mul_ex_mult_76_n49, mul_ex_mult_76_n48, mul_ex_mult_76_n47,
         mul_ex_mult_76_n45, mul_ex_mult_76_n44, mul_ex_mult_76_n43,
         mul_ex_mult_76_n42, mul_ex_mult_76_n41, mul_ex_mult_76_n40,
         mul_ex_mult_76_n39, mul_ex_mult_76_n38, mul_ex_mult_76_n37,
         mul_ex_mult_76_n36, mul_ex_mult_76_n35, mul_ex_mult_76_n34,
         mul_ex_mult_76_n33, mul_ex_mult_76_n32, mul_ex_mult_76_n31,
         mul_ex_mult_76_n30, mul_ex_mult_76_n29, mul_ex_mult_76_n28,
         mul_ex_mult_76_n27, mul_ex_mult_76_n26, mul_ex_mult_76_n25,
         mul_ex_mult_76_n24, mul_ex_mult_76_n23, mul_ex_mult_76_n22,
         mul_ex_mult_76_n21, mul_ex_mult_76_n20, mul_ex_mult_76_n19,
         mul_ex_mult_76_n18, mul_ex_mult_76_n17, mul_ex_mult_76_n16,
         mul_ex_mult_76_n15, mul_ex_mult_76_n14, mul_ex_mult_76_n13,
         mul_ex_mult_76_n12, mul_ex_mult_76_n11, mul_ex_mult_76_n10,
         mul_ex_mult_76_n9, mul_ex_mult_76_n8, mul_ex_mult_76_n7,
         mul_ex_mult_76_n6, mul_ex_mult_76_n5, mul_ex_mult_76_n4,
         mul_ex_mult_76_n3, mul_ex_mult_76_A1_0_, mul_ex_mult_76_A1_1_,
         mul_ex_mult_76_A1_2_, mul_ex_mult_76_A1_3_, mul_ex_mult_76_A1_4_,
         mul_ex_mult_76_A1_5_, mul_ex_mult_76_A1_6_, mul_ex_mult_76_A1_7_,
         mul_ex_mult_76_A1_8_, mul_ex_mult_76_A1_9_, mul_ex_mult_76_A1_10_,
         mul_ex_mult_76_A1_11_, mul_ex_mult_76_A1_12_,
         mul_ex_mult_76_SUMB_2__1_, mul_ex_mult_76_SUMB_2__2_,
         mul_ex_mult_76_SUMB_2__3_, mul_ex_mult_76_SUMB_2__4_,
         mul_ex_mult_76_SUMB_2__5_, mul_ex_mult_76_SUMB_2__6_,
         mul_ex_mult_76_SUMB_2__7_, mul_ex_mult_76_SUMB_2__8_,
         mul_ex_mult_76_SUMB_2__9_, mul_ex_mult_76_SUMB_2__10_,
         mul_ex_mult_76_SUMB_2__11_, mul_ex_mult_76_SUMB_2__12_,
         mul_ex_mult_76_SUMB_2__13_, mul_ex_mult_76_SUMB_2__14_,
         mul_ex_mult_76_SUMB_3__1_, mul_ex_mult_76_SUMB_3__2_,
         mul_ex_mult_76_SUMB_3__3_, mul_ex_mult_76_SUMB_3__4_,
         mul_ex_mult_76_SUMB_3__5_, mul_ex_mult_76_SUMB_3__6_,
         mul_ex_mult_76_SUMB_3__7_, mul_ex_mult_76_SUMB_3__8_,
         mul_ex_mult_76_SUMB_3__9_, mul_ex_mult_76_SUMB_3__10_,
         mul_ex_mult_76_SUMB_3__11_, mul_ex_mult_76_SUMB_3__12_,
         mul_ex_mult_76_SUMB_3__13_, mul_ex_mult_76_SUMB_3__14_,
         mul_ex_mult_76_SUMB_4__1_, mul_ex_mult_76_SUMB_4__2_,
         mul_ex_mult_76_SUMB_4__3_, mul_ex_mult_76_SUMB_4__4_,
         mul_ex_mult_76_SUMB_4__5_, mul_ex_mult_76_SUMB_4__6_,
         mul_ex_mult_76_SUMB_4__7_, mul_ex_mult_76_SUMB_4__8_,
         mul_ex_mult_76_SUMB_4__9_, mul_ex_mult_76_SUMB_4__10_,
         mul_ex_mult_76_SUMB_4__11_, mul_ex_mult_76_SUMB_4__12_,
         mul_ex_mult_76_SUMB_4__13_, mul_ex_mult_76_SUMB_4__14_,
         mul_ex_mult_76_SUMB_5__1_, mul_ex_mult_76_SUMB_5__2_,
         mul_ex_mult_76_SUMB_5__3_, mul_ex_mult_76_SUMB_5__4_,
         mul_ex_mult_76_SUMB_5__5_, mul_ex_mult_76_SUMB_5__6_,
         mul_ex_mult_76_SUMB_5__7_, mul_ex_mult_76_SUMB_5__8_,
         mul_ex_mult_76_SUMB_5__9_, mul_ex_mult_76_SUMB_5__10_,
         mul_ex_mult_76_SUMB_5__11_, mul_ex_mult_76_SUMB_5__12_,
         mul_ex_mult_76_SUMB_5__13_, mul_ex_mult_76_SUMB_5__14_,
         mul_ex_mult_76_SUMB_6__1_, mul_ex_mult_76_SUMB_6__2_,
         mul_ex_mult_76_SUMB_6__3_, mul_ex_mult_76_SUMB_6__4_,
         mul_ex_mult_76_SUMB_6__5_, mul_ex_mult_76_SUMB_6__6_,
         mul_ex_mult_76_SUMB_6__7_, mul_ex_mult_76_SUMB_6__8_,
         mul_ex_mult_76_SUMB_6__9_, mul_ex_mult_76_SUMB_6__10_,
         mul_ex_mult_76_SUMB_6__11_, mul_ex_mult_76_SUMB_6__12_,
         mul_ex_mult_76_SUMB_6__13_, mul_ex_mult_76_SUMB_6__14_,
         mul_ex_mult_76_SUMB_7__1_, mul_ex_mult_76_SUMB_7__2_,
         mul_ex_mult_76_SUMB_7__3_, mul_ex_mult_76_SUMB_7__4_,
         mul_ex_mult_76_SUMB_7__5_, mul_ex_mult_76_SUMB_7__6_,
         mul_ex_mult_76_SUMB_7__7_, mul_ex_mult_76_SUMB_7__8_,
         mul_ex_mult_76_SUMB_7__9_, mul_ex_mult_76_SUMB_7__10_,
         mul_ex_mult_76_SUMB_7__11_, mul_ex_mult_76_SUMB_7__12_,
         mul_ex_mult_76_SUMB_7__13_, mul_ex_mult_76_SUMB_7__14_,
         mul_ex_mult_76_SUMB_8__1_, mul_ex_mult_76_SUMB_8__2_,
         mul_ex_mult_76_SUMB_8__3_, mul_ex_mult_76_SUMB_8__4_,
         mul_ex_mult_76_SUMB_8__5_, mul_ex_mult_76_SUMB_8__6_,
         mul_ex_mult_76_SUMB_8__7_, mul_ex_mult_76_SUMB_8__8_,
         mul_ex_mult_76_SUMB_8__9_, mul_ex_mult_76_SUMB_8__10_,
         mul_ex_mult_76_SUMB_8__11_, mul_ex_mult_76_SUMB_8__12_,
         mul_ex_mult_76_SUMB_8__13_, mul_ex_mult_76_SUMB_8__14_,
         mul_ex_mult_76_SUMB_9__1_, mul_ex_mult_76_SUMB_9__2_,
         mul_ex_mult_76_SUMB_9__3_, mul_ex_mult_76_SUMB_9__4_,
         mul_ex_mult_76_SUMB_9__5_, mul_ex_mult_76_SUMB_9__6_,
         mul_ex_mult_76_SUMB_9__7_, mul_ex_mult_76_SUMB_9__8_,
         mul_ex_mult_76_SUMB_9__9_, mul_ex_mult_76_SUMB_9__10_,
         mul_ex_mult_76_SUMB_9__11_, mul_ex_mult_76_SUMB_9__12_,
         mul_ex_mult_76_SUMB_9__13_, mul_ex_mult_76_SUMB_9__14_,
         mul_ex_mult_76_SUMB_10__1_, mul_ex_mult_76_SUMB_10__2_,
         mul_ex_mult_76_SUMB_10__3_, mul_ex_mult_76_SUMB_10__4_,
         mul_ex_mult_76_SUMB_10__5_, mul_ex_mult_76_SUMB_10__6_,
         mul_ex_mult_76_SUMB_10__7_, mul_ex_mult_76_SUMB_10__8_,
         mul_ex_mult_76_SUMB_10__9_, mul_ex_mult_76_SUMB_10__10_,
         mul_ex_mult_76_SUMB_10__11_, mul_ex_mult_76_SUMB_10__12_,
         mul_ex_mult_76_SUMB_10__13_, mul_ex_mult_76_SUMB_10__14_,
         mul_ex_mult_76_SUMB_11__1_, mul_ex_mult_76_SUMB_11__2_,
         mul_ex_mult_76_SUMB_11__3_, mul_ex_mult_76_SUMB_11__4_,
         mul_ex_mult_76_SUMB_11__5_, mul_ex_mult_76_SUMB_11__6_,
         mul_ex_mult_76_SUMB_11__7_, mul_ex_mult_76_SUMB_11__8_,
         mul_ex_mult_76_SUMB_11__9_, mul_ex_mult_76_SUMB_11__10_,
         mul_ex_mult_76_SUMB_11__11_, mul_ex_mult_76_SUMB_11__12_,
         mul_ex_mult_76_SUMB_11__13_, mul_ex_mult_76_SUMB_11__14_,
         mul_ex_mult_76_SUMB_12__1_, mul_ex_mult_76_SUMB_12__2_,
         mul_ex_mult_76_SUMB_12__3_, mul_ex_mult_76_SUMB_12__4_,
         mul_ex_mult_76_SUMB_12__5_, mul_ex_mult_76_SUMB_12__6_,
         mul_ex_mult_76_SUMB_12__7_, mul_ex_mult_76_SUMB_12__8_,
         mul_ex_mult_76_SUMB_12__9_, mul_ex_mult_76_SUMB_12__10_,
         mul_ex_mult_76_SUMB_12__11_, mul_ex_mult_76_SUMB_12__12_,
         mul_ex_mult_76_SUMB_12__13_, mul_ex_mult_76_SUMB_12__14_,
         mul_ex_mult_76_SUMB_13__1_, mul_ex_mult_76_SUMB_13__2_,
         mul_ex_mult_76_SUMB_13__3_, mul_ex_mult_76_SUMB_13__4_,
         mul_ex_mult_76_SUMB_13__5_, mul_ex_mult_76_SUMB_13__6_,
         mul_ex_mult_76_SUMB_13__7_, mul_ex_mult_76_SUMB_13__8_,
         mul_ex_mult_76_SUMB_13__9_, mul_ex_mult_76_SUMB_13__10_,
         mul_ex_mult_76_SUMB_13__11_, mul_ex_mult_76_SUMB_13__12_,
         mul_ex_mult_76_SUMB_13__13_, mul_ex_mult_76_SUMB_13__14_,
         mul_ex_mult_76_SUMB_14__1_, mul_ex_mult_76_SUMB_14__2_,
         mul_ex_mult_76_SUMB_14__3_, mul_ex_mult_76_SUMB_14__4_,
         mul_ex_mult_76_SUMB_14__5_, mul_ex_mult_76_SUMB_14__6_,
         mul_ex_mult_76_SUMB_14__7_, mul_ex_mult_76_SUMB_14__8_,
         mul_ex_mult_76_SUMB_14__9_, mul_ex_mult_76_SUMB_14__10_,
         mul_ex_mult_76_SUMB_14__11_, mul_ex_mult_76_SUMB_14__12_,
         mul_ex_mult_76_SUMB_14__13_, mul_ex_mult_76_SUMB_14__14_,
         mul_ex_mult_76_SUMB_15__0_, mul_ex_mult_76_SUMB_15__1_,
         mul_ex_mult_76_SUMB_15__2_, mul_ex_mult_76_SUMB_15__3_,
         mul_ex_mult_76_SUMB_15__4_, mul_ex_mult_76_SUMB_15__5_,
         mul_ex_mult_76_SUMB_15__6_, mul_ex_mult_76_SUMB_15__7_,
         mul_ex_mult_76_SUMB_15__8_, mul_ex_mult_76_SUMB_15__9_,
         mul_ex_mult_76_SUMB_15__10_, mul_ex_mult_76_SUMB_15__11_,
         mul_ex_mult_76_SUMB_15__12_, mul_ex_mult_76_SUMB_15__13_,
         mul_ex_mult_76_SUMB_15__14_, mul_ex_mult_76_CARRYB_2__0_,
         mul_ex_mult_76_CARRYB_2__1_, mul_ex_mult_76_CARRYB_2__2_,
         mul_ex_mult_76_CARRYB_2__3_, mul_ex_mult_76_CARRYB_2__4_,
         mul_ex_mult_76_CARRYB_2__5_, mul_ex_mult_76_CARRYB_2__6_,
         mul_ex_mult_76_CARRYB_2__7_, mul_ex_mult_76_CARRYB_2__8_,
         mul_ex_mult_76_CARRYB_2__9_, mul_ex_mult_76_CARRYB_2__10_,
         mul_ex_mult_76_CARRYB_2__11_, mul_ex_mult_76_CARRYB_2__12_,
         mul_ex_mult_76_CARRYB_2__13_, mul_ex_mult_76_CARRYB_2__14_,
         mul_ex_mult_76_CARRYB_3__0_, mul_ex_mult_76_CARRYB_3__1_,
         mul_ex_mult_76_CARRYB_3__2_, mul_ex_mult_76_CARRYB_3__3_,
         mul_ex_mult_76_CARRYB_3__4_, mul_ex_mult_76_CARRYB_3__5_,
         mul_ex_mult_76_CARRYB_3__6_, mul_ex_mult_76_CARRYB_3__7_,
         mul_ex_mult_76_CARRYB_3__8_, mul_ex_mult_76_CARRYB_3__9_,
         mul_ex_mult_76_CARRYB_3__10_, mul_ex_mult_76_CARRYB_3__11_,
         mul_ex_mult_76_CARRYB_3__12_, mul_ex_mult_76_CARRYB_3__13_,
         mul_ex_mult_76_CARRYB_3__14_, mul_ex_mult_76_CARRYB_4__0_,
         mul_ex_mult_76_CARRYB_4__1_, mul_ex_mult_76_CARRYB_4__2_,
         mul_ex_mult_76_CARRYB_4__3_, mul_ex_mult_76_CARRYB_4__4_,
         mul_ex_mult_76_CARRYB_4__5_, mul_ex_mult_76_CARRYB_4__6_,
         mul_ex_mult_76_CARRYB_4__7_, mul_ex_mult_76_CARRYB_4__8_,
         mul_ex_mult_76_CARRYB_4__9_, mul_ex_mult_76_CARRYB_4__10_,
         mul_ex_mult_76_CARRYB_4__11_, mul_ex_mult_76_CARRYB_4__12_,
         mul_ex_mult_76_CARRYB_4__13_, mul_ex_mult_76_CARRYB_4__14_,
         mul_ex_mult_76_CARRYB_5__0_, mul_ex_mult_76_CARRYB_5__1_,
         mul_ex_mult_76_CARRYB_5__2_, mul_ex_mult_76_CARRYB_5__3_,
         mul_ex_mult_76_CARRYB_5__4_, mul_ex_mult_76_CARRYB_5__5_,
         mul_ex_mult_76_CARRYB_5__6_, mul_ex_mult_76_CARRYB_5__7_,
         mul_ex_mult_76_CARRYB_5__8_, mul_ex_mult_76_CARRYB_5__9_,
         mul_ex_mult_76_CARRYB_5__10_, mul_ex_mult_76_CARRYB_5__11_,
         mul_ex_mult_76_CARRYB_5__12_, mul_ex_mult_76_CARRYB_5__13_,
         mul_ex_mult_76_CARRYB_5__14_, mul_ex_mult_76_CARRYB_6__0_,
         mul_ex_mult_76_CARRYB_6__1_, mul_ex_mult_76_CARRYB_6__2_,
         mul_ex_mult_76_CARRYB_6__3_, mul_ex_mult_76_CARRYB_6__4_,
         mul_ex_mult_76_CARRYB_6__5_, mul_ex_mult_76_CARRYB_6__6_,
         mul_ex_mult_76_CARRYB_6__7_, mul_ex_mult_76_CARRYB_6__8_,
         mul_ex_mult_76_CARRYB_6__9_, mul_ex_mult_76_CARRYB_6__10_,
         mul_ex_mult_76_CARRYB_6__11_, mul_ex_mult_76_CARRYB_6__12_,
         mul_ex_mult_76_CARRYB_6__13_, mul_ex_mult_76_CARRYB_6__14_,
         mul_ex_mult_76_CARRYB_7__0_, mul_ex_mult_76_CARRYB_7__1_,
         mul_ex_mult_76_CARRYB_7__2_, mul_ex_mult_76_CARRYB_7__3_,
         mul_ex_mult_76_CARRYB_7__4_, mul_ex_mult_76_CARRYB_7__5_,
         mul_ex_mult_76_CARRYB_7__6_, mul_ex_mult_76_CARRYB_7__7_,
         mul_ex_mult_76_CARRYB_7__8_, mul_ex_mult_76_CARRYB_7__9_,
         mul_ex_mult_76_CARRYB_7__10_, mul_ex_mult_76_CARRYB_7__11_,
         mul_ex_mult_76_CARRYB_7__12_, mul_ex_mult_76_CARRYB_7__13_,
         mul_ex_mult_76_CARRYB_7__14_, mul_ex_mult_76_CARRYB_8__0_,
         mul_ex_mult_76_CARRYB_8__1_, mul_ex_mult_76_CARRYB_8__2_,
         mul_ex_mult_76_CARRYB_8__3_, mul_ex_mult_76_CARRYB_8__4_,
         mul_ex_mult_76_CARRYB_8__5_, mul_ex_mult_76_CARRYB_8__6_,
         mul_ex_mult_76_CARRYB_8__7_, mul_ex_mult_76_CARRYB_8__8_,
         mul_ex_mult_76_CARRYB_8__9_, mul_ex_mult_76_CARRYB_8__10_,
         mul_ex_mult_76_CARRYB_8__11_, mul_ex_mult_76_CARRYB_8__12_,
         mul_ex_mult_76_CARRYB_8__13_, mul_ex_mult_76_CARRYB_8__14_,
         mul_ex_mult_76_CARRYB_9__0_, mul_ex_mult_76_CARRYB_9__1_,
         mul_ex_mult_76_CARRYB_9__2_, mul_ex_mult_76_CARRYB_9__3_,
         mul_ex_mult_76_CARRYB_9__4_, mul_ex_mult_76_CARRYB_9__5_,
         mul_ex_mult_76_CARRYB_9__6_, mul_ex_mult_76_CARRYB_9__7_,
         mul_ex_mult_76_CARRYB_9__8_, mul_ex_mult_76_CARRYB_9__9_,
         mul_ex_mult_76_CARRYB_9__10_, mul_ex_mult_76_CARRYB_9__11_,
         mul_ex_mult_76_CARRYB_9__12_, mul_ex_mult_76_CARRYB_9__13_,
         mul_ex_mult_76_CARRYB_9__14_, mul_ex_mult_76_CARRYB_10__0_,
         mul_ex_mult_76_CARRYB_10__1_, mul_ex_mult_76_CARRYB_10__2_,
         mul_ex_mult_76_CARRYB_10__3_, mul_ex_mult_76_CARRYB_10__4_,
         mul_ex_mult_76_CARRYB_10__5_, mul_ex_mult_76_CARRYB_10__6_,
         mul_ex_mult_76_CARRYB_10__7_, mul_ex_mult_76_CARRYB_10__8_,
         mul_ex_mult_76_CARRYB_10__9_, mul_ex_mult_76_CARRYB_10__10_,
         mul_ex_mult_76_CARRYB_10__11_, mul_ex_mult_76_CARRYB_10__12_,
         mul_ex_mult_76_CARRYB_10__13_, mul_ex_mult_76_CARRYB_10__14_,
         mul_ex_mult_76_CARRYB_11__0_, mul_ex_mult_76_CARRYB_11__1_,
         mul_ex_mult_76_CARRYB_11__2_, mul_ex_mult_76_CARRYB_11__3_,
         mul_ex_mult_76_CARRYB_11__4_, mul_ex_mult_76_CARRYB_11__5_,
         mul_ex_mult_76_CARRYB_11__6_, mul_ex_mult_76_CARRYB_11__7_,
         mul_ex_mult_76_CARRYB_11__8_, mul_ex_mult_76_CARRYB_11__9_,
         mul_ex_mult_76_CARRYB_11__10_, mul_ex_mult_76_CARRYB_11__11_,
         mul_ex_mult_76_CARRYB_11__12_, mul_ex_mult_76_CARRYB_11__13_,
         mul_ex_mult_76_CARRYB_11__14_, mul_ex_mult_76_CARRYB_12__0_,
         mul_ex_mult_76_CARRYB_12__1_, mul_ex_mult_76_CARRYB_12__2_,
         mul_ex_mult_76_CARRYB_12__3_, mul_ex_mult_76_CARRYB_12__4_,
         mul_ex_mult_76_CARRYB_12__5_, mul_ex_mult_76_CARRYB_12__6_,
         mul_ex_mult_76_CARRYB_12__7_, mul_ex_mult_76_CARRYB_12__8_,
         mul_ex_mult_76_CARRYB_12__9_, mul_ex_mult_76_CARRYB_12__10_,
         mul_ex_mult_76_CARRYB_12__11_, mul_ex_mult_76_CARRYB_12__12_,
         mul_ex_mult_76_CARRYB_12__13_, mul_ex_mult_76_CARRYB_12__14_,
         mul_ex_mult_76_CARRYB_13__0_, mul_ex_mult_76_CARRYB_13__1_,
         mul_ex_mult_76_CARRYB_13__2_, mul_ex_mult_76_CARRYB_13__3_,
         mul_ex_mult_76_CARRYB_13__4_, mul_ex_mult_76_CARRYB_13__5_,
         mul_ex_mult_76_CARRYB_13__6_, mul_ex_mult_76_CARRYB_13__7_,
         mul_ex_mult_76_CARRYB_13__8_, mul_ex_mult_76_CARRYB_13__9_,
         mul_ex_mult_76_CARRYB_13__10_, mul_ex_mult_76_CARRYB_13__11_,
         mul_ex_mult_76_CARRYB_13__12_, mul_ex_mult_76_CARRYB_13__13_,
         mul_ex_mult_76_CARRYB_13__14_, mul_ex_mult_76_CARRYB_14__0_,
         mul_ex_mult_76_CARRYB_14__1_, mul_ex_mult_76_CARRYB_14__2_,
         mul_ex_mult_76_CARRYB_14__3_, mul_ex_mult_76_CARRYB_14__4_,
         mul_ex_mult_76_CARRYB_14__5_, mul_ex_mult_76_CARRYB_14__6_,
         mul_ex_mult_76_CARRYB_14__7_, mul_ex_mult_76_CARRYB_14__8_,
         mul_ex_mult_76_CARRYB_14__9_, mul_ex_mult_76_CARRYB_14__10_,
         mul_ex_mult_76_CARRYB_14__11_, mul_ex_mult_76_CARRYB_14__12_,
         mul_ex_mult_76_CARRYB_14__13_, mul_ex_mult_76_CARRYB_14__14_,
         mul_ex_mult_76_CARRYB_15__0_, mul_ex_mult_76_CARRYB_15__1_,
         mul_ex_mult_76_CARRYB_15__2_, mul_ex_mult_76_CARRYB_15__3_,
         mul_ex_mult_76_CARRYB_15__4_, mul_ex_mult_76_CARRYB_15__5_,
         mul_ex_mult_76_CARRYB_15__6_, mul_ex_mult_76_CARRYB_15__7_,
         mul_ex_mult_76_CARRYB_15__8_, mul_ex_mult_76_CARRYB_15__9_,
         mul_ex_mult_76_CARRYB_15__10_, mul_ex_mult_76_CARRYB_15__11_,
         mul_ex_mult_76_CARRYB_15__12_, mul_ex_mult_76_CARRYB_15__13_,
         mul_ex_mult_76_CARRYB_15__14_, mul_ex_mult_76_ab_0__1_,
         mul_ex_mult_76_ab_0__2_, mul_ex_mult_76_ab_0__3_,
         mul_ex_mult_76_ab_0__4_, mul_ex_mult_76_ab_0__5_,
         mul_ex_mult_76_ab_0__6_, mul_ex_mult_76_ab_0__7_,
         mul_ex_mult_76_ab_0__8_, mul_ex_mult_76_ab_0__9_,
         mul_ex_mult_76_ab_0__10_, mul_ex_mult_76_ab_0__11_,
         mul_ex_mult_76_ab_0__12_, mul_ex_mult_76_ab_0__13_,
         mul_ex_mult_76_ab_0__14_, mul_ex_mult_76_ab_0__15_,
         mul_ex_mult_76_ab_1__0_, mul_ex_mult_76_ab_1__1_,
         mul_ex_mult_76_ab_1__2_, mul_ex_mult_76_ab_1__3_,
         mul_ex_mult_76_ab_1__4_, mul_ex_mult_76_ab_1__5_,
         mul_ex_mult_76_ab_1__6_, mul_ex_mult_76_ab_1__7_,
         mul_ex_mult_76_ab_1__8_, mul_ex_mult_76_ab_1__9_,
         mul_ex_mult_76_ab_1__10_, mul_ex_mult_76_ab_1__11_,
         mul_ex_mult_76_ab_1__12_, mul_ex_mult_76_ab_1__13_,
         mul_ex_mult_76_ab_1__14_, mul_ex_mult_76_ab_1__15_,
         mul_ex_mult_76_ab_2__0_, mul_ex_mult_76_ab_2__1_,
         mul_ex_mult_76_ab_2__2_, mul_ex_mult_76_ab_2__3_,
         mul_ex_mult_76_ab_2__4_, mul_ex_mult_76_ab_2__5_,
         mul_ex_mult_76_ab_2__6_, mul_ex_mult_76_ab_2__7_,
         mul_ex_mult_76_ab_2__8_, mul_ex_mult_76_ab_2__9_,
         mul_ex_mult_76_ab_2__10_, mul_ex_mult_76_ab_2__11_,
         mul_ex_mult_76_ab_2__12_, mul_ex_mult_76_ab_2__13_,
         mul_ex_mult_76_ab_2__14_, mul_ex_mult_76_ab_2__15_,
         mul_ex_mult_76_ab_3__0_, mul_ex_mult_76_ab_3__1_,
         mul_ex_mult_76_ab_3__2_, mul_ex_mult_76_ab_3__3_,
         mul_ex_mult_76_ab_3__4_, mul_ex_mult_76_ab_3__5_,
         mul_ex_mult_76_ab_3__6_, mul_ex_mult_76_ab_3__7_,
         mul_ex_mult_76_ab_3__8_, mul_ex_mult_76_ab_3__9_,
         mul_ex_mult_76_ab_3__10_, mul_ex_mult_76_ab_3__11_,
         mul_ex_mult_76_ab_3__12_, mul_ex_mult_76_ab_3__13_,
         mul_ex_mult_76_ab_3__14_, mul_ex_mult_76_ab_3__15_,
         mul_ex_mult_76_ab_4__0_, mul_ex_mult_76_ab_4__1_,
         mul_ex_mult_76_ab_4__2_, mul_ex_mult_76_ab_4__3_,
         mul_ex_mult_76_ab_4__4_, mul_ex_mult_76_ab_4__5_,
         mul_ex_mult_76_ab_4__6_, mul_ex_mult_76_ab_4__7_,
         mul_ex_mult_76_ab_4__8_, mul_ex_mult_76_ab_4__9_,
         mul_ex_mult_76_ab_4__10_, mul_ex_mult_76_ab_4__11_,
         mul_ex_mult_76_ab_4__12_, mul_ex_mult_76_ab_4__13_,
         mul_ex_mult_76_ab_4__14_, mul_ex_mult_76_ab_4__15_,
         mul_ex_mult_76_ab_5__0_, mul_ex_mult_76_ab_5__1_,
         mul_ex_mult_76_ab_5__2_, mul_ex_mult_76_ab_5__3_,
         mul_ex_mult_76_ab_5__4_, mul_ex_mult_76_ab_5__5_,
         mul_ex_mult_76_ab_5__6_, mul_ex_mult_76_ab_5__7_,
         mul_ex_mult_76_ab_5__8_, mul_ex_mult_76_ab_5__9_,
         mul_ex_mult_76_ab_5__10_, mul_ex_mult_76_ab_5__11_,
         mul_ex_mult_76_ab_5__12_, mul_ex_mult_76_ab_5__13_,
         mul_ex_mult_76_ab_5__14_, mul_ex_mult_76_ab_5__15_,
         mul_ex_mult_76_ab_6__0_, mul_ex_mult_76_ab_6__1_,
         mul_ex_mult_76_ab_6__2_, mul_ex_mult_76_ab_6__3_,
         mul_ex_mult_76_ab_6__4_, mul_ex_mult_76_ab_6__5_,
         mul_ex_mult_76_ab_6__6_, mul_ex_mult_76_ab_6__7_,
         mul_ex_mult_76_ab_6__8_, mul_ex_mult_76_ab_6__9_,
         mul_ex_mult_76_ab_6__10_, mul_ex_mult_76_ab_6__11_,
         mul_ex_mult_76_ab_6__12_, mul_ex_mult_76_ab_6__13_,
         mul_ex_mult_76_ab_6__14_, mul_ex_mult_76_ab_6__15_,
         mul_ex_mult_76_ab_7__0_, mul_ex_mult_76_ab_7__1_,
         mul_ex_mult_76_ab_7__2_, mul_ex_mult_76_ab_7__3_,
         mul_ex_mult_76_ab_7__4_, mul_ex_mult_76_ab_7__5_,
         mul_ex_mult_76_ab_7__6_, mul_ex_mult_76_ab_7__7_,
         mul_ex_mult_76_ab_7__8_, mul_ex_mult_76_ab_7__9_,
         mul_ex_mult_76_ab_7__10_, mul_ex_mult_76_ab_7__11_,
         mul_ex_mult_76_ab_7__12_, mul_ex_mult_76_ab_7__13_,
         mul_ex_mult_76_ab_7__14_, mul_ex_mult_76_ab_7__15_,
         mul_ex_mult_76_ab_8__0_, mul_ex_mult_76_ab_8__1_,
         mul_ex_mult_76_ab_8__2_, mul_ex_mult_76_ab_8__3_,
         mul_ex_mult_76_ab_8__4_, mul_ex_mult_76_ab_8__5_,
         mul_ex_mult_76_ab_8__6_, mul_ex_mult_76_ab_8__7_,
         mul_ex_mult_76_ab_8__8_, mul_ex_mult_76_ab_8__9_,
         mul_ex_mult_76_ab_8__10_, mul_ex_mult_76_ab_8__11_,
         mul_ex_mult_76_ab_8__12_, mul_ex_mult_76_ab_8__13_,
         mul_ex_mult_76_ab_8__14_, mul_ex_mult_76_ab_8__15_,
         mul_ex_mult_76_ab_9__0_, mul_ex_mult_76_ab_9__1_,
         mul_ex_mult_76_ab_9__2_, mul_ex_mult_76_ab_9__3_,
         mul_ex_mult_76_ab_9__4_, mul_ex_mult_76_ab_9__5_,
         mul_ex_mult_76_ab_9__6_, mul_ex_mult_76_ab_9__7_,
         mul_ex_mult_76_ab_9__8_, mul_ex_mult_76_ab_9__9_,
         mul_ex_mult_76_ab_9__10_, mul_ex_mult_76_ab_9__11_,
         mul_ex_mult_76_ab_9__12_, mul_ex_mult_76_ab_9__13_,
         mul_ex_mult_76_ab_9__14_, mul_ex_mult_76_ab_9__15_,
         mul_ex_mult_76_ab_10__0_, mul_ex_mult_76_ab_10__1_,
         mul_ex_mult_76_ab_10__2_, mul_ex_mult_76_ab_10__3_,
         mul_ex_mult_76_ab_10__4_, mul_ex_mult_76_ab_10__5_,
         mul_ex_mult_76_ab_10__6_, mul_ex_mult_76_ab_10__7_,
         mul_ex_mult_76_ab_10__8_, mul_ex_mult_76_ab_10__9_,
         mul_ex_mult_76_ab_10__10_, mul_ex_mult_76_ab_10__11_,
         mul_ex_mult_76_ab_10__12_, mul_ex_mult_76_ab_10__13_,
         mul_ex_mult_76_ab_10__14_, mul_ex_mult_76_ab_10__15_,
         mul_ex_mult_76_ab_11__0_, mul_ex_mult_76_ab_11__1_,
         mul_ex_mult_76_ab_11__2_, mul_ex_mult_76_ab_11__3_,
         mul_ex_mult_76_ab_11__4_, mul_ex_mult_76_ab_11__5_,
         mul_ex_mult_76_ab_11__6_, mul_ex_mult_76_ab_11__7_,
         mul_ex_mult_76_ab_11__8_, mul_ex_mult_76_ab_11__9_,
         mul_ex_mult_76_ab_11__10_, mul_ex_mult_76_ab_11__11_,
         mul_ex_mult_76_ab_11__12_, mul_ex_mult_76_ab_11__13_,
         mul_ex_mult_76_ab_11__14_, mul_ex_mult_76_ab_11__15_,
         mul_ex_mult_76_ab_12__0_, mul_ex_mult_76_ab_12__1_,
         mul_ex_mult_76_ab_12__2_, mul_ex_mult_76_ab_12__3_,
         mul_ex_mult_76_ab_12__4_, mul_ex_mult_76_ab_12__5_,
         mul_ex_mult_76_ab_12__6_, mul_ex_mult_76_ab_12__7_,
         mul_ex_mult_76_ab_12__8_, mul_ex_mult_76_ab_12__9_,
         mul_ex_mult_76_ab_12__10_, mul_ex_mult_76_ab_12__11_,
         mul_ex_mult_76_ab_12__12_, mul_ex_mult_76_ab_12__13_,
         mul_ex_mult_76_ab_12__14_, mul_ex_mult_76_ab_12__15_,
         mul_ex_mult_76_ab_13__0_, mul_ex_mult_76_ab_13__1_,
         mul_ex_mult_76_ab_13__2_, mul_ex_mult_76_ab_13__3_,
         mul_ex_mult_76_ab_13__4_, mul_ex_mult_76_ab_13__5_,
         mul_ex_mult_76_ab_13__6_, mul_ex_mult_76_ab_13__7_,
         mul_ex_mult_76_ab_13__8_, mul_ex_mult_76_ab_13__9_,
         mul_ex_mult_76_ab_13__10_, mul_ex_mult_76_ab_13__11_,
         mul_ex_mult_76_ab_13__12_, mul_ex_mult_76_ab_13__13_,
         mul_ex_mult_76_ab_13__14_, mul_ex_mult_76_ab_13__15_,
         mul_ex_mult_76_ab_14__0_, mul_ex_mult_76_ab_14__1_,
         mul_ex_mult_76_ab_14__2_, mul_ex_mult_76_ab_14__3_,
         mul_ex_mult_76_ab_14__4_, mul_ex_mult_76_ab_14__5_,
         mul_ex_mult_76_ab_14__6_, mul_ex_mult_76_ab_14__7_,
         mul_ex_mult_76_ab_14__8_, mul_ex_mult_76_ab_14__9_,
         mul_ex_mult_76_ab_14__10_, mul_ex_mult_76_ab_14__11_,
         mul_ex_mult_76_ab_14__12_, mul_ex_mult_76_ab_14__13_,
         mul_ex_mult_76_ab_14__14_, mul_ex_mult_76_ab_14__15_,
         mul_ex_mult_76_ab_15__0_, mul_ex_mult_76_ab_15__1_,
         mul_ex_mult_76_ab_15__2_, mul_ex_mult_76_ab_15__3_,
         mul_ex_mult_76_ab_15__4_, mul_ex_mult_76_ab_15__5_,
         mul_ex_mult_76_ab_15__6_, mul_ex_mult_76_ab_15__7_,
         mul_ex_mult_76_ab_15__8_, mul_ex_mult_76_ab_15__9_,
         mul_ex_mult_76_ab_15__10_, mul_ex_mult_76_ab_15__11_,
         mul_ex_mult_76_ab_15__12_, mul_ex_mult_76_ab_15__13_,
         mul_ex_mult_76_ab_15__14_, mul_ex_mult_76_ab_15__15_,
         mul_ex_mult_76_FS_1_n70, mul_ex_mult_76_FS_1_n69,
         mul_ex_mult_76_FS_1_n68, mul_ex_mult_76_FS_1_n67,
         mul_ex_mult_76_FS_1_n66, mul_ex_mult_76_FS_1_n65,
         mul_ex_mult_76_FS_1_n64, mul_ex_mult_76_FS_1_n63,
         mul_ex_mult_76_FS_1_n62, mul_ex_mult_76_FS_1_n61,
         mul_ex_mult_76_FS_1_n60, mul_ex_mult_76_FS_1_n59,
         mul_ex_mult_76_FS_1_n58, mul_ex_mult_76_FS_1_n57,
         mul_ex_mult_76_FS_1_n56, mul_ex_mult_76_FS_1_n55,
         mul_ex_mult_76_FS_1_n54, mul_ex_mult_76_FS_1_n53,
         mul_ex_mult_76_FS_1_n52, mul_ex_mult_76_FS_1_n51,
         mul_ex_mult_76_FS_1_n50, mul_ex_mult_76_FS_1_n49,
         mul_ex_mult_76_FS_1_n48, mul_ex_mult_76_FS_1_n47,
         mul_ex_mult_76_FS_1_n46, mul_ex_mult_76_FS_1_n45,
         mul_ex_mult_76_FS_1_n44, mul_ex_mult_76_FS_1_n43,
         mul_ex_mult_76_FS_1_n42, mul_ex_mult_76_FS_1_n41,
         mul_ex_mult_76_FS_1_n40, mul_ex_mult_76_FS_1_n39,
         mul_ex_mult_76_FS_1_n38, mul_ex_mult_76_FS_1_n37,
         mul_ex_mult_76_FS_1_n36, mul_ex_mult_76_FS_1_n35,
         mul_ex_mult_76_FS_1_n34, mul_ex_mult_76_FS_1_n33,
         mul_ex_mult_76_FS_1_n32, mul_ex_mult_76_FS_1_n31,
         mul_ex_mult_76_FS_1_n30, mul_ex_mult_76_FS_1_n29,
         mul_ex_mult_76_FS_1_n28, mul_ex_mult_76_FS_1_n27,
         mul_ex_mult_76_FS_1_n26, mul_ex_mult_76_FS_1_n25,
         mul_ex_mult_76_FS_1_n24, mul_ex_mult_76_FS_1_n23,
         mul_ex_mult_76_FS_1_n22, mul_ex_mult_76_FS_1_n21,
         mul_ex_mult_76_FS_1_n20, mul_ex_mult_76_FS_1_n19,
         mul_ex_mult_76_FS_1_n18, mul_ex_mult_76_FS_1_n17,
         mul_ex_mult_76_FS_1_n16, mul_ex_mult_76_FS_1_n15,
         mul_ex_mult_76_FS_1_n14, mul_ex_mult_76_FS_1_n13,
         mul_ex_mult_76_FS_1_n12, mul_ex_mult_76_FS_1_n11,
         mul_ex_mult_76_FS_1_n10, mul_ex_mult_76_FS_1_n9,
         mul_ex_mult_76_FS_1_n8, mul_ex_mult_76_FS_1_n7,
         mul_ex_mult_76_FS_1_n6, mul_ex_mult_76_FS_1_n5,
         mul_ex_mult_76_FS_1_n4, mul_ex_mult_76_FS_1_n3,
         mul_ex_mult_76_FS_1_n1, mul_ex_mult_86_n94, mul_ex_mult_86_n93,
         mul_ex_mult_86_n92, mul_ex_mult_86_n91, mul_ex_mult_86_n90,
         mul_ex_mult_86_n89, mul_ex_mult_86_n88, mul_ex_mult_86_n87,
         mul_ex_mult_86_n86, mul_ex_mult_86_n85, mul_ex_mult_86_n84,
         mul_ex_mult_86_n83, mul_ex_mult_86_n82, mul_ex_mult_86_n81,
         mul_ex_mult_86_n80, mul_ex_mult_86_n79, mul_ex_mult_86_n78,
         mul_ex_mult_86_n77, mul_ex_mult_86_n76, mul_ex_mult_86_n75,
         mul_ex_mult_86_n74, mul_ex_mult_86_n73, mul_ex_mult_86_n72,
         mul_ex_mult_86_n71, mul_ex_mult_86_n70, mul_ex_mult_86_n69,
         mul_ex_mult_86_n68, mul_ex_mult_86_n67, mul_ex_mult_86_n66,
         mul_ex_mult_86_n65, mul_ex_mult_86_n64, mul_ex_mult_86_n63,
         mul_ex_mult_86_n62, mul_ex_mult_86_n61, mul_ex_mult_86_n59,
         mul_ex_mult_86_n58, mul_ex_mult_86_n57, mul_ex_mult_86_n56,
         mul_ex_mult_86_n55, mul_ex_mult_86_n54, mul_ex_mult_86_n53,
         mul_ex_mult_86_n52, mul_ex_mult_86_n51, mul_ex_mult_86_n50,
         mul_ex_mult_86_n49, mul_ex_mult_86_n48, mul_ex_mult_86_n47,
         mul_ex_mult_86_n46, mul_ex_mult_86_n45, mul_ex_mult_86_n44,
         mul_ex_mult_86_n43, mul_ex_mult_86_n42, mul_ex_mult_86_n41,
         mul_ex_mult_86_n40, mul_ex_mult_86_n39, mul_ex_mult_86_n38,
         mul_ex_mult_86_n37, mul_ex_mult_86_n36, mul_ex_mult_86_n35,
         mul_ex_mult_86_n34, mul_ex_mult_86_n33, mul_ex_mult_86_n32,
         mul_ex_mult_86_n31, mul_ex_mult_86_n30, mul_ex_mult_86_n29,
         mul_ex_mult_86_n28, mul_ex_mult_86_n27, mul_ex_mult_86_n26,
         mul_ex_mult_86_n25, mul_ex_mult_86_n24, mul_ex_mult_86_n23,
         mul_ex_mult_86_n22, mul_ex_mult_86_n21, mul_ex_mult_86_n20,
         mul_ex_mult_86_n19, mul_ex_mult_86_n18, mul_ex_mult_86_n17,
         mul_ex_mult_86_n16, mul_ex_mult_86_n15, mul_ex_mult_86_n14,
         mul_ex_mult_86_n13, mul_ex_mult_86_n12, mul_ex_mult_86_n11,
         mul_ex_mult_86_n10, mul_ex_mult_86_n9, mul_ex_mult_86_n8,
         mul_ex_mult_86_n7, mul_ex_mult_86_n6, mul_ex_mult_86_n5,
         mul_ex_mult_86_n4, mul_ex_mult_86_n3, mul_ex_mult_86_A1_0_,
         mul_ex_mult_86_A1_1_, mul_ex_mult_86_A1_2_, mul_ex_mult_86_A1_3_,
         mul_ex_mult_86_A1_4_, mul_ex_mult_86_A1_5_, mul_ex_mult_86_A1_6_,
         mul_ex_mult_86_A1_7_, mul_ex_mult_86_A1_8_, mul_ex_mult_86_A1_9_,
         mul_ex_mult_86_A1_10_, mul_ex_mult_86_A1_11_, mul_ex_mult_86_A1_12_,
         mul_ex_mult_86_SUMB_2__1_, mul_ex_mult_86_SUMB_2__2_,
         mul_ex_mult_86_SUMB_2__3_, mul_ex_mult_86_SUMB_2__4_,
         mul_ex_mult_86_SUMB_2__5_, mul_ex_mult_86_SUMB_2__6_,
         mul_ex_mult_86_SUMB_2__7_, mul_ex_mult_86_SUMB_2__8_,
         mul_ex_mult_86_SUMB_2__9_, mul_ex_mult_86_SUMB_2__10_,
         mul_ex_mult_86_SUMB_2__11_, mul_ex_mult_86_SUMB_2__12_,
         mul_ex_mult_86_SUMB_2__13_, mul_ex_mult_86_SUMB_2__14_,
         mul_ex_mult_86_SUMB_3__1_, mul_ex_mult_86_SUMB_3__2_,
         mul_ex_mult_86_SUMB_3__3_, mul_ex_mult_86_SUMB_3__4_,
         mul_ex_mult_86_SUMB_3__5_, mul_ex_mult_86_SUMB_3__6_,
         mul_ex_mult_86_SUMB_3__7_, mul_ex_mult_86_SUMB_3__8_,
         mul_ex_mult_86_SUMB_3__9_, mul_ex_mult_86_SUMB_3__10_,
         mul_ex_mult_86_SUMB_3__11_, mul_ex_mult_86_SUMB_3__12_,
         mul_ex_mult_86_SUMB_3__13_, mul_ex_mult_86_SUMB_3__14_,
         mul_ex_mult_86_SUMB_4__1_, mul_ex_mult_86_SUMB_4__2_,
         mul_ex_mult_86_SUMB_4__3_, mul_ex_mult_86_SUMB_4__4_,
         mul_ex_mult_86_SUMB_4__5_, mul_ex_mult_86_SUMB_4__6_,
         mul_ex_mult_86_SUMB_4__7_, mul_ex_mult_86_SUMB_4__8_,
         mul_ex_mult_86_SUMB_4__9_, mul_ex_mult_86_SUMB_4__10_,
         mul_ex_mult_86_SUMB_4__11_, mul_ex_mult_86_SUMB_4__12_,
         mul_ex_mult_86_SUMB_4__13_, mul_ex_mult_86_SUMB_4__14_,
         mul_ex_mult_86_SUMB_5__1_, mul_ex_mult_86_SUMB_5__2_,
         mul_ex_mult_86_SUMB_5__3_, mul_ex_mult_86_SUMB_5__4_,
         mul_ex_mult_86_SUMB_5__5_, mul_ex_mult_86_SUMB_5__6_,
         mul_ex_mult_86_SUMB_5__7_, mul_ex_mult_86_SUMB_5__8_,
         mul_ex_mult_86_SUMB_5__9_, mul_ex_mult_86_SUMB_5__10_,
         mul_ex_mult_86_SUMB_5__11_, mul_ex_mult_86_SUMB_5__12_,
         mul_ex_mult_86_SUMB_5__13_, mul_ex_mult_86_SUMB_5__14_,
         mul_ex_mult_86_SUMB_6__1_, mul_ex_mult_86_SUMB_6__2_,
         mul_ex_mult_86_SUMB_6__3_, mul_ex_mult_86_SUMB_6__4_,
         mul_ex_mult_86_SUMB_6__5_, mul_ex_mult_86_SUMB_6__6_,
         mul_ex_mult_86_SUMB_6__7_, mul_ex_mult_86_SUMB_6__8_,
         mul_ex_mult_86_SUMB_6__9_, mul_ex_mult_86_SUMB_6__10_,
         mul_ex_mult_86_SUMB_6__11_, mul_ex_mult_86_SUMB_6__12_,
         mul_ex_mult_86_SUMB_6__13_, mul_ex_mult_86_SUMB_6__14_,
         mul_ex_mult_86_SUMB_7__1_, mul_ex_mult_86_SUMB_7__2_,
         mul_ex_mult_86_SUMB_7__3_, mul_ex_mult_86_SUMB_7__4_,
         mul_ex_mult_86_SUMB_7__5_, mul_ex_mult_86_SUMB_7__6_,
         mul_ex_mult_86_SUMB_7__7_, mul_ex_mult_86_SUMB_7__8_,
         mul_ex_mult_86_SUMB_7__9_, mul_ex_mult_86_SUMB_7__10_,
         mul_ex_mult_86_SUMB_7__11_, mul_ex_mult_86_SUMB_7__12_,
         mul_ex_mult_86_SUMB_7__13_, mul_ex_mult_86_SUMB_7__14_,
         mul_ex_mult_86_SUMB_8__1_, mul_ex_mult_86_SUMB_8__2_,
         mul_ex_mult_86_SUMB_8__3_, mul_ex_mult_86_SUMB_8__4_,
         mul_ex_mult_86_SUMB_8__5_, mul_ex_mult_86_SUMB_8__6_,
         mul_ex_mult_86_SUMB_8__7_, mul_ex_mult_86_SUMB_8__8_,
         mul_ex_mult_86_SUMB_8__9_, mul_ex_mult_86_SUMB_8__10_,
         mul_ex_mult_86_SUMB_8__11_, mul_ex_mult_86_SUMB_8__12_,
         mul_ex_mult_86_SUMB_8__13_, mul_ex_mult_86_SUMB_8__14_,
         mul_ex_mult_86_SUMB_9__1_, mul_ex_mult_86_SUMB_9__2_,
         mul_ex_mult_86_SUMB_9__3_, mul_ex_mult_86_SUMB_9__4_,
         mul_ex_mult_86_SUMB_9__5_, mul_ex_mult_86_SUMB_9__6_,
         mul_ex_mult_86_SUMB_9__7_, mul_ex_mult_86_SUMB_9__8_,
         mul_ex_mult_86_SUMB_9__9_, mul_ex_mult_86_SUMB_9__10_,
         mul_ex_mult_86_SUMB_9__11_, mul_ex_mult_86_SUMB_9__12_,
         mul_ex_mult_86_SUMB_9__13_, mul_ex_mult_86_SUMB_9__14_,
         mul_ex_mult_86_SUMB_10__1_, mul_ex_mult_86_SUMB_10__2_,
         mul_ex_mult_86_SUMB_10__3_, mul_ex_mult_86_SUMB_10__4_,
         mul_ex_mult_86_SUMB_10__5_, mul_ex_mult_86_SUMB_10__6_,
         mul_ex_mult_86_SUMB_10__7_, mul_ex_mult_86_SUMB_10__8_,
         mul_ex_mult_86_SUMB_10__9_, mul_ex_mult_86_SUMB_10__10_,
         mul_ex_mult_86_SUMB_10__11_, mul_ex_mult_86_SUMB_10__12_,
         mul_ex_mult_86_SUMB_10__13_, mul_ex_mult_86_SUMB_10__14_,
         mul_ex_mult_86_SUMB_11__1_, mul_ex_mult_86_SUMB_11__2_,
         mul_ex_mult_86_SUMB_11__3_, mul_ex_mult_86_SUMB_11__4_,
         mul_ex_mult_86_SUMB_11__5_, mul_ex_mult_86_SUMB_11__6_,
         mul_ex_mult_86_SUMB_11__7_, mul_ex_mult_86_SUMB_11__8_,
         mul_ex_mult_86_SUMB_11__9_, mul_ex_mult_86_SUMB_11__10_,
         mul_ex_mult_86_SUMB_11__11_, mul_ex_mult_86_SUMB_11__12_,
         mul_ex_mult_86_SUMB_11__13_, mul_ex_mult_86_SUMB_11__14_,
         mul_ex_mult_86_SUMB_12__1_, mul_ex_mult_86_SUMB_12__2_,
         mul_ex_mult_86_SUMB_12__3_, mul_ex_mult_86_SUMB_12__4_,
         mul_ex_mult_86_SUMB_12__5_, mul_ex_mult_86_SUMB_12__6_,
         mul_ex_mult_86_SUMB_12__7_, mul_ex_mult_86_SUMB_12__8_,
         mul_ex_mult_86_SUMB_12__9_, mul_ex_mult_86_SUMB_12__10_,
         mul_ex_mult_86_SUMB_12__11_, mul_ex_mult_86_SUMB_12__12_,
         mul_ex_mult_86_SUMB_12__13_, mul_ex_mult_86_SUMB_12__14_,
         mul_ex_mult_86_SUMB_13__1_, mul_ex_mult_86_SUMB_13__2_,
         mul_ex_mult_86_SUMB_13__3_, mul_ex_mult_86_SUMB_13__4_,
         mul_ex_mult_86_SUMB_13__5_, mul_ex_mult_86_SUMB_13__6_,
         mul_ex_mult_86_SUMB_13__7_, mul_ex_mult_86_SUMB_13__8_,
         mul_ex_mult_86_SUMB_13__9_, mul_ex_mult_86_SUMB_13__10_,
         mul_ex_mult_86_SUMB_13__11_, mul_ex_mult_86_SUMB_13__12_,
         mul_ex_mult_86_SUMB_13__13_, mul_ex_mult_86_SUMB_13__14_,
         mul_ex_mult_86_SUMB_14__1_, mul_ex_mult_86_SUMB_14__2_,
         mul_ex_mult_86_SUMB_14__3_, mul_ex_mult_86_SUMB_14__4_,
         mul_ex_mult_86_SUMB_14__5_, mul_ex_mult_86_SUMB_14__6_,
         mul_ex_mult_86_SUMB_14__7_, mul_ex_mult_86_SUMB_14__8_,
         mul_ex_mult_86_SUMB_14__9_, mul_ex_mult_86_SUMB_14__10_,
         mul_ex_mult_86_SUMB_14__11_, mul_ex_mult_86_SUMB_14__12_,
         mul_ex_mult_86_SUMB_14__13_, mul_ex_mult_86_SUMB_14__14_,
         mul_ex_mult_86_SUMB_15__0_, mul_ex_mult_86_SUMB_15__1_,
         mul_ex_mult_86_SUMB_15__2_, mul_ex_mult_86_SUMB_15__3_,
         mul_ex_mult_86_SUMB_15__4_, mul_ex_mult_86_SUMB_15__5_,
         mul_ex_mult_86_SUMB_15__6_, mul_ex_mult_86_SUMB_15__7_,
         mul_ex_mult_86_SUMB_15__8_, mul_ex_mult_86_SUMB_15__9_,
         mul_ex_mult_86_SUMB_15__10_, mul_ex_mult_86_SUMB_15__11_,
         mul_ex_mult_86_SUMB_15__12_, mul_ex_mult_86_SUMB_15__13_,
         mul_ex_mult_86_SUMB_15__14_, mul_ex_mult_86_CARRYB_2__0_,
         mul_ex_mult_86_CARRYB_2__1_, mul_ex_mult_86_CARRYB_2__2_,
         mul_ex_mult_86_CARRYB_2__3_, mul_ex_mult_86_CARRYB_2__4_,
         mul_ex_mult_86_CARRYB_2__5_, mul_ex_mult_86_CARRYB_2__6_,
         mul_ex_mult_86_CARRYB_2__7_, mul_ex_mult_86_CARRYB_2__8_,
         mul_ex_mult_86_CARRYB_2__9_, mul_ex_mult_86_CARRYB_2__10_,
         mul_ex_mult_86_CARRYB_2__11_, mul_ex_mult_86_CARRYB_2__12_,
         mul_ex_mult_86_CARRYB_2__13_, mul_ex_mult_86_CARRYB_2__14_,
         mul_ex_mult_86_CARRYB_3__0_, mul_ex_mult_86_CARRYB_3__1_,
         mul_ex_mult_86_CARRYB_3__2_, mul_ex_mult_86_CARRYB_3__3_,
         mul_ex_mult_86_CARRYB_3__4_, mul_ex_mult_86_CARRYB_3__5_,
         mul_ex_mult_86_CARRYB_3__6_, mul_ex_mult_86_CARRYB_3__7_,
         mul_ex_mult_86_CARRYB_3__8_, mul_ex_mult_86_CARRYB_3__9_,
         mul_ex_mult_86_CARRYB_3__10_, mul_ex_mult_86_CARRYB_3__11_,
         mul_ex_mult_86_CARRYB_3__12_, mul_ex_mult_86_CARRYB_3__13_,
         mul_ex_mult_86_CARRYB_3__14_, mul_ex_mult_86_CARRYB_4__0_,
         mul_ex_mult_86_CARRYB_4__1_, mul_ex_mult_86_CARRYB_4__2_,
         mul_ex_mult_86_CARRYB_4__3_, mul_ex_mult_86_CARRYB_4__4_,
         mul_ex_mult_86_CARRYB_4__5_, mul_ex_mult_86_CARRYB_4__6_,
         mul_ex_mult_86_CARRYB_4__7_, mul_ex_mult_86_CARRYB_4__8_,
         mul_ex_mult_86_CARRYB_4__9_, mul_ex_mult_86_CARRYB_4__10_,
         mul_ex_mult_86_CARRYB_4__11_, mul_ex_mult_86_CARRYB_4__12_,
         mul_ex_mult_86_CARRYB_4__13_, mul_ex_mult_86_CARRYB_4__14_,
         mul_ex_mult_86_CARRYB_5__0_, mul_ex_mult_86_CARRYB_5__1_,
         mul_ex_mult_86_CARRYB_5__2_, mul_ex_mult_86_CARRYB_5__3_,
         mul_ex_mult_86_CARRYB_5__4_, mul_ex_mult_86_CARRYB_5__5_,
         mul_ex_mult_86_CARRYB_5__6_, mul_ex_mult_86_CARRYB_5__7_,
         mul_ex_mult_86_CARRYB_5__8_, mul_ex_mult_86_CARRYB_5__9_,
         mul_ex_mult_86_CARRYB_5__10_, mul_ex_mult_86_CARRYB_5__11_,
         mul_ex_mult_86_CARRYB_5__12_, mul_ex_mult_86_CARRYB_5__13_,
         mul_ex_mult_86_CARRYB_5__14_, mul_ex_mult_86_CARRYB_6__0_,
         mul_ex_mult_86_CARRYB_6__1_, mul_ex_mult_86_CARRYB_6__2_,
         mul_ex_mult_86_CARRYB_6__3_, mul_ex_mult_86_CARRYB_6__4_,
         mul_ex_mult_86_CARRYB_6__5_, mul_ex_mult_86_CARRYB_6__6_,
         mul_ex_mult_86_CARRYB_6__7_, mul_ex_mult_86_CARRYB_6__8_,
         mul_ex_mult_86_CARRYB_6__9_, mul_ex_mult_86_CARRYB_6__10_,
         mul_ex_mult_86_CARRYB_6__11_, mul_ex_mult_86_CARRYB_6__12_,
         mul_ex_mult_86_CARRYB_6__13_, mul_ex_mult_86_CARRYB_6__14_,
         mul_ex_mult_86_CARRYB_7__0_, mul_ex_mult_86_CARRYB_7__1_,
         mul_ex_mult_86_CARRYB_7__2_, mul_ex_mult_86_CARRYB_7__3_,
         mul_ex_mult_86_CARRYB_7__4_, mul_ex_mult_86_CARRYB_7__5_,
         mul_ex_mult_86_CARRYB_7__6_, mul_ex_mult_86_CARRYB_7__7_,
         mul_ex_mult_86_CARRYB_7__8_, mul_ex_mult_86_CARRYB_7__9_,
         mul_ex_mult_86_CARRYB_7__10_, mul_ex_mult_86_CARRYB_7__11_,
         mul_ex_mult_86_CARRYB_7__12_, mul_ex_mult_86_CARRYB_7__13_,
         mul_ex_mult_86_CARRYB_7__14_, mul_ex_mult_86_CARRYB_8__0_,
         mul_ex_mult_86_CARRYB_8__1_, mul_ex_mult_86_CARRYB_8__2_,
         mul_ex_mult_86_CARRYB_8__3_, mul_ex_mult_86_CARRYB_8__4_,
         mul_ex_mult_86_CARRYB_8__5_, mul_ex_mult_86_CARRYB_8__6_,
         mul_ex_mult_86_CARRYB_8__7_, mul_ex_mult_86_CARRYB_8__8_,
         mul_ex_mult_86_CARRYB_8__9_, mul_ex_mult_86_CARRYB_8__10_,
         mul_ex_mult_86_CARRYB_8__11_, mul_ex_mult_86_CARRYB_8__12_,
         mul_ex_mult_86_CARRYB_8__13_, mul_ex_mult_86_CARRYB_8__14_,
         mul_ex_mult_86_CARRYB_9__0_, mul_ex_mult_86_CARRYB_9__1_,
         mul_ex_mult_86_CARRYB_9__2_, mul_ex_mult_86_CARRYB_9__3_,
         mul_ex_mult_86_CARRYB_9__4_, mul_ex_mult_86_CARRYB_9__5_,
         mul_ex_mult_86_CARRYB_9__6_, mul_ex_mult_86_CARRYB_9__7_,
         mul_ex_mult_86_CARRYB_9__8_, mul_ex_mult_86_CARRYB_9__9_,
         mul_ex_mult_86_CARRYB_9__10_, mul_ex_mult_86_CARRYB_9__11_,
         mul_ex_mult_86_CARRYB_9__12_, mul_ex_mult_86_CARRYB_9__13_,
         mul_ex_mult_86_CARRYB_9__14_, mul_ex_mult_86_CARRYB_10__0_,
         mul_ex_mult_86_CARRYB_10__1_, mul_ex_mult_86_CARRYB_10__2_,
         mul_ex_mult_86_CARRYB_10__3_, mul_ex_mult_86_CARRYB_10__4_,
         mul_ex_mult_86_CARRYB_10__5_, mul_ex_mult_86_CARRYB_10__6_,
         mul_ex_mult_86_CARRYB_10__7_, mul_ex_mult_86_CARRYB_10__8_,
         mul_ex_mult_86_CARRYB_10__9_, mul_ex_mult_86_CARRYB_10__10_,
         mul_ex_mult_86_CARRYB_10__11_, mul_ex_mult_86_CARRYB_10__12_,
         mul_ex_mult_86_CARRYB_10__13_, mul_ex_mult_86_CARRYB_10__14_,
         mul_ex_mult_86_CARRYB_11__0_, mul_ex_mult_86_CARRYB_11__1_,
         mul_ex_mult_86_CARRYB_11__2_, mul_ex_mult_86_CARRYB_11__3_,
         mul_ex_mult_86_CARRYB_11__4_, mul_ex_mult_86_CARRYB_11__5_,
         mul_ex_mult_86_CARRYB_11__6_, mul_ex_mult_86_CARRYB_11__7_,
         mul_ex_mult_86_CARRYB_11__8_, mul_ex_mult_86_CARRYB_11__9_,
         mul_ex_mult_86_CARRYB_11__10_, mul_ex_mult_86_CARRYB_11__11_,
         mul_ex_mult_86_CARRYB_11__12_, mul_ex_mult_86_CARRYB_11__13_,
         mul_ex_mult_86_CARRYB_11__14_, mul_ex_mult_86_CARRYB_12__0_,
         mul_ex_mult_86_CARRYB_12__1_, mul_ex_mult_86_CARRYB_12__2_,
         mul_ex_mult_86_CARRYB_12__3_, mul_ex_mult_86_CARRYB_12__4_,
         mul_ex_mult_86_CARRYB_12__5_, mul_ex_mult_86_CARRYB_12__6_,
         mul_ex_mult_86_CARRYB_12__7_, mul_ex_mult_86_CARRYB_12__8_,
         mul_ex_mult_86_CARRYB_12__9_, mul_ex_mult_86_CARRYB_12__10_,
         mul_ex_mult_86_CARRYB_12__11_, mul_ex_mult_86_CARRYB_12__12_,
         mul_ex_mult_86_CARRYB_12__13_, mul_ex_mult_86_CARRYB_12__14_,
         mul_ex_mult_86_CARRYB_13__0_, mul_ex_mult_86_CARRYB_13__1_,
         mul_ex_mult_86_CARRYB_13__2_, mul_ex_mult_86_CARRYB_13__3_,
         mul_ex_mult_86_CARRYB_13__4_, mul_ex_mult_86_CARRYB_13__5_,
         mul_ex_mult_86_CARRYB_13__6_, mul_ex_mult_86_CARRYB_13__7_,
         mul_ex_mult_86_CARRYB_13__8_, mul_ex_mult_86_CARRYB_13__9_,
         mul_ex_mult_86_CARRYB_13__10_, mul_ex_mult_86_CARRYB_13__11_,
         mul_ex_mult_86_CARRYB_13__12_, mul_ex_mult_86_CARRYB_13__13_,
         mul_ex_mult_86_CARRYB_13__14_, mul_ex_mult_86_CARRYB_14__0_,
         mul_ex_mult_86_CARRYB_14__1_, mul_ex_mult_86_CARRYB_14__2_,
         mul_ex_mult_86_CARRYB_14__3_, mul_ex_mult_86_CARRYB_14__4_,
         mul_ex_mult_86_CARRYB_14__5_, mul_ex_mult_86_CARRYB_14__6_,
         mul_ex_mult_86_CARRYB_14__7_, mul_ex_mult_86_CARRYB_14__8_,
         mul_ex_mult_86_CARRYB_14__9_, mul_ex_mult_86_CARRYB_14__10_,
         mul_ex_mult_86_CARRYB_14__11_, mul_ex_mult_86_CARRYB_14__12_,
         mul_ex_mult_86_CARRYB_14__13_, mul_ex_mult_86_CARRYB_14__14_,
         mul_ex_mult_86_CARRYB_15__0_, mul_ex_mult_86_CARRYB_15__1_,
         mul_ex_mult_86_CARRYB_15__2_, mul_ex_mult_86_CARRYB_15__3_,
         mul_ex_mult_86_CARRYB_15__4_, mul_ex_mult_86_CARRYB_15__5_,
         mul_ex_mult_86_CARRYB_15__6_, mul_ex_mult_86_CARRYB_15__7_,
         mul_ex_mult_86_CARRYB_15__8_, mul_ex_mult_86_CARRYB_15__9_,
         mul_ex_mult_86_CARRYB_15__10_, mul_ex_mult_86_CARRYB_15__11_,
         mul_ex_mult_86_CARRYB_15__12_, mul_ex_mult_86_CARRYB_15__13_,
         mul_ex_mult_86_CARRYB_15__14_, mul_ex_mult_86_ab_0__1_,
         mul_ex_mult_86_ab_0__2_, mul_ex_mult_86_ab_0__3_,
         mul_ex_mult_86_ab_0__4_, mul_ex_mult_86_ab_0__5_,
         mul_ex_mult_86_ab_0__6_, mul_ex_mult_86_ab_0__7_,
         mul_ex_mult_86_ab_0__8_, mul_ex_mult_86_ab_0__9_,
         mul_ex_mult_86_ab_0__10_, mul_ex_mult_86_ab_0__11_,
         mul_ex_mult_86_ab_0__12_, mul_ex_mult_86_ab_0__13_,
         mul_ex_mult_86_ab_0__14_, mul_ex_mult_86_ab_0__15_,
         mul_ex_mult_86_ab_1__0_, mul_ex_mult_86_ab_1__1_,
         mul_ex_mult_86_ab_1__2_, mul_ex_mult_86_ab_1__3_,
         mul_ex_mult_86_ab_1__4_, mul_ex_mult_86_ab_1__5_,
         mul_ex_mult_86_ab_1__6_, mul_ex_mult_86_ab_1__7_,
         mul_ex_mult_86_ab_1__8_, mul_ex_mult_86_ab_1__9_,
         mul_ex_mult_86_ab_1__10_, mul_ex_mult_86_ab_1__11_,
         mul_ex_mult_86_ab_1__12_, mul_ex_mult_86_ab_1__13_,
         mul_ex_mult_86_ab_1__14_, mul_ex_mult_86_ab_1__15_,
         mul_ex_mult_86_ab_2__0_, mul_ex_mult_86_ab_2__1_,
         mul_ex_mult_86_ab_2__2_, mul_ex_mult_86_ab_2__3_,
         mul_ex_mult_86_ab_2__4_, mul_ex_mult_86_ab_2__5_,
         mul_ex_mult_86_ab_2__6_, mul_ex_mult_86_ab_2__7_,
         mul_ex_mult_86_ab_2__8_, mul_ex_mult_86_ab_2__9_,
         mul_ex_mult_86_ab_2__10_, mul_ex_mult_86_ab_2__11_,
         mul_ex_mult_86_ab_2__12_, mul_ex_mult_86_ab_2__13_,
         mul_ex_mult_86_ab_2__14_, mul_ex_mult_86_ab_2__15_,
         mul_ex_mult_86_ab_3__0_, mul_ex_mult_86_ab_3__1_,
         mul_ex_mult_86_ab_3__2_, mul_ex_mult_86_ab_3__3_,
         mul_ex_mult_86_ab_3__4_, mul_ex_mult_86_ab_3__5_,
         mul_ex_mult_86_ab_3__6_, mul_ex_mult_86_ab_3__7_,
         mul_ex_mult_86_ab_3__8_, mul_ex_mult_86_ab_3__9_,
         mul_ex_mult_86_ab_3__10_, mul_ex_mult_86_ab_3__11_,
         mul_ex_mult_86_ab_3__12_, mul_ex_mult_86_ab_3__13_,
         mul_ex_mult_86_ab_3__14_, mul_ex_mult_86_ab_3__15_,
         mul_ex_mult_86_ab_4__0_, mul_ex_mult_86_ab_4__1_,
         mul_ex_mult_86_ab_4__2_, mul_ex_mult_86_ab_4__3_,
         mul_ex_mult_86_ab_4__4_, mul_ex_mult_86_ab_4__5_,
         mul_ex_mult_86_ab_4__6_, mul_ex_mult_86_ab_4__7_,
         mul_ex_mult_86_ab_4__8_, mul_ex_mult_86_ab_4__9_,
         mul_ex_mult_86_ab_4__10_, mul_ex_mult_86_ab_4__11_,
         mul_ex_mult_86_ab_4__12_, mul_ex_mult_86_ab_4__13_,
         mul_ex_mult_86_ab_4__14_, mul_ex_mult_86_ab_4__15_,
         mul_ex_mult_86_ab_5__0_, mul_ex_mult_86_ab_5__1_,
         mul_ex_mult_86_ab_5__2_, mul_ex_mult_86_ab_5__3_,
         mul_ex_mult_86_ab_5__4_, mul_ex_mult_86_ab_5__5_,
         mul_ex_mult_86_ab_5__6_, mul_ex_mult_86_ab_5__7_,
         mul_ex_mult_86_ab_5__8_, mul_ex_mult_86_ab_5__9_,
         mul_ex_mult_86_ab_5__10_, mul_ex_mult_86_ab_5__11_,
         mul_ex_mult_86_ab_5__12_, mul_ex_mult_86_ab_5__13_,
         mul_ex_mult_86_ab_5__14_, mul_ex_mult_86_ab_5__15_,
         mul_ex_mult_86_ab_6__0_, mul_ex_mult_86_ab_6__1_,
         mul_ex_mult_86_ab_6__2_, mul_ex_mult_86_ab_6__3_,
         mul_ex_mult_86_ab_6__4_, mul_ex_mult_86_ab_6__5_,
         mul_ex_mult_86_ab_6__6_, mul_ex_mult_86_ab_6__7_,
         mul_ex_mult_86_ab_6__8_, mul_ex_mult_86_ab_6__9_,
         mul_ex_mult_86_ab_6__10_, mul_ex_mult_86_ab_6__11_,
         mul_ex_mult_86_ab_6__12_, mul_ex_mult_86_ab_6__13_,
         mul_ex_mult_86_ab_6__14_, mul_ex_mult_86_ab_6__15_,
         mul_ex_mult_86_ab_7__0_, mul_ex_mult_86_ab_7__1_,
         mul_ex_mult_86_ab_7__2_, mul_ex_mult_86_ab_7__3_,
         mul_ex_mult_86_ab_7__4_, mul_ex_mult_86_ab_7__5_,
         mul_ex_mult_86_ab_7__6_, mul_ex_mult_86_ab_7__7_,
         mul_ex_mult_86_ab_7__8_, mul_ex_mult_86_ab_7__9_,
         mul_ex_mult_86_ab_7__10_, mul_ex_mult_86_ab_7__11_,
         mul_ex_mult_86_ab_7__12_, mul_ex_mult_86_ab_7__13_,
         mul_ex_mult_86_ab_7__14_, mul_ex_mult_86_ab_7__15_,
         mul_ex_mult_86_ab_8__0_, mul_ex_mult_86_ab_8__1_,
         mul_ex_mult_86_ab_8__2_, mul_ex_mult_86_ab_8__3_,
         mul_ex_mult_86_ab_8__4_, mul_ex_mult_86_ab_8__5_,
         mul_ex_mult_86_ab_8__6_, mul_ex_mult_86_ab_8__7_,
         mul_ex_mult_86_ab_8__8_, mul_ex_mult_86_ab_8__9_,
         mul_ex_mult_86_ab_8__10_, mul_ex_mult_86_ab_8__11_,
         mul_ex_mult_86_ab_8__12_, mul_ex_mult_86_ab_8__13_,
         mul_ex_mult_86_ab_8__14_, mul_ex_mult_86_ab_8__15_,
         mul_ex_mult_86_ab_9__0_, mul_ex_mult_86_ab_9__1_,
         mul_ex_mult_86_ab_9__2_, mul_ex_mult_86_ab_9__3_,
         mul_ex_mult_86_ab_9__4_, mul_ex_mult_86_ab_9__5_,
         mul_ex_mult_86_ab_9__6_, mul_ex_mult_86_ab_9__7_,
         mul_ex_mult_86_ab_9__8_, mul_ex_mult_86_ab_9__9_,
         mul_ex_mult_86_ab_9__10_, mul_ex_mult_86_ab_9__11_,
         mul_ex_mult_86_ab_9__12_, mul_ex_mult_86_ab_9__13_,
         mul_ex_mult_86_ab_9__14_, mul_ex_mult_86_ab_9__15_,
         mul_ex_mult_86_ab_10__0_, mul_ex_mult_86_ab_10__1_,
         mul_ex_mult_86_ab_10__2_, mul_ex_mult_86_ab_10__3_,
         mul_ex_mult_86_ab_10__4_, mul_ex_mult_86_ab_10__5_,
         mul_ex_mult_86_ab_10__6_, mul_ex_mult_86_ab_10__7_,
         mul_ex_mult_86_ab_10__8_, mul_ex_mult_86_ab_10__9_,
         mul_ex_mult_86_ab_10__10_, mul_ex_mult_86_ab_10__11_,
         mul_ex_mult_86_ab_10__12_, mul_ex_mult_86_ab_10__13_,
         mul_ex_mult_86_ab_10__14_, mul_ex_mult_86_ab_10__15_,
         mul_ex_mult_86_ab_11__0_, mul_ex_mult_86_ab_11__1_,
         mul_ex_mult_86_ab_11__2_, mul_ex_mult_86_ab_11__3_,
         mul_ex_mult_86_ab_11__4_, mul_ex_mult_86_ab_11__5_,
         mul_ex_mult_86_ab_11__6_, mul_ex_mult_86_ab_11__7_,
         mul_ex_mult_86_ab_11__8_, mul_ex_mult_86_ab_11__9_,
         mul_ex_mult_86_ab_11__10_, mul_ex_mult_86_ab_11__11_,
         mul_ex_mult_86_ab_11__12_, mul_ex_mult_86_ab_11__13_,
         mul_ex_mult_86_ab_11__14_, mul_ex_mult_86_ab_11__15_,
         mul_ex_mult_86_ab_12__0_, mul_ex_mult_86_ab_12__1_,
         mul_ex_mult_86_ab_12__2_, mul_ex_mult_86_ab_12__3_,
         mul_ex_mult_86_ab_12__4_, mul_ex_mult_86_ab_12__5_,
         mul_ex_mult_86_ab_12__6_, mul_ex_mult_86_ab_12__7_,
         mul_ex_mult_86_ab_12__8_, mul_ex_mult_86_ab_12__9_,
         mul_ex_mult_86_ab_12__10_, mul_ex_mult_86_ab_12__11_,
         mul_ex_mult_86_ab_12__12_, mul_ex_mult_86_ab_12__13_,
         mul_ex_mult_86_ab_12__14_, mul_ex_mult_86_ab_12__15_,
         mul_ex_mult_86_ab_13__0_, mul_ex_mult_86_ab_13__1_,
         mul_ex_mult_86_ab_13__2_, mul_ex_mult_86_ab_13__3_,
         mul_ex_mult_86_ab_13__4_, mul_ex_mult_86_ab_13__5_,
         mul_ex_mult_86_ab_13__6_, mul_ex_mult_86_ab_13__7_,
         mul_ex_mult_86_ab_13__8_, mul_ex_mult_86_ab_13__9_,
         mul_ex_mult_86_ab_13__10_, mul_ex_mult_86_ab_13__11_,
         mul_ex_mult_86_ab_13__12_, mul_ex_mult_86_ab_13__13_,
         mul_ex_mult_86_ab_13__14_, mul_ex_mult_86_ab_13__15_,
         mul_ex_mult_86_ab_14__0_, mul_ex_mult_86_ab_14__1_,
         mul_ex_mult_86_ab_14__2_, mul_ex_mult_86_ab_14__3_,
         mul_ex_mult_86_ab_14__4_, mul_ex_mult_86_ab_14__5_,
         mul_ex_mult_86_ab_14__6_, mul_ex_mult_86_ab_14__7_,
         mul_ex_mult_86_ab_14__8_, mul_ex_mult_86_ab_14__9_,
         mul_ex_mult_86_ab_14__10_, mul_ex_mult_86_ab_14__11_,
         mul_ex_mult_86_ab_14__12_, mul_ex_mult_86_ab_14__13_,
         mul_ex_mult_86_ab_14__14_, mul_ex_mult_86_ab_14__15_,
         mul_ex_mult_86_ab_15__0_, mul_ex_mult_86_ab_15__1_,
         mul_ex_mult_86_ab_15__2_, mul_ex_mult_86_ab_15__3_,
         mul_ex_mult_86_ab_15__4_, mul_ex_mult_86_ab_15__5_,
         mul_ex_mult_86_ab_15__6_, mul_ex_mult_86_ab_15__7_,
         mul_ex_mult_86_ab_15__8_, mul_ex_mult_86_ab_15__9_,
         mul_ex_mult_86_ab_15__10_, mul_ex_mult_86_ab_15__11_,
         mul_ex_mult_86_ab_15__12_, mul_ex_mult_86_ab_15__13_,
         mul_ex_mult_86_ab_15__14_, mul_ex_mult_86_ab_15__15_,
         mul_ex_mult_86_FS_1_n70, mul_ex_mult_86_FS_1_n69,
         mul_ex_mult_86_FS_1_n68, mul_ex_mult_86_FS_1_n67,
         mul_ex_mult_86_FS_1_n66, mul_ex_mult_86_FS_1_n65,
         mul_ex_mult_86_FS_1_n64, mul_ex_mult_86_FS_1_n63,
         mul_ex_mult_86_FS_1_n62, mul_ex_mult_86_FS_1_n61,
         mul_ex_mult_86_FS_1_n60, mul_ex_mult_86_FS_1_n59,
         mul_ex_mult_86_FS_1_n58, mul_ex_mult_86_FS_1_n57,
         mul_ex_mult_86_FS_1_n56, mul_ex_mult_86_FS_1_n55,
         mul_ex_mult_86_FS_1_n54, mul_ex_mult_86_FS_1_n53,
         mul_ex_mult_86_FS_1_n52, mul_ex_mult_86_FS_1_n51,
         mul_ex_mult_86_FS_1_n50, mul_ex_mult_86_FS_1_n49,
         mul_ex_mult_86_FS_1_n48, mul_ex_mult_86_FS_1_n47,
         mul_ex_mult_86_FS_1_n46, mul_ex_mult_86_FS_1_n45,
         mul_ex_mult_86_FS_1_n44, mul_ex_mult_86_FS_1_n43,
         mul_ex_mult_86_FS_1_n42, mul_ex_mult_86_FS_1_n41,
         mul_ex_mult_86_FS_1_n40, mul_ex_mult_86_FS_1_n39,
         mul_ex_mult_86_FS_1_n38, mul_ex_mult_86_FS_1_n37,
         mul_ex_mult_86_FS_1_n36, mul_ex_mult_86_FS_1_n35,
         mul_ex_mult_86_FS_1_n34, mul_ex_mult_86_FS_1_n33,
         mul_ex_mult_86_FS_1_n32, mul_ex_mult_86_FS_1_n31,
         mul_ex_mult_86_FS_1_n30, mul_ex_mult_86_FS_1_n29,
         mul_ex_mult_86_FS_1_n28, mul_ex_mult_86_FS_1_n27,
         mul_ex_mult_86_FS_1_n26, mul_ex_mult_86_FS_1_n25,
         mul_ex_mult_86_FS_1_n24, mul_ex_mult_86_FS_1_n23,
         mul_ex_mult_86_FS_1_n22, mul_ex_mult_86_FS_1_n21,
         mul_ex_mult_86_FS_1_n20, mul_ex_mult_86_FS_1_n19,
         mul_ex_mult_86_FS_1_n18, mul_ex_mult_86_FS_1_n17,
         mul_ex_mult_86_FS_1_n16, mul_ex_mult_86_FS_1_n15,
         mul_ex_mult_86_FS_1_n14, mul_ex_mult_86_FS_1_n13,
         mul_ex_mult_86_FS_1_n12, mul_ex_mult_86_FS_1_n11,
         mul_ex_mult_86_FS_1_n10, mul_ex_mult_86_FS_1_n9,
         mul_ex_mult_86_FS_1_n8, mul_ex_mult_86_FS_1_n7,
         mul_ex_mult_86_FS_1_n6, mul_ex_mult_86_FS_1_n5,
         mul_ex_mult_86_FS_1_n4, mul_ex_mult_86_FS_1_n3,
         mul_ex_mult_86_FS_1_n1, CHOOSE_MULT_OR_INT_n8, CHOOSE_MULT_OR_INT_n7,
         CHOOSE_MULT_OR_INT_n6, CHOOSE_MULT_OR_INT_n5, CHOOSE_MULT_OR_INT_n4,
         CHOOSE_MULT_OR_INT_n3, CHOOSE_MULT_OR_INT_n2, CHOOSE_MULT_OR_INT_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_0__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_1__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_2__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_3__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_4__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_5__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_6__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_7__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_8__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_9__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_10__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_11__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_12__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_13__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_14__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_15__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_16__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_17__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_18__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_19__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_20__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_21__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_22__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_23__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_24__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_25__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_26__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_27__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_28__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_29__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_30__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_31__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_32__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_32__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_33__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_33__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_34__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_34__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_35__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_35__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_36__MUX_n5,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_36__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_36__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_37__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_37__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_38__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_38__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_39__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_39__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_40__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_40__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_41__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_41__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_42__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_42__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_43__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_43__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_44__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_44__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_45__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_45__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_46__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_46__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_47__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_47__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_48__MUX_n5,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_48__MUX_n2,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_48__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_49__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_49__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_50__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_50__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_51__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_51__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_52__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_52__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_53__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_53__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_54__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_54__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_55__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_55__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_56__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_56__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_57__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_57__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_58__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_58__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_59__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_59__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_60__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_60__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_61__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_61__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_62__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_62__MUX_n1,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_63__MUX_n4,
         CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_63__MUX_n1, decide_if_leap_n3,
         decide_if_leap_n2, decide_if_leap_zeroBit, decide_if_leap_ZERO_A_n10,
         decide_if_leap_ZERO_A_n9, decide_if_leap_ZERO_A_n8,
         decide_if_leap_ZERO_A_n7, decide_if_leap_ZERO_A_n6,
         decide_if_leap_ZERO_A_n5, decide_if_leap_ZERO_A_n4,
         decide_if_leap_ZERO_A_n3, decide_if_leap_ZERO_A_n2,
         decide_if_leap_ZERO_A_n1, EXTEND_IMM16_n18, CHOOSE_IMMEDIATE_n3,
         CHOOSE_IMMEDIATE_n2, CHOOSE_IMMEDIATE_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_0__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_0__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_1__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_1__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_2__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_2__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_3__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_3__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_4__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_4__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_5__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_5__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_6__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_6__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_7__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_7__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_8__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_8__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_9__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_9__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_10__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_10__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_11__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_11__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_12__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_12__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_13__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_13__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_14__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_14__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_15__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_15__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_16__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_16__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_17__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_17__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_18__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_18__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_19__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_19__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_20__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_20__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_21__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_21__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_22__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_22__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_23__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_23__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_24__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_24__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_25__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_25__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_26__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_26__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_27__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_27__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_28__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_28__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_29__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_29__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_30__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_30__MUX_n1,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_31__MUX_n4,
         CHOOSE_IMMEDIATE_MUX2TO1_32BIT_31__MUX_n1;
  wire   [0:31] not_mul_result;
  wire   [0:63] mul_result_long;
  wire   [0:31] imm16_32;
  wire   [0:31] imm26_32;
  wire   [0:31] alu_ex_add_sub_in;
  wire   [0:31] alu_ex_b_not;
  wire   [0:31] alu_ex_xor_out;
  wire   [0:31] alu_ex_or_out;
  wire   [1:31] alu_ex_FULL_ADDER_carry;
  wire   [0:31] alu_ex_SHIFTER_rtemp4;
  wire   [0:31] alu_ex_SHIFTER_ltemp4;
  wire   [0:31] alu_ex_SET_FLAGS_b_not;
  wire   [0:31] alu_ex_FINAL_MUX_bus2;
  wire   [0:31] alu_ex_FINAL_MUX_bus1;
  wire   [0:31] alu_ex_FINAL_MUX_MUX_BUS1_bus2;
  wire   [0:31] alu_ex_FINAL_MUX_MUX_BUS1_bus1;
  wire   [0:31] alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1;
  wire   [0:31] alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2;
  wire   [0:31] alu_ex_FINAL_MUX_MUX_BUS2_bus2;
  wire   [0:31] alu_ex_FINAL_MUX_MUX_BUS2_bus1;
  wire   [0:31] alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2;
  wire   [0:31] alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1;
  wire   [0:31] alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2;
  wire   [0:31] alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1;
  wire   [0:31] mul_ex_P2;
  wire   [0:31] mul_ex_P;
  wire   [0:31] mul_ex_P1;
  wire   [0:31] mul_ex_H;
  wire   [15:2] mul_ex_add_85_carry;
  wire   [15:2] mul_ex_add_77_carry;
  wire   [31:1] mul_ex_sub_1_root_sub_0_root_sub_94_2_carry;
  wire   [31:1] mul_ex_sub_0_root_sub_0_root_sub_94_2_carry;

  NOR2_X2 U5 ( .A1(mul_done), .A2(n2), .ZN(stall_out) );
  INV_X4 U6 ( .A(mul_in), .ZN(n2) );
  BUF_X32 U8 ( .A(mul_in), .Z(mul_out) );
  BUF_X32 U9 ( .A(FPRegWrite_in), .Z(FPRegWrite_out) );
  BUF_X32 U10 ( .A(fDestReg_in[4]), .Z(fDestReg_out[4]) );
  BUF_X32 U11 ( .A(fDestReg_in[3]), .Z(fDestReg_out[3]) );
  BUF_X32 U12 ( .A(fDestReg_in[2]), .Z(fDestReg_out[2]) );
  BUF_X32 U13 ( .A(fDestReg_in[1]), .Z(fDestReg_out[1]) );
  BUF_X32 U14 ( .A(fDestReg_in[0]), .Z(fDestReg_out[0]) );
  BUF_X32 U15 ( .A(memVal_in[31]), .Z(memVal_out[31]) );
  BUF_X32 U16 ( .A(memVal_in[30]), .Z(memVal_out[30]) );
  BUF_X32 U17 ( .A(memVal_in[29]), .Z(memVal_out[29]) );
  BUF_X32 U18 ( .A(memVal_in[28]), .Z(memVal_out[28]) );
  BUF_X32 U19 ( .A(memVal_in[27]), .Z(memVal_out[27]) );
  BUF_X32 U20 ( .A(memVal_in[26]), .Z(memVal_out[26]) );
  BUF_X32 U21 ( .A(memVal_in[25]), .Z(memVal_out[25]) );
  BUF_X32 U22 ( .A(memVal_in[24]), .Z(memVal_out[24]) );
  BUF_X32 U23 ( .A(memVal_in[23]), .Z(memVal_out[23]) );
  BUF_X32 U24 ( .A(memVal_in[22]), .Z(memVal_out[22]) );
  BUF_X32 U25 ( .A(memVal_in[21]), .Z(memVal_out[21]) );
  BUF_X32 U26 ( .A(memVal_in[20]), .Z(memVal_out[20]) );
  BUF_X32 U27 ( .A(memVal_in[19]), .Z(memVal_out[19]) );
  BUF_X32 U28 ( .A(memVal_in[18]), .Z(memVal_out[18]) );
  BUF_X32 U29 ( .A(memVal_in[17]), .Z(memVal_out[17]) );
  BUF_X32 U30 ( .A(memVal_in[16]), .Z(memVal_out[16]) );
  BUF_X32 U31 ( .A(memVal_in[15]), .Z(memVal_out[15]) );
  BUF_X32 U32 ( .A(memVal_in[14]), .Z(memVal_out[14]) );
  BUF_X32 U33 ( .A(memVal_in[13]), .Z(memVal_out[13]) );
  BUF_X32 U34 ( .A(memVal_in[12]), .Z(memVal_out[12]) );
  BUF_X32 U35 ( .A(memVal_in[11]), .Z(memVal_out[11]) );
  BUF_X32 U36 ( .A(memVal_in[10]), .Z(memVal_out[10]) );
  BUF_X32 U37 ( .A(memVal_in[9]), .Z(memVal_out[9]) );
  BUF_X32 U38 ( .A(memVal_in[8]), .Z(memVal_out[8]) );
  BUF_X32 U39 ( .A(memVal_in[7]), .Z(memVal_out[7]) );
  BUF_X32 U40 ( .A(memVal_in[6]), .Z(memVal_out[6]) );
  BUF_X32 U41 ( .A(memVal_in[5]), .Z(memVal_out[5]) );
  BUF_X32 U42 ( .A(memVal_in[4]), .Z(memVal_out[4]) );
  BUF_X32 U43 ( .A(memVal_in[3]), .Z(memVal_out[3]) );
  BUF_X32 U44 ( .A(memVal_in[2]), .Z(memVal_out[2]) );
  BUF_X32 U45 ( .A(memVal_in[1]), .Z(memVal_out[1]) );
  BUF_X32 U46 ( .A(memVal_in[0]), .Z(memVal_out[0]) );
  BUF_X32 U47 ( .A(DSize_in[1]), .Z(DSize_out[1]) );
  BUF_X32 U48 ( .A(DSize_in[0]), .Z(DSize_out[0]) );
  BUF_X32 U49 ( .A(loadSign_in), .Z(loadSign_out) );
  BUF_X32 U50 ( .A(MemWrite_in), .Z(MemWrite_out) );
  BUF_X32 U51 ( .A(MemToReg_in), .Z(MemToReg_out) );
  BUF_X32 U52 ( .A(RegWrite_in), .Z(RegWrite_out) );
  BUF_X32 U53 ( .A(RegToPC_in), .Z(RegToPC_out) );
  BUF_X32 U54 ( .A(PCtoReg_in), .Z(PCtoReg_out) );
  BUF_X32 U55 ( .A(destReg_in[4]), .Z(destReg_out[4]) );
  BUF_X32 U56 ( .A(destReg_in[3]), .Z(destReg_out[3]) );
  BUF_X32 U57 ( .A(destReg_in[2]), .Z(destReg_out[2]) );
  BUF_X32 U58 ( .A(destReg_in[1]), .Z(destReg_out[1]) );
  BUF_X32 U59 ( .A(destReg_in[0]), .Z(destReg_out[0]) );
  BUF_X32 U60 ( .A(nextPC_in[31]), .Z(nextPC_out[31]) );
  BUF_X32 U61 ( .A(nextPC_in[30]), .Z(nextPC_out[30]) );
  BUF_X32 U62 ( .A(nextPC_in[29]), .Z(nextPC_out[29]) );
  BUF_X32 U63 ( .A(nextPC_in[28]), .Z(nextPC_out[28]) );
  BUF_X32 U64 ( .A(nextPC_in[27]), .Z(nextPC_out[27]) );
  BUF_X32 U65 ( .A(nextPC_in[26]), .Z(nextPC_out[26]) );
  BUF_X32 U66 ( .A(nextPC_in[25]), .Z(nextPC_out[25]) );
  BUF_X32 U67 ( .A(nextPC_in[24]), .Z(nextPC_out[24]) );
  BUF_X32 U68 ( .A(nextPC_in[23]), .Z(nextPC_out[23]) );
  BUF_X32 U69 ( .A(nextPC_in[22]), .Z(nextPC_out[22]) );
  BUF_X32 U70 ( .A(nextPC_in[21]), .Z(nextPC_out[21]) );
  BUF_X32 U71 ( .A(nextPC_in[20]), .Z(nextPC_out[20]) );
  BUF_X32 U72 ( .A(nextPC_in[19]), .Z(nextPC_out[19]) );
  BUF_X32 U73 ( .A(nextPC_in[18]), .Z(nextPC_out[18]) );
  BUF_X32 U74 ( .A(nextPC_in[17]), .Z(nextPC_out[17]) );
  BUF_X32 U75 ( .A(nextPC_in[16]), .Z(nextPC_out[16]) );
  BUF_X32 U76 ( .A(nextPC_in[15]), .Z(nextPC_out[15]) );
  BUF_X32 U77 ( .A(nextPC_in[14]), .Z(nextPC_out[14]) );
  BUF_X32 U78 ( .A(nextPC_in[13]), .Z(nextPC_out[13]) );
  BUF_X32 U79 ( .A(nextPC_in[12]), .Z(nextPC_out[12]) );
  BUF_X32 U80 ( .A(nextPC_in[11]), .Z(nextPC_out[11]) );
  BUF_X32 U81 ( .A(nextPC_in[10]), .Z(nextPC_out[10]) );
  BUF_X32 U82 ( .A(nextPC_in[9]), .Z(nextPC_out[9]) );
  BUF_X32 U83 ( .A(nextPC_in[8]), .Z(nextPC_out[8]) );
  BUF_X32 U84 ( .A(nextPC_in[7]), .Z(nextPC_out[7]) );
  BUF_X32 U85 ( .A(nextPC_in[6]), .Z(nextPC_out[6]) );
  BUF_X32 U86 ( .A(nextPC_in[5]), .Z(nextPC_out[5]) );
  BUF_X32 U87 ( .A(nextPC_in[4]), .Z(nextPC_out[4]) );
  BUF_X32 U88 ( .A(nextPC_in[3]), .Z(nextPC_out[3]) );
  BUF_X32 U89 ( .A(nextPC_in[2]), .Z(nextPC_out[2]) );
  BUF_X32 U90 ( .A(nextPC_in[1]), .Z(nextPC_out[1]) );
  BUF_X32 U91 ( .A(nextPC_in[0]), .Z(nextPC_out[0]) );
  BUF_X4 alu_ex_U4 ( .A(opB_in[31]), .Z(alu_ex_n4) );
  BUF_X4 alu_ex_U2 ( .A(opB_in[30]), .Z(alu_ex_n1) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_0__AND_1_U1 ( .A1(opB_in[0]), .A2(opA_in[0]), 
        .ZN(alu_ex_and_out_0_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_1__AND_1_U1 ( .A1(opB_in[1]), .A2(opA_in[1]), 
        .ZN(alu_ex_and_out_1_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_2__AND_1_U1 ( .A1(opB_in[2]), .A2(opA_in[2]), 
        .ZN(alu_ex_and_out_2_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_3__AND_1_U1 ( .A1(opB_in[3]), .A2(opA_in[3]), 
        .ZN(alu_ex_and_out_3_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_4__AND_1_U1 ( .A1(opB_in[4]), .A2(opA_in[4]), 
        .ZN(alu_ex_and_out_4_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_5__AND_1_U1 ( .A1(opB_in[5]), .A2(opA_in[5]), 
        .ZN(alu_ex_and_out_5_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_6__AND_1_U1 ( .A1(opB_in[6]), .A2(opA_in[6]), 
        .ZN(alu_ex_and_out_6_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_7__AND_1_U1 ( .A1(opB_in[7]), .A2(opA_in[7]), 
        .ZN(alu_ex_and_out_7_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_8__AND_1_U1 ( .A1(opB_in[8]), .A2(opA_in[8]), 
        .ZN(alu_ex_and_out_8_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_9__AND_1_U1 ( .A1(opB_in[9]), .A2(opA_in[9]), 
        .ZN(alu_ex_and_out_9_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_10__AND_1_U1 ( .A1(opB_in[10]), .A2(
        opA_in[10]), .ZN(alu_ex_and_out_10_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_11__AND_1_U1 ( .A1(opB_in[11]), .A2(
        opA_in[11]), .ZN(alu_ex_and_out_11_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_12__AND_1_U1 ( .A1(opB_in[12]), .A2(
        opA_in[12]), .ZN(alu_ex_and_out_12_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_13__AND_1_U1 ( .A1(opB_in[13]), .A2(
        opA_in[13]), .ZN(alu_ex_and_out_13_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_14__AND_1_U1 ( .A1(opB_in[14]), .A2(
        opA_in[14]), .ZN(alu_ex_and_out_14_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_15__AND_1_U1 ( .A1(opB_in[15]), .A2(
        opA_in[15]), .ZN(alu_ex_and_out_15_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_16__AND_1_U1 ( .A1(opB_in[16]), .A2(
        opA_in[16]), .ZN(alu_ex_and_out_16_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_17__AND_1_U1 ( .A1(opB_in[17]), .A2(
        opA_in[17]), .ZN(alu_ex_and_out_17_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_18__AND_1_U1 ( .A1(opB_in[18]), .A2(
        opA_in[18]), .ZN(alu_ex_and_out_18_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_19__AND_1_U1 ( .A1(opB_in[19]), .A2(
        opA_in[19]), .ZN(alu_ex_and_out_19_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_20__AND_1_U1 ( .A1(opB_in[20]), .A2(
        opA_in[20]), .ZN(alu_ex_and_out_20_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_21__AND_1_U1 ( .A1(opB_in[21]), .A2(
        opA_in[21]), .ZN(alu_ex_and_out_21_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_22__AND_1_U1 ( .A1(opB_in[22]), .A2(
        opA_in[22]), .ZN(alu_ex_and_out_22_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_23__AND_1_U1 ( .A1(opB_in[23]), .A2(
        opA_in[23]), .ZN(alu_ex_and_out_23_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_24__AND_1_U1 ( .A1(opB_in[24]), .A2(
        opA_in[24]), .ZN(alu_ex_and_out_24_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_25__AND_1_U1 ( .A1(opB_in[25]), .A2(
        opA_in[25]), .ZN(alu_ex_and_out_25_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_26__AND_1_U1 ( .A1(opB_in[26]), .A2(
        opA_in[26]), .ZN(alu_ex_and_out_26_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_27__AND_1_U1 ( .A1(opB_in[27]), .A2(
        opA_in[27]), .ZN(alu_ex_and_out_27_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_28__AND_1_U1 ( .A1(opB_in[28]), .A2(
        opA_in[28]), .ZN(alu_ex_and_out_28_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_29__AND_1_U1 ( .A1(opB_in[29]), .A2(
        opA_in[29]), .ZN(alu_ex_and_out_29_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_30__AND_1_U1 ( .A1(alu_ex_n1), .A2(
        opA_in[30]), .ZN(alu_ex_and_out_30_) );
  AND2_X2 alu_ex_AND_32_AND_32BIT_31__AND_1_U1 ( .A1(alu_ex_n4), .A2(
        opA_in[31]), .ZN(alu_ex_and_out_31_) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_0__OR_1_U1 ( .A1(opA_in[0]), .A2(opB_in[0]), 
        .ZN(alu_ex_or_out[0]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_1__OR_1_U1 ( .A1(opA_in[1]), .A2(opB_in[1]), 
        .ZN(alu_ex_or_out[1]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_2__OR_1_U1 ( .A1(opA_in[2]), .A2(opB_in[2]), 
        .ZN(alu_ex_or_out[2]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_3__OR_1_U1 ( .A1(opA_in[3]), .A2(opB_in[3]), 
        .ZN(alu_ex_or_out[3]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_4__OR_1_U1 ( .A1(opA_in[4]), .A2(opB_in[4]), 
        .ZN(alu_ex_or_out[4]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_5__OR_1_U1 ( .A1(opA_in[5]), .A2(opB_in[5]), 
        .ZN(alu_ex_or_out[5]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_6__OR_1_U1 ( .A1(opA_in[6]), .A2(opB_in[6]), 
        .ZN(alu_ex_or_out[6]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_7__OR_1_U1 ( .A1(opA_in[7]), .A2(opB_in[7]), 
        .ZN(alu_ex_or_out[7]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_8__OR_1_U1 ( .A1(opA_in[8]), .A2(opB_in[8]), 
        .ZN(alu_ex_or_out[8]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_9__OR_1_U1 ( .A1(opA_in[9]), .A2(opB_in[9]), 
        .ZN(alu_ex_or_out[9]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_10__OR_1_U1 ( .A1(opA_in[10]), .A2(opB_in[10]), 
        .ZN(alu_ex_or_out[10]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_11__OR_1_U1 ( .A1(opA_in[11]), .A2(opB_in[11]), 
        .ZN(alu_ex_or_out[11]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_12__OR_1_U1 ( .A1(opA_in[12]), .A2(opB_in[12]), 
        .ZN(alu_ex_or_out[12]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_13__OR_1_U1 ( .A1(opA_in[13]), .A2(opB_in[13]), 
        .ZN(alu_ex_or_out[13]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_14__OR_1_U1 ( .A1(opA_in[14]), .A2(opB_in[14]), 
        .ZN(alu_ex_or_out[14]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_15__OR_1_U1 ( .A1(opA_in[15]), .A2(opB_in[15]), 
        .ZN(alu_ex_or_out[15]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_16__OR_1_U1 ( .A1(opA_in[16]), .A2(opB_in[16]), 
        .ZN(alu_ex_or_out[16]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_17__OR_1_U1 ( .A1(opA_in[17]), .A2(opB_in[17]), 
        .ZN(alu_ex_or_out[17]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_18__OR_1_U1 ( .A1(opA_in[18]), .A2(opB_in[18]), 
        .ZN(alu_ex_or_out[18]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_19__OR_1_U1 ( .A1(opA_in[19]), .A2(opB_in[19]), 
        .ZN(alu_ex_or_out[19]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_20__OR_1_U1 ( .A1(opA_in[20]), .A2(opB_in[20]), 
        .ZN(alu_ex_or_out[20]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_21__OR_1_U1 ( .A1(opA_in[21]), .A2(opB_in[21]), 
        .ZN(alu_ex_or_out[21]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_22__OR_1_U1 ( .A1(opA_in[22]), .A2(opB_in[22]), 
        .ZN(alu_ex_or_out[22]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_23__OR_1_U1 ( .A1(opA_in[23]), .A2(opB_in[23]), 
        .ZN(alu_ex_or_out[23]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_24__OR_1_U1 ( .A1(opA_in[24]), .A2(opB_in[24]), 
        .ZN(alu_ex_or_out[24]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_25__OR_1_U1 ( .A1(opA_in[25]), .A2(opB_in[25]), 
        .ZN(alu_ex_or_out[25]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_26__OR_1_U1 ( .A1(opA_in[26]), .A2(opB_in[26]), 
        .ZN(alu_ex_or_out[26]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_27__OR_1_U1 ( .A1(opA_in[27]), .A2(opB_in[27]), 
        .ZN(alu_ex_or_out[27]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_28__OR_1_U1 ( .A1(opA_in[28]), .A2(opB_in[28]), 
        .ZN(alu_ex_or_out[28]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_29__OR_1_U1 ( .A1(opA_in[29]), .A2(opB_in[29]), 
        .ZN(alu_ex_or_out[29]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_30__OR_1_U1 ( .A1(opA_in[30]), .A2(alu_ex_n1), 
        .ZN(alu_ex_or_out[30]) );
  OR2_X2 alu_ex_OR_32_OR_32BIT_31__OR_1_U1 ( .A1(opA_in[31]), .A2(alu_ex_n4), 
        .ZN(alu_ex_or_out[31]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_0__XOR_1_U1 ( .A(opB_in[0]), .B(opA_in[0]), 
        .Z(alu_ex_xor_out[0]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_1__XOR_1_U1 ( .A(opB_in[1]), .B(opA_in[1]), 
        .Z(alu_ex_xor_out[1]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_2__XOR_1_U1 ( .A(opB_in[2]), .B(opA_in[2]), 
        .Z(alu_ex_xor_out[2]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_3__XOR_1_U1 ( .A(opB_in[3]), .B(opA_in[3]), 
        .Z(alu_ex_xor_out[3]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_4__XOR_1_U1 ( .A(opB_in[4]), .B(opA_in[4]), 
        .Z(alu_ex_xor_out[4]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_5__XOR_1_U1 ( .A(opB_in[5]), .B(opA_in[5]), 
        .Z(alu_ex_xor_out[5]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_6__XOR_1_U1 ( .A(opB_in[6]), .B(opA_in[6]), 
        .Z(alu_ex_xor_out[6]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_7__XOR_1_U1 ( .A(opB_in[7]), .B(opA_in[7]), 
        .Z(alu_ex_xor_out[7]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_8__XOR_1_U1 ( .A(opB_in[8]), .B(opA_in[8]), 
        .Z(alu_ex_xor_out[8]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_9__XOR_1_U1 ( .A(opB_in[9]), .B(opA_in[9]), 
        .Z(alu_ex_xor_out[9]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_10__XOR_1_U1 ( .A(opB_in[10]), .B(opA_in[10]), .Z(alu_ex_xor_out[10]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_11__XOR_1_U1 ( .A(opB_in[11]), .B(opA_in[11]), .Z(alu_ex_xor_out[11]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_12__XOR_1_U1 ( .A(opB_in[12]), .B(opA_in[12]), .Z(alu_ex_xor_out[12]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_13__XOR_1_U1 ( .A(opB_in[13]), .B(opA_in[13]), .Z(alu_ex_xor_out[13]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_14__XOR_1_U1 ( .A(opB_in[14]), .B(opA_in[14]), .Z(alu_ex_xor_out[14]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_15__XOR_1_U1 ( .A(opB_in[15]), .B(opA_in[15]), .Z(alu_ex_xor_out[15]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_16__XOR_1_U1 ( .A(opB_in[16]), .B(opA_in[16]), .Z(alu_ex_xor_out[16]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_17__XOR_1_U1 ( .A(opB_in[17]), .B(opA_in[17]), .Z(alu_ex_xor_out[17]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_18__XOR_1_U1 ( .A(opB_in[18]), .B(opA_in[18]), .Z(alu_ex_xor_out[18]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_19__XOR_1_U1 ( .A(opB_in[19]), .B(opA_in[19]), .Z(alu_ex_xor_out[19]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_20__XOR_1_U1 ( .A(opB_in[20]), .B(opA_in[20]), .Z(alu_ex_xor_out[20]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_21__XOR_1_U1 ( .A(opB_in[21]), .B(opA_in[21]), .Z(alu_ex_xor_out[21]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_22__XOR_1_U1 ( .A(opB_in[22]), .B(opA_in[22]), .Z(alu_ex_xor_out[22]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_23__XOR_1_U1 ( .A(opB_in[23]), .B(opA_in[23]), .Z(alu_ex_xor_out[23]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_24__XOR_1_U1 ( .A(opB_in[24]), .B(opA_in[24]), .Z(alu_ex_xor_out[24]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_25__XOR_1_U1 ( .A(opB_in[25]), .B(opA_in[25]), .Z(alu_ex_xor_out[25]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_26__XOR_1_U1 ( .A(opB_in[26]), .B(opA_in[26]), .Z(alu_ex_xor_out[26]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_27__XOR_1_U1 ( .A(opB_in[27]), .B(opA_in[27]), .Z(alu_ex_xor_out[27]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_28__XOR_1_U1 ( .A(opB_in[28]), .B(opA_in[28]), .Z(alu_ex_xor_out[28]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_29__XOR_1_U1 ( .A(opB_in[29]), .B(opA_in[29]), .Z(alu_ex_xor_out[29]) );
  XOR2_X1 alu_ex_XOR_32_XOR_32BIT_30__XOR_1_U1 ( .A(alu_ex_n1), .B(opA_in[30]), 
        .Z(alu_ex_xor_out[30]) );
  XOR2_X2 alu_ex_XOR_32_XOR_32BIT_31__XOR_1_U1 ( .A(alu_ex_n4), .B(opA_in[31]), 
        .Z(alu_ex_xor_out[31]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_0__NOT_1_U1 ( .A(opB_in[0]), .ZN(
        alu_ex_b_not[0]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_1__NOT_1_U1 ( .A(opB_in[1]), .ZN(
        alu_ex_b_not[1]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_2__NOT_1_U1 ( .A(opB_in[2]), .ZN(
        alu_ex_b_not[2]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_3__NOT_1_U1 ( .A(opB_in[3]), .ZN(
        alu_ex_b_not[3]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_4__NOT_1_U1 ( .A(opB_in[4]), .ZN(
        alu_ex_b_not[4]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_5__NOT_1_U1 ( .A(opB_in[5]), .ZN(
        alu_ex_b_not[5]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_6__NOT_1_U1 ( .A(opB_in[6]), .ZN(
        alu_ex_b_not[6]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_7__NOT_1_U1 ( .A(opB_in[7]), .ZN(
        alu_ex_b_not[7]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_8__NOT_1_U1 ( .A(opB_in[8]), .ZN(
        alu_ex_b_not[8]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_9__NOT_1_U1 ( .A(opB_in[9]), .ZN(
        alu_ex_b_not[9]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_10__NOT_1_U1 ( .A(opB_in[10]), .ZN(
        alu_ex_b_not[10]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_11__NOT_1_U1 ( .A(opB_in[11]), .ZN(
        alu_ex_b_not[11]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_12__NOT_1_U1 ( .A(opB_in[12]), .ZN(
        alu_ex_b_not[12]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_13__NOT_1_U1 ( .A(opB_in[13]), .ZN(
        alu_ex_b_not[13]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_14__NOT_1_U1 ( .A(opB_in[14]), .ZN(
        alu_ex_b_not[14]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_15__NOT_1_U1 ( .A(opB_in[15]), .ZN(
        alu_ex_b_not[15]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_16__NOT_1_U1 ( .A(opB_in[16]), .ZN(
        alu_ex_b_not[16]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_17__NOT_1_U1 ( .A(opB_in[17]), .ZN(
        alu_ex_b_not[17]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_18__NOT_1_U1 ( .A(opB_in[18]), .ZN(
        alu_ex_b_not[18]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_19__NOT_1_U1 ( .A(opB_in[19]), .ZN(
        alu_ex_b_not[19]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_20__NOT_1_U1 ( .A(opB_in[20]), .ZN(
        alu_ex_b_not[20]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_21__NOT_1_U1 ( .A(opB_in[21]), .ZN(
        alu_ex_b_not[21]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_22__NOT_1_U1 ( .A(opB_in[22]), .ZN(
        alu_ex_b_not[22]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_23__NOT_1_U1 ( .A(opB_in[23]), .ZN(
        alu_ex_b_not[23]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_24__NOT_1_U1 ( .A(opB_in[24]), .ZN(
        alu_ex_b_not[24]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_25__NOT_1_U1 ( .A(opB_in[25]), .ZN(
        alu_ex_b_not[25]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_26__NOT_1_U1 ( .A(opB_in[26]), .ZN(
        alu_ex_b_not[26]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_27__NOT_1_U1 ( .A(opB_in[27]), .ZN(
        alu_ex_b_not[27]) );
  INV_X1 alu_ex_NEGATE_B_NOT_32BIT_28__NOT_1_U1 ( .A(opB_in[28]), .ZN(
        alu_ex_b_not[28]) );
  INV_X1 alu_ex_NEGATE_B_NOT_32BIT_29__NOT_1_U1 ( .A(opB_in[29]), .ZN(
        alu_ex_b_not[29]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_30__NOT_1_U1 ( .A(opB_in[30]), .ZN(
        alu_ex_b_not[30]) );
  INV_X4 alu_ex_NEGATE_B_NOT_32BIT_31__NOT_1_U1 ( .A(opB_in[31]), .ZN(
        alu_ex_b_not[31]) );
  INV_X4 alu_ex_ADD_OR_SUB_U4 ( .A(alu_ex_ADD_OR_SUB_n4), .ZN(
        alu_ex_ADD_OR_SUB_n3) );
  INV_X4 alu_ex_ADD_OR_SUB_U3 ( .A(alu_ex_ADD_OR_SUB_n4), .ZN(
        alu_ex_ADD_OR_SUB_n2) );
  INV_X4 alu_ex_ADD_OR_SUB_U2 ( .A(alu_ex_ADD_OR_SUB_n4), .ZN(
        alu_ex_ADD_OR_SUB_n1) );
  INV_X4 alu_ex_ADD_OR_SUB_U1 ( .A(ALUCtrl_in[3]), .ZN(alu_ex_ADD_OR_SUB_n4)
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_0__MUX_U3 ( .A(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_0__MUX_n4), .ZN(alu_ex_add_sub_in[0])
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_0__MUX_U2 ( .A(alu_ex_ADD_OR_SUB_n3), 
        .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_0__MUX_U1 ( .A1(opB_in[0]), .A2(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_0__MUX_n1), .B1(alu_ex_b_not[0]), .B2(
        alu_ex_ADD_OR_SUB_n3), .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_0__MUX_n4)
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_1__MUX_n4), .ZN(alu_ex_add_sub_in[1])
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_1__MUX_U2 ( .A(alu_ex_ADD_OR_SUB_n2), 
        .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_1__MUX_U1 ( .A1(opB_in[1]), .A2(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_1__MUX_n1), .B1(alu_ex_b_not[1]), .B2(
        alu_ex_ADD_OR_SUB_n2), .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_1__MUX_n4)
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_2__MUX_U3 ( .A(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_2__MUX_n4), .ZN(alu_ex_add_sub_in[2])
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_2__MUX_U2 ( .A(alu_ex_ADD_OR_SUB_n1), 
        .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_2__MUX_U1 ( .A1(opB_in[2]), .A2(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_2__MUX_n1), .B1(alu_ex_b_not[2]), .B2(
        alu_ex_ADD_OR_SUB_n1), .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_2__MUX_n4)
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_3__MUX_U3 ( .A(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_3__MUX_n4), .ZN(alu_ex_add_sub_in[3])
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_3__MUX_U2 ( .A(alu_ex_ADD_OR_SUB_n3), 
        .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_3__MUX_U1 ( .A1(opB_in[3]), .A2(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_3__MUX_n1), .B1(alu_ex_b_not[3]), .B2(
        alu_ex_ADD_OR_SUB_n3), .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_3__MUX_n4)
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_4__MUX_U3 ( .A(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_4__MUX_n4), .ZN(alu_ex_add_sub_in[4])
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_4__MUX_U2 ( .A(alu_ex_ADD_OR_SUB_n2), 
        .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_4__MUX_U1 ( .A1(opB_in[4]), .A2(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_4__MUX_n1), .B1(alu_ex_b_not[4]), .B2(
        alu_ex_ADD_OR_SUB_n2), .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_4__MUX_n4)
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_5__MUX_U3 ( .A(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_5__MUX_n4), .ZN(alu_ex_add_sub_in[5])
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_5__MUX_U2 ( .A(alu_ex_ADD_OR_SUB_n1), 
        .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_5__MUX_U1 ( .A1(opB_in[5]), .A2(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_5__MUX_n1), .B1(alu_ex_b_not[5]), .B2(
        alu_ex_ADD_OR_SUB_n1), .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_5__MUX_n4)
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_6__MUX_U3 ( .A(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_6__MUX_n4), .ZN(alu_ex_add_sub_in[6])
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_6__MUX_U2 ( .A(alu_ex_ADD_OR_SUB_n3), 
        .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_6__MUX_U1 ( .A1(opB_in[6]), .A2(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_6__MUX_n1), .B1(alu_ex_b_not[6]), .B2(
        alu_ex_ADD_OR_SUB_n3), .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_6__MUX_n4)
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_7__MUX_U3 ( .A(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_7__MUX_n4), .ZN(alu_ex_add_sub_in[7])
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_7__MUX_U2 ( .A(alu_ex_ADD_OR_SUB_n2), 
        .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_7__MUX_U1 ( .A1(opB_in[7]), .A2(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_7__MUX_n1), .B1(alu_ex_b_not[7]), .B2(
        alu_ex_ADD_OR_SUB_n2), .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_7__MUX_n4)
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_8__MUX_U3 ( .A(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_8__MUX_n4), .ZN(alu_ex_add_sub_in[8])
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_8__MUX_U2 ( .A(alu_ex_ADD_OR_SUB_n1), 
        .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_8__MUX_U1 ( .A1(opB_in[8]), .A2(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_8__MUX_n1), .B1(alu_ex_b_not[8]), .B2(
        alu_ex_ADD_OR_SUB_n1), .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_8__MUX_n4)
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_9__MUX_U3 ( .A(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_9__MUX_n4), .ZN(alu_ex_add_sub_in[9])
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_9__MUX_U2 ( .A(alu_ex_ADD_OR_SUB_n3), 
        .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_9__MUX_U1 ( .A1(opB_in[9]), .A2(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_9__MUX_n1), .B1(alu_ex_b_not[9]), .B2(
        alu_ex_ADD_OR_SUB_n3), .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_9__MUX_n4)
         );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_10__MUX_U3 ( .A(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_10__MUX_n4), .ZN(alu_ex_add_sub_in[10]) );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_10__MUX_U2 ( .A(alu_ex_ADD_OR_SUB_n2), 
        .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_10__MUX_n1) );
  AOI22_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_10__MUX_U1 ( .A1(opB_in[10]), .A2(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_10__MUX_n1), .B1(alu_ex_b_not[10]), 
        .B2(alu_ex_ADD_OR_SUB_n2), .ZN(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_10__MUX_n4) );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_11__MUX_U3 ( .A(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_11__MUX_n4), .ZN(alu_ex_add_sub_in[11]) );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_11__MUX_U2 ( .A(alu_ex_ADD_OR_SUB_n1), 
        .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_11__MUX_n1) );
  AOI22_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_11__MUX_U1 ( .A1(opB_in[11]), .A2(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_11__MUX_n1), .B1(alu_ex_b_not[11]), 
        .B2(alu_ex_ADD_OR_SUB_n1), .ZN(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_11__MUX_n4) );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_12__MUX_U3 ( .A(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_12__MUX_n4), .ZN(alu_ex_add_sub_in[12]) );
  INV_X1 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_12__MUX_U2 ( .A(alu_ex_ADD_OR_SUB_n3), 
        .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_12__MUX_n1) );
  AOI22_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_12__MUX_U1 ( .A1(opB_in[12]), .A2(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_12__MUX_n1), .B1(alu_ex_b_not[12]), 
        .B2(alu_ex_ADD_OR_SUB_n3), .ZN(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_12__MUX_n4) );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_13__MUX_U1 ( .A(opB_in[13]), .B(
        alu_ex_b_not[13]), .S(alu_ex_ADD_OR_SUB_n3), .Z(alu_ex_add_sub_in[13])
         );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_14__MUX_U1 ( .A(opB_in[14]), .B(
        alu_ex_b_not[14]), .S(alu_ex_ADD_OR_SUB_n2), .Z(alu_ex_add_sub_in[14])
         );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_15__MUX_U1 ( .A(opB_in[15]), .B(
        alu_ex_b_not[15]), .S(alu_ex_ADD_OR_SUB_n1), .Z(alu_ex_add_sub_in[15])
         );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_16__MUX_U1 ( .A(opB_in[16]), .B(
        alu_ex_b_not[16]), .S(ALUCtrl_in[3]), .Z(alu_ex_add_sub_in[16]) );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_17__MUX_U1 ( .A(opB_in[17]), .B(
        alu_ex_b_not[17]), .S(ALUCtrl_in[3]), .Z(alu_ex_add_sub_in[17]) );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_18__MUX_U1 ( .A(opB_in[18]), .B(
        alu_ex_b_not[18]), .S(ALUCtrl_in[3]), .Z(alu_ex_add_sub_in[18]) );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_19__MUX_U1 ( .A(opB_in[19]), .B(
        alu_ex_b_not[19]), .S(ALUCtrl_in[3]), .Z(alu_ex_add_sub_in[19]) );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_20__MUX_U1 ( .A(opB_in[20]), .B(
        alu_ex_b_not[20]), .S(ALUCtrl_in[3]), .Z(alu_ex_add_sub_in[20]) );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_21__MUX_U1 ( .A(opB_in[21]), .B(
        alu_ex_b_not[21]), .S(ALUCtrl_in[3]), .Z(alu_ex_add_sub_in[21]) );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_22__MUX_U1 ( .A(opB_in[22]), .B(
        alu_ex_b_not[22]), .S(ALUCtrl_in[3]), .Z(alu_ex_add_sub_in[22]) );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_23__MUX_U1 ( .A(opB_in[23]), .B(
        alu_ex_b_not[23]), .S(ALUCtrl_in[3]), .Z(alu_ex_add_sub_in[23]) );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_24__MUX_U1 ( .A(opB_in[24]), .B(
        alu_ex_b_not[24]), .S(ALUCtrl_in[3]), .Z(alu_ex_add_sub_in[24]) );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_25__MUX_U1 ( .A(opB_in[25]), .B(
        alu_ex_b_not[25]), .S(ALUCtrl_in[3]), .Z(alu_ex_add_sub_in[25]) );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_26__MUX_U1 ( .A(opB_in[26]), .B(
        alu_ex_b_not[26]), .S(ALUCtrl_in[3]), .Z(alu_ex_add_sub_in[26]) );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_27__MUX_U1 ( .A(opB_in[27]), .B(
        alu_ex_b_not[27]), .S(ALUCtrl_in[3]), .Z(alu_ex_add_sub_in[27]) );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_28__MUX_U1 ( .A(opB_in[28]), .B(
        alu_ex_b_not[28]), .S(ALUCtrl_in[3]), .Z(alu_ex_add_sub_in[28]) );
  MUX2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_29__MUX_U1 ( .A(opB_in[29]), .B(
        alu_ex_b_not[29]), .S(ALUCtrl_in[3]), .Z(alu_ex_add_sub_in[29]) );
  NAND2_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_30__MUX_U4 ( .A1(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_30__MUX_n2), .A2(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_30__MUX_n3), .ZN(alu_ex_add_sub_in[30]) );
  NAND2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_30__MUX_U3 ( .A1(alu_ex_b_not[30]), 
        .A2(ALUCtrl_in[3]), .ZN(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_30__MUX_n3) );
  INV_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_30__MUX_U2 ( .A(ALUCtrl_in[3]), .ZN(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_30__MUX_n1) );
  NAND2_X2 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_30__MUX_U1 ( .A1(opB_in[30]), .A2(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_30__MUX_n1), .ZN(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_30__MUX_n2) );
  OAI21_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_31__MUX_U3 ( .B1(alu_ex_b_not[31]), 
        .B2(ALUCtrl_in[3]), .A(alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_31__MUX_n3), 
        .ZN(alu_ex_add_sub_in[31]) );
  NAND2_X4 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_31__MUX_U2 ( .A1(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_31__MUX_n2), .A2(ALUCtrl_in[3]), .ZN(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_31__MUX_n3) );
  INV_X16 alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_31__MUX_U1 ( .A(opB_in[31]), .ZN(
        alu_ex_ADD_OR_SUB_MUX2TO1_32BIT_31__MUX_n2) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_0__FA_U2 ( .A(alu_ex_FULL_ADDER_carry[1]), 
        .B(alu_ex_FULL_ADDER_FA_NBIT_0__FA_n1), .ZN(alu_ex_add_sub_out_0_) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_0__FA_U1 ( .A(alu_ex_add_sub_in[0]), .B(
        opA_in[0]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_0__FA_n1) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_1__FA_U6 ( .A(alu_ex_FULL_ADDER_carry[2]), 
        .B(alu_ex_FULL_ADDER_FA_NBIT_1__FA_n4), .ZN(alu_ex_add_sub_out_1_) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_1__FA_U5 ( .A1(alu_ex_add_sub_in[1]), 
        .A2(opA_in[1]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_1__FA_n2) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_1__FA_U4 ( .A1(alu_ex_FULL_ADDER_carry[2]), .A2(alu_ex_FULL_ADDER_FA_NBIT_1__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_1__FA_n3) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_1__FA_U3 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_1__FA_n4), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_1__FA_n1) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_1__FA_U2 ( .A(alu_ex_add_sub_in[1]), .B(
        opA_in[1]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_1__FA_n4) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_1__FA_U1 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_1__FA_n3), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_1__FA_n2), .ZN(alu_ex_FULL_ADDER_carry[1])
         );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_2__FA_U6 ( .A(alu_ex_FULL_ADDER_carry[3]), 
        .B(alu_ex_FULL_ADDER_FA_NBIT_2__FA_n4), .ZN(alu_ex_add_sub_out_2_) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_2__FA_U5 ( .A1(alu_ex_add_sub_in[2]), 
        .A2(opA_in[2]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_2__FA_n2) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_2__FA_U4 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_2__FA_n4), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_2__FA_n1) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_2__FA_U3 ( .A(alu_ex_add_sub_in[2]), .B(
        opA_in[2]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_2__FA_n4) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_2__FA_U2 ( .A1(alu_ex_FULL_ADDER_carry[3]), .A2(alu_ex_FULL_ADDER_FA_NBIT_2__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_2__FA_n3) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_2__FA_U1 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_2__FA_n3), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_2__FA_n2), .ZN(alu_ex_FULL_ADDER_carry[2])
         );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_3__FA_U6 ( .A(alu_ex_FULL_ADDER_carry[4]), 
        .B(alu_ex_FULL_ADDER_FA_NBIT_3__FA_n4), .ZN(alu_ex_add_sub_out_3_) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_3__FA_U5 ( .A1(alu_ex_add_sub_in[3]), 
        .A2(opA_in[3]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_3__FA_n2) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_3__FA_U4 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_3__FA_n4), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_3__FA_n1) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_3__FA_U3 ( .A(alu_ex_add_sub_in[3]), .B(
        opA_in[3]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_3__FA_n4) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_3__FA_U2 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_3__FA_n3), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_3__FA_n2), .ZN(alu_ex_FULL_ADDER_carry[3])
         );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_3__FA_U1 ( .A1(alu_ex_FULL_ADDER_carry[4]), .A2(alu_ex_FULL_ADDER_FA_NBIT_3__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_3__FA_n3) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_4__FA_U6 ( .A1(alu_ex_add_sub_in[4]), 
        .A2(opA_in[4]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_4__FA_n2) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_4__FA_U5 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_4__FA_n4), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_4__FA_n1) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_4__FA_U4 ( .A(alu_ex_add_sub_in[4]), .B(
        opA_in[4]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_4__FA_n4) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_4__FA_U3 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_4__FA_n3), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_4__FA_n2), .ZN(alu_ex_FULL_ADDER_carry[4])
         );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_4__FA_U2 ( .A1(alu_ex_FULL_ADDER_carry[5]), .A2(alu_ex_FULL_ADDER_FA_NBIT_4__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_4__FA_n3) );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_4__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[5]), 
        .B(alu_ex_FULL_ADDER_FA_NBIT_4__FA_n4), .ZN(alu_ex_add_sub_out_4_) );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_5__FA_U2 ( .A(alu_ex_FULL_ADDER_carry[6]), 
        .B(alu_ex_FULL_ADDER_FA_NBIT_5__FA_n6), .ZN(alu_ex_add_sub_out_5_) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_5__FA_U8 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_5__FA_n6), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_5__FA_n5) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_5__FA_U7 ( .A(alu_ex_add_sub_in[5]), .B(
        opA_in[5]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_5__FA_n6) );
  INV_X8 alu_ex_FULL_ADDER_FA_NBIT_5__FA_U6 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_5__FA_n4), .ZN(alu_ex_FULL_ADDER_carry[5])
         );
  AOI21_X4 alu_ex_FULL_ADDER_FA_NBIT_5__FA_U5 ( .B1(alu_ex_FULL_ADDER_carry[6]), .B2(alu_ex_FULL_ADDER_FA_NBIT_5__FA_n5), .A(
        alu_ex_FULL_ADDER_FA_NBIT_5__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_5__FA_n4) );
  AND2_X4 alu_ex_FULL_ADDER_FA_NBIT_5__FA_U1 ( .A1(alu_ex_add_sub_in[5]), .A2(
        opA_in[5]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_5__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_6__FA_U8 ( .A1(alu_ex_add_sub_in[6]), 
        .A2(opA_in[6]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_6__FA_n4) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_6__FA_U7 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_6__FA_n6), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_6__FA_n3) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_6__FA_U6 ( .A(alu_ex_add_sub_in[6]), .B(
        opA_in[6]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_6__FA_n6) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_6__FA_U5 ( .A1(alu_ex_FULL_ADDER_carry[7]), .A2(alu_ex_FULL_ADDER_FA_NBIT_6__FA_n3), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_6__FA_n5) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_6__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_6__FA_n5), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_6__FA_n4), .ZN(alu_ex_FULL_ADDER_carry[6])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_6__FA_U3 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_6__FA_n2), .B(
        alu_ex_FULL_ADDER_FA_NBIT_6__FA_n6), .ZN(alu_ex_add_sub_out_6_) );
  INV_X2 alu_ex_FULL_ADDER_FA_NBIT_6__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_6__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_6__FA_n2) );
  INV_X1 alu_ex_FULL_ADDER_FA_NBIT_6__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[7]), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_6__FA_n1) );
  BUF_X8 alu_ex_FULL_ADDER_FA_NBIT_7__FA_U9 ( .A(alu_ex_FULL_ADDER_carry[8]), 
        .Z(alu_ex_FULL_ADDER_FA_NBIT_7__FA_n8) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_7__FA_U8 ( .A1(alu_ex_add_sub_in[7]), 
        .A2(opA_in[7]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_7__FA_n4) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_7__FA_U7 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_7__FA_n6), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_7__FA_n3) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_7__FA_U6 ( .A(alu_ex_add_sub_in[7]), .B(
        opA_in[7]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_7__FA_n6) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_7__FA_U5 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_7__FA_n5), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_7__FA_n4), .ZN(alu_ex_FULL_ADDER_carry[7])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_7__FA_U4 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_7__FA_n2), .B(
        alu_ex_FULL_ADDER_FA_NBIT_7__FA_n6), .ZN(alu_ex_add_sub_out_7_) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_7__FA_U3 ( .A1(alu_ex_FULL_ADDER_carry[8]), .A2(alu_ex_FULL_ADDER_FA_NBIT_7__FA_n3), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_7__FA_n5) );
  INV_X2 alu_ex_FULL_ADDER_FA_NBIT_7__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_7__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_7__FA_n2) );
  INV_X1 alu_ex_FULL_ADDER_FA_NBIT_7__FA_U1 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_7__FA_n8), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_7__FA_n1) );
  BUF_X16 alu_ex_FULL_ADDER_FA_NBIT_8__FA_U9 ( .A(alu_ex_FULL_ADDER_carry[9]), 
        .Z(alu_ex_FULL_ADDER_FA_NBIT_8__FA_n8) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_8__FA_U8 ( .A1(alu_ex_add_sub_in[8]), 
        .A2(opA_in[8]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_8__FA_n4) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_8__FA_U7 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_8__FA_n6), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_8__FA_n3) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_8__FA_U6 ( .A(alu_ex_add_sub_in[8]), .B(
        opA_in[8]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_8__FA_n6) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_8__FA_U5 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_8__FA_n5), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_8__FA_n4), .ZN(alu_ex_FULL_ADDER_carry[8])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_8__FA_U4 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_8__FA_n2), .B(
        alu_ex_FULL_ADDER_FA_NBIT_8__FA_n6), .ZN(alu_ex_add_sub_out_8_) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_8__FA_U3 ( .A1(alu_ex_FULL_ADDER_carry[9]), .A2(alu_ex_FULL_ADDER_FA_NBIT_8__FA_n3), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_8__FA_n5) );
  INV_X2 alu_ex_FULL_ADDER_FA_NBIT_8__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_8__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_8__FA_n2) );
  INV_X1 alu_ex_FULL_ADDER_FA_NBIT_8__FA_U1 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_8__FA_n8), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_8__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_9__FA_U8 ( .A1(alu_ex_add_sub_in[9]), 
        .A2(opA_in[9]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_9__FA_n4) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_9__FA_U7 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_9__FA_n6), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_9__FA_n3) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_9__FA_U6 ( .A(alu_ex_add_sub_in[9]), .B(
        opA_in[9]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_9__FA_n6) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_9__FA_U5 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_9__FA_n5), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_9__FA_n4), .ZN(alu_ex_FULL_ADDER_carry[9])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_9__FA_U4 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_9__FA_n2), .B(
        alu_ex_FULL_ADDER_FA_NBIT_9__FA_n6), .ZN(alu_ex_add_sub_out_9_) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_9__FA_U3 ( .A1(
        alu_ex_FULL_ADDER_carry[10]), .A2(alu_ex_FULL_ADDER_FA_NBIT_9__FA_n3), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_9__FA_n5) );
  INV_X2 alu_ex_FULL_ADDER_FA_NBIT_9__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_9__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_9__FA_n2) );
  INV_X1 alu_ex_FULL_ADDER_FA_NBIT_9__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[10]), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_9__FA_n1) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_10__FA_U9 ( .A(alu_ex_FULL_ADDER_carry[11]), .Z(alu_ex_FULL_ADDER_FA_NBIT_10__FA_n8) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_10__FA_U8 ( .A1(alu_ex_add_sub_in[10]), 
        .A2(opA_in[10]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_10__FA_n4) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_10__FA_U7 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_10__FA_n6), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_10__FA_n3) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_10__FA_U6 ( .A(alu_ex_add_sub_in[10]), 
        .B(opA_in[10]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_10__FA_n6) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_10__FA_U5 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_10__FA_n5), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_10__FA_n4), .ZN(alu_ex_FULL_ADDER_carry[10])
         );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_10__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_carry[11]), .A2(alu_ex_FULL_ADDER_FA_NBIT_10__FA_n3), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_10__FA_n5) );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_10__FA_U3 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_10__FA_n2), .B(
        alu_ex_FULL_ADDER_FA_NBIT_10__FA_n6), .ZN(alu_ex_add_sub_out_10_) );
  INV_X2 alu_ex_FULL_ADDER_FA_NBIT_10__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_10__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_10__FA_n2) );
  INV_X1 alu_ex_FULL_ADDER_FA_NBIT_10__FA_U1 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_10__FA_n8), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_10__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_11__FA_U7 ( .A1(alu_ex_add_sub_in[11]), 
        .A2(opA_in[11]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_11__FA_n3) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_11__FA_U6 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_11__FA_n5), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_11__FA_n2) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_11__FA_U5 ( .A(alu_ex_add_sub_in[11]), 
        .B(opA_in[11]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_11__FA_n5) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_11__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_carry[12]), .A2(alu_ex_FULL_ADDER_FA_NBIT_11__FA_n2), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_11__FA_n4) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_11__FA_U3 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_11__FA_n4), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_11__FA_n3), .ZN(alu_ex_FULL_ADDER_carry[11])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_11__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_11__FA_n1), .B(
        alu_ex_FULL_ADDER_FA_NBIT_11__FA_n5), .ZN(alu_ex_add_sub_out_11_) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_11__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[12]), .Z(alu_ex_FULL_ADDER_FA_NBIT_11__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_12__FA_U7 ( .A1(alu_ex_add_sub_in[12]), 
        .A2(opA_in[12]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_12__FA_n3) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_12__FA_U6 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_12__FA_n5), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_12__FA_n2) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_12__FA_U5 ( .A(alu_ex_add_sub_in[12]), 
        .B(opA_in[12]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_12__FA_n5) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_12__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_12__FA_n4), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_12__FA_n3), .ZN(alu_ex_FULL_ADDER_carry[12])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_12__FA_U3 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_12__FA_n1), .B(
        alu_ex_FULL_ADDER_FA_NBIT_12__FA_n5), .ZN(alu_ex_add_sub_out_12_) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_12__FA_U2 ( .A1(
        alu_ex_FULL_ADDER_carry[13]), .A2(alu_ex_FULL_ADDER_FA_NBIT_12__FA_n2), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_12__FA_n4) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_12__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[13]), .Z(alu_ex_FULL_ADDER_FA_NBIT_12__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_13__FA_U7 ( .A1(alu_ex_add_sub_in[13]), 
        .A2(opA_in[13]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_13__FA_n3) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_13__FA_U6 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_13__FA_n5), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_13__FA_n2) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_13__FA_U5 ( .A(alu_ex_add_sub_in[13]), 
        .B(opA_in[13]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_13__FA_n5) );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_13__FA_U4 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_13__FA_n1), .B(
        alu_ex_FULL_ADDER_FA_NBIT_13__FA_n5), .ZN(alu_ex_add_sub_out_13_) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_13__FA_U3 ( .A1(
        alu_ex_FULL_ADDER_carry[14]), .A2(alu_ex_FULL_ADDER_FA_NBIT_13__FA_n2), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_13__FA_n4) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_13__FA_U2 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_13__FA_n4), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_13__FA_n3), .ZN(alu_ex_FULL_ADDER_carry[13])
         );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_13__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[14]), .Z(alu_ex_FULL_ADDER_FA_NBIT_13__FA_n1) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_14__FA_U9 ( .A(alu_ex_FULL_ADDER_carry[15]), .Z(alu_ex_FULL_ADDER_FA_NBIT_14__FA_n8) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_14__FA_U8 ( .A1(alu_ex_add_sub_in[14]), 
        .A2(opA_in[14]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_14__FA_n4) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_14__FA_U7 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_14__FA_n6), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_14__FA_n3) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_14__FA_U6 ( .A(alu_ex_add_sub_in[14]), 
        .B(opA_in[14]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_14__FA_n6) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_14__FA_U5 ( .A1(
        alu_ex_FULL_ADDER_carry[15]), .A2(alu_ex_FULL_ADDER_FA_NBIT_14__FA_n3), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_14__FA_n5) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_14__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_14__FA_n5), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_14__FA_n4), .ZN(alu_ex_FULL_ADDER_carry[14])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_14__FA_U3 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_14__FA_n2), .B(
        alu_ex_FULL_ADDER_FA_NBIT_14__FA_n6), .ZN(alu_ex_add_sub_out_14_) );
  INV_X2 alu_ex_FULL_ADDER_FA_NBIT_14__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_14__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_14__FA_n2) );
  INV_X1 alu_ex_FULL_ADDER_FA_NBIT_14__FA_U1 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_14__FA_n8), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_14__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_15__FA_U7 ( .A1(alu_ex_add_sub_in[15]), 
        .A2(opA_in[15]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_15__FA_n3) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_15__FA_U6 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_15__FA_n5), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_15__FA_n2) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_15__FA_U5 ( .A(alu_ex_add_sub_in[15]), 
        .B(opA_in[15]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_15__FA_n5) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_15__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_carry[16]), .A2(alu_ex_FULL_ADDER_FA_NBIT_15__FA_n2), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_15__FA_n4) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_15__FA_U3 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_15__FA_n4), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_15__FA_n3), .ZN(alu_ex_FULL_ADDER_carry[15])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_15__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_15__FA_n1), .B(
        alu_ex_FULL_ADDER_FA_NBIT_15__FA_n5), .ZN(alu_ex_add_sub_out_15_) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_15__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[16]), .Z(alu_ex_FULL_ADDER_FA_NBIT_15__FA_n1) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_16__FA_U9 ( .A(alu_ex_FULL_ADDER_carry[17]), .Z(alu_ex_FULL_ADDER_FA_NBIT_16__FA_n8) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_16__FA_U8 ( .A1(alu_ex_add_sub_in[16]), 
        .A2(opA_in[16]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_16__FA_n4) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_16__FA_U7 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_16__FA_n6), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_16__FA_n3) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_16__FA_U6 ( .A(alu_ex_add_sub_in[16]), 
        .B(opA_in[16]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_16__FA_n6) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_16__FA_U5 ( .A1(
        alu_ex_FULL_ADDER_carry[17]), .A2(alu_ex_FULL_ADDER_FA_NBIT_16__FA_n3), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_16__FA_n5) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_16__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_16__FA_n5), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_16__FA_n4), .ZN(alu_ex_FULL_ADDER_carry[16])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_16__FA_U3 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_16__FA_n2), .B(
        alu_ex_FULL_ADDER_FA_NBIT_16__FA_n6), .ZN(alu_ex_add_sub_out_16_) );
  INV_X2 alu_ex_FULL_ADDER_FA_NBIT_16__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_16__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_16__FA_n2) );
  INV_X1 alu_ex_FULL_ADDER_FA_NBIT_16__FA_U1 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_16__FA_n8), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_16__FA_n1) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_17__FA_U9 ( .A(alu_ex_FULL_ADDER_carry[18]), .Z(alu_ex_FULL_ADDER_FA_NBIT_17__FA_n8) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_17__FA_U8 ( .A1(alu_ex_add_sub_in[17]), 
        .A2(opA_in[17]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_17__FA_n4) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_17__FA_U7 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_17__FA_n6), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_17__FA_n3) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_17__FA_U6 ( .A(alu_ex_add_sub_in[17]), 
        .B(opA_in[17]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_17__FA_n6) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_17__FA_U5 ( .A1(
        alu_ex_FULL_ADDER_carry[18]), .A2(alu_ex_FULL_ADDER_FA_NBIT_17__FA_n3), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_17__FA_n5) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_17__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_17__FA_n5), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_17__FA_n4), .ZN(alu_ex_FULL_ADDER_carry[17])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_17__FA_U3 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_17__FA_n2), .B(
        alu_ex_FULL_ADDER_FA_NBIT_17__FA_n6), .ZN(alu_ex_add_sub_out_17_) );
  INV_X2 alu_ex_FULL_ADDER_FA_NBIT_17__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_17__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_17__FA_n2) );
  INV_X1 alu_ex_FULL_ADDER_FA_NBIT_17__FA_U1 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_17__FA_n8), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_17__FA_n1) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_18__FA_U9 ( .A(alu_ex_FULL_ADDER_carry[19]), .Z(alu_ex_FULL_ADDER_FA_NBIT_18__FA_n8) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_18__FA_U8 ( .A1(alu_ex_add_sub_in[18]), 
        .A2(opA_in[18]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_18__FA_n4) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_18__FA_U7 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_18__FA_n6), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_18__FA_n3) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_18__FA_U6 ( .A(alu_ex_add_sub_in[18]), 
        .B(opA_in[18]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_18__FA_n6) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_18__FA_U5 ( .A1(
        alu_ex_FULL_ADDER_carry[19]), .A2(alu_ex_FULL_ADDER_FA_NBIT_18__FA_n3), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_18__FA_n5) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_18__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_18__FA_n5), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_18__FA_n4), .ZN(alu_ex_FULL_ADDER_carry[18])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_18__FA_U3 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_18__FA_n2), .B(
        alu_ex_FULL_ADDER_FA_NBIT_18__FA_n6), .ZN(alu_ex_add_sub_out_18_) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_18__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_18__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_18__FA_n2) );
  INV_X1 alu_ex_FULL_ADDER_FA_NBIT_18__FA_U1 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_18__FA_n8), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_18__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_19__FA_U7 ( .A1(alu_ex_add_sub_in[19]), 
        .A2(opA_in[19]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_19__FA_n3) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_19__FA_U6 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_19__FA_n5), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_19__FA_n2) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_19__FA_U5 ( .A(alu_ex_add_sub_in[19]), 
        .B(opA_in[19]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_19__FA_n5) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_19__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_19__FA_n4), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_19__FA_n3), .ZN(alu_ex_FULL_ADDER_carry[19])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_19__FA_U3 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_19__FA_n1), .B(
        alu_ex_FULL_ADDER_FA_NBIT_19__FA_n5), .ZN(alu_ex_add_sub_out_19_) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_19__FA_U2 ( .A1(
        alu_ex_FULL_ADDER_carry[20]), .A2(alu_ex_FULL_ADDER_FA_NBIT_19__FA_n2), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_19__FA_n4) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_19__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[20]), .Z(alu_ex_FULL_ADDER_FA_NBIT_19__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_20__FA_U7 ( .A1(alu_ex_add_sub_in[20]), 
        .A2(opA_in[20]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_20__FA_n3) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_20__FA_U6 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_20__FA_n5), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_20__FA_n2) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_20__FA_U5 ( .A(alu_ex_add_sub_in[20]), 
        .B(opA_in[20]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_20__FA_n5) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_20__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_20__FA_n4), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_20__FA_n3), .ZN(alu_ex_FULL_ADDER_carry[20])
         );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_20__FA_U3 ( .A1(
        alu_ex_FULL_ADDER_carry[21]), .A2(alu_ex_FULL_ADDER_FA_NBIT_20__FA_n2), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_20__FA_n4) );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_20__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_20__FA_n1), .B(
        alu_ex_FULL_ADDER_FA_NBIT_20__FA_n5), .ZN(alu_ex_add_sub_out_20_) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_20__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[21]), .Z(alu_ex_FULL_ADDER_FA_NBIT_20__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_21__FA_U9 ( .A1(alu_ex_add_sub_in[21]), 
        .A2(opA_in[21]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_21__FA_n5) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_21__FA_U8 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_21__FA_n7), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_21__FA_n4) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_21__FA_U7 ( .A(alu_ex_add_sub_in[21]), 
        .B(opA_in[21]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_21__FA_n7) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_21__FA_U6 ( .A1(
        alu_ex_FULL_ADDER_carry[22]), .A2(alu_ex_FULL_ADDER_FA_NBIT_21__FA_n4), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_21__FA_n6) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_21__FA_U5 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_21__FA_n6), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_21__FA_n5), .ZN(alu_ex_FULL_ADDER_carry[21])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_21__FA_U4 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_21__FA_n3), .B(
        alu_ex_FULL_ADDER_FA_NBIT_21__FA_n7), .ZN(alu_ex_add_sub_out_21_) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_21__FA_U3 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_21__FA_n2), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_21__FA_n3) );
  INV_X1 alu_ex_FULL_ADDER_FA_NBIT_21__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_21__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_21__FA_n2) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_21__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[22]), .Z(alu_ex_FULL_ADDER_FA_NBIT_21__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_22__FA_U7 ( .A1(alu_ex_add_sub_in[22]), 
        .A2(opA_in[22]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_22__FA_n3) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_22__FA_U6 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_22__FA_n5), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_22__FA_n2) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_22__FA_U5 ( .A(alu_ex_add_sub_in[22]), 
        .B(opA_in[22]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_22__FA_n5) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_22__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_22__FA_n4), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_22__FA_n3), .ZN(alu_ex_FULL_ADDER_carry[22])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_22__FA_U3 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_22__FA_n1), .B(
        alu_ex_FULL_ADDER_FA_NBIT_22__FA_n5), .ZN(alu_ex_add_sub_out_22_) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_22__FA_U2 ( .A1(
        alu_ex_FULL_ADDER_carry[23]), .A2(alu_ex_FULL_ADDER_FA_NBIT_22__FA_n2), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_22__FA_n4) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_22__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[23]), .Z(alu_ex_FULL_ADDER_FA_NBIT_22__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_23__FA_U7 ( .A1(alu_ex_add_sub_in[23]), 
        .A2(opA_in[23]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_23__FA_n3) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_23__FA_U6 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_23__FA_n5), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_23__FA_n2) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_23__FA_U5 ( .A(alu_ex_add_sub_in[23]), 
        .B(opA_in[23]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_23__FA_n5) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_23__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_carry[24]), .A2(alu_ex_FULL_ADDER_FA_NBIT_23__FA_n2), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_23__FA_n4) );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_23__FA_U3 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_23__FA_n1), .B(
        alu_ex_FULL_ADDER_FA_NBIT_23__FA_n5), .ZN(alu_ex_add_sub_out_23_) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_23__FA_U2 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_23__FA_n4), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_23__FA_n3), .ZN(alu_ex_FULL_ADDER_carry[23])
         );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_23__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[24]), .Z(alu_ex_FULL_ADDER_FA_NBIT_23__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_24__FA_U7 ( .A1(alu_ex_add_sub_in[24]), 
        .A2(opA_in[24]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_24__FA_n3) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_24__FA_U6 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_24__FA_n5), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_24__FA_n2) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_24__FA_U5 ( .A(alu_ex_add_sub_in[24]), 
        .B(opA_in[24]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_24__FA_n5) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_24__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_24__FA_n4), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_24__FA_n3), .ZN(alu_ex_FULL_ADDER_carry[24])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_24__FA_U3 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_24__FA_n1), .B(
        alu_ex_FULL_ADDER_FA_NBIT_24__FA_n5), .ZN(alu_ex_add_sub_out_24_) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_24__FA_U2 ( .A1(
        alu_ex_FULL_ADDER_carry[25]), .A2(alu_ex_FULL_ADDER_FA_NBIT_24__FA_n2), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_24__FA_n4) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_24__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[25]), .Z(alu_ex_FULL_ADDER_FA_NBIT_24__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_25__FA_U7 ( .A1(alu_ex_add_sub_in[25]), 
        .A2(opA_in[25]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_25__FA_n3) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_25__FA_U6 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_25__FA_n5), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_25__FA_n2) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_25__FA_U5 ( .A(alu_ex_add_sub_in[25]), 
        .B(opA_in[25]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_25__FA_n5) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_25__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_25__FA_n4), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_25__FA_n3), .ZN(alu_ex_FULL_ADDER_carry[25])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_25__FA_U3 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_25__FA_n1), .B(
        alu_ex_FULL_ADDER_FA_NBIT_25__FA_n5), .ZN(alu_ex_add_sub_out_25_) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_25__FA_U2 ( .A1(
        alu_ex_FULL_ADDER_carry[26]), .A2(alu_ex_FULL_ADDER_FA_NBIT_25__FA_n2), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_25__FA_n4) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_25__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[26]), .Z(alu_ex_FULL_ADDER_FA_NBIT_25__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_26__FA_U7 ( .A1(alu_ex_add_sub_in[26]), 
        .A2(opA_in[26]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_26__FA_n3) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_26__FA_U6 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_26__FA_n5), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_26__FA_n2) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_26__FA_U5 ( .A(alu_ex_add_sub_in[26]), 
        .B(opA_in[26]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_26__FA_n5) );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_26__FA_U4 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_26__FA_n1), .B(
        alu_ex_FULL_ADDER_FA_NBIT_26__FA_n5), .ZN(alu_ex_add_sub_out_26_) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_26__FA_U3 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_26__FA_n4), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_26__FA_n3), .ZN(alu_ex_FULL_ADDER_carry[26])
         );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_26__FA_U2 ( .A1(
        alu_ex_FULL_ADDER_carry[27]), .A2(alu_ex_FULL_ADDER_FA_NBIT_26__FA_n2), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_26__FA_n4) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_26__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[27]), .Z(alu_ex_FULL_ADDER_FA_NBIT_26__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_27__FA_U7 ( .A1(alu_ex_add_sub_in[27]), 
        .A2(opA_in[27]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_27__FA_n3) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_27__FA_U6 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_27__FA_n5), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_27__FA_n2) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_27__FA_U5 ( .A(alu_ex_add_sub_in[27]), 
        .B(opA_in[27]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_27__FA_n5) );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_27__FA_U4 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_27__FA_n1), .B(
        alu_ex_FULL_ADDER_FA_NBIT_27__FA_n5), .ZN(alu_ex_add_sub_out_27_) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_27__FA_U3 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_27__FA_n4), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_27__FA_n3), .ZN(alu_ex_FULL_ADDER_carry[27])
         );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_27__FA_U2 ( .A1(
        alu_ex_FULL_ADDER_carry[28]), .A2(alu_ex_FULL_ADDER_FA_NBIT_27__FA_n2), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_27__FA_n4) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_27__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[28]), .Z(alu_ex_FULL_ADDER_FA_NBIT_27__FA_n1) );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_28__FA_U7 ( .A1(alu_ex_add_sub_in[28]), 
        .A2(opA_in[28]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_28__FA_n3) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_28__FA_U6 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_28__FA_n5), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_28__FA_n2) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_28__FA_U5 ( .A(alu_ex_add_sub_in[28]), 
        .B(opA_in[28]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_28__FA_n5) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_28__FA_U4 ( .A1(
        alu_ex_FULL_ADDER_carry[29]), .A2(alu_ex_FULL_ADDER_FA_NBIT_28__FA_n2), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_28__FA_n4) );
  NAND2_X4 alu_ex_FULL_ADDER_FA_NBIT_28__FA_U3 ( .A1(
        alu_ex_FULL_ADDER_FA_NBIT_28__FA_n4), .A2(
        alu_ex_FULL_ADDER_FA_NBIT_28__FA_n3), .ZN(alu_ex_FULL_ADDER_carry[28])
         );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_28__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_28__FA_n1), .B(
        alu_ex_FULL_ADDER_FA_NBIT_28__FA_n5), .ZN(alu_ex_add_sub_out_28_) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_28__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[29]), .Z(alu_ex_FULL_ADDER_FA_NBIT_28__FA_n1) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_29__FA_U8 ( .A(alu_ex_add_sub_in[29]), 
        .B(opA_in[29]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_29__FA_n6) );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_29__FA_U7 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_29__FA_n2), .B(
        alu_ex_FULL_ADDER_FA_NBIT_29__FA_n3), .ZN(alu_ex_add_sub_out_29_) );
  OAI21_X4 alu_ex_FULL_ADDER_FA_NBIT_29__FA_U6 ( .B1(
        alu_ex_FULL_ADDER_FA_NBIT_29__FA_n6), .B2(
        alu_ex_FULL_ADDER_FA_NBIT_29__FA_n4), .A(
        alu_ex_FULL_ADDER_FA_NBIT_29__FA_n5), .ZN(alu_ex_FULL_ADDER_carry[29])
         );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_29__FA_U5 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_29__FA_n6), .Z(
        alu_ex_FULL_ADDER_FA_NBIT_29__FA_n3) );
  NAND2_X1 alu_ex_FULL_ADDER_FA_NBIT_29__FA_U4 ( .A1(alu_ex_add_sub_in[29]), 
        .A2(opA_in[29]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_29__FA_n5) );
  INV_X8 alu_ex_FULL_ADDER_FA_NBIT_29__FA_U3 ( .A(alu_ex_FULL_ADDER_carry[30]), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_29__FA_n4) );
  INV_X1 alu_ex_FULL_ADDER_FA_NBIT_29__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_29__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_29__FA_n2) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_29__FA_U1 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_29__FA_n4), .Z(
        alu_ex_FULL_ADDER_FA_NBIT_29__FA_n1) );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_30__FA_U7 ( .A(alu_ex_add_sub_in[30]), 
        .B(opA_in[30]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_30__FA_n5) );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_30__FA_U6 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_30__FA_n2), .B(
        alu_ex_FULL_ADDER_FA_NBIT_30__FA_n5), .ZN(alu_ex_add_sub_out_30_) );
  OAI21_X4 alu_ex_FULL_ADDER_FA_NBIT_30__FA_U5 ( .B1(
        alu_ex_FULL_ADDER_FA_NBIT_30__FA_n4), .B2(
        alu_ex_FULL_ADDER_FA_NBIT_30__FA_n5), .A(
        alu_ex_FULL_ADDER_FA_NBIT_30__FA_n3), .ZN(alu_ex_FULL_ADDER_carry[30])
         );
  NAND2_X2 alu_ex_FULL_ADDER_FA_NBIT_30__FA_U4 ( .A1(alu_ex_add_sub_in[30]), 
        .A2(opA_in[30]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_30__FA_n3) );
  INV_X1 alu_ex_FULL_ADDER_FA_NBIT_30__FA_U3 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_30__FA_n1), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_30__FA_n2) );
  BUF_X32 alu_ex_FULL_ADDER_FA_NBIT_30__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_30__FA_n4), .Z(
        alu_ex_FULL_ADDER_FA_NBIT_30__FA_n1) );
  INV_X4 alu_ex_FULL_ADDER_FA_NBIT_30__FA_U1 ( .A(alu_ex_FULL_ADDER_carry[31]), 
        .ZN(alu_ex_FULL_ADDER_FA_NBIT_30__FA_n4) );
  OAI21_X4 alu_ex_FULL_ADDER_FA_NBIT_31__FA_U7 ( .B1(
        alu_ex_FULL_ADDER_FA_NBIT_31__FA_n5), .B2(
        alu_ex_FULL_ADDER_FA_NBIT_31__FA_n3), .A(
        alu_ex_FULL_ADDER_FA_NBIT_31__FA_n4), .ZN(alu_ex_FULL_ADDER_carry[31])
         );
  XNOR2_X2 alu_ex_FULL_ADDER_FA_NBIT_31__FA_U6 ( .A(alu_ex_add_sub_in[31]), 
        .B(opA_in[31]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_31__FA_n5) );
  INV_X1 alu_ex_FULL_ADDER_FA_NBIT_31__FA_U5 ( .A(ALUCtrl_in[3]), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_31__FA_n3) );
  XOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_31__FA_U4 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_31__FA_n2), .B(
        alu_ex_FULL_ADDER_FA_NBIT_31__FA_n3), .Z(alu_ex_add_sub_out_31_) );
  NAND2_X1 alu_ex_FULL_ADDER_FA_NBIT_31__FA_U3 ( .A1(opA_in[31]), .A2(
        alu_ex_add_sub_in[31]), .ZN(alu_ex_FULL_ADDER_FA_NBIT_31__FA_n4) );
  XNOR2_X1 alu_ex_FULL_ADDER_FA_NBIT_31__FA_U2 ( .A(
        alu_ex_FULL_ADDER_FA_NBIT_31__FA_n1), .B(opA_in[31]), .ZN(
        alu_ex_FULL_ADDER_FA_NBIT_31__FA_n2) );
  BUF_X8 alu_ex_FULL_ADDER_FA_NBIT_31__FA_U1 ( .A(alu_ex_add_sub_in[31]), .Z(
        alu_ex_FULL_ADDER_FA_NBIT_31__FA_n1) );
  INV_X4 alu_ex_SHIFTER_U13 ( .A(opB_in[31]), .ZN(alu_ex_SHIFTER_n6) );
  INV_X4 alu_ex_SHIFTER_U12 ( .A(alu_ex_SHIFTER_n6), .ZN(alu_ex_SHIFTER_n5) );
  NAND2_X2 alu_ex_SHIFTER_U11 ( .A1(ALUCtrl_in[1]), .A2(opA_in[0]), .ZN(
        alu_ex_SHIFTER_n1) );
  INV_X4 alu_ex_SHIFTER_U10 ( .A(alu_ex_SHIFTER_n1), .ZN(alu_ex_SHIFTER_n4) );
  INV_X1 alu_ex_SHIFTER_U9 ( .A(opB_in[29]), .ZN(alu_ex_SHIFTER_n8) );
  INV_X4 alu_ex_SHIFTER_U8 ( .A(alu_ex_SHIFTER_n8), .ZN(alu_ex_SHIFTER_n7) );
  INV_X1 alu_ex_SHIFTER_U7 ( .A(opB_in[28]), .ZN(alu_ex_SHIFTER_n10) );
  INV_X4 alu_ex_SHIFTER_U6 ( .A(alu_ex_SHIFTER_n10), .ZN(alu_ex_SHIFTER_n9) );
  INV_X4 alu_ex_SHIFTER_U5 ( .A(opB_in[27]), .ZN(alu_ex_SHIFTER_n12) );
  INV_X4 alu_ex_SHIFTER_U4 ( .A(alu_ex_SHIFTER_n12), .ZN(alu_ex_SHIFTER_n11)
         );
  INV_X4 alu_ex_SHIFTER_U3 ( .A(alu_ex_SHIFTER_n1), .ZN(alu_ex_SHIFTER_n3) );
  INV_X4 alu_ex_SHIFTER_U2 ( .A(alu_ex_SHIFTER_n1), .ZN(alu_ex_SHIFTER_n2) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_U4 ( .A(alu_ex_SHIFTER_n11), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_U3 ( .A(alu_ex_SHIFTER_SHIFTLEFT16_n4), 
        .ZN(alu_ex_SHIFTER_SHIFTLEFT16_n3) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_U2 ( .A(alu_ex_SHIFTER_SHIFTLEFT16_n4), 
        .ZN(alu_ex_SHIFTER_SHIFTLEFT16_n1) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_U1 ( .A(alu_ex_SHIFTER_SHIFTLEFT16_n4), 
        .ZN(alu_ex_SHIFTER_SHIFTLEFT16_n2) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_0__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_0__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_0_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_0__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_0__MUX_U1 ( .A1(opA_in[0]), 
        .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_0__MUX_n1), .B1(
        opA_in[16]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_0__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_1__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_1_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_1__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_1__MUX_U1 ( .A1(opA_in[1]), 
        .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_1__MUX_n1), .B1(
        opA_in[17]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_1__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_2__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_2__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_2_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_2__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_2__MUX_U1 ( .A1(opA_in[2]), 
        .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_2__MUX_n1), .B1(
        opA_in[18]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_2__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_3__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_3__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_3_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_3__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_3__MUX_U1 ( .A1(opA_in[3]), 
        .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_3__MUX_n1), .B1(
        opA_in[19]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_3__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_4__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_4__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_4_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_4__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_4__MUX_U1 ( .A1(opA_in[4]), 
        .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_4__MUX_n1), .B1(
        opA_in[20]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_4__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_5__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_5__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_5_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_5__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_5__MUX_U1 ( .A1(opA_in[5]), 
        .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_5__MUX_n1), .B1(
        opA_in[21]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_5__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_6__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_6__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_6_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_6__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_6__MUX_U1 ( .A1(opA_in[6]), 
        .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_6__MUX_n1), .B1(
        opA_in[22]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_6__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_7__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_7__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_7_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_7__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_7__MUX_U1 ( .A1(opA_in[7]), 
        .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_7__MUX_n1), .B1(
        opA_in[23]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_7__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_8__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_8__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_8_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_8__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_8__MUX_U1 ( .A1(opA_in[8]), 
        .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_8__MUX_n1), .B1(
        opA_in[24]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_8__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_9__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_9__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_9_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_9__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_9__MUX_U1 ( .A1(opA_in[9]), 
        .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_9__MUX_n1), .B1(
        opA_in[25]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_9__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_10__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_10__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_10_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_10__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_10__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_10__MUX_U1 ( .A1(
        opA_in[10]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_10__MUX_n1), 
        .B1(opA_in[26]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_10__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_11__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_11__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_11_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_11__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_11__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_11__MUX_U1 ( .A1(
        opA_in[11]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_11__MUX_n1), 
        .B1(opA_in[27]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_11__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_12__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_12__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_12_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_12__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_12__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_12__MUX_U1 ( .A1(
        opA_in[12]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_12__MUX_n1), 
        .B1(opA_in[28]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_12__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_13__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_13__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_13_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_13__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_13__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_13__MUX_U1 ( .A1(
        opA_in[13]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_13__MUX_n1), 
        .B1(opA_in[29]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_13__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_14__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_14__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_14_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_14__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_14__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_14__MUX_U1 ( .A1(
        opA_in[14]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_14__MUX_n1), 
        .B1(opA_in[30]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_14__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_15__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_15__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp0_15_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_15__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_15__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_15__MUX_U1 ( .A1(
        opA_in[15]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_15__MUX_n1), 
        .B1(opA_in[31]), .B2(alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_15__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_16__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_16__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_16__MUX_U1 ( .A1(opA_in[16]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_16__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_16_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_17__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_17__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_17__MUX_U1 ( .A1(opA_in[17]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_17__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_17_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_18__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_18__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_18__MUX_U1 ( .A1(opA_in[18]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_18__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_18_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_19__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_19__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_19__MUX_U1 ( .A1(opA_in[19]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_19__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_19_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_20__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_20__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_20__MUX_U1 ( .A1(opA_in[20]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_20__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_20_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_21__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_21__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_21__MUX_U1 ( .A1(opA_in[21]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_21__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_21_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_22__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_22__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_22__MUX_U1 ( .A1(opA_in[22]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_22__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_22_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_23__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_23__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_23__MUX_U1 ( .A1(opA_in[23]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_23__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_23_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_24__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_24__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_24__MUX_U1 ( .A1(opA_in[24]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_24__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_24_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_25__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_25__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_25__MUX_U1 ( .A1(opA_in[25]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_25__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_25_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_26__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_26__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_26__MUX_U1 ( .A1(opA_in[26]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_26__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_26_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_27__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_27__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_27__MUX_U1 ( .A1(opA_in[27]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_27__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_27_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_28__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_28__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_28__MUX_U1 ( .A1(opA_in[28]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_28__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_28_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_29__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_29__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_29__MUX_U1 ( .A1(opA_in[29]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_29__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_29_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_30__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_30__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_30__MUX_U1 ( .A1(opA_in[30]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_30__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_30_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_31__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT16_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_31__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_31__MUX_U1 ( .A1(opA_in[31]), .A2(alu_ex_SHIFTER_SHIFTLEFT16_MUX2TO1_32BIT_31__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp0_31_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_U3 ( .A(alu_ex_SHIFTER_n9), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_n3) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_U2 ( .A(alu_ex_SHIFTER_SHIFTLEFT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_n1) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_U1 ( .A(alu_ex_SHIFTER_SHIFTLEFT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_n2) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_0__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_0__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_0_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_0__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_0__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_0_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_0__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_8_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_0__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_1__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_1_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_1__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_1__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_1_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_1__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_9_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_1__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_2__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_2__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_2_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_2__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_2__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_2_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_2__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_10_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_2__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_3__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_3__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_3_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_3__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_3__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_3_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_3__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_11_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_3__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_4__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_4__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_4_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_4__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_4__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_4_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_4__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_12_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_4__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_5__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_5__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_5_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_5__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_5__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_5_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_5__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_13_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_5__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_6__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_6__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_6_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_6__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_6__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_6_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_6__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_14_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_6__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_7__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_7__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_7_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_7__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_7__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_7_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_7__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_15_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_7__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_8__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_8__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_8_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_8__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_8__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_8_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_8__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_16_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_8__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_9__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_9__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_9_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_9__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_9__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_9_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_9__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_17_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_9__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_10__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_10__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_10_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_10__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_10__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_10__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_10_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_10__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_18_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_10__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_11__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_11__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_11_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_11__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_11__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_11__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_11_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_11__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_19_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_11__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_12__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_12__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_12_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_12__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_12__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_12__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_12_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_12__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_20_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_12__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_13__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_13__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_13_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_13__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_13__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_13__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_13_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_13__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_21_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_13__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_14__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_14__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_14_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_14__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_14__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_14__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_14_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_14__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_22_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_14__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_15__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_15__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_15_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_15__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_15__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_15__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_15_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_15__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_23_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_15__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_16__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_16__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_16_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_16__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_16__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_16__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_16_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_16__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_24_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_16__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_17__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_17__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_17_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_17__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_17__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_17__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_17_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_17__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_25_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_17__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_18__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_18__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_18_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_18__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_18__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_18__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_18_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_18__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_26_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_18__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_19__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_19__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_19_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_19__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_19__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_19__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_19_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_19__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_27_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_19__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_20__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_20__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_20_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_20__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_20__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_20__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_20_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_20__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_28_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_20__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_21__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_21__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_21_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_21__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_21__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_21__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_21_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_21__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_29_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_21__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_22__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_22__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_22_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_22__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_22__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_22__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_22_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_22__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_30_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_22__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_23__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_23__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp1_23_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_23__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_23__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_23__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_23_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_23__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp0_31_), .B2(alu_ex_SHIFTER_SHIFTLEFT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_23__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_24__MUX_U2 ( .A(
        alu_ex_SHIFTER_n9), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_24__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_24__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_24_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_24__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp1_24_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_25__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_25__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_25__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_25_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_25__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp1_25_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_26__MUX_U2 ( .A(
        alu_ex_SHIFTER_n9), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_26__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_26__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_26_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_26__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp1_26_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_27__MUX_U2 ( .A(
        alu_ex_SHIFTER_n9), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_27__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_27__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_27_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_27__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp1_27_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_28__MUX_U2 ( .A(
        alu_ex_SHIFTER_n9), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_28__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_28__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_28_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_28__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp1_28_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_29__MUX_U2 ( .A(
        alu_ex_SHIFTER_n9), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_29__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_29__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_29_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_29__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp1_29_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_30__MUX_U2 ( .A(
        alu_ex_SHIFTER_n9), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_30__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_30__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_30_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_30__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp1_30_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_31__MUX_U2 ( .A(
        alu_ex_SHIFTER_n9), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_31__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_31__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp0_31_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT8_MUX2TO1_32BIT_31__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp1_31_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_U3 ( .A(alu_ex_SHIFTER_n7), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_n3) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_U2 ( .A(alu_ex_SHIFTER_SHIFTLEFT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_n1) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_U1 ( .A(alu_ex_SHIFTER_SHIFTLEFT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_n2) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_0__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_0__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_0_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_0__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_0__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_0_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_0__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_4_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_0__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_1__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_1_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_1__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_1__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_1_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_1__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_5_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_1__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_2__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_2__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_2_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_2__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_2__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_2_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_2__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_6_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_2__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_3__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_3__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_3_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_3__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_3__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_3_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_3__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_7_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_3__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_4__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_4__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_4_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_4__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_4__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_4_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_4__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_8_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_4__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_5__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_5__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_5_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_5__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_5__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_5_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_5__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_9_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_5__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_6__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_6__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_6_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_6__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_6__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_6_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_6__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_10_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_6__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_7__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_7__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_7_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_7__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_7__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_7_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_7__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_11_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_7__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_8__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_8__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_8_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_8__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_8__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_8_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_8__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_12_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_8__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_9__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_9__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_9_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_9__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_9__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_9_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_9__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_13_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_9__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_10__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_10__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_10_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_10__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_10__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_10__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_10_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_10__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_14_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_10__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_11__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_11__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_11_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_11__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_11__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_11__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_11_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_11__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_15_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_11__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_12__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_12__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_12_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_12__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_12__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_12__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_12_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_12__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_16_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_12__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_13__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_13__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_13_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_13__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_13__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_13__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_13_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_13__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_17_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_13__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_14__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_14__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_14_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_14__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_14__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_14__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_14_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_14__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_18_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_14__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_15__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_15__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_15_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_15__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_15__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_15__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_15_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_15__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_19_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_15__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_16__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_16__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_16_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_16__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_16__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_16__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_16_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_16__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_20_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_16__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_17__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_17__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_17_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_17__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_17__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_17__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_17_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_17__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_21_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_17__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_18__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_18__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_18_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_18__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_18__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_18__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_18_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_18__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_22_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_18__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_19__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_19__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_19_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_19__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_19__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_19__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_19_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_19__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_23_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_19__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_20__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_20__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_20_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_20__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_20__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_20__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_20_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_20__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_24_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_20__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_21__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_21__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_21_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_21__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_21__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_21__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_21_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_21__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_25_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_21__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_22__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_22__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_22_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_22__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_22__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_22__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_22_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_22__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_26_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_22__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_23__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_23__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_23_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_23__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_23__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_23__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_23_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_23__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_27_), .B2(alu_ex_SHIFTER_SHIFTLEFT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_23__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_24__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_24__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_24_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_24__MUX_U2 ( .A(
        alu_ex_SHIFTER_n7), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_24__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_24__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_24_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_24__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_28_), .B2(alu_ex_SHIFTER_n7), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_24__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_25__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_25__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_25_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_25__MUX_U2 ( .A(
        alu_ex_SHIFTER_n7), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_25__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_25__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_25_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_25__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_29_), .B2(alu_ex_SHIFTER_n7), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_25__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_26__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_26__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_26_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_26__MUX_U2 ( .A(
        alu_ex_SHIFTER_n7), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_26__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_26__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_26_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_26__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_30_), .B2(alu_ex_SHIFTER_n7), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_26__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_27__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_27__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp2_27_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_27__MUX_U2 ( .A(
        alu_ex_SHIFTER_n7), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_27__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_27__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_27_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_27__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp1_31_), .B2(alu_ex_SHIFTER_n7), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_27__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_28__MUX_U2 ( .A(
        alu_ex_SHIFTER_n7), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_28__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_28__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_28_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_28__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp2_28_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_29__MUX_U2 ( .A(
        alu_ex_SHIFTER_n7), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_29__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_29__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_29_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_29__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp2_29_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_30__MUX_U2 ( .A(
        alu_ex_SHIFTER_n7), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_30__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_30__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_30_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_30__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp2_30_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_31__MUX_U2 ( .A(
        alu_ex_SHIFTER_n7), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_31__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_31__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp1_31_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT4_MUX2TO1_32BIT_31__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp2_31_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_U4 ( .A(opB_in[30]), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_U3 ( .A(alu_ex_SHIFTER_SHIFTLEFT2_n4), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_n3) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_U2 ( .A(alu_ex_SHIFTER_SHIFTLEFT2_n4), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_n1) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_U1 ( .A(alu_ex_SHIFTER_SHIFTLEFT2_n4), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_n2) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_0__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_0__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_0_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_0__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_0__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_0_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_0__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_2_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_0__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_1__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_1_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_1__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_1__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_1_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_1__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_3_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_1__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_2__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_2__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_2_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_2__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_2__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_2_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_2__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_4_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_2__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_3__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_3__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_3_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_3__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_3__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_3_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_3__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_5_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_3__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_4__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_4__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_4_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_4__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_4__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_4_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_4__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_6_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_4__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_5__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_5__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_5_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_5__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_5__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_5_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_5__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_7_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_5__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_6__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_6__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_6_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_6__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_6__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_6_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_6__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_8_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_6__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_7__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_7__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_7_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_7__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_7__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_7_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_7__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_9_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_7__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_8__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_8__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_8_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_8__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_8__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_8_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_8__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_10_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_8__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_9__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_9__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_9_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_9__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_9__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_9_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_9__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_11_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_9__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_10__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_10__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_10_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_10__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_10__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_10__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_10_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_10__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_12_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_10__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_11__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_11__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_11_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_11__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_11__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_11__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_11_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_11__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_13_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_11__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_12__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_12__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_12_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_12__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_12__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_12__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_12_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_12__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_14_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_12__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_13__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_13__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_13_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_13__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_13__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_13__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_13_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_13__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_15_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_13__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_14__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_14__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_14_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_14__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_14__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_14__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_14_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_14__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_16_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_14__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_15__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_15__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_15_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_15__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_15__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_15__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_15_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_15__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_17_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_15__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_16__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_16__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_16_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_16__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_16__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_16__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_16_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_16__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_18_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_16__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_17__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_17__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_17_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_17__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_17__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_17__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_17_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_17__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_19_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_17__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_18__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_18__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_18_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_18__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_18__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_18__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_18_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_18__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_20_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_18__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_19__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_19__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_19_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_19__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_19__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_19__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_19_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_19__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_21_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_19__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_20__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_20__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_20_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_20__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_20__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_20__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_20_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_20__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_22_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_20__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_21__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_21__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_21_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_21__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_21__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_21__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_21_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_21__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_23_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_21__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_22__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_22__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_22_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_22__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_22__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_22__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_22_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_22__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_24_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_22__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_23__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_23__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_23_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_23__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_23__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_23__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_23_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_23__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_25_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_23__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_24__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_24__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_24_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_24__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_24__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_24__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_24_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_24__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_26_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_24__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_25__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_25__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_25_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_25__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_25__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_25__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_25_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_25__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_27_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_25__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_26__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_26__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_26_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_26__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_26__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_26__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_26_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_26__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_28_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_26__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_27__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_27__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_27_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_27__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_27__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_27__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_27_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_27__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_29_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_27__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_28__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_28__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_28_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_28__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_28__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_28__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_28_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_28__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_30_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_28__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_29__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_29__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp3_29_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_29__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_29__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_29__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_29_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_29__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp2_31_), .B2(alu_ex_SHIFTER_SHIFTLEFT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_29__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_30__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_30__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_30__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_30_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_30__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp3_30_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_31__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_31__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_31__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp2_31_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT2_MUX2TO1_32BIT_31__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp3_31_) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_U3 ( .A(alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_n3) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_U2 ( .A(alu_ex_SHIFTER_SHIFTLEFT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_n1) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_U1 ( .A(alu_ex_SHIFTER_SHIFTLEFT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_n2) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_0__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_0__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[0]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_0__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_0__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_0_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_0__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_1_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_0__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_1__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[1]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_1__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_1__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_1_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_1__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_2_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_1__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_2__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_2__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[2]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_2__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_2__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_2_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_2__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_3_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_2__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_3__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_3__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[3]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_3__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_3__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_3_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_3__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_4_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_3__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_4__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_4__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[4]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_4__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_4__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_4_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_4__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_5_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_4__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_5__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_5__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[5]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_5__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_5__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_5_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_5__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_6_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_5__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_6__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_6__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[6]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_6__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_6__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_6_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_6__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_7_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_6__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_7__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_7__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[7]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_7__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_7__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_7_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_7__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_8_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_7__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_8__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_8__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[8]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_8__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_8__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_8_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_8__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_9_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_8__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_9__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_9__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[9]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_9__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_9__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_9_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_9__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_10_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_9__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_10__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_10__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[10]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_10__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_10__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_10__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_10_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_10__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_11_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_10__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_11__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_11__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[11]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_11__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_11__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_11__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_11_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_11__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_12_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_11__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_12__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_12__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[12]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_12__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_12__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_12__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_12_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_12__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_13_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_12__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_13__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_13__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[13]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_13__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_13__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_13__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_13_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_13__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_14_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_13__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_14__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_14__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[14]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_14__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_14__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_14__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_14_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_14__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_15_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_14__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_15__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_15__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[15]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_15__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_15__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_15__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_15_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_15__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_16_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_15__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_16__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_16__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[16]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_16__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_16__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_16__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_16_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_16__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_17_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_16__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_17__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_17__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[17]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_17__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_17__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_17__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_17_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_17__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_18_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_17__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_18__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_18__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[18]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_18__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_18__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_18__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_18_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_18__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_19_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_18__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_19__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_19__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[19]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_19__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_19__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_19__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_19_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_19__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_20_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_19__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_20__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_20__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[20]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_20__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_20__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_20__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_20_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_20__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_21_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_20__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_21__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_21__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[21]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_21__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_21__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_21__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_21_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_21__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_22_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_21__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_22__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_22__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[22]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_22__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_22__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_22__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_22_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_22__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_23_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_22__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_23__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_23__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[23]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_23__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_23__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_23__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_23_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_23__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_24_), .B2(alu_ex_SHIFTER_SHIFTLEFT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_23__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_24__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_24__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[24]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_24__MUX_U2 ( .A(
        alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_24__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_24__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_24_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_24__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_25_), .B2(alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_24__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_25__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_25__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[25]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_25__MUX_U2 ( .A(
        alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_25__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_25__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_25_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_25__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_26_), .B2(alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_25__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_26__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_26__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[26]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_26__MUX_U2 ( .A(
        alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_26__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_26__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_26_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_26__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_27_), .B2(alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_26__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_27__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_27__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[27]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_27__MUX_U2 ( .A(
        alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_27__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_27__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_27_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_27__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_28_), .B2(alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_27__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_28__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_28__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[28]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_28__MUX_U2 ( .A(
        alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_28__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_28__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_28_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_28__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_29_), .B2(alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_28__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_29__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_29__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[29]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_29__MUX_U2 ( .A(
        alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_29__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_29__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_29_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_29__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_30_), .B2(alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_29__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_30__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_30__MUX_n4), .ZN(
        alu_ex_SHIFTER_ltemp4[30]) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_30__MUX_U2 ( .A(
        alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_30__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_30__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_30_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_30__MUX_n1), .B1(
        alu_ex_SHIFTER_ltemp3_31_), .B2(alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_30__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_31__MUX_U2 ( .A(
        alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_31__MUX_n2) );
  AND2_X4 alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_31__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp3_31_), .A2(
        alu_ex_SHIFTER_SHIFTLEFT1_MUX2TO1_32BIT_31__MUX_n2), .ZN(
        alu_ex_SHIFTER_ltemp4[31]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_U3 ( .A(alu_ex_SHIFTER_n11), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_n3) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_U2 ( .A(alu_ex_SHIFTER_SHIFTRIGHT16_n3), 
        .ZN(alu_ex_SHIFTER_SHIFTRIGHT16_n1) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_U1 ( .A(alu_ex_SHIFTER_SHIFTRIGHT16_n3), 
        .ZN(alu_ex_SHIFTER_SHIFTRIGHT16_n2) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_0__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_0__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_0_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_0__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_0__MUX_U1 ( .A1(opA_in[0]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_0__MUX_n1), .B1(
        alu_ex_SHIFTER_n3), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_0__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_1__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_1_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_1__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_1__MUX_U1 ( .A1(opA_in[1]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_1__MUX_n1), .B1(
        alu_ex_SHIFTER_n3), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_1__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_2__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_2__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_2_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_2__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_2__MUX_U1 ( .A1(opA_in[2]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_2__MUX_n1), .B1(
        alu_ex_SHIFTER_n3), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_2__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_3__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_3__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_3_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_3__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_3__MUX_U1 ( .A1(opA_in[3]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_3__MUX_n1), .B1(
        alu_ex_SHIFTER_n3), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_3__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_4__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_4__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_4_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_4__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_4__MUX_U1 ( .A1(opA_in[4]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_4__MUX_n1), .B1(
        alu_ex_SHIFTER_n2), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_4__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_5__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_5__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_5_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_5__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_5__MUX_U1 ( .A1(opA_in[5]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_5__MUX_n1), .B1(
        alu_ex_SHIFTER_n2), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_5__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_6__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_6__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_6_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_6__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_6__MUX_U1 ( .A1(opA_in[6]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_6__MUX_n1), .B1(
        alu_ex_SHIFTER_n2), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_6__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_7__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_7__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_7_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_7__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_7__MUX_U1 ( .A1(opA_in[7]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_7__MUX_n1), .B1(
        alu_ex_SHIFTER_n2), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_7__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_8__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_8__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_8_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_8__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_8__MUX_U1 ( .A1(opA_in[8]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_8__MUX_n1), .B1(
        alu_ex_SHIFTER_n2), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_8__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_9__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_9__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_9_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_9__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_9__MUX_U1 ( .A1(opA_in[9]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_9__MUX_n1), .B1(
        alu_ex_SHIFTER_n2), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_9__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_10__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_10__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_10_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_10__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_10__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_10__MUX_U1 ( .A1(
        opA_in[10]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_10__MUX_n1), 
        .B1(alu_ex_SHIFTER_n2), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_10__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_11__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_11__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_11_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_11__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_11__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_11__MUX_U1 ( .A1(
        opA_in[11]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_11__MUX_n1), 
        .B1(alu_ex_SHIFTER_n2), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_11__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_12__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_12__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_12_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_12__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_12__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_12__MUX_U1 ( .A1(
        opA_in[12]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_12__MUX_n1), 
        .B1(alu_ex_SHIFTER_n2), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_12__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_13__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_13__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_13_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_13__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_13__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_13__MUX_U1 ( .A1(
        opA_in[13]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_13__MUX_n1), 
        .B1(alu_ex_SHIFTER_n2), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_13__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_14__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_14__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_14_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_14__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_14__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_14__MUX_U1 ( .A1(
        opA_in[14]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_14__MUX_n1), 
        .B1(alu_ex_SHIFTER_n2), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_14__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_15__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_15__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_15_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_15__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_15__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_15__MUX_U1 ( .A1(
        opA_in[15]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_15__MUX_n1), 
        .B1(alu_ex_SHIFTER_n2), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_15__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_16__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_16__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_16_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_16__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_16__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_16__MUX_U1 ( .A1(
        opA_in[16]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_16__MUX_n1), 
        .B1(opA_in[0]), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_16__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_17__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_17__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_17_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_17__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_17__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_17__MUX_U1 ( .A1(
        opA_in[17]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_17__MUX_n1), 
        .B1(opA_in[1]), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_17__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_18__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_18__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_18_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_18__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_18__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_18__MUX_U1 ( .A1(
        opA_in[18]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_18__MUX_n1), 
        .B1(opA_in[2]), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_18__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_19__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_19__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_19_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_19__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_19__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_19__MUX_U1 ( .A1(
        opA_in[19]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_19__MUX_n1), 
        .B1(opA_in[3]), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_19__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_20__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_20__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_20_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_20__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_20__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_20__MUX_U1 ( .A1(
        opA_in[20]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_20__MUX_n1), 
        .B1(opA_in[4]), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_20__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_21__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_21__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_21_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_21__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_21__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_21__MUX_U1 ( .A1(
        opA_in[21]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_21__MUX_n1), 
        .B1(opA_in[5]), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_21__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_22__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_22__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_22_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_22__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_22__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_22__MUX_U1 ( .A1(
        opA_in[22]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_22__MUX_n1), 
        .B1(opA_in[6]), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_22__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_23__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_23__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_23_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_23__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_23__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_23__MUX_U1 ( .A1(
        opA_in[23]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_23__MUX_n1), 
        .B1(opA_in[7]), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_23__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_24__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_24__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_24_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_24__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_24__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_24__MUX_U1 ( .A1(
        opA_in[24]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_24__MUX_n1), 
        .B1(opA_in[8]), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_24__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_25__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_25__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_25_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_25__MUX_U2 ( .A(
        alu_ex_SHIFTER_n11), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_25__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_25__MUX_U1 ( .A1(
        opA_in[25]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_25__MUX_n1), 
        .B1(opA_in[9]), .B2(alu_ex_SHIFTER_n11), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_25__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_26__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_26__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_26_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_26__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_26__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_26__MUX_U1 ( .A1(
        opA_in[26]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_26__MUX_n1), 
        .B1(opA_in[10]), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_26__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_27__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_27__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_27_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_27__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_27__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_27__MUX_U1 ( .A1(
        opA_in[27]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_27__MUX_n1), 
        .B1(opA_in[11]), .B2(alu_ex_SHIFTER_SHIFTRIGHT16_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_27__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_28__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_28__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_28_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_28__MUX_U2 ( .A(
        alu_ex_SHIFTER_n11), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_28__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_28__MUX_U1 ( .A1(
        opA_in[28]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_28__MUX_n1), 
        .B1(opA_in[12]), .B2(alu_ex_SHIFTER_n11), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_28__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_29__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_29__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_29_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_29__MUX_U2 ( .A(
        alu_ex_SHIFTER_n11), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_29__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_29__MUX_U1 ( .A1(
        opA_in[29]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_29__MUX_n1), 
        .B1(opA_in[13]), .B2(alu_ex_SHIFTER_n11), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_29__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_30__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_30__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_30_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_30__MUX_U2 ( .A(
        alu_ex_SHIFTER_n11), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_30__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_30__MUX_U1 ( .A1(
        opA_in[30]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_30__MUX_n1), 
        .B1(opA_in[14]), .B2(alu_ex_SHIFTER_n11), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_30__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_31__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_31__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp0_31_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_31__MUX_U2 ( .A(
        alu_ex_SHIFTER_n11), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_31__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_31__MUX_U1 ( .A1(
        opA_in[31]), .A2(alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_31__MUX_n1), 
        .B1(opA_in[15]), .B2(alu_ex_SHIFTER_n11), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT16_MUX2TO1_32BIT_31__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_U4 ( .A(alu_ex_SHIFTER_n9), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_U3 ( .A(alu_ex_SHIFTER_SHIFTRIGHT8_n4), 
        .ZN(alu_ex_SHIFTER_SHIFTRIGHT8_n3) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_U2 ( .A(alu_ex_SHIFTER_SHIFTRIGHT8_n4), 
        .ZN(alu_ex_SHIFTER_SHIFTRIGHT8_n1) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_U1 ( .A(alu_ex_SHIFTER_SHIFTRIGHT8_n4), 
        .ZN(alu_ex_SHIFTER_SHIFTRIGHT8_n2) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_0__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_0__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_0_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_0__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_0__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_0_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_0__MUX_n1), .B1(
        alu_ex_SHIFTER_n3), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_0__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_1__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_1_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_1__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_1__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_1_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_1__MUX_n1), .B1(
        alu_ex_SHIFTER_n3), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_1__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_2__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_2__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_2_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_2__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_2__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_2_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_2__MUX_n1), .B1(
        alu_ex_SHIFTER_n3), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_2__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_3__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_3__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_3_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_3__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_3__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_3_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_3__MUX_n1), .B1(
        alu_ex_SHIFTER_n3), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_3__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_4__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_4__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_4_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_4__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_4__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_4_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_4__MUX_n1), .B1(
        alu_ex_SHIFTER_n3), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_4__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_5__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_5__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_5_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_5__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_5__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_5_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_5__MUX_n1), .B1(
        alu_ex_SHIFTER_n3), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_5__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_6__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_6__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_6_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_6__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_6__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_6_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_6__MUX_n1), .B1(
        alu_ex_SHIFTER_n3), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_6__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_7__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_7__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_7_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_7__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_7__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_7_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_7__MUX_n1), .B1(
        alu_ex_SHIFTER_n3), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_7__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_8__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_8__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_8_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_8__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_8__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_8_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_8__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_0_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_8__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_9__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_9__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_9_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_9__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_9__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_9_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_9__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_1_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_9__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_10__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_10__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_10_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_10__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_10__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_10__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_10_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_10__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_2_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_10__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_11__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_11__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_11_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_11__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_11__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_11__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_11_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_11__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_3_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_11__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_12__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_12__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_12_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_12__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_12__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_12__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_12_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_12__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_4_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_12__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_13__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_13__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_13_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_13__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_13__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_13__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_13_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_13__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_5_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_13__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_14__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_14__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_14_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_14__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_14__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_14__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_14_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_14__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_6_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_14__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_15__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_15__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_15_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_15__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_15__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_15__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_15_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_15__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_7_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_15__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_16__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_16__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_16_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_16__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_16__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_16__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_16_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_16__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_8_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_16__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_17__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_17__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_17_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_17__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_17__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_17__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_17_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_17__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_9_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_17__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_18__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_18__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_18_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_18__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_18__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_18__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_18_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_18__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_10_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_18__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_19__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_19__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_19_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_19__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_19__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_19__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_19_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_19__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_11_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_19__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_20__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_20__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_20_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_20__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_20__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_20__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_20_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_20__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_12_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_20__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_21__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_21__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_21_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_21__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_21__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_21__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_21_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_21__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_13_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_21__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_22__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_22__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_22_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_22__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_22__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_22__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_22_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_22__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_14_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_22__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_23__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_23__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_23_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_23__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_23__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_23__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_23_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_23__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_15_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_23__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_24__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_24__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_24_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_24__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_24__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_24__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_24_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_24__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_16_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_24__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_25__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_25__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_25_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_25__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_25__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_25__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_25_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_25__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_17_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_25__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_26__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_26__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_26_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_26__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_26__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_26__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_26_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_26__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_18_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_26__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_27__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_27__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_27_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_27__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_27__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_27__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_27_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_27__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_19_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_27__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_28__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_28__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_28_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_28__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_28__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_28__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_28_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_28__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_20_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_28__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_29__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_29__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_29_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_29__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_29__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_29__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_29_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_29__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_21_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_29__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_30__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_30__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_30_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_30__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_30__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_30__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_30_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_30__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_22_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_30__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_31__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_31__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp1_31_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_31__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_31__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_31__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp0_31_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_31__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp0_23_), .B2(alu_ex_SHIFTER_SHIFTRIGHT8_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT8_MUX2TO1_32BIT_31__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_U4 ( .A(alu_ex_SHIFTER_n7), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_U3 ( .A(alu_ex_SHIFTER_SHIFTRIGHT4_n4), 
        .ZN(alu_ex_SHIFTER_SHIFTRIGHT4_n3) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_U2 ( .A(alu_ex_SHIFTER_SHIFTRIGHT4_n4), 
        .ZN(alu_ex_SHIFTER_SHIFTRIGHT4_n1) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_U1 ( .A(alu_ex_SHIFTER_SHIFTRIGHT4_n4), 
        .ZN(alu_ex_SHIFTER_SHIFTRIGHT4_n2) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_0__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_0__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_0_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_0__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_0__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_0_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_0__MUX_n1), .B1(
        alu_ex_SHIFTER_n4), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_0__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_1__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_1_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_1__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_1__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_1_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_1__MUX_n1), .B1(
        alu_ex_SHIFTER_n4), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_1__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_2__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_2__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_2_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_2__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_2__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_2_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_2__MUX_n1), .B1(
        alu_ex_SHIFTER_n4), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_2__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_3__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_3__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_3_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_3__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_3__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_3_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_3__MUX_n1), .B1(
        alu_ex_SHIFTER_n4), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_3__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_4__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_4__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_4_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_4__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_4__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_4_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_4__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_0_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_4__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_5__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_5__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_5_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_5__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_5__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_5_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_5__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_1_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_5__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_6__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_6__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_6_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_6__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_6__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_6_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_6__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_2_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_6__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_7__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_7__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_7_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_7__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_7__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_7_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_7__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_3_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_7__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_8__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_8__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_8_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_8__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_8__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_8_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_8__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_4_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_8__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_9__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_9__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_9_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_9__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_9__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_9_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_9__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_5_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_9__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_10__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_10__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_10_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_10__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_10__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_10__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_10_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_10__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_6_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_10__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_11__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_11__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_11_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_11__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_11__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_11__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_11_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_11__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_7_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_11__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_12__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_12__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_12_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_12__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_12__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_12__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_12_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_12__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_8_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_12__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_13__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_13__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_13_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_13__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_13__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_13__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_13_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_13__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_9_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_13__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_14__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_14__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_14_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_14__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_14__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_14__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_14_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_14__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_10_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_14__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_15__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_15__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_15_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_15__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_15__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_15__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_15_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_15__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_11_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_15__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_16__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_16__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_16_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_16__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_16__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_16__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_16_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_16__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_12_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_16__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_17__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_17__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_17_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_17__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_17__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_17__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_17_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_17__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_13_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_17__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_18__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_18__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_18_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_18__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_18__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_18__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_18_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_18__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_14_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_18__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_19__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_19__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_19_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_19__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_19__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_19__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_19_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_19__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_15_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_19__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_20__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_20__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_20_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_20__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_20__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_20__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_20_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_20__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_16_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_20__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_21__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_21__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_21_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_21__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_21__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_21__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_21_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_21__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_17_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_21__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_22__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_22__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_22_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_22__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_22__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_22__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_22_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_22__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_18_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_22__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_23__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_23__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_23_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_23__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_23__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_23__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_23_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_23__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_19_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_23__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_24__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_24__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_24_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_24__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_24__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_24__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_24_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_24__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_20_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_24__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_25__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_25__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_25_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_25__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_25__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_25__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_25_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_25__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_21_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_25__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_26__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_26__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_26_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_26__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_26__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_26__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_26_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_26__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_22_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_26__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_27__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_27__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_27_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_27__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_27__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_27__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_27_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_27__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_23_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_27__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_28__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_28__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_28_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_28__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_28__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_28__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_28_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_28__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_24_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_28__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_29__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_29__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_29_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_29__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_29__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_29__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_29_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_29__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_25_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_29__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_30__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_30__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_30_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_30__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_30__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_30__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_30_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_30__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_26_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_30__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_31__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_31__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp2_31_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_31__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_31__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_31__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp1_31_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_31__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp1_27_), .B2(alu_ex_SHIFTER_SHIFTRIGHT4_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT4_MUX2TO1_32BIT_31__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_U4 ( .A(opB_in[30]), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_U3 ( .A(alu_ex_SHIFTER_SHIFTRIGHT2_n4), 
        .ZN(alu_ex_SHIFTER_SHIFTRIGHT2_n3) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_U2 ( .A(alu_ex_SHIFTER_SHIFTRIGHT2_n4), 
        .ZN(alu_ex_SHIFTER_SHIFTRIGHT2_n1) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_U1 ( .A(alu_ex_SHIFTER_SHIFTRIGHT2_n4), 
        .ZN(alu_ex_SHIFTER_SHIFTRIGHT2_n2) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_0__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_0__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_0_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_0__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_0__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_0_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_0__MUX_n1), .B1(
        alu_ex_SHIFTER_n4), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_0__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_1__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_1_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_1__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_1__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_1_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_1__MUX_n1), .B1(
        alu_ex_SHIFTER_n4), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_1__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_2__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_2__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_2_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_2__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_2__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_2_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_2__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_0_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_2__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_3__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_3__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_3_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_3__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_3__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_3_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_3__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_1_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_3__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_4__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_4__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_4_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_4__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_4__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_4_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_4__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_2_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_4__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_5__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_5__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_5_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_5__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_5__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_5_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_5__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_3_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_5__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_6__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_6__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_6_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_6__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_6__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_6_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_6__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_4_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_6__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_7__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_7__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_7_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_7__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_7__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_7_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_7__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_5_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_7__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_8__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_8__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_8_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_8__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_8__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_8_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_8__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_6_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_8__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_9__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_9__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_9_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_9__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_9__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_9_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_9__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_7_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_9__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_10__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_10__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_10_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_10__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_10__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_10__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_10_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_10__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_8_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_10__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_11__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_11__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_11_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_11__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_11__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_11__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_11_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_11__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_9_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_11__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_12__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_12__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_12_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_12__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_12__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_12__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_12_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_12__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_10_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_12__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_13__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_13__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_13_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_13__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_13__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_13__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_13_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_13__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_11_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_13__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_14__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_14__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_14_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_14__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_14__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_14__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_14_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_14__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_12_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_14__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_15__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_15__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_15_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_15__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_15__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_15__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_15_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_15__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_13_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_15__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_16__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_16__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_16_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_16__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_16__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_16__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_16_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_16__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_14_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_16__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_17__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_17__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_17_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_17__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_17__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_17__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_17_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_17__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_15_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_17__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_18__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_18__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_18_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_18__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_18__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_18__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_18_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_18__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_16_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_18__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_19__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_19__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_19_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_19__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_19__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_19__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_19_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_19__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_17_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_19__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_20__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_20__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_20_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_20__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_20__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_20__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_20_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_20__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_18_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_20__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_21__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_21__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_21_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_21__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_21__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_21__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_21_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_21__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_19_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_21__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_22__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_22__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_22_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_22__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_22__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_22__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_22_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_22__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_20_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_22__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_23__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_23__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_23_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_23__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_23__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_23__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_23_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_23__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_21_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_23__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_24__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_24__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_24_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_24__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_24__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_24__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_24_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_24__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_22_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_24__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_25__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_25__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_25_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_25__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_25__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_25__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_25_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_25__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_23_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_25__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_26__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_26__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_26_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_26__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_26__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_26__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_26_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_26__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_24_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_26__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_27__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_27__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_27_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_27__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_27__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_27__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_27_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_27__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_25_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_27__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_28__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_28__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_28_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_28__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_28__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_28__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_28_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_28__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_26_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_28__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_29__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_29__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_29_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_29__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_29__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_29__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_29_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_29__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_27_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_29__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_30__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_30__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_30_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_30__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_30__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_30__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_30_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_30__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_28_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_30__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_31__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_31__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp3_31_) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_31__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_31__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_31__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp2_31_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_31__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp2_29_), .B2(alu_ex_SHIFTER_SHIFTRIGHT2_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT2_MUX2TO1_32BIT_31__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_U4 ( .A(alu_ex_SHIFTER_n5), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_U3 ( .A(alu_ex_SHIFTER_SHIFTRIGHT1_n4), 
        .ZN(alu_ex_SHIFTER_SHIFTRIGHT1_n3) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_U2 ( .A(alu_ex_SHIFTER_SHIFTRIGHT1_n4), 
        .ZN(alu_ex_SHIFTER_SHIFTRIGHT1_n1) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_U1 ( .A(alu_ex_SHIFTER_SHIFTRIGHT1_n4), 
        .ZN(alu_ex_SHIFTER_SHIFTRIGHT1_n2) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_0__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_0__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[0]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_0__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_0__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_0_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_0__MUX_n1), .B1(
        alu_ex_SHIFTER_n4), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_0__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_1__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[1]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_1__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_1__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_1_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_1__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_0_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_1__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_2__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_2__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[2]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_2__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_2__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_2_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_2__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_1_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_2__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_3__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_3__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[3]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_3__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_3__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_3_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_3__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_2_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_3__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_4__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_4__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[4]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_4__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_4__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_4_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_4__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_3_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_4__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_5__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_5__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[5]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_5__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_5__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_5_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_5__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_4_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_5__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_6__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_6__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[6]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_6__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_6__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_6_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_6__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_5_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_6__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_7__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_7__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[7]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_7__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_7__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_7_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_7__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_6_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_7__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_8__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_8__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[8]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_8__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_8__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_8_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_8__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_7_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_8__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_9__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_9__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[9]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_9__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_9__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_9_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_9__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_8_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_9__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_10__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_10__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[10]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_10__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_10__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_10__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_10_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_10__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_9_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_10__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_11__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_11__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[11]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_11__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_11__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_11__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_11_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_11__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_10_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n1), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_11__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_12__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_12__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[12]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_12__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_12__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_12__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_12_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_12__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_11_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_12__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_13__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_13__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[13]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_13__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_13__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_13__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_13_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_13__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_12_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_13__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_14__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_14__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[14]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_14__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_14__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_14__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_14_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_14__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_13_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_14__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_15__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_15__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[15]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_15__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_15__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_15__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_15_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_15__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_14_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_15__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_16__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_16__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[16]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_16__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_16__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_16__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_16_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_16__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_15_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_16__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_17__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_17__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[17]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_17__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_17__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_17__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_17_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_17__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_16_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_17__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_18__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_18__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[18]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_18__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_18__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_18__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_18_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_18__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_17_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_18__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_19__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_19__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[19]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_19__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_19__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_19__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_19_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_19__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_18_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_19__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_20__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_20__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[20]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_20__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_20__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_20__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_20_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_20__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_19_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_20__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_21__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_21__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[21]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_21__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_21__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_21__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_21_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_21__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_20_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_21__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_22__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_22__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[22]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_22__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_22__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_22__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_22_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_22__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_21_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_22__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_23__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_23__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[23]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_23__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_23__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_23__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_23_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_23__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_22_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n2), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_23__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_24__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_24__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[24]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_24__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_24__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_24__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_24_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_24__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_23_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_24__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_25__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_25__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[25]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_25__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_25__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_25__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_25_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_25__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_24_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_25__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_26__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_26__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[26]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_26__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_26__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_26__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_26_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_26__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_25_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_26__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_27__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_27__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[27]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_27__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_27__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_27__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_27_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_27__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_26_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_27__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_28__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_28__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[28]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_28__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_28__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_28__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_28_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_28__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_27_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_28__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_29__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_29__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[29]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_29__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_29__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_29__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_29_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_29__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_28_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_29__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_30__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_30__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[30]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_30__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_30__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_30__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_30_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_30__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_29_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_30__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_31__MUX_U3 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_31__MUX_n4), .ZN(
        alu_ex_SHIFTER_rtemp4[31]) );
  INV_X4 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_31__MUX_U2 ( .A(
        alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_31__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_31__MUX_U1 ( .A1(
        alu_ex_SHIFTER_rtemp3_31_), .A2(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_31__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp3_30_), .B2(alu_ex_SHIFTER_SHIFTRIGHT1_n3), .ZN(
        alu_ex_SHIFTER_SHIFTRIGHT1_MUX2TO1_32BIT_31__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_U4 ( .A(ALUCtrl_in[2]), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_U3 ( .A(alu_ex_SHIFTER_LEFTORRIGHT_n4), 
        .ZN(alu_ex_SHIFTER_LEFTORRIGHT_n3) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_U2 ( .A(alu_ex_SHIFTER_LEFTORRIGHT_n4), 
        .ZN(alu_ex_SHIFTER_LEFTORRIGHT_n1) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_U1 ( .A(alu_ex_SHIFTER_LEFTORRIGHT_n4), 
        .ZN(alu_ex_SHIFTER_LEFTORRIGHT_n2) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_0__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_0__MUX_n4), .ZN(
        alu_ex_shift_out_0_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_0__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_0__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[0]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_0__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[0]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_0__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_1__MUX_n4), .ZN(
        alu_ex_shift_out_1_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_1__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_1__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[1]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_1__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[1]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_1__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_2__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_2__MUX_n4), .ZN(
        alu_ex_shift_out_2_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_2__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_2__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[2]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_2__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[2]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_2__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_3__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_3__MUX_n4), .ZN(
        alu_ex_shift_out_3_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_3__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_3__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[3]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_3__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[3]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_3__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_4__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_4__MUX_n4), .ZN(
        alu_ex_shift_out_4_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_4__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_4__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[4]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_4__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[4]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_4__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_5__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_5__MUX_n4), .ZN(
        alu_ex_shift_out_5_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_5__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_5__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[5]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_5__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[5]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_5__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_6__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_6__MUX_n4), .ZN(
        alu_ex_shift_out_6_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_6__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_6__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[6]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_6__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[6]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_6__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_7__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_7__MUX_n4), .ZN(
        alu_ex_shift_out_7_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_7__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_7__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[7]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_7__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[7]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_7__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_8__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_8__MUX_n4), .ZN(
        alu_ex_shift_out_8_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_8__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_8__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[8]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_8__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[8]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_8__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_9__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_9__MUX_n4), .ZN(
        alu_ex_shift_out_9_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_9__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_9__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[9]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_9__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[9]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_9__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_10__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_10__MUX_n4), .ZN(
        alu_ex_shift_out_10_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_10__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_10__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_10__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[10]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_10__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[10]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_10__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_11__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_11__MUX_n4), .ZN(
        alu_ex_shift_out_11_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_11__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_11__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_11__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[11]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_11__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[11]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n1), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_11__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_12__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_12__MUX_n4), .ZN(
        alu_ex_shift_out_12_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_12__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_12__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_12__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[12]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_12__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[12]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_12__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_13__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_13__MUX_n4), .ZN(
        alu_ex_shift_out_13_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_13__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_13__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_13__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[13]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_13__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[13]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_13__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_14__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_14__MUX_n4), .ZN(
        alu_ex_shift_out_14_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_14__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_14__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_14__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[14]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_14__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[14]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_14__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_15__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_15__MUX_n4), .ZN(
        alu_ex_shift_out_15_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_15__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_15__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_15__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[15]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_15__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[15]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_15__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_16__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_16__MUX_n4), .ZN(
        alu_ex_shift_out_16_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_16__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_16__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_16__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[16]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_16__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[16]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_16__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_17__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_17__MUX_n4), .ZN(
        alu_ex_shift_out_17_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_17__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_17__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_17__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[17]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_17__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[17]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_17__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_18__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_18__MUX_n4), .ZN(
        alu_ex_shift_out_18_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_18__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_18__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_18__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[18]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_18__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[18]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_18__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_19__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_19__MUX_n4), .ZN(
        alu_ex_shift_out_19_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_19__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_19__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_19__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[19]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_19__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[19]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_19__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_20__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_20__MUX_n4), .ZN(
        alu_ex_shift_out_20_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_20__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_20__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_20__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[20]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_20__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[20]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_20__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_21__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_21__MUX_n4), .ZN(
        alu_ex_shift_out_21_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_21__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_21__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_21__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[21]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_21__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[21]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_21__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_22__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_22__MUX_n4), .ZN(
        alu_ex_shift_out_22_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_22__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_22__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_22__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[22]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_22__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[22]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_22__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_23__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_23__MUX_n4), .ZN(
        alu_ex_shift_out_23_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_23__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_23__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_23__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[23]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_23__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[23]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n2), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_23__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_24__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_24__MUX_n4), .ZN(
        alu_ex_shift_out_24_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_24__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_24__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_24__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[24]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_24__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[24]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_24__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_25__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_25__MUX_n4), .ZN(
        alu_ex_shift_out_25_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_25__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_25__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_25__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[25]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_25__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[25]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_25__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_26__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_26__MUX_n4), .ZN(
        alu_ex_shift_out_26_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_26__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_26__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_26__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[26]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_26__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[26]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_26__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_27__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_27__MUX_n4), .ZN(
        alu_ex_shift_out_27_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_27__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_27__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_27__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[27]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_27__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[27]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_27__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_28__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_28__MUX_n4), .ZN(
        alu_ex_shift_out_28_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_28__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_28__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_28__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[28]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_28__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[28]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_28__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_29__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_29__MUX_n4), .ZN(
        alu_ex_shift_out_29_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_29__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_29__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_29__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[29]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_29__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[29]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_29__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_30__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_30__MUX_n4), .ZN(
        alu_ex_shift_out_30_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_30__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_30__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_30__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[30]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_30__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[30]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_30__MUX_n4) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_31__MUX_U3 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_31__MUX_n4), .ZN(
        alu_ex_shift_out_31_) );
  INV_X4 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_31__MUX_U2 ( .A(
        alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_31__MUX_n1) );
  AOI22_X2 alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_31__MUX_U1 ( .A1(
        alu_ex_SHIFTER_ltemp4[31]), .A2(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_31__MUX_n1), .B1(
        alu_ex_SHIFTER_rtemp4[31]), .B2(alu_ex_SHIFTER_LEFTORRIGHT_n3), .ZN(
        alu_ex_SHIFTER_LEFTORRIGHT_MUX2TO1_32BIT_31__MUX_n4) );
  INV_X4 alu_ex_SET_FLAGS_U13 ( .A(alu_ex_n3), .ZN(alu_ex_sne_1bit) );
  BUF_X4 alu_ex_SET_FLAGS_U11 ( .A(alu_ex_sne_1bit), .Z(alu_ex_SET_FLAGS_n2)
         );
  NAND2_X2 alu_ex_SET_FLAGS_U8 ( .A1(alu_ex_SET_FLAGS_n2), .A2(alu_ex_sge_1bit), .ZN(alu_ex_sle_1bit) );
  NAND2_X2 alu_ex_SET_FLAGS_U7 ( .A1(alu_ex_SET_FLAGS_n5), .A2(
        alu_ex_SET_FLAGS_n6), .ZN(alu_ex_sge_1bit) );
  NAND2_X2 alu_ex_SET_FLAGS_U3 ( .A1(alu_ex_SET_FLAGS_difference_0_), .A2(
        alu_ex_SET_FLAGS_sub_of), .ZN(alu_ex_SET_FLAGS_n5) );
  NAND2_X4 alu_ex_SET_FLAGS_U12 ( .A1(alu_ex_SET_FLAGS_n5), .A2(
        alu_ex_SET_FLAGS_n6), .ZN(alu_ex_SET_FLAGS_n12) );
  NAND2_X4 alu_ex_SET_FLAGS_U10 ( .A1(alu_ex_SET_FLAGS_n3), .A2(
        alu_ex_SET_FLAGS_n4), .ZN(alu_ex_SET_FLAGS_n6) );
  NOR2_X4 alu_ex_SET_FLAGS_U9 ( .A1(alu_ex_slt_1bit), .A2(alu_ex_SET_FLAGS_n1), 
        .ZN(alu_ex_sgt_1bit) );
  INV_X4 alu_ex_SET_FLAGS_U6 ( .A(alu_ex_SET_FLAGS_sub_of), .ZN(
        alu_ex_SET_FLAGS_n3) );
  INV_X8 alu_ex_SET_FLAGS_U5 ( .A(alu_ex_SET_FLAGS_n12), .ZN(alu_ex_slt_1bit)
         );
  INV_X1 alu_ex_SET_FLAGS_U4 ( .A(alu_ex_sne_1bit), .ZN(alu_ex_SET_FLAGS_n1)
         );
  INV_X2 alu_ex_SET_FLAGS_U2 ( .A(alu_ex_SET_FLAGS_difference_0_), .ZN(
        alu_ex_SET_FLAGS_n4) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_0__NOT_1_U1 ( .A(opB_in[0]), .ZN(
        alu_ex_SET_FLAGS_b_not[0]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_1__NOT_1_U1 ( .A(opB_in[1]), .ZN(
        alu_ex_SET_FLAGS_b_not[1]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_2__NOT_1_U1 ( .A(opB_in[2]), .ZN(
        alu_ex_SET_FLAGS_b_not[2]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_3__NOT_1_U1 ( .A(opB_in[3]), .ZN(
        alu_ex_SET_FLAGS_b_not[3]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_4__NOT_1_U1 ( .A(opB_in[4]), .ZN(
        alu_ex_SET_FLAGS_b_not[4]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_5__NOT_1_U1 ( .A(opB_in[5]), .ZN(
        alu_ex_SET_FLAGS_b_not[5]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_6__NOT_1_U1 ( .A(opB_in[6]), .ZN(
        alu_ex_SET_FLAGS_b_not[6]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_7__NOT_1_U1 ( .A(opB_in[7]), .ZN(
        alu_ex_SET_FLAGS_b_not[7]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_8__NOT_1_U1 ( .A(opB_in[8]), .ZN(
        alu_ex_SET_FLAGS_b_not[8]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_9__NOT_1_U1 ( .A(opB_in[9]), .ZN(
        alu_ex_SET_FLAGS_b_not[9]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_10__NOT_1_U1 ( .A(opB_in[10]), 
        .ZN(alu_ex_SET_FLAGS_b_not[10]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_11__NOT_1_U1 ( .A(opB_in[11]), 
        .ZN(alu_ex_SET_FLAGS_b_not[11]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_12__NOT_1_U1 ( .A(opB_in[12]), 
        .ZN(alu_ex_SET_FLAGS_b_not[12]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_13__NOT_1_U1 ( .A(opB_in[13]), 
        .ZN(alu_ex_SET_FLAGS_b_not[13]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_14__NOT_1_U1 ( .A(opB_in[14]), 
        .ZN(alu_ex_SET_FLAGS_b_not[14]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_15__NOT_1_U1 ( .A(opB_in[15]), 
        .ZN(alu_ex_SET_FLAGS_b_not[15]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_16__NOT_1_U1 ( .A(opB_in[16]), 
        .ZN(alu_ex_SET_FLAGS_b_not[16]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_17__NOT_1_U1 ( .A(opB_in[17]), 
        .ZN(alu_ex_SET_FLAGS_b_not[17]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_18__NOT_1_U1 ( .A(opB_in[18]), 
        .ZN(alu_ex_SET_FLAGS_b_not[18]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_19__NOT_1_U1 ( .A(opB_in[19]), 
        .ZN(alu_ex_SET_FLAGS_b_not[19]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_20__NOT_1_U1 ( .A(opB_in[20]), 
        .ZN(alu_ex_SET_FLAGS_b_not[20]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_21__NOT_1_U1 ( .A(opB_in[21]), 
        .ZN(alu_ex_SET_FLAGS_b_not[21]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_22__NOT_1_U1 ( .A(opB_in[22]), 
        .ZN(alu_ex_SET_FLAGS_b_not[22]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_23__NOT_1_U1 ( .A(opB_in[23]), 
        .ZN(alu_ex_SET_FLAGS_b_not[23]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_24__NOT_1_U1 ( .A(opB_in[24]), 
        .ZN(alu_ex_SET_FLAGS_b_not[24]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_25__NOT_1_U1 ( .A(opB_in[25]), 
        .ZN(alu_ex_SET_FLAGS_b_not[25]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_26__NOT_1_U1 ( .A(opB_in[26]), 
        .ZN(alu_ex_SET_FLAGS_b_not[26]) );
  INV_X4 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_27__NOT_1_U1 ( .A(opB_in[27]), 
        .ZN(alu_ex_SET_FLAGS_b_not[27]) );
  INV_X32 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_28__NOT_1_U1 ( .A(opB_in[28]), 
        .ZN(alu_ex_SET_FLAGS_b_not[28]) );
  INV_X32 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_29__NOT_1_U1 ( .A(opB_in[29]), 
        .ZN(alu_ex_SET_FLAGS_b_not[29]) );
  INV_X32 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_30__NOT_1_U1 ( .A(opB_in[30]), 
        .ZN(alu_ex_SET_FLAGS_b_not[30]) );
  INV_X32 alu_ex_SET_FLAGS_NEGATE_B_NOT_32BIT_31__NOT_1_U1 ( .A(opB_in[31]), 
        .ZN(alu_ex_SET_FLAGS_b_not[31]) );
  INV_X2 alu_ex_SET_FLAGS_FULL_ADDER_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_1_), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_n1) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_U6 ( .A(alu_ex_SET_FLAGS_FULL_ADDER_n1), 
        .ZN(alu_ex_SET_FLAGS_FULL_ADDER_n5) );
  INV_X8 alu_ex_SET_FLAGS_FULL_ADDER_U5 ( .A(alu_ex_SET_FLAGS_FULL_ADDER_n3), 
        .ZN(alu_ex_SET_FLAGS_FULL_ADDER_n4) );
  NAND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_U4 ( .A1(alu_ex_SET_FLAGS_FULL_ADDER_n6), .A2(alu_ex_SET_FLAGS_FULL_ADDER_n7), .ZN(alu_ex_SET_FLAGS_sub_of) );
  NAND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_U2 ( .A1(alu_ex_SET_FLAGS_FULL_ADDER_n4), .A2(alu_ex_SET_FLAGS_FULL_ADDER_n5), .ZN(alu_ex_SET_FLAGS_FULL_ADDER_n7) );
  NAND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_U1 ( .A1(alu_ex_SET_FLAGS_FULL_ADDER_n3), .A2(alu_ex_SET_FLAGS_FULL_ADDER_n1), .ZN(alu_ex_SET_FLAGS_FULL_ADDER_n6) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_U13 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n15), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n5) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_U6 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n10), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n14) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_U5 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n3), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n14), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n15) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_U4 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n10), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n12) );
  AOI21_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_U3 ( .B1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_1_), .B2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n12), .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n7), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n13) );
  INV_X8 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n13), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_n3) );
  INV_X8 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_U1 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_1_), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_U12 ( .A(
        alu_ex_SET_FLAGS_b_not[0]), .B(opA_in[0]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n10) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_U11 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n8), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n7) );
  NAND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_U10 ( .A1(
        alu_ex_SET_FLAGS_b_not[0]), .A2(opA_in[0]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n8) );
  INV_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_U9 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n10), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n4) );
  NAND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_0_) );
  NAND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_U7 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n3), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_0__FA_n6) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_U7 ( .A(
        alu_ex_SET_FLAGS_b_not[1]), .B(opA_in[1]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n5) );
  NAND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_U6 ( .A1(
        alu_ex_SET_FLAGS_b_not[1]), .A2(opA_in[1]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n4) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_2_), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n5), .ZN(
        alu_ex_SET_FLAGS_difference_1_) );
  INV_X8 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_U4 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n2), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_1_) );
  OAI21_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_U3 ( .B1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_2_), .B2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n3), .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n2) );
  NAND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_U2 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n1) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_U1 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_1__FA_n3) );
  INV_X8 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_U8 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n2) );
  INV_X8 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n8), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_2_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n7) );
  OAI21_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_U2 ( .B1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_3_), .B2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n2), .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n7), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n8) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_U1 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_3_), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n5), .ZN(
        alu_ex_SET_FLAGS_difference_2_) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_U6 ( .A(
        alu_ex_SET_FLAGS_b_not[2]), .B(opA_in[2]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n5) );
  NAND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_b_not[2]), .A2(opA_in[2]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n3) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_2__FA_n1) );
  INV_X8 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_U9 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n3) );
  INV_X8 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_U8 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n9), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_3_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_U6 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n2), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n8) );
  OAI21_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_U5 ( .B1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_4_), .B2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n3), .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n8), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n9) );
  BUF_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_4_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n1) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_U7 ( .A(
        alu_ex_SET_FLAGS_b_not[3]), .B(opA_in[3]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n6) );
  NAND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_b_not[3]), .A2(opA_in[3]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n4) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n6), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n2) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_U1 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n1), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_3__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_3_) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_U9 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n6), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_4_) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_U8 ( .A(
        alu_ex_SET_FLAGS_b_not[4]), .B(opA_in[4]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n7) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n5), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n4) );
  NAND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_U6 ( .A1(
        alu_ex_SET_FLAGS_b_not[4]), .A2(opA_in[4]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n5) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n7), .ZN(
        alu_ex_SET_FLAGS_difference_4_) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n7), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n5), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n3) );
  INV_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_U3 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n2) );
  INV_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_5_), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_5_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_4__FA_n6) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n2), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_5_) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_U7 ( .A(
        alu_ex_SET_FLAGS_b_not[5]), .B(opA_in[5]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n6) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_U6 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_6_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n5) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n3) );
  NAND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_b_not[5]), .A2(opA_in[5]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n4) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_U3 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n1), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_5_) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_U2 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n6), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n2) );
  BUF_X16 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_U1 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_6_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_5__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n2), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_6_) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_U7 ( .A(
        alu_ex_SET_FLAGS_b_not[6]), .B(opA_in[6]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n6) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_U6 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_7_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n5) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n3) );
  NAND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_b_not[6]), .A2(opA_in[6]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n4) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n6), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n2) );
  BUF_X16 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_7_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n1) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_U1 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n1), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_6__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_6_) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_U10 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n10), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_7_) );
  INV_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_U9 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n9), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n10) );
  INV_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n8), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n9) );
  BUF_X16 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_U1 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_8_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n8) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n2), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_7_) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_U7 ( .A(
        alu_ex_SET_FLAGS_b_not[7]), .B(opA_in[7]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n6) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_U6 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_8_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n5) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n3) );
  NAND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_b_not[7]), .A2(opA_in[7]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n4) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n6), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_7__FA_n2) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_U8 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n9) );
  INV_X8 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_U6 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n3) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_U3 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n8), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_8_) );
  AOI21_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_U2 ( .B1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_9_), .B2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n9), .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n8) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_U7 ( .A(
        alu_ex_SET_FLAGS_b_not[8]), .B(opA_in[8]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n6) );
  NAND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_U5 ( .A1(
        alu_ex_SET_FLAGS_b_not[8]), .A2(opA_in[8]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n4) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_U4 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n1), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_8_) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_U1 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_9_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_8__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n2), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_9_) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_U7 ( .A(
        alu_ex_SET_FLAGS_b_not[9]), .B(opA_in[9]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n6) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_U6 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n3) );
  NAND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_U5 ( .A1(
        alu_ex_SET_FLAGS_b_not[9]), .A2(opA_in[9]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n4) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_U4 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n1), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_9_) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n6), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n2) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_U2 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_10_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n5) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_U1 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_10_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_9__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n2), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_10_) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_U7 ( .A(
        alu_ex_SET_FLAGS_b_not[10]), .B(opA_in[10]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n6) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_U6 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_11_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n5) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n3) );
  NAND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_b_not[10]), .A2(opA_in[10]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n4) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_U3 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n1), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_10_) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_U2 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n6), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n2) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_U1 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_11_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_10__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_11_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_U6 ( .A(
        alu_ex_SET_FLAGS_b_not[11]), .B(opA_in[11]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n6) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_U5 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_12_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n5) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_U4 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_11_) );
  NOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n4) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_12_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n2) );
  AND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[11]), .A2(opA_in[11]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_11__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_12_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_U6 ( .A(
        alu_ex_SET_FLAGS_b_not[12]), .B(opA_in[12]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n6) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_U5 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_13_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n5) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_U4 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_12_) );
  NOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n4) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_13_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n2) );
  AND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[12]), .A2(opA_in[12]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_12__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_13_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_U6 ( .A(
        alu_ex_SET_FLAGS_b_not[13]), .B(opA_in[13]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n6) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_U5 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_14_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n5) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_U4 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_13_) );
  NOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n4) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_14_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n2) );
  AND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[13]), .A2(opA_in[13]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_13__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_14_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_U6 ( .A(
        alu_ex_SET_FLAGS_b_not[14]), .B(opA_in[14]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n6) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_U5 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_15_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n5) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_U4 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_14_) );
  NOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n4) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_15_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n2) );
  AND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[14]), .A2(opA_in[14]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_14__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_U9 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n6), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n5), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_15_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_U8 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n7), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n4) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_U7 ( .A(
        alu_ex_SET_FLAGS_b_not[15]), .B(opA_in[15]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n7) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_U6 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_16_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n6) );
  INV_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n2), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n3) );
  XOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_U4 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n3), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n7), .Z(
        alu_ex_SET_FLAGS_difference_15_) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_U3 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_16_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n2) );
  AND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_U2 ( .A1(
        alu_ex_SET_FLAGS_b_not[15]), .A2(opA_in[15]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n1) );
  NOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_15__FA_n5) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_16_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_U6 ( .A(
        alu_ex_SET_FLAGS_b_not[16]), .B(opA_in[16]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n6) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_16_) );
  NOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n4) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_17_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n5) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_17_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n2) );
  AND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[16]), .A2(opA_in[16]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_16__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_17_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_U6 ( .A(
        alu_ex_SET_FLAGS_b_not[17]), .B(opA_in[17]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n6) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_17_) );
  NOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n4) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_18_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n5) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_18_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n2) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[17]), .A2(opA_in[17]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_17__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_18_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_U6 ( .A(
        alu_ex_SET_FLAGS_b_not[18]), .B(opA_in[18]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n6) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_18_) );
  NOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n4) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_19_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n5) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_19_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n2) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[18]), .A2(opA_in[18]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_18__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_19_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_U6 ( .A(
        alu_ex_SET_FLAGS_b_not[19]), .B(opA_in[19]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n6) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_19_) );
  NOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n4) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_20_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n5) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_20_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n2) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[19]), .A2(opA_in[19]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_19__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_20_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_U6 ( .A(
        alu_ex_SET_FLAGS_b_not[20]), .B(opA_in[20]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n6) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_20_) );
  NOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n4) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_21_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n5) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_21_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n2) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[20]), .A2(opA_in[20]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_20__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_21_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_U6 ( .A(
        alu_ex_SET_FLAGS_b_not[21]), .B(opA_in[21]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n6) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_21_) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n4) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_22_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n5) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_22_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n2) );
  AND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[21]), .A2(opA_in[21]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_21__FA_n1) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_U8 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_U7 ( .A(
        alu_ex_SET_FLAGS_b_not[22]), .B(opA_in[22]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n6) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_U6 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_22_) );
  NOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_U5 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n4) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_23_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n5) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_22_) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_23_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n2) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[22]), .A2(opA_in[22]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_22__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_23_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_U6 ( .A(
        alu_ex_SET_FLAGS_b_not[23]), .B(opA_in[23]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n6) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_23_) );
  NOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n4) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_24_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n5) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_24_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n2) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[23]), .A2(opA_in[23]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_23__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_24_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_U6 ( .A(
        alu_ex_SET_FLAGS_b_not[24]), .B(opA_in[24]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n6) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_24_) );
  NOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n4) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_25_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n5) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_25_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n2) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[24]), .A2(opA_in[24]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_24__FA_n1) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_U8 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_U7 ( .A(
        alu_ex_SET_FLAGS_b_not[25]), .B(opA_in[25]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n6) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_U6 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_25_) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_U5 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n4) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_25_) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_26_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n5) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_26_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n2) );
  AND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[25]), .A2(opA_in[25]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_25__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_26_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_U6 ( .A(
        alu_ex_SET_FLAGS_b_not[26]), .B(opA_in[26]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n6) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_26_) );
  NOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n4) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_27_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n5) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_27_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n2) );
  AND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[26]), .A2(opA_in[26]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_26__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_27_) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_U6 ( .A(
        alu_ex_SET_FLAGS_b_not[27]), .B(opA_in[27]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n6) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_27_) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n4) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_28_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n5) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_28_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n2) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[27]), .A2(opA_in[27]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_27__FA_n1) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_U5 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n1), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n4) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_U8 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n3) );
  XNOR2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_U7 ( .A(
        alu_ex_SET_FLAGS_b_not[28]), .B(opA_in[28]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n6) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_U6 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n6), .ZN(
        alu_ex_SET_FLAGS_difference_28_) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_29_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n5) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n4), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_28_) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_29_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n2) );
  AND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[28]), .A2(opA_in[28]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_28__FA_n1) );
  INV_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_U9 ( .A(opA_in[29]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n7) );
  INV_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_U3 ( .A(
        alu_ex_SET_FLAGS_b_not[29]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n3) );
  AND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_U2 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n3), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n7), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n8) );
  AND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_U1 ( .A1(
        alu_ex_SET_FLAGS_b_not[29]), .A2(opA_in[29]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n1) );
  XNOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_U12 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n2), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n10), .ZN(
        alu_ex_SET_FLAGS_difference_29_) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_U11 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_30_), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n1), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n9) );
  INV_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_U10 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n6), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n10) );
  NAND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_U8 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n3), .A2(opA_in[29]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n5) );
  NAND2_X2 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_U7 ( .A1(
        alu_ex_SET_FLAGS_b_not[29]), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n7), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n4) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_U6 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n9), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n8), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_29_) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_30_), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n2) );
  NAND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n4), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n5), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_29__FA_n6) );
  OAI21_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_U10 ( .B1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n8), .B2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n13), .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n9), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_30_) );
  INV_X8 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_U9 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_31_), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n8) );
  INV_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_U7 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n12), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n14) );
  NAND2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_U6 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n6), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n9), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n10) );
  NOR2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_U4 ( .A1(
        alu_ex_SET_FLAGS_b_not[30]), .A2(opA_in[30]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n13) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_U2 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n8), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n12) );
  INV_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_U1 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n13), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n6) );
  INV_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_U11 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n3), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n7) );
  XOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_U8 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n14), .B(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n7), .Z(
        alu_ex_SET_FLAGS_difference_30_) );
  BUF_X32 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_U5 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n10), .Z(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n3) );
  NAND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_U3 ( .A1(
        alu_ex_SET_FLAGS_b_not[30]), .A2(opA_in[30]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_30__FA_n9) );
  NAND2_X4 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_31__FA_U5 ( .A1(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_31__FA_n5), .A2(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_31__FA_n2), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_carry_31_) );
  XOR2_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_31__FA_U4 ( .A(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_31__FA_n1), .B(opA_in[31]), .Z(
        alu_ex_SET_FLAGS_difference_31_) );
  INV_X1 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_31__FA_U3 ( .A(
        alu_ex_SET_FLAGS_b_not[31]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_31__FA_n1) );
  INV_X16 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_31__FA_U2 ( .A(
        alu_ex_SET_FLAGS_b_not[31]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_31__FA_n5) );
  INV_X8 alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_31__FA_U1 ( .A(opA_in[31]), .ZN(
        alu_ex_SET_FLAGS_FULL_ADDER_FA_NBIT_31__FA_n2) );
  NOR2_X2 alu_ex_SET_FLAGS_CHECK_EQ_U16 ( .A1(alu_ex_SET_FLAGS_difference_3_), 
        .A2(alu_ex_SET_FLAGS_difference_4_), .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n9)
         );
  NAND4_X2 alu_ex_SET_FLAGS_CHECK_EQ_U2 ( .A1(alu_ex_SET_FLAGS_CHECK_EQ_n9), 
        .A2(alu_ex_SET_FLAGS_CHECK_EQ_n8), .A3(alu_ex_SET_FLAGS_CHECK_EQ_n7), 
        .A4(alu_ex_SET_FLAGS_CHECK_EQ_n6), .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n16)
         );
  NAND4_X2 alu_ex_SET_FLAGS_CHECK_EQ_U20 ( .A1(alu_ex_SET_FLAGS_CHECK_EQ_n14), 
        .A2(alu_ex_SET_FLAGS_CHECK_EQ_n13), .A3(alu_ex_SET_FLAGS_CHECK_EQ_n12), 
        .A4(alu_ex_SET_FLAGS_CHECK_EQ_n11), .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n15)
         );
  NOR4_X2 alu_ex_SET_FLAGS_CHECK_EQ_U19 ( .A1(alu_ex_SET_FLAGS_CHECK_EQ_n10), 
        .A2(alu_ex_SET_FLAGS_CHECK_EQ_n4), .A3(alu_ex_SET_FLAGS_difference_24_), .A4(alu_ex_SET_FLAGS_difference_25_), .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n11) );
  NOR4_X2 alu_ex_SET_FLAGS_CHECK_EQ_U18 ( .A1(alu_ex_SET_FLAGS_difference_20_), 
        .A2(alu_ex_SET_FLAGS_difference_21_), .A3(
        alu_ex_SET_FLAGS_difference_22_), .A4(alu_ex_SET_FLAGS_difference_23_), 
        .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n12) );
  INV_X4 alu_ex_SET_FLAGS_CHECK_EQ_U17 ( .A(alu_ex_SET_FLAGS_difference_17_), 
        .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n13) );
  NOR4_X2 alu_ex_SET_FLAGS_CHECK_EQ_U15 ( .A1(alu_ex_SET_FLAGS_CHECK_EQ_n5), 
        .A2(alu_ex_SET_FLAGS_CHECK_EQ_n2), .A3(alu_ex_SET_FLAGS_difference_9_), 
        .A4(alu_ex_SET_FLAGS_difference_10_), .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n6) );
  INV_X2 alu_ex_SET_FLAGS_CHECK_EQ_U14 ( .A(alu_ex_SET_FLAGS_difference_2_), 
        .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n8) );
  INV_X2 alu_ex_SET_FLAGS_CHECK_EQ_U13 ( .A(alu_ex_SET_FLAGS_difference_1_), 
        .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n17) );
  OR2_X2 alu_ex_SET_FLAGS_CHECK_EQ_U12 ( .A1(alu_ex_SET_FLAGS_difference_26_), 
        .A2(alu_ex_SET_FLAGS_difference_27_), .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n4) );
  OR2_X4 alu_ex_SET_FLAGS_CHECK_EQ_U11 ( .A1(alu_ex_SET_FLAGS_difference_30_), 
        .A2(alu_ex_SET_FLAGS_difference_31_), .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n3) );
  OR3_X2 alu_ex_SET_FLAGS_CHECK_EQ_U10 ( .A1(alu_ex_SET_FLAGS_difference_29_), 
        .A2(alu_ex_SET_FLAGS_difference_28_), .A3(alu_ex_SET_FLAGS_CHECK_EQ_n3), .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n10) );
  OR2_X2 alu_ex_SET_FLAGS_CHECK_EQ_U9 ( .A1(alu_ex_SET_FLAGS_difference_11_), 
        .A2(alu_ex_SET_FLAGS_difference_12_), .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n2) );
  OR2_X4 alu_ex_SET_FLAGS_CHECK_EQ_U8 ( .A1(alu_ex_SET_FLAGS_difference_15_), 
        .A2(alu_ex_SET_FLAGS_difference_16_), .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n1) );
  OR3_X2 alu_ex_SET_FLAGS_CHECK_EQ_U7 ( .A1(alu_ex_SET_FLAGS_difference_14_), 
        .A2(alu_ex_SET_FLAGS_difference_13_), .A3(alu_ex_SET_FLAGS_CHECK_EQ_n1), .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n5) );
  NOR2_X2 alu_ex_SET_FLAGS_CHECK_EQ_U6 ( .A1(alu_ex_SET_FLAGS_difference_18_), 
        .A2(alu_ex_SET_FLAGS_difference_19_), .ZN(
        alu_ex_SET_FLAGS_CHECK_EQ_n14) );
  NOR2_X4 alu_ex_SET_FLAGS_CHECK_EQ_U5 ( .A1(alu_ex_SET_FLAGS_difference_0_), 
        .A2(alu_ex_SET_FLAGS_CHECK_EQ_n19), .ZN(alu_ex_n3) );
  NOR2_X4 alu_ex_SET_FLAGS_CHECK_EQ_U4 ( .A1(alu_ex_SET_FLAGS_CHECK_EQ_n16), 
        .A2(alu_ex_SET_FLAGS_CHECK_EQ_n15), .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n18)
         );
  NAND2_X4 alu_ex_SET_FLAGS_CHECK_EQ_U3 ( .A1(alu_ex_SET_FLAGS_CHECK_EQ_n18), 
        .A2(alu_ex_SET_FLAGS_CHECK_EQ_n17), .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n19)
         );
  NOR4_X2 alu_ex_SET_FLAGS_CHECK_EQ_U1 ( .A1(alu_ex_SET_FLAGS_difference_5_), 
        .A2(alu_ex_SET_FLAGS_difference_6_), .A3(
        alu_ex_SET_FLAGS_difference_7_), .A4(alu_ex_SET_FLAGS_difference_8_), 
        .ZN(alu_ex_SET_FLAGS_CHECK_EQ_n7) );
  INV_X8 alu_ex_EXTEND_SEQ_U2 ( .A(alu_ex_n3), .ZN(alu_ex_EXTEND_SEQ_n1) );
  INV_X4 alu_ex_EXTEND_SEQ_U1 ( .A(alu_ex_EXTEND_SEQ_n1), .ZN(
        alu_ex_seq_out_31_) );
  INV_X2 alu_ex_EXTEND_SNE_U2 ( .A(alu_ex_EXTEND_SNE_n1), .ZN(
        alu_ex_sne_out_31_) );
  INV_X2 alu_ex_EXTEND_SNE_U1 ( .A(alu_ex_sne_1bit), .ZN(alu_ex_EXTEND_SNE_n1)
         );
  INV_X4 alu_ex_EXTEND_SLE_U2 ( .A(alu_ex_sle_1bit), .ZN(alu_ex_EXTEND_SLE_n1)
         );
  INV_X4 alu_ex_EXTEND_SLE_U1 ( .A(alu_ex_EXTEND_SLE_n1), .ZN(
        alu_ex_sle_out_31_) );
  INV_X4 alu_ex_EXTEND_SLT_U2 ( .A(alu_ex_slt_1bit), .ZN(alu_ex_EXTEND_SLT_n1)
         );
  INV_X4 alu_ex_EXTEND_SLT_U1 ( .A(alu_ex_EXTEND_SLT_n1), .ZN(
        alu_ex_slt_out_31_) );
  INV_X2 alu_ex_EXTEND_SGE_U2 ( .A(alu_ex_EXTEND_SGE_n1), .ZN(
        alu_ex_sge_out_31_) );
  INV_X1 alu_ex_EXTEND_SGE_U1 ( .A(alu_ex_sge_1bit), .ZN(alu_ex_EXTEND_SGE_n1)
         );
  INV_X4 alu_ex_EXTEND_SGT_U2 ( .A(alu_ex_sgt_1bit), .ZN(alu_ex_EXTEND_SGT_n1)
         );
  INV_X8 alu_ex_EXTEND_SGT_U1 ( .A(alu_ex_EXTEND_SGT_n1), .ZN(
        alu_ex_sgt_out_31_) );
  INV_X1 alu_ex_FINAL_MUX_U2 ( .A(ALUCtrl_in[3]), .ZN(alu_ex_FINAL_MUX_n2) );
  INV_X4 alu_ex_FINAL_MUX_U1 ( .A(alu_ex_FINAL_MUX_n2), .ZN(
        alu_ex_FINAL_MUX_n1) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_U4 ( .A(
        alu_ex_FINAL_MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n2) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1) );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_U4 ( 
        .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_n3), 
        .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[0]) );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_U3 ( 
        .A1(alu_ex_add_sub_out_0_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_n1), 
        .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_n2)
         );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n2), .A2(
        alu_ex_add_sub_out_0_), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_n3)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_n1)
         );
  MUX2_X1 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_1__MUX_U1 ( 
        .A(alu_ex_add_sub_out_1_), .B(alu_ex_add_sub_out_1_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[1]) );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_U4 ( 
        .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_n3), 
        .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[2]) );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_U3 ( 
        .A1(alu_ex_add_sub_out_2_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_n1), 
        .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_n2)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_n1)
         );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_U1 ( 
        .A1(alu_ex_add_sub_out_2_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_n3)
         );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_3__MUX_U1 ( 
        .A(alu_ex_add_sub_out_3_), .B(alu_ex_add_sub_out_3_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[3]) );
  MUX2_X1 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_4__MUX_U1 ( 
        .A(alu_ex_add_sub_out_4_), .B(alu_ex_add_sub_out_4_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[4]) );
  MUX2_X1 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_5__MUX_U1 ( 
        .A(alu_ex_add_sub_out_5_), .B(alu_ex_add_sub_out_5_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[5]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_6__MUX_U1 ( 
        .A(alu_ex_add_sub_out_6_), .B(alu_ex_add_sub_out_6_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[6]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_7__MUX_U1 ( 
        .A(alu_ex_add_sub_out_7_), .B(alu_ex_add_sub_out_7_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[7]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_8__MUX_U1 ( 
        .A(alu_ex_add_sub_out_8_), .B(alu_ex_add_sub_out_8_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[8]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_9__MUX_U1 ( 
        .A(alu_ex_add_sub_out_9_), .B(alu_ex_add_sub_out_9_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[9]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_10__MUX_U1 ( 
        .A(alu_ex_add_sub_out_10_), .B(alu_ex_add_sub_out_10_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[10]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_11__MUX_U1 ( 
        .A(alu_ex_add_sub_out_11_), .B(alu_ex_add_sub_out_11_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[11]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_12__MUX_U1 ( 
        .A(alu_ex_add_sub_out_12_), .B(alu_ex_add_sub_out_12_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[12]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_13__MUX_U1 ( 
        .A(alu_ex_add_sub_out_13_), .B(alu_ex_add_sub_out_13_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[13]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_14__MUX_U1 ( 
        .A(alu_ex_add_sub_out_14_), .B(alu_ex_add_sub_out_14_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[14]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_15__MUX_U1 ( 
        .A(alu_ex_add_sub_out_15_), .B(alu_ex_add_sub_out_15_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[15]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_16__MUX_U1 ( 
        .A(alu_ex_add_sub_out_16_), .B(alu_ex_add_sub_out_16_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[16]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_17__MUX_U1 ( 
        .A(alu_ex_add_sub_out_17_), .B(alu_ex_add_sub_out_17_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[17]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_18__MUX_U1 ( 
        .A(alu_ex_add_sub_out_18_), .B(alu_ex_add_sub_out_18_), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[18]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[19]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_U1 ( 
        .A1(alu_ex_add_sub_out_19_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_n1), 
        .B1(alu_ex_add_sub_out_19_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[20]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_U1 ( 
        .A1(alu_ex_add_sub_out_20_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_n1), 
        .B1(alu_ex_add_sub_out_20_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[21]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_U1 ( 
        .A1(alu_ex_add_sub_out_21_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_n1), 
        .B1(alu_ex_add_sub_out_21_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[22]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_U1 ( 
        .A1(alu_ex_add_sub_out_22_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_n1), 
        .B1(alu_ex_add_sub_out_22_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[23]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_U1 ( 
        .A1(alu_ex_add_sub_out_23_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_n1), 
        .B1(alu_ex_add_sub_out_23_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[24]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_U1 ( 
        .A1(alu_ex_add_sub_out_24_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_n1), 
        .B1(alu_ex_add_sub_out_24_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[25]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_U1 ( 
        .A1(alu_ex_add_sub_out_25_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_n1), 
        .B1(alu_ex_add_sub_out_25_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[26]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_U1 ( 
        .A1(alu_ex_add_sub_out_26_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_n1), 
        .B1(alu_ex_add_sub_out_26_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[27]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_U1 ( 
        .A1(alu_ex_add_sub_out_27_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_n1), 
        .B1(alu_ex_add_sub_out_27_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[28]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_U1 ( 
        .A1(alu_ex_add_sub_out_28_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_n1), 
        .B1(alu_ex_add_sub_out_28_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[29]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_U1 ( 
        .A1(alu_ex_add_sub_out_29_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_n1), 
        .B1(alu_ex_add_sub_out_29_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[30]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_U1 ( 
        .A1(alu_ex_add_sub_out_30_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_n1), 
        .B1(alu_ex_add_sub_out_30_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[31]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_U1 ( 
        .A1(alu_ex_add_sub_out_31_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n1), 
        .B1(alu_ex_add_sub_out_31_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n4)
         );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_U4 ( 
        .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n3), 
        .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus2_31_) );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_U1 ( 
        .A1(alu_ex_sle_out_31_), .A2(alu_ex_FINAL_MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n3)
         );
  NAND2_X1 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_U3 ( 
        .A1(alu_ex_slt_out_31_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n1), 
        .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n2)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n1)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_U6 ( .A(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n6) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_U5 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n6), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n5) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_U4 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n6), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n6), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n6), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n2) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n6), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n1) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_n2) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[0]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[0]) );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[1]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[1]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1) );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_2__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[2]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_2__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[2]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_2__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n5), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_2__MUX_n1) );
  NOR2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_3__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_3__MUX_n1), .A2(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[3]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_3__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[3]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_3__MUX_n1) );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_4__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[4]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_4__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[4]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_4__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_4__MUX_n1) );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_5__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[5]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_5__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[5]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_5__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_5__MUX_n1) );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_6__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[6]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_6__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[6]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_6__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n5), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_6__MUX_n1) );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_7__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[7]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_7__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[7]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_7__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_7__MUX_n1) );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_8__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[8]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_8__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[8]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_8__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_8__MUX_n1) );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_9__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[9]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_9__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[9]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_9__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n5), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_9__MUX_n1) );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_10__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[10]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_10__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[10]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_10__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_10__MUX_n1)
         );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_11__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[11]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_11__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[11]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_11__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_11__MUX_n1)
         );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_12__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[12]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_12__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[12]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_12__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n5), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_12__MUX_n1)
         );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_13__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[13]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_13__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[13]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_13__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_13__MUX_n1)
         );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_14__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[14]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_14__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[14]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_14__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_14__MUX_n1)
         );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_15__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[15]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_15__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[15]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_15__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n5), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_15__MUX_n1)
         );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_16__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[16]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_16__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[16]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_16__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_16__MUX_n1)
         );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_17__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[17]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_17__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[17]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_17__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_17__MUX_n1)
         );
  AND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_18__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[18]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_18__MUX_n1), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[18]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_18__MUX_U1 ( 
        .A(ALUCtrl_in[2]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_18__MUX_n1)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[19]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[19]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[20]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[20]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[21]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[21]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[22]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[22]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[23]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[23]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[24]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[24]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[25]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[25]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[26]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[26]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[27]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[27]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[28]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[28]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[29]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[29]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[30]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[30]) );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus2_31_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n3)
         );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_U4 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_bus1[31]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n1), 
        .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n2)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n1)
         );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_U2 ( 
        .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n3), 
        .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus1[31]) );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_U2 ( 
        .A1(alu_ex_sge_out_31_), .A2(alu_ex_FINAL_MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n2)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_U4 ( 
        .A(alu_ex_FINAL_MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n1)
         );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_U3 ( 
        .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n3), 
        .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus1_31_) );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_U1 ( 
        .A1(alu_ex_sgt_out_31_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n1), 
        .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n3)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_U4 ( .A(
        alu_ex_FINAL_MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[0]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_U1 ( 
        .A1(alu_ex_and_out_0_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_n1), 
        .B1(alu_ex_shift_out_0_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[1]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_U1 ( 
        .A1(alu_ex_and_out_1_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_n1), 
        .B1(alu_ex_shift_out_1_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[2]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_U1 ( 
        .A1(alu_ex_and_out_2_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_n1), 
        .B1(alu_ex_shift_out_2_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[3]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_U1 ( 
        .A1(alu_ex_and_out_3_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_n1), 
        .B1(alu_ex_shift_out_3_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[4]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_U1 ( 
        .A1(alu_ex_and_out_4_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_n1), 
        .B1(alu_ex_shift_out_4_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[5]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_U1 ( 
        .A1(alu_ex_and_out_5_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_n1), 
        .B1(alu_ex_shift_out_5_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[6]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_U1 ( 
        .A1(alu_ex_and_out_6_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_n1), 
        .B1(alu_ex_shift_out_6_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[7]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_U1 ( 
        .A1(alu_ex_and_out_7_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_n1), 
        .B1(alu_ex_shift_out_7_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[8]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_U1 ( 
        .A1(alu_ex_and_out_8_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_n1), 
        .B1(alu_ex_shift_out_8_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[9]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_U1 ( 
        .A1(alu_ex_and_out_9_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_n1), 
        .B1(alu_ex_shift_out_9_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[10]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_U1 ( 
        .A1(alu_ex_and_out_10_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_n1), 
        .B1(alu_ex_shift_out_10_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[11]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_U1 ( 
        .A1(alu_ex_and_out_11_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_n1), 
        .B1(alu_ex_shift_out_11_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[12]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_U1 ( 
        .A1(alu_ex_and_out_12_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_n1), 
        .B1(alu_ex_shift_out_12_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[13]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_U1 ( 
        .A1(alu_ex_and_out_13_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_n1), 
        .B1(alu_ex_shift_out_13_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[14]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_U1 ( 
        .A1(alu_ex_and_out_14_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_n1), 
        .B1(alu_ex_shift_out_14_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[15]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_U1 ( 
        .A1(alu_ex_and_out_15_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_n1), 
        .B1(alu_ex_shift_out_15_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[16]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_U1 ( 
        .A1(alu_ex_and_out_16_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_n1), 
        .B1(alu_ex_shift_out_16_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[17]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_U1 ( 
        .A1(alu_ex_and_out_17_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_n1), 
        .B1(alu_ex_shift_out_17_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[18]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_U1 ( 
        .A1(alu_ex_and_out_18_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_n1), 
        .B1(alu_ex_shift_out_18_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[19]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_U1 ( 
        .A1(alu_ex_and_out_19_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_n1), 
        .B1(alu_ex_shift_out_19_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[20]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_U1 ( 
        .A1(alu_ex_and_out_20_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_n1), 
        .B1(alu_ex_shift_out_20_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[21]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_U1 ( 
        .A1(alu_ex_and_out_21_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_n1), 
        .B1(alu_ex_shift_out_21_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[22]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_U1 ( 
        .A1(alu_ex_and_out_22_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_n1), 
        .B1(alu_ex_shift_out_22_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[23]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_U1 ( 
        .A1(alu_ex_and_out_23_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_n1), 
        .B1(alu_ex_shift_out_23_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[24]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_U1 ( 
        .A1(alu_ex_and_out_24_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_n1), 
        .B1(alu_ex_shift_out_24_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[25]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_U1 ( 
        .A1(alu_ex_and_out_25_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_n1), 
        .B1(alu_ex_shift_out_25_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[26]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_U1 ( 
        .A1(alu_ex_and_out_26_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_n1), 
        .B1(alu_ex_shift_out_26_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[27]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_U1 ( 
        .A1(alu_ex_and_out_27_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_n1), 
        .B1(alu_ex_shift_out_27_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[28]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_U1 ( 
        .A1(alu_ex_and_out_28_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_n1), 
        .B1(alu_ex_shift_out_28_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[29]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_U1 ( 
        .A1(alu_ex_and_out_29_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_n1), 
        .B1(alu_ex_shift_out_29_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[30]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_U1 ( 
        .A1(alu_ex_and_out_30_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_n1), 
        .B1(alu_ex_shift_out_30_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[31]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_U1 ( 
        .A1(alu_ex_and_out_31_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n1), 
        .B1(alu_ex_shift_out_31_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n4)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[0]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[0]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[1]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[1]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[2]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[2]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[3]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[3]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[4]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[4]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[5]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[5]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[6]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[6]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[7]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[7]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[8]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[8]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[9]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[9]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[10]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[10]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[11]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[11]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[12]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[12]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[13]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[13]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[14]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[14]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[15]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[15]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[16]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[16]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[17]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[17]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[18]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[18]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[19]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[19]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[20]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[20]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[21]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[21]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[22]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[22]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[23]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[23]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[24]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[24]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[25]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[25]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[26]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[26]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[27]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[27]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[28]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[28]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[29]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[29]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[30]), .A2(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[30]) );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_U4 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus2[31]), .A2(ALUCtrl_in[2]), 
        .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n2)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_U3 ( 
        .A(ALUCtrl_in[2]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n1)
         );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_U2 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_bus1_31_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n1), 
        .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n3)
         );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_U1 ( 
        .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n3), 
        .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS1_bus2[31]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_U4 ( .A(ALUCtrl_in[1]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1) );
  OAI21_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_U3 ( .B1(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_n2), .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_n1), .ZN(
        alu_ex_FINAL_MUX_bus1[0]) );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_U2 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[0]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_n1) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[0]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_n2) );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_U4 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[1]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1) );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_U2 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[1]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n2) );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n3), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n2), .ZN(
        alu_ex_FINAL_MUX_bus1[1]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_2__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[2]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[2]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[2]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_3__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[3]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[3]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[3]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_4__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[4]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[4]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[4]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_5__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[5]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[5]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[5]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_6__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[6]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[6]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[6]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_7__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[7]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[7]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[7]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_8__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[8]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[8]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[8]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_9__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[9]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[9]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[9]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_10__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[10]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[10]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[10])
         );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_11__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[11]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[11]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[11])
         );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_12__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[12]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[12]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[12])
         );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_13__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[13]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[13]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[13])
         );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_14__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[14]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[14]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[14])
         );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_15__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[15]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[15]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[15])
         );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_16__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[16]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[16]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[16])
         );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_17__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[17]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[17]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[17])
         );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_18__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[18]), .B(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[18]), .S(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n3), .Z(alu_ex_FINAL_MUX_bus1[18])
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus1[19]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[19]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[19]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus1[20]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[20]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[20]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus1[21]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[21]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[21]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus1[22]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[22]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[22]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus1[23]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[23]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[23]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus1[24]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[24]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[24]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus1[25]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[25]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[25]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus1[26]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[26]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[26]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus1[27]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[27]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[27]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus1[28]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[28]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[28]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus1[29]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[29]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[29]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus1[30]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[30]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[30]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_n4) );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_U2 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus2[31]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n2) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_U4 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n1) );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_U3 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n3), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n2), .ZN(
        alu_ex_FINAL_MUX_bus1[31]) );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS1_bus1[31]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_U4 ( .A(
        alu_ex_FINAL_MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[0]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_U1 ( 
        .A1(alu_ex_and_out_0_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_n1), 
        .B1(alu_ex_shift_out_0_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_0__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_1__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_1__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[1]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_1__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_1__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_1__MUX_U1 ( 
        .A1(alu_ex_and_out_1_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_1__MUX_n1), 
        .B1(alu_ex_shift_out_1_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_1__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[2]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_U1 ( 
        .A1(alu_ex_and_out_2_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_n1), 
        .B1(alu_ex_shift_out_2_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_2__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_3__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_3__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[3]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_3__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_3__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_3__MUX_U1 ( 
        .A1(alu_ex_and_out_3_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_3__MUX_n1), 
        .B1(alu_ex_shift_out_3_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_3__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_4__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_4__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[4]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_4__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_4__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_4__MUX_U1 ( 
        .A1(alu_ex_and_out_4_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_4__MUX_n1), 
        .B1(alu_ex_shift_out_4_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_4__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_5__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_5__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[5]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_5__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_5__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_5__MUX_U1 ( 
        .A1(alu_ex_and_out_5_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_5__MUX_n1), 
        .B1(alu_ex_shift_out_5_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_5__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_6__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_6__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[6]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_6__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_6__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_6__MUX_U1 ( 
        .A1(alu_ex_and_out_6_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_6__MUX_n1), 
        .B1(alu_ex_shift_out_6_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_6__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_7__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_7__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[7]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_7__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_7__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_7__MUX_U1 ( 
        .A1(alu_ex_and_out_7_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_7__MUX_n1), 
        .B1(alu_ex_shift_out_7_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_7__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_8__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_8__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[8]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_8__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_8__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_8__MUX_U1 ( 
        .A1(alu_ex_and_out_8_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_8__MUX_n1), 
        .B1(alu_ex_shift_out_8_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_8__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_9__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_9__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[9]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_9__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_9__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_9__MUX_U1 ( 
        .A1(alu_ex_and_out_9_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_9__MUX_n1), 
        .B1(alu_ex_shift_out_9_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_9__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_10__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_10__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[10]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_10__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_10__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_10__MUX_U1 ( 
        .A1(alu_ex_and_out_10_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_10__MUX_n1), 
        .B1(alu_ex_shift_out_10_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_10__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_11__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_11__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[11]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_11__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_11__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_11__MUX_U1 ( 
        .A1(alu_ex_and_out_11_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_11__MUX_n1), 
        .B1(alu_ex_shift_out_11_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_11__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_12__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_12__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[12]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_12__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_12__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_12__MUX_U1 ( 
        .A1(alu_ex_and_out_12_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_12__MUX_n1), 
        .B1(alu_ex_shift_out_12_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_12__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_13__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_13__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[13]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_13__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_13__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_13__MUX_U1 ( 
        .A1(alu_ex_and_out_13_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_13__MUX_n1), 
        .B1(alu_ex_shift_out_13_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_13__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_14__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_14__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[14]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_14__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_14__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_14__MUX_U1 ( 
        .A1(alu_ex_and_out_14_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_14__MUX_n1), 
        .B1(alu_ex_shift_out_14_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_14__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_15__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_15__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[15]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_15__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_15__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_15__MUX_U1 ( 
        .A1(alu_ex_and_out_15_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_15__MUX_n1), 
        .B1(alu_ex_shift_out_15_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_15__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_16__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_16__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[16]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_16__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_16__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_16__MUX_U1 ( 
        .A1(alu_ex_and_out_16_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_16__MUX_n1), 
        .B1(alu_ex_shift_out_16_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_16__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_17__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_17__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[17]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_17__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_17__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_17__MUX_U1 ( 
        .A1(alu_ex_and_out_17_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_17__MUX_n1), 
        .B1(alu_ex_shift_out_17_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_17__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_18__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_18__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[18]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_18__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_18__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_18__MUX_U1 ( 
        .A1(alu_ex_and_out_18_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_18__MUX_n1), 
        .B1(alu_ex_shift_out_18_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_18__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[19]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_U1 ( 
        .A1(alu_ex_and_out_19_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_n1), 
        .B1(alu_ex_shift_out_19_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_19__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[20]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_U1 ( 
        .A1(alu_ex_and_out_20_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_n1), 
        .B1(alu_ex_shift_out_20_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_20__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[21]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_U1 ( 
        .A1(alu_ex_and_out_21_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_n1), 
        .B1(alu_ex_shift_out_21_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_21__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[22]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_U1 ( 
        .A1(alu_ex_and_out_22_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_n1), 
        .B1(alu_ex_shift_out_22_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_22__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[23]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_U1 ( 
        .A1(alu_ex_and_out_23_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_n1), 
        .B1(alu_ex_shift_out_23_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_23__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[24]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_U1 ( 
        .A1(alu_ex_and_out_24_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_n1), 
        .B1(alu_ex_shift_out_24_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_24__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[25]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_U1 ( 
        .A1(alu_ex_and_out_25_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_n1), 
        .B1(alu_ex_shift_out_25_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_25__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[26]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_U1 ( 
        .A1(alu_ex_and_out_26_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_n1), 
        .B1(alu_ex_shift_out_26_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_26__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[27]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_U1 ( 
        .A1(alu_ex_and_out_27_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_n1), 
        .B1(alu_ex_shift_out_27_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_27__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[28]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_U1 ( 
        .A1(alu_ex_and_out_28_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_n1), 
        .B1(alu_ex_shift_out_28_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_28__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[29]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_U1 ( 
        .A1(alu_ex_and_out_29_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_n1), 
        .B1(alu_ex_shift_out_29_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_29__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[30]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_U1 ( 
        .A1(alu_ex_and_out_30_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_n1), 
        .B1(alu_ex_shift_out_30_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_30__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[31]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_U1 ( 
        .A1(alu_ex_and_out_31_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n1), 
        .B1(alu_ex_shift_out_31_), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_U4 ( .A(
        alu_ex_FINAL_MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n1) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n2) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_0__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_0__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_0__MUX_U1 ( 
        .A1(alu_ex_shift_out_0_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_0__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[0]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_1__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_1__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_1__MUX_U1 ( 
        .A1(alu_ex_shift_out_1_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_1__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[1]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_2__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_2__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_2__MUX_U1 ( 
        .A1(alu_ex_shift_out_2_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_2__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[2]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_3__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_3__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_3__MUX_U1 ( 
        .A1(alu_ex_shift_out_3_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_3__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[3]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_4__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_4__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_4__MUX_U1 ( 
        .A1(alu_ex_shift_out_4_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_4__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[4]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_5__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_5__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_5__MUX_U1 ( 
        .A1(alu_ex_shift_out_5_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_5__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[5]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_6__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_6__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_6__MUX_U1 ( 
        .A1(alu_ex_shift_out_6_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_6__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[6]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_7__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_7__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_7__MUX_U1 ( 
        .A1(alu_ex_shift_out_7_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_7__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[7]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_8__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_8__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_8__MUX_U1 ( 
        .A1(alu_ex_shift_out_8_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_8__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[8]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_9__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_9__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_9__MUX_U1 ( 
        .A1(alu_ex_shift_out_9_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_9__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[9]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_10__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_10__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_10__MUX_U1 ( 
        .A1(alu_ex_shift_out_10_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_10__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[10]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_11__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_11__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_11__MUX_U1 ( 
        .A1(alu_ex_shift_out_11_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_11__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[11]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_12__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_12__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_12__MUX_U1 ( 
        .A1(alu_ex_shift_out_12_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_12__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[12]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_13__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_13__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_13__MUX_U1 ( 
        .A1(alu_ex_shift_out_13_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_13__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[13]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_14__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_14__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_14__MUX_U1 ( 
        .A1(alu_ex_shift_out_14_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_14__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[14]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_15__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_15__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_15__MUX_U1 ( 
        .A1(alu_ex_shift_out_15_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_15__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[15]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_16__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_16__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_16__MUX_U1 ( 
        .A1(alu_ex_shift_out_16_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_16__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[16]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_17__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_17__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_17__MUX_U1 ( 
        .A1(alu_ex_shift_out_17_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_17__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[17]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_18__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_18__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_18__MUX_U1 ( 
        .A1(alu_ex_shift_out_18_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_18__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[18]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_19__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_19__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_19__MUX_U1 ( 
        .A1(alu_ex_shift_out_19_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_19__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[19]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_20__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_20__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_20__MUX_U1 ( 
        .A1(alu_ex_shift_out_20_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_20__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[20]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_21__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_21__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_21__MUX_U1 ( 
        .A1(alu_ex_shift_out_21_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_21__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[21]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_22__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_22__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_22__MUX_U1 ( 
        .A1(alu_ex_shift_out_22_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_22__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[22]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_23__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_23__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_23__MUX_U1 ( 
        .A1(alu_ex_shift_out_23_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_23__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[23]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_24__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_24__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_24__MUX_U1 ( 
        .A1(alu_ex_shift_out_24_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_24__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[24]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_25__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_25__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_25__MUX_U1 ( 
        .A1(alu_ex_shift_out_25_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_25__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[25]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_26__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_26__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_26__MUX_U1 ( 
        .A1(alu_ex_shift_out_26_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_26__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[26]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_27__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_27__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_27__MUX_U1 ( 
        .A1(alu_ex_shift_out_27_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_27__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[27]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_28__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_28__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_28__MUX_U1 ( 
        .A1(alu_ex_shift_out_28_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_28__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[28]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_29__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_29__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_29__MUX_U1 ( 
        .A1(alu_ex_shift_out_29_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_29__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[29]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_30__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_30__MUX_n2)
         );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_30__MUX_U1 ( 
        .A1(alu_ex_shift_out_30_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_30__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[30]) );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_U1 ( 
        .A1(alu_ex_seq_out_31_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n1)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_U4 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n3)
         );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_U3 ( 
        .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n1), 
        .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n2), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[31]) );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_U2 ( 
        .A1(alu_ex_shift_out_31_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n3), 
        .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n2)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_U4 ( .A(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[0]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[0]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[0]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_0__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[1]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[1]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[1]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_1__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_2__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_2__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[2]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_2__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_2__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[2]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_2__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[2]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_2__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_3__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_3__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[3]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_3__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_3__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[3]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_3__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[3]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_3__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_4__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_4__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[4]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_4__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_4__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[4]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_4__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[4]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_4__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_5__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_5__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[5]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_5__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_5__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[5]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_5__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[5]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_5__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_6__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_6__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[6]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_6__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_6__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[6]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_6__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[6]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_6__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_7__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_7__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[7]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_7__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_7__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[7]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_7__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[7]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_7__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_8__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_8__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[8]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_8__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_8__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[8]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_8__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[8]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_8__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_9__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_9__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[9]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_9__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_9__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[9]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_9__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[9]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_9__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_10__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_10__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[10]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_10__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_10__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_10__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[10]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_10__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[10]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_10__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_11__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_11__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[11]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_11__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_11__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_11__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[11]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_11__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[11]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_11__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_12__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_12__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[12]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_12__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_12__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_12__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[12]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_12__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[12]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_12__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_13__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_13__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[13]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_13__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_13__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_13__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[13]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_13__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[13]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_13__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_14__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_14__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[14]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_14__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_14__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_14__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[14]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_14__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[14]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_14__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_15__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_15__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[15]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_15__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_15__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_15__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[15]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_15__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[15]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_15__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_16__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_16__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[16]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_16__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_16__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_16__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[16]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_16__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[16]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_16__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_17__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_17__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[17]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_17__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_17__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_17__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[17]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_17__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[17]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_17__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_18__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_18__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[18]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_18__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_18__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_18__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[18]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_18__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[18]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_18__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[19]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[19]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[19]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_19__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[20]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[20]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[20]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_20__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[21]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[21]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[21]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_21__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[22]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[22]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[22]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_22__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[23]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[23]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[23]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_23__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[24]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[24]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[24]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_24__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[25]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[25]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[25]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_25__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[26]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[26]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[26]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_26__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[27]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[27]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[27]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_27__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[28]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[28]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[28]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_28__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[29]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[29]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[29]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_29__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus1[30]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[30]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[30]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_30__MUX_n4)
         );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_MUX2TO1_32BIT_31__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus1[31]), .B(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_bus2[31]), .S(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS1_MUX_OUT_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[31]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_U3 ( .A(
        alu_ex_FINAL_MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_0__MUX_U1 ( 
        .A1(alu_ex_and_out_0_), .A2(alu_ex_FINAL_MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[0]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_1__MUX_U1 ( 
        .A1(alu_ex_and_out_1_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[1]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_2__MUX_U1 ( 
        .A1(alu_ex_and_out_2_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[2]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_3__MUX_U1 ( 
        .A1(alu_ex_and_out_3_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[3]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_4__MUX_U1 ( 
        .A1(alu_ex_and_out_4_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[4]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_5__MUX_U1 ( 
        .A1(alu_ex_and_out_5_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[5]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_6__MUX_U1 ( 
        .A1(alu_ex_and_out_6_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[6]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_7__MUX_U1 ( 
        .A1(alu_ex_and_out_7_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[7]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_8__MUX_U1 ( 
        .A1(alu_ex_and_out_8_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[8]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_9__MUX_U1 ( 
        .A1(alu_ex_and_out_9_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[9]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_10__MUX_U1 ( 
        .A1(alu_ex_and_out_10_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[10]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_11__MUX_U1 ( 
        .A1(alu_ex_and_out_11_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[11]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_12__MUX_U1 ( 
        .A1(alu_ex_and_out_12_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[12]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_13__MUX_U1 ( 
        .A1(alu_ex_and_out_13_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[13]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_14__MUX_U1 ( 
        .A1(alu_ex_and_out_14_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[14]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_15__MUX_U1 ( 
        .A1(alu_ex_and_out_15_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[15]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_16__MUX_U1 ( 
        .A1(alu_ex_and_out_16_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[16]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_17__MUX_U1 ( 
        .A1(alu_ex_and_out_17_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[17]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_18__MUX_U1 ( 
        .A1(alu_ex_and_out_18_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[18]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_19__MUX_U1 ( 
        .A1(alu_ex_and_out_19_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[19]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_20__MUX_U1 ( 
        .A1(alu_ex_and_out_20_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[20]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_21__MUX_U1 ( 
        .A1(alu_ex_and_out_21_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[21]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_22__MUX_U1 ( 
        .A1(alu_ex_and_out_22_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[22]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_23__MUX_U1 ( 
        .A1(alu_ex_and_out_23_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[23]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_24__MUX_U1 ( 
        .A1(alu_ex_and_out_24_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[24]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_25__MUX_U1 ( 
        .A1(alu_ex_and_out_25_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[25]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_26__MUX_U1 ( 
        .A1(alu_ex_and_out_26_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[26]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_27__MUX_U1 ( 
        .A1(alu_ex_and_out_27_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[27]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_28__MUX_U1 ( 
        .A1(alu_ex_and_out_28_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[28]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_29__MUX_U1 ( 
        .A1(alu_ex_and_out_29_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[29]) );
  AND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_30__MUX_U1 ( 
        .A1(alu_ex_and_out_30_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[30]) );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_U3 ( 
        .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n2), 
        .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n3), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[31]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_U4 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n1)
         );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_U2 ( 
        .A1(alu_ex_and_out_31_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n3)
         );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_U1 ( 
        .A1(alu_ex_sne_out_31_), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n1), 
        .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS1_MUX2TO1_32BIT_31__MUX_n2)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_U4 ( .A(
        alu_ex_FINAL_MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[0]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_U1 ( 
        .A1(alu_ex_or_out[0]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_n1), 
        .B1(alu_ex_xor_out[0]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_0__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[1]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_U1 ( 
        .A1(alu_ex_or_out[1]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_n1), 
        .B1(alu_ex_xor_out[1]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_1__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[2]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_U1 ( 
        .A1(alu_ex_or_out[2]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_n1), 
        .B1(alu_ex_xor_out[2]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_2__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[3]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_U1 ( 
        .A1(alu_ex_or_out[3]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_n1), 
        .B1(alu_ex_xor_out[3]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_3__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[4]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_U1 ( 
        .A1(alu_ex_or_out[4]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_n1), 
        .B1(alu_ex_xor_out[4]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_4__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[5]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_U1 ( 
        .A1(alu_ex_or_out[5]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_n1), 
        .B1(alu_ex_xor_out[5]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_5__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[6]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_U1 ( 
        .A1(alu_ex_or_out[6]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_n1), 
        .B1(alu_ex_xor_out[6]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_6__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[7]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_U1 ( 
        .A1(alu_ex_or_out[7]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_n1), 
        .B1(alu_ex_xor_out[7]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_7__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[8]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_U1 ( 
        .A1(alu_ex_or_out[8]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_n1), 
        .B1(alu_ex_xor_out[8]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_8__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[9]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_U1 ( 
        .A1(alu_ex_or_out[9]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_n1), 
        .B1(alu_ex_xor_out[9]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_9__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[10]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_U1 ( 
        .A1(alu_ex_or_out[10]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_n1), 
        .B1(alu_ex_xor_out[10]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_10__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[11]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_U1 ( 
        .A1(alu_ex_or_out[11]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_n1), 
        .B1(alu_ex_xor_out[11]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_11__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[12]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_U1 ( 
        .A1(alu_ex_or_out[12]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_n1), 
        .B1(alu_ex_xor_out[12]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_12__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[13]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_U1 ( 
        .A1(alu_ex_or_out[13]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_n1), 
        .B1(alu_ex_xor_out[13]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_13__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[14]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_U1 ( 
        .A1(alu_ex_or_out[14]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_n1), 
        .B1(alu_ex_xor_out[14]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_14__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[15]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_U1 ( 
        .A1(alu_ex_or_out[15]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_n1), 
        .B1(alu_ex_xor_out[15]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_15__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[16]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_U1 ( 
        .A1(alu_ex_or_out[16]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_n1), 
        .B1(alu_ex_xor_out[16]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_16__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[17]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_U1 ( 
        .A1(alu_ex_or_out[17]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_n1), 
        .B1(alu_ex_xor_out[17]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_17__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[18]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_U1 ( 
        .A1(alu_ex_or_out[18]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_n1), 
        .B1(alu_ex_xor_out[18]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_18__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[19]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_U1 ( 
        .A1(alu_ex_or_out[19]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_n1), 
        .B1(alu_ex_xor_out[19]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_19__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[20]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_U1 ( 
        .A1(alu_ex_or_out[20]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_n1), 
        .B1(alu_ex_xor_out[20]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_20__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[21]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_U1 ( 
        .A1(alu_ex_or_out[21]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_n1), 
        .B1(alu_ex_xor_out[21]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_21__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[22]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_U1 ( 
        .A1(alu_ex_or_out[22]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_n1), 
        .B1(alu_ex_xor_out[22]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_22__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[23]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_U1 ( 
        .A1(alu_ex_or_out[23]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_n1), 
        .B1(alu_ex_xor_out[23]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_23__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[24]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_U1 ( 
        .A1(alu_ex_or_out[24]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_n1), 
        .B1(alu_ex_xor_out[24]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_24__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[25]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_U1 ( 
        .A1(alu_ex_or_out[25]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_n1), 
        .B1(alu_ex_xor_out[25]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_25__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[26]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_U1 ( 
        .A1(alu_ex_or_out[26]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_n1), 
        .B1(alu_ex_xor_out[26]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_26__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[27]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_U1 ( 
        .A1(alu_ex_or_out[27]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_n1), 
        .B1(alu_ex_xor_out[27]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_27__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[28]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_U1 ( 
        .A1(alu_ex_or_out[28]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_n1), 
        .B1(alu_ex_xor_out[28]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_28__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[29]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_U1 ( 
        .A1(alu_ex_or_out[29]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_n1), 
        .B1(alu_ex_xor_out[29]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_29__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[30]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_U1 ( 
        .A1(alu_ex_or_out[30]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_n1), 
        .B1(alu_ex_xor_out[30]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_30__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_U3 ( 
        .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[31]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_U1 ( 
        .A1(alu_ex_or_out[31]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n1), 
        .B1(alu_ex_xor_out[31]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_BUS2_MUX2TO1_32BIT_31__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_U4 ( .A(ALUCtrl_in[2]), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[0]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[0]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[0]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[1]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[1]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[1]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[2]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[2]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[2]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[3]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[3]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[3]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[4]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[4]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[4]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[5]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[5]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[5]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[6]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[6]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[6]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[7]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[7]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[7]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[8]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[8]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[8]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_n4), 
        .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[9]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[9]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[9]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[10]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[10]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[10]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[11]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[11]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[11]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[12]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[12]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[12]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[13]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[13]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[13]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[14]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[14]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[14]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[15]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[15]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[15]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[16]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[16]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[16]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[17]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[17]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[17]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[18]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[18]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[18]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[19]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[19]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[19]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[20]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[20]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[20]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[21]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[21]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[21]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[22]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[22]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[22]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[23]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[23]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[23]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[24]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[24]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[24]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[25]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[25]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[25]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[26]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[26]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[26]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[27]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[27]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[27]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[28]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[28]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[28]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[29]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[29]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[29]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_n4)
         );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_U3 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_n4), .ZN(alu_ex_FINAL_MUX_MUX_BUS2_bus2[30]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_U2 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_n1)
         );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_U1 ( 
        .A1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[30]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_n1), 
        .B1(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[30]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_n4)
         );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_U1 ( 
        .A(alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus1[31]), .B(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_bus2[31]), .S(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_BUS2_MUX_OUT_n3), .Z(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[31]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_U6 ( .A(ALUCtrl_in[1]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n6) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_U5 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n6), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n5) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_U4 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n6), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n6), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n6), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n6), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n1) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[0]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n5), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[0]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[0]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n5), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_0__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[1]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n5), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[1]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[1]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n5), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_1__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[2]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n5), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[2]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[2]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n5), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_2__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[3]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n5), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[3]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[3]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n5), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_3__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[4]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[4]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[4]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_4__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[5]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[5]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[5]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_5__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[6]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_U2 ( .A(
        ALUCtrl_in[1]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[6]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[6]), .B2(ALUCtrl_in[1]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_6__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[7]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[7]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[7]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_7__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[8]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[8]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[8]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_8__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[9]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_U2 ( .A(
        ALUCtrl_in[1]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[9]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[9]), .B2(ALUCtrl_in[1]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_9__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[10]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[10]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[10]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_10__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[11]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[11]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[11]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_11__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[12]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_U2 ( .A(
        ALUCtrl_in[1]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[12]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[12]), .B2(ALUCtrl_in[1]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_12__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[13]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[13]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[13]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_13__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[14]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[14]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[14]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_14__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[15]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_U2 ( .A(
        ALUCtrl_in[1]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[15]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[15]), .B2(ALUCtrl_in[1]), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_15__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[16]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[16]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[16]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_16__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[17]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[17]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[17]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_17__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[18]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n5), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[18]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[18]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n5), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_18__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[19]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[19]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[19]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_19__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[20]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[20]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[20]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_20__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[21]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[21]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[21]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_21__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[22]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[22]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[22]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_22__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[23]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[23]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[23]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_23__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[24]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[24]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[24]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_24__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[25]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[25]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[25]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_25__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[26]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[26]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[26]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_26__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[27]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[27]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[27]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_27__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[28]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[28]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[28]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_28__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[29]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[29]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[29]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_29__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_n4), .ZN(
        alu_ex_FINAL_MUX_bus2[30]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[30]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_n1), .B1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[30]), .B2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_30__MUX_n4) );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_U4 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n3), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n2), .ZN(
        alu_ex_FINAL_MUX_bus2[31]) );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_U3 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus2[31]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n2) );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_U2 ( .A1(
        alu_ex_FINAL_MUX_MUX_BUS2_bus1[31]), .A2(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_BUS2_MUX_OUT_MUX2TO1_32BIT_31__MUX_n1) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_U4 ( .A(ALUCtrl_in[0]), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_U3 ( .A(alu_ex_FINAL_MUX_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_U2 ( .A(alu_ex_FINAL_MUX_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_n2) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_U1 ( .A(alu_ex_FINAL_MUX_MUX_OUT_n4), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_n1) );
  OAI21_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_0__MUX_U3 ( .B1(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_0__MUX_n2), .B2(
        alu_ex_FINAL_MUX_MUX_OUT_n3), .A(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_0__MUX_n1), .ZN(
        not_mul_result[0]) );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_0__MUX_U2 ( .A1(
        alu_ex_FINAL_MUX_MUX_OUT_n3), .A2(alu_ex_FINAL_MUX_bus2[0]), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_0__MUX_n1) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_0__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[0]), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_0__MUX_n2) );
  NAND2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_1__MUX_U4 ( .A1(
        alu_ex_FINAL_MUX_MUX_OUT_n1), .A2(alu_ex_FINAL_MUX_bus2[1]), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_1__MUX_n3) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1) );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_1__MUX_U2 ( .A1(
        alu_ex_FINAL_MUX_bus1[1]), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_1__MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_1__MUX_n2) );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_1__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_1__MUX_n2), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_1__MUX_n3), .ZN(
        not_mul_result[1]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_2__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[2]), .B(alu_ex_FINAL_MUX_bus2[2]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[2]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_3__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[3]), .B(alu_ex_FINAL_MUX_bus2[3]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[3]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_4__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[4]), .B(alu_ex_FINAL_MUX_bus2[4]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[4]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_5__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[5]), .B(alu_ex_FINAL_MUX_bus2[5]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[5]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_6__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[6]), .B(alu_ex_FINAL_MUX_bus2[6]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[6]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_7__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[7]), .B(alu_ex_FINAL_MUX_bus2[7]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[7]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_8__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[8]), .B(alu_ex_FINAL_MUX_bus2[8]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[8]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_9__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[9]), .B(alu_ex_FINAL_MUX_bus2[9]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[9]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_10__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[10]), .B(alu_ex_FINAL_MUX_bus2[10]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[10]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_11__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[11]), .B(alu_ex_FINAL_MUX_bus2[11]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[11]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_12__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[12]), .B(alu_ex_FINAL_MUX_bus2[12]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[12]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_13__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[13]), .B(alu_ex_FINAL_MUX_bus2[13]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[13]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_14__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[14]), .B(alu_ex_FINAL_MUX_bus2[14]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[14]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_15__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[15]), .B(alu_ex_FINAL_MUX_bus2[15]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[15]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_16__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[16]), .B(alu_ex_FINAL_MUX_bus2[16]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[16]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_17__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[17]), .B(alu_ex_FINAL_MUX_bus2[17]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[17]) );
  MUX2_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_18__MUX_U1 ( .A(
        alu_ex_FINAL_MUX_bus1[18]), .B(alu_ex_FINAL_MUX_bus2[18]), .S(
        ALUCtrl_in[0]), .Z(not_mul_result[18]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_19__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_19__MUX_n4), .ZN(
        not_mul_result[19]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_19__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_19__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_19__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_bus1[19]), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_19__MUX_n1), .B1(
        alu_ex_FINAL_MUX_bus2[19]), .B2(alu_ex_FINAL_MUX_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_19__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_20__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_20__MUX_n4), .ZN(
        not_mul_result[20]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_20__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_20__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_20__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_bus1[20]), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_20__MUX_n1), .B1(
        alu_ex_FINAL_MUX_bus2[20]), .B2(alu_ex_FINAL_MUX_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_20__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_21__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_21__MUX_n4), .ZN(
        not_mul_result[21]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_21__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_21__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_21__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_bus1[21]), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_21__MUX_n1), .B1(
        alu_ex_FINAL_MUX_bus2[21]), .B2(alu_ex_FINAL_MUX_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_21__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_22__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_22__MUX_n4), .ZN(
        not_mul_result[22]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_22__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_22__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_22__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_bus1[22]), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_22__MUX_n1), .B1(
        alu_ex_FINAL_MUX_bus2[22]), .B2(alu_ex_FINAL_MUX_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_22__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_23__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_23__MUX_n4), .ZN(
        not_mul_result[23]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_23__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_23__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_23__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_bus1[23]), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_23__MUX_n1), .B1(
        alu_ex_FINAL_MUX_bus2[23]), .B2(alu_ex_FINAL_MUX_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_23__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_24__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_24__MUX_n4), .ZN(
        not_mul_result[24]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_24__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_24__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_24__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_bus1[24]), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_24__MUX_n1), .B1(
        alu_ex_FINAL_MUX_bus2[24]), .B2(alu_ex_FINAL_MUX_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_24__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_25__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_25__MUX_n4), .ZN(
        not_mul_result[25]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_25__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_25__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_25__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_bus1[25]), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_25__MUX_n1), .B1(
        alu_ex_FINAL_MUX_bus2[25]), .B2(alu_ex_FINAL_MUX_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_25__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_26__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_26__MUX_n4), .ZN(
        not_mul_result[26]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_26__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_26__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_26__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_bus1[26]), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_26__MUX_n1), .B1(
        alu_ex_FINAL_MUX_bus2[26]), .B2(alu_ex_FINAL_MUX_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_26__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_27__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_27__MUX_n4), .ZN(
        not_mul_result[27]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_27__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_27__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_27__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_bus1[27]), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_27__MUX_n1), .B1(
        alu_ex_FINAL_MUX_bus2[27]), .B2(alu_ex_FINAL_MUX_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_27__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_28__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_28__MUX_n4), .ZN(
        not_mul_result[28]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_28__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_28__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_28__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_bus1[28]), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_28__MUX_n1), .B1(
        alu_ex_FINAL_MUX_bus2[28]), .B2(alu_ex_FINAL_MUX_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_28__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_29__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_29__MUX_n4), .ZN(
        not_mul_result[29]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_29__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_29__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_29__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_bus1[29]), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_29__MUX_n1), .B1(
        alu_ex_FINAL_MUX_bus2[29]), .B2(alu_ex_FINAL_MUX_MUX_OUT_n2), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_29__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_30__MUX_U3 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_30__MUX_n4), .ZN(
        not_mul_result[30]) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_30__MUX_U2 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_30__MUX_n1) );
  AOI22_X2 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_30__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_bus1[30]), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_30__MUX_n1), .B1(
        alu_ex_FINAL_MUX_bus2[30]), .B2(alu_ex_FINAL_MUX_MUX_OUT_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_30__MUX_n4) );
  INV_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_31__MUX_U4 ( .A(
        alu_ex_FINAL_MUX_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_31__MUX_n1) );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_31__MUX_U3 ( .A1(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_31__MUX_n3), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_31__MUX_n2), .ZN(
        not_mul_result[31]) );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_31__MUX_U2 ( .A1(
        alu_ex_FINAL_MUX_bus1[31]), .A2(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_31__MUX_n1), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_31__MUX_n3) );
  NAND2_X4 alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_31__MUX_U1 ( .A1(
        alu_ex_FINAL_MUX_bus2[31]), .A2(alu_ex_FINAL_MUX_MUX_OUT_n3), .ZN(
        alu_ex_FINAL_MUX_MUX_OUT_MUX2TO1_32BIT_31__MUX_n2) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_U3 ( .A(movfp2i_in), .ZN(CHOOSE_FP_OR_NOTMUL_n3)
         );
  INV_X4 CHOOSE_FP_OR_NOTMUL_U2 ( .A(CHOOSE_FP_OR_NOTMUL_n3), .ZN(
        CHOOSE_FP_OR_NOTMUL_n2) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_U1 ( .A(CHOOSE_FP_OR_NOTMUL_n3), .ZN(
        CHOOSE_FP_OR_NOTMUL_n1) );
  AOI21_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_0__MUX_U4 ( .B1(not_mul_result[0]), .B2(CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_0__MUX_n2), .A(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_0__MUX_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_0__MUX_n3) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_0__MUX_U3 ( .A(
        CHOOSE_FP_OR_NOTMUL_n2), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_0__MUX_n2) );
  INV_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_0__MUX_U2 ( .A(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_0__MUX_n3), .ZN(aluResult_out[0]) );
  AND2_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_0__MUX_U1 ( .A1(
        CHOOSE_FP_OR_NOTMUL_n2), .A2(f1_in[0]), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_0__MUX_n1) );
  MUX2_X1 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_1__MUX_U1 ( .A(not_mul_result[1]), 
        .B(f1_in[1]), .S(movfp2i_in), .Z(aluResult_out[1]) );
  MUX2_X1 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_2__MUX_U1 ( .A(not_mul_result[2]), 
        .B(f1_in[2]), .S(movfp2i_in), .Z(aluResult_out[2]) );
  MUX2_X1 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_3__MUX_U1 ( .A(not_mul_result[3]), 
        .B(f1_in[3]), .S(movfp2i_in), .Z(aluResult_out[3]) );
  MUX2_X1 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_4__MUX_U1 ( .A(not_mul_result[4]), 
        .B(f1_in[4]), .S(movfp2i_in), .Z(aluResult_out[4]) );
  MUX2_X1 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_5__MUX_U1 ( .A(not_mul_result[5]), 
        .B(f1_in[5]), .S(movfp2i_in), .Z(aluResult_out[5]) );
  MUX2_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_6__MUX_U1 ( .A(not_mul_result[6]), 
        .B(f1_in[6]), .S(movfp2i_in), .Z(aluResult_out[6]) );
  MUX2_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_7__MUX_U1 ( .A(not_mul_result[7]), 
        .B(f1_in[7]), .S(movfp2i_in), .Z(aluResult_out[7]) );
  MUX2_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_8__MUX_U1 ( .A(not_mul_result[8]), 
        .B(f1_in[8]), .S(movfp2i_in), .Z(aluResult_out[8]) );
  MUX2_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_9__MUX_U1 ( .A(not_mul_result[9]), 
        .B(f1_in[9]), .S(movfp2i_in), .Z(aluResult_out[9]) );
  MUX2_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_10__MUX_U1 ( .A(not_mul_result[10]), .B(f1_in[10]), .S(movfp2i_in), .Z(aluResult_out[10]) );
  MUX2_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_11__MUX_U1 ( .A(not_mul_result[11]), .B(f1_in[11]), .S(movfp2i_in), .Z(aluResult_out[11]) );
  MUX2_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_12__MUX_U1 ( .A(not_mul_result[12]), .B(f1_in[12]), .S(movfp2i_in), .Z(aluResult_out[12]) );
  MUX2_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_13__MUX_U1 ( .A(not_mul_result[13]), .B(f1_in[13]), .S(movfp2i_in), .Z(aluResult_out[13]) );
  MUX2_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_14__MUX_U1 ( .A(not_mul_result[14]), .B(f1_in[14]), .S(movfp2i_in), .Z(aluResult_out[14]) );
  MUX2_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_15__MUX_U1 ( .A(not_mul_result[15]), .B(f1_in[15]), .S(movfp2i_in), .Z(aluResult_out[15]) );
  MUX2_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_16__MUX_U1 ( .A(not_mul_result[16]), .B(f1_in[16]), .S(movfp2i_in), .Z(aluResult_out[16]) );
  MUX2_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_17__MUX_U1 ( .A(not_mul_result[17]), .B(f1_in[17]), .S(movfp2i_in), .Z(aluResult_out[17]) );
  MUX2_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_18__MUX_U1 ( .A(not_mul_result[18]), .B(f1_in[18]), .S(movfp2i_in), .Z(aluResult_out[18]) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_19__MUX_U3 ( .A(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_19__MUX_n4), .ZN(aluResult_out[19])
         );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_19__MUX_U2 ( .A(
        CHOOSE_FP_OR_NOTMUL_n2), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_19__MUX_n1) );
  AOI22_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_19__MUX_U1 ( .A1(
        not_mul_result[19]), .A2(CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_19__MUX_n1), 
        .B1(f1_in[19]), .B2(CHOOSE_FP_OR_NOTMUL_n2), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_19__MUX_n4) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_20__MUX_U3 ( .A(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_20__MUX_n4), .ZN(aluResult_out[20])
         );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_20__MUX_U2 ( .A(
        CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_20__MUX_n1) );
  AOI22_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_20__MUX_U1 ( .A1(
        not_mul_result[20]), .A2(CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_20__MUX_n1), 
        .B1(f1_in[20]), .B2(CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_20__MUX_n4) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_21__MUX_U3 ( .A(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_21__MUX_n4), .ZN(aluResult_out[21])
         );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_21__MUX_U2 ( .A(
        CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_21__MUX_n1) );
  AOI22_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_21__MUX_U1 ( .A1(
        not_mul_result[21]), .A2(CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_21__MUX_n1), 
        .B1(f1_in[21]), .B2(CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_21__MUX_n4) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_22__MUX_U3 ( .A(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_22__MUX_n4), .ZN(aluResult_out[22])
         );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_22__MUX_U2 ( .A(
        CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_22__MUX_n1) );
  AOI22_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_22__MUX_U1 ( .A1(
        not_mul_result[22]), .A2(CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_22__MUX_n1), 
        .B1(f1_in[22]), .B2(CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_22__MUX_n4) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_23__MUX_U3 ( .A(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_23__MUX_n4), .ZN(aluResult_out[23])
         );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_23__MUX_U2 ( .A(
        CHOOSE_FP_OR_NOTMUL_n2), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_23__MUX_n1) );
  AOI22_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_23__MUX_U1 ( .A1(
        not_mul_result[23]), .A2(CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_23__MUX_n1), 
        .B1(f1_in[23]), .B2(CHOOSE_FP_OR_NOTMUL_n2), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_23__MUX_n4) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_24__MUX_U3 ( .A(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_24__MUX_n4), .ZN(aluResult_out[24])
         );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_24__MUX_U2 ( .A(
        CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_24__MUX_n1) );
  AOI22_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_24__MUX_U1 ( .A1(
        not_mul_result[24]), .A2(CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_24__MUX_n1), 
        .B1(f1_in[24]), .B2(CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_24__MUX_n4) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_25__MUX_U3 ( .A(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_25__MUX_n4), .ZN(aluResult_out[25])
         );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_25__MUX_U2 ( .A(
        CHOOSE_FP_OR_NOTMUL_n2), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_25__MUX_n1) );
  AOI22_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_25__MUX_U1 ( .A1(
        not_mul_result[25]), .A2(CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_25__MUX_n1), 
        .B1(f1_in[25]), .B2(CHOOSE_FP_OR_NOTMUL_n2), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_25__MUX_n4) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_26__MUX_U3 ( .A(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_26__MUX_n4), .ZN(aluResult_out[26])
         );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_26__MUX_U2 ( .A(
        CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_26__MUX_n1) );
  AOI22_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_26__MUX_U1 ( .A1(
        not_mul_result[26]), .A2(CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_26__MUX_n1), 
        .B1(f1_in[26]), .B2(CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_26__MUX_n4) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_27__MUX_U3 ( .A(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_27__MUX_n4), .ZN(aluResult_out[27])
         );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_27__MUX_U2 ( .A(
        CHOOSE_FP_OR_NOTMUL_n2), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_27__MUX_n1) );
  AOI22_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_27__MUX_U1 ( .A1(
        not_mul_result[27]), .A2(CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_27__MUX_n1), 
        .B1(f1_in[27]), .B2(CHOOSE_FP_OR_NOTMUL_n2), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_27__MUX_n4) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_28__MUX_U3 ( .A(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_28__MUX_n4), .ZN(aluResult_out[28])
         );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_28__MUX_U2 ( .A(
        CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_28__MUX_n1) );
  AOI22_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_28__MUX_U1 ( .A1(
        not_mul_result[28]), .A2(CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_28__MUX_n1), 
        .B1(f1_in[28]), .B2(CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_28__MUX_n4) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_29__MUX_U3 ( .A(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_29__MUX_n4), .ZN(aluResult_out[29])
         );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_29__MUX_U2 ( .A(
        CHOOSE_FP_OR_NOTMUL_n2), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_29__MUX_n1) );
  AOI22_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_29__MUX_U1 ( .A1(
        not_mul_result[29]), .A2(CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_29__MUX_n1), 
        .B1(f1_in[29]), .B2(CHOOSE_FP_OR_NOTMUL_n2), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_29__MUX_n4) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_30__MUX_U3 ( .A(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_30__MUX_n4), .ZN(aluResult_out[30])
         );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_30__MUX_U2 ( .A(
        CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_30__MUX_n1) );
  AOI22_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_30__MUX_U1 ( .A1(
        not_mul_result[30]), .A2(CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_30__MUX_n1), 
        .B1(f1_in[30]), .B2(CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_30__MUX_n4) );
  NAND2_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_31__MUX_U4 ( .A1(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_31__MUX_n3), .A2(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_31__MUX_n2), .ZN(aluResult_out[31])
         );
  NAND2_X2 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_31__MUX_U3 ( .A1(f1_in[31]), .A2(
        CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_31__MUX_n2) );
  INV_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_31__MUX_U2 ( .A(
        CHOOSE_FP_OR_NOTMUL_n1), .ZN(
        CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_31__MUX_n1) );
  NAND2_X4 CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_31__MUX_U1 ( .A1(
        not_mul_result[31]), .A2(CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_31__MUX_n1), 
        .ZN(CHOOSE_FP_OR_NOTMUL_MUX2TO1_32BIT_31__MUX_n3) );
  INV_X4 mul_ex_U169 ( .A(reset), .ZN(mul_ex_n40) );
  INV_X4 mul_ex_U168 ( .A(mul_ex_n35), .ZN(mul_ex_n39) );
  NOR3_X2 mul_ex_U137 ( .A1(mul_ex_CurrentState_1_), .A2(
        mul_ex_CurrentState_2_), .A3(mul_ex_CurrentState_0_), .ZN(mul_ex_N43)
         );
  NAND3_X2 mul_ex_U136 ( .A1(mul_ex_n5), .A2(mul_ex_n4), .A3(
        mul_ex_CurrentState_1_), .ZN(mul_ex_n35) );
  NAND3_X2 mul_ex_U135 ( .A1(mul_ex_n5), .A2(mul_ex_n4), .A3(mul_in), .ZN(
        mul_ex_n36) );
  AOI21_X2 mul_ex_U134 ( .B1(mul_ex_n35), .B2(mul_ex_n36), .A(mul_ex_n40), 
        .ZN(mul_ex_N14) );
  NAND3_X2 mul_ex_U133 ( .A1(mul_ex_CurrentState_2_), .A2(mul_ex_n5), .A3(
        mul_ex_CurrentState_1_), .ZN(mul_ex_n33) );
  INV_X4 mul_ex_U132 ( .A(mul_ex_n6), .ZN(mul_ex_n18) );
  INV_X4 mul_ex_U131 ( .A(mul_ex_N43), .ZN(mul_ex_n37) );
  INV_X4 mul_ex_U130 ( .A(mul_ex_n37), .ZN(mul_ex_n31) );
  INV_X4 mul_ex_U129 ( .A(mul_ex_n37), .ZN(mul_ex_n32) );
  AND2_X2 mul_ex_U128 ( .A1(mul_ex_n37), .A2(mul_ex_n35), .ZN(mul_ex_n10) );
  AND2_X2 mul_ex_U127 ( .A1(mul_ex_n37), .A2(mul_ex_n33), .ZN(mul_ex_n9) );
  INV_X4 mul_ex_U126 ( .A(mul_ex_n3), .ZN(mul_ex_n15) );
  NOR2_X2 mul_ex_U125 ( .A1(mul_ex_n15), .A2(mul_ex_n11), .ZN(mul_ex_n34) );
  NOR2_X2 mul_ex_U124 ( .A1(mul_ex_n34), .A2(mul_ex_n40), .ZN(mul_ex_N15) );
  NOR2_X2 mul_ex_U123 ( .A1(mul_ex_n33), .A2(mul_ex_n40), .ZN(mul_ex_N16) );
  INV_X4 mul_ex_U122 ( .A(mul_ex_n3), .ZN(mul_ex_n17) );
  OR2_X2 mul_ex_U121 ( .A1(mul_ex_n18), .A2(mul_ex_n31), .ZN(mul_ex_n8) );
  INV_X4 mul_ex_U120 ( .A(mul_ex_n33), .ZN(mul_ex_n14) );
  INV_X4 mul_ex_U119 ( .A(mul_ex_n33), .ZN(mul_ex_n12) );
  INV_X4 mul_ex_U118 ( .A(mul_ex_n33), .ZN(mul_ex_n13) );
  INV_X4 mul_ex_U117 ( .A(mul_ex_n10), .ZN(mul_ex_n24) );
  INV_X4 mul_ex_U116 ( .A(mul_ex_n9), .ZN(mul_ex_n27) );
  INV_X4 mul_ex_U115 ( .A(mul_ex_n10), .ZN(mul_ex_n22) );
  INV_X4 mul_ex_U114 ( .A(mul_ex_n10), .ZN(mul_ex_n23) );
  INV_X4 mul_ex_U113 ( .A(mul_ex_n9), .ZN(mul_ex_n25) );
  INV_X4 mul_ex_U112 ( .A(mul_ex_n9), .ZN(mul_ex_n26) );
  INV_X4 mul_ex_U111 ( .A(mul_ex_n6), .ZN(mul_ex_n21) );
  INV_X4 mul_ex_U110 ( .A(mul_ex_n3), .ZN(mul_ex_n16) );
  INV_X4 mul_ex_U109 ( .A(mul_ex_n6), .ZN(mul_ex_n20) );
  INV_X4 mul_ex_U108 ( .A(mul_ex_n6), .ZN(mul_ex_n19) );
  INV_X4 mul_ex_U107 ( .A(mul_ex_n35), .ZN(mul_ex_n11) );
  INV_X4 mul_ex_U74 ( .A(mul_ex_n7), .ZN(mul_ex_n30) );
  INV_X4 mul_ex_U41 ( .A(mul_ex_n7), .ZN(mul_ex_n28) );
  INV_X4 mul_ex_U6 ( .A(mul_ex_n7), .ZN(mul_ex_n29) );
  NOR2_X2 mul_ex_U5 ( .A1(mul_ex_N43), .A2(mul_ex_n17), .ZN(mul_ex_n7) );
  OR3_X4 mul_ex_U4 ( .A1(mul_ex_CurrentState_1_), .A2(mul_ex_CurrentState_2_), 
        .A3(mul_ex_n5), .ZN(mul_ex_n6) );
  OR3_X4 mul_ex_U3 ( .A1(mul_ex_CurrentState_0_), .A2(mul_ex_CurrentState_1_), 
        .A3(mul_ex_n4), .ZN(mul_ex_n3) );
  DLH_X2 mul_ex_H_reg_31_ ( .G(mul_ex_n31), .D(mul_ex_N56), .Q(mul_ex_H[31])
         );
  DLH_X2 mul_ex_H_reg_30_ ( .G(mul_ex_n31), .D(mul_ex_N57), .Q(mul_ex_H[30])
         );
  DLH_X2 mul_ex_H_reg_29_ ( .G(mul_ex_n31), .D(mul_ex_N58), .Q(mul_ex_H[29])
         );
  DLH_X2 mul_ex_H_reg_28_ ( .G(mul_ex_n31), .D(mul_ex_N59), .Q(mul_ex_H[28])
         );
  DLH_X2 mul_ex_H_reg_27_ ( .G(mul_ex_n31), .D(mul_ex_N60), .Q(mul_ex_H[27])
         );
  DLH_X2 mul_ex_H_reg_26_ ( .G(mul_ex_n31), .D(mul_ex_N61), .Q(mul_ex_H[26])
         );
  DLH_X2 mul_ex_H_reg_25_ ( .G(mul_ex_n31), .D(mul_ex_N62), .Q(mul_ex_H[25])
         );
  DLH_X2 mul_ex_H_reg_24_ ( .G(mul_ex_n31), .D(mul_ex_N63), .Q(mul_ex_H[24])
         );
  DLH_X2 mul_ex_H_reg_23_ ( .G(mul_ex_n31), .D(mul_ex_N64), .Q(mul_ex_H[23])
         );
  DLH_X2 mul_ex_H_reg_22_ ( .G(mul_ex_n31), .D(mul_ex_N65), .Q(mul_ex_H[22])
         );
  DLH_X2 mul_ex_H_reg_21_ ( .G(mul_ex_n31), .D(mul_ex_N66), .Q(mul_ex_H[21])
         );
  DLH_X2 mul_ex_H_reg_20_ ( .G(mul_ex_n31), .D(mul_ex_N67), .Q(mul_ex_H[20])
         );
  DLH_X2 mul_ex_H_reg_19_ ( .G(mul_ex_n31), .D(mul_ex_N68), .Q(mul_ex_H[19])
         );
  DLH_X2 mul_ex_H_reg_18_ ( .G(mul_ex_n31), .D(mul_ex_N69), .Q(mul_ex_H[18])
         );
  DLH_X2 mul_ex_H_reg_17_ ( .G(mul_ex_n32), .D(mul_ex_N70), .Q(mul_ex_H[17])
         );
  DLH_X2 mul_ex_H_reg_16_ ( .G(mul_ex_n31), .D(mul_ex_N71), .Q(mul_ex_H[16])
         );
  DLH_X2 mul_ex_H_reg_15_ ( .G(mul_ex_n31), .D(mul_ex_N72), .Q(mul_ex_H[15])
         );
  DLH_X2 mul_ex_H_reg_14_ ( .G(mul_ex_n32), .D(mul_ex_N73), .Q(mul_ex_H[14])
         );
  DLH_X2 mul_ex_H_reg_13_ ( .G(mul_ex_n32), .D(mul_ex_N74), .Q(mul_ex_H[13])
         );
  DLH_X2 mul_ex_H_reg_12_ ( .G(mul_ex_n32), .D(mul_ex_N75), .Q(mul_ex_H[12])
         );
  DLH_X2 mul_ex_H_reg_11_ ( .G(mul_ex_n32), .D(mul_ex_N76), .Q(mul_ex_H[11])
         );
  DLH_X2 mul_ex_H_reg_10_ ( .G(mul_ex_n32), .D(mul_ex_N77), .Q(mul_ex_H[10])
         );
  DLH_X2 mul_ex_H_reg_9_ ( .G(mul_ex_n32), .D(mul_ex_N78), .Q(mul_ex_H[9]) );
  DLH_X2 mul_ex_H_reg_8_ ( .G(mul_ex_n32), .D(mul_ex_N79), .Q(mul_ex_H[8]) );
  DLH_X2 mul_ex_H_reg_7_ ( .G(mul_ex_n32), .D(mul_ex_N80), .Q(mul_ex_H[7]) );
  DLH_X2 mul_ex_H_reg_6_ ( .G(mul_ex_n32), .D(mul_ex_N81), .Q(mul_ex_H[6]) );
  DLH_X2 mul_ex_H_reg_5_ ( .G(mul_ex_n32), .D(mul_ex_N82), .Q(mul_ex_H[5]) );
  DLH_X2 mul_ex_H_reg_4_ ( .G(mul_ex_n32), .D(mul_ex_N83), .Q(mul_ex_H[4]) );
  DLH_X2 mul_ex_H_reg_3_ ( .G(mul_ex_n32), .D(mul_ex_N84), .Q(mul_ex_H[3]) );
  DLH_X2 mul_ex_H_reg_2_ ( .G(mul_ex_n32), .D(mul_ex_N85), .Q(mul_ex_H[2]) );
  DLH_X2 mul_ex_H_reg_1_ ( .G(mul_ex_n32), .D(mul_ex_N86), .Q(mul_ex_H[1]) );
  DLH_X2 mul_ex_H_reg_0_ ( .G(mul_ex_n32), .D(mul_ex_N87), .Q(mul_ex_H[0]) );
  DLH_X2 mul_ex_result_reg_63_ ( .G(mul_ex_n18), .D(mul_ex_N314), .Q(
        mul_result_long[63]) );
  DLH_X2 mul_ex_result_reg_62_ ( .G(mul_ex_n18), .D(mul_ex_N315), .Q(
        mul_result_long[62]) );
  DLH_X2 mul_ex_result_reg_61_ ( .G(mul_ex_n18), .D(mul_ex_N316), .Q(
        mul_result_long[61]) );
  DLH_X2 mul_ex_result_reg_60_ ( .G(mul_ex_n18), .D(mul_ex_N317), .Q(
        mul_result_long[60]) );
  DLH_X2 mul_ex_result_reg_59_ ( .G(mul_ex_n18), .D(mul_ex_N318), .Q(
        mul_result_long[59]) );
  DLH_X2 mul_ex_result_reg_58_ ( .G(mul_ex_n18), .D(mul_ex_N319), .Q(
        mul_result_long[58]) );
  DLH_X2 mul_ex_result_reg_57_ ( .G(mul_ex_n18), .D(mul_ex_N320), .Q(
        mul_result_long[57]) );
  DLH_X2 mul_ex_result_reg_56_ ( .G(mul_ex_n18), .D(mul_ex_N321), .Q(
        mul_result_long[56]) );
  DLH_X2 mul_ex_result_reg_55_ ( .G(mul_ex_n18), .D(mul_ex_N322), .Q(
        mul_result_long[55]) );
  DLH_X2 mul_ex_result_reg_54_ ( .G(mul_ex_n18), .D(mul_ex_N323), .Q(
        mul_result_long[54]) );
  DLH_X2 mul_ex_result_reg_53_ ( .G(mul_ex_n18), .D(mul_ex_N324), .Q(
        mul_result_long[53]) );
  DLH_X2 mul_ex_result_reg_52_ ( .G(mul_ex_n18), .D(mul_ex_N325), .Q(
        mul_result_long[52]) );
  DLH_X2 mul_ex_result_reg_51_ ( .G(mul_ex_n18), .D(mul_ex_N326), .Q(
        mul_result_long[51]) );
  DLH_X2 mul_ex_result_reg_50_ ( .G(mul_ex_n18), .D(mul_ex_N327), .Q(
        mul_result_long[50]) );
  DLH_X2 mul_ex_result_reg_49_ ( .G(mul_ex_n19), .D(mul_ex_N328), .Q(
        mul_result_long[49]) );
  DLH_X2 mul_ex_result_reg_48_ ( .G(mul_ex_n19), .D(mul_ex_N329), .Q(
        mul_result_long[48]) );
  DLH_X2 mul_ex_result_reg_47_ ( .G(mul_ex_n19), .D(mul_ex_N330), .Q(
        mul_result_long[47]) );
  DLH_X2 mul_ex_result_reg_46_ ( .G(mul_ex_n19), .D(mul_ex_N331), .Q(
        mul_result_long[46]) );
  DLH_X2 mul_ex_result_reg_45_ ( .G(mul_ex_n19), .D(mul_ex_N332), .Q(
        mul_result_long[45]) );
  DLH_X2 mul_ex_result_reg_44_ ( .G(mul_ex_n19), .D(mul_ex_N333), .Q(
        mul_result_long[44]) );
  DLH_X2 mul_ex_result_reg_43_ ( .G(mul_ex_n19), .D(mul_ex_N334), .Q(
        mul_result_long[43]) );
  DLH_X2 mul_ex_result_reg_42_ ( .G(mul_ex_n19), .D(mul_ex_N335), .Q(
        mul_result_long[42]) );
  DLH_X2 mul_ex_result_reg_41_ ( .G(mul_ex_n19), .D(mul_ex_N336), .Q(
        mul_result_long[41]) );
  DLH_X2 mul_ex_result_reg_40_ ( .G(mul_ex_n19), .D(mul_ex_N337), .Q(
        mul_result_long[40]) );
  DLH_X2 mul_ex_result_reg_39_ ( .G(mul_ex_n19), .D(mul_ex_N338), .Q(
        mul_result_long[39]) );
  DLH_X2 mul_ex_result_reg_38_ ( .G(mul_ex_n19), .D(mul_ex_N339), .Q(
        mul_result_long[38]) );
  DLH_X2 mul_ex_result_reg_37_ ( .G(mul_ex_n19), .D(mul_ex_N340), .Q(
        mul_result_long[37]) );
  DLH_X2 mul_ex_result_reg_36_ ( .G(mul_ex_n19), .D(mul_ex_N341), .Q(
        mul_result_long[36]) );
  DLH_X2 mul_ex_result_reg_35_ ( .G(mul_ex_n19), .D(mul_ex_N342), .Q(
        mul_result_long[35]) );
  DLH_X2 mul_ex_result_reg_34_ ( .G(mul_ex_n19), .D(mul_ex_N343), .Q(
        mul_result_long[34]) );
  DLH_X2 mul_ex_result_reg_33_ ( .G(mul_ex_n19), .D(mul_ex_N344), .Q(
        mul_result_long[33]) );
  DLH_X2 mul_ex_result_reg_32_ ( .G(mul_ex_n20), .D(mul_ex_N345), .Q(
        mul_result_long[32]) );
  DLH_X2 mul_ex_result_reg_31_ ( .G(mul_ex_n20), .D(mul_ex_N346), .Q(
        mul_result_long[31]) );
  DLH_X2 mul_ex_result_reg_30_ ( .G(mul_ex_n20), .D(mul_ex_N347), .Q(
        mul_result_long[30]) );
  DLH_X2 mul_ex_result_reg_29_ ( .G(mul_ex_n20), .D(mul_ex_N348), .Q(
        mul_result_long[29]) );
  DLH_X2 mul_ex_result_reg_28_ ( .G(mul_ex_n20), .D(mul_ex_N349), .Q(
        mul_result_long[28]) );
  DLH_X2 mul_ex_result_reg_27_ ( .G(mul_ex_n20), .D(mul_ex_N350), .Q(
        mul_result_long[27]) );
  DLH_X2 mul_ex_result_reg_26_ ( .G(mul_ex_n20), .D(mul_ex_N351), .Q(
        mul_result_long[26]) );
  DLH_X2 mul_ex_result_reg_25_ ( .G(mul_ex_n20), .D(mul_ex_N352), .Q(
        mul_result_long[25]) );
  DLH_X2 mul_ex_result_reg_24_ ( .G(mul_ex_n20), .D(mul_ex_N353), .Q(
        mul_result_long[24]) );
  DLH_X2 mul_ex_result_reg_23_ ( .G(mul_ex_n20), .D(mul_ex_N354), .Q(
        mul_result_long[23]) );
  DLH_X2 mul_ex_result_reg_22_ ( .G(mul_ex_n20), .D(mul_ex_N355), .Q(
        mul_result_long[22]) );
  DLH_X2 mul_ex_result_reg_21_ ( .G(mul_ex_n20), .D(mul_ex_N356), .Q(
        mul_result_long[21]) );
  DLH_X2 mul_ex_result_reg_20_ ( .G(mul_ex_n20), .D(mul_ex_N357), .Q(
        mul_result_long[20]) );
  DLH_X2 mul_ex_result_reg_19_ ( .G(mul_ex_n20), .D(mul_ex_N358), .Q(
        mul_result_long[19]) );
  DLH_X2 mul_ex_result_reg_18_ ( .G(mul_ex_n20), .D(mul_ex_N359), .Q(
        mul_result_long[18]) );
  DLH_X2 mul_ex_result_reg_17_ ( .G(mul_ex_n20), .D(mul_ex_N360), .Q(
        mul_result_long[17]) );
  DLH_X2 mul_ex_result_reg_16_ ( .G(mul_ex_n20), .D(mul_ex_N361), .Q(
        mul_result_long[16]) );
  DLH_X2 mul_ex_result_reg_15_ ( .G(mul_ex_n21), .D(mul_ex_N362), .Q(
        mul_result_long[15]) );
  DLH_X2 mul_ex_result_reg_14_ ( .G(mul_ex_n21), .D(mul_ex_N363), .Q(
        mul_result_long[14]) );
  DLH_X2 mul_ex_result_reg_13_ ( .G(mul_ex_n21), .D(mul_ex_N364), .Q(
        mul_result_long[13]) );
  DLH_X2 mul_ex_result_reg_12_ ( .G(mul_ex_n21), .D(mul_ex_N365), .Q(
        mul_result_long[12]) );
  DLH_X2 mul_ex_result_reg_11_ ( .G(mul_ex_n21), .D(mul_ex_N366), .Q(
        mul_result_long[11]) );
  DLH_X2 mul_ex_result_reg_10_ ( .G(mul_ex_n21), .D(mul_ex_N367), .Q(
        mul_result_long[10]) );
  DLH_X2 mul_ex_result_reg_9_ ( .G(mul_ex_n21), .D(mul_ex_N368), .Q(
        mul_result_long[9]) );
  DLH_X2 mul_ex_result_reg_8_ ( .G(mul_ex_n21), .D(mul_ex_N369), .Q(
        mul_result_long[8]) );
  DLH_X2 mul_ex_result_reg_7_ ( .G(mul_ex_n21), .D(mul_ex_N370), .Q(
        mul_result_long[7]) );
  DLH_X2 mul_ex_result_reg_6_ ( .G(mul_ex_n21), .D(mul_ex_N371), .Q(
        mul_result_long[6]) );
  DLH_X2 mul_ex_result_reg_5_ ( .G(mul_ex_n21), .D(mul_ex_N372), .Q(
        mul_result_long[5]) );
  DLH_X2 mul_ex_result_reg_4_ ( .G(mul_ex_n21), .D(mul_ex_N373), .Q(
        mul_result_long[4]) );
  DLH_X2 mul_ex_result_reg_3_ ( .G(mul_ex_n21), .D(mul_ex_N374), .Q(
        mul_result_long[3]) );
  DLH_X2 mul_ex_result_reg_2_ ( .G(mul_ex_n21), .D(mul_ex_N375), .Q(
        mul_result_long[2]) );
  DLH_X2 mul_ex_result_reg_1_ ( .G(mul_ex_n21), .D(mul_ex_N376), .Q(
        mul_result_long[1]) );
  DLH_X2 mul_ex_result_reg_0_ ( .G(mul_ex_n18), .D(mul_ex_N377), .Q(
        mul_result_long[0]) );
  DLH_X2 mul_ex_Z_reg_31_ ( .G(mul_ex_n27), .D(mul_ex_N412), .Q(mul_ex_Z_31_)
         );
  DLH_X2 mul_ex_Z_reg_30_ ( .G(mul_ex_n27), .D(mul_ex_N413), .Q(mul_ex_Z_30_)
         );
  DLH_X2 mul_ex_Z_reg_29_ ( .G(mul_ex_n27), .D(mul_ex_N414), .Q(mul_ex_Z_29_)
         );
  DLH_X2 mul_ex_Z_reg_28_ ( .G(mul_ex_n27), .D(mul_ex_N415), .Q(mul_ex_Z_28_)
         );
  DLH_X2 mul_ex_Z_reg_27_ ( .G(mul_ex_n27), .D(mul_ex_N416), .Q(mul_ex_Z_27_)
         );
  DLH_X2 mul_ex_Z_reg_26_ ( .G(mul_ex_n27), .D(mul_ex_N417), .Q(mul_ex_Z_26_)
         );
  DLH_X2 mul_ex_Z_reg_25_ ( .G(mul_ex_n27), .D(mul_ex_N418), .Q(mul_ex_Z_25_)
         );
  DLH_X2 mul_ex_Z_reg_24_ ( .G(mul_ex_n27), .D(mul_ex_N419), .Q(mul_ex_Z_24_)
         );
  DLH_X2 mul_ex_Z_reg_23_ ( .G(mul_ex_n27), .D(mul_ex_N420), .Q(mul_ex_Z_23_)
         );
  DLH_X2 mul_ex_Z_reg_22_ ( .G(mul_ex_n27), .D(mul_ex_N421), .Q(mul_ex_Z_22_)
         );
  DLH_X2 mul_ex_Z_reg_21_ ( .G(mul_ex_n26), .D(mul_ex_N422), .Q(mul_ex_Z_21_)
         );
  DLH_X2 mul_ex_Z_reg_20_ ( .G(mul_ex_n26), .D(mul_ex_N423), .Q(mul_ex_Z_20_)
         );
  DLH_X2 mul_ex_Z_reg_19_ ( .G(mul_ex_n26), .D(mul_ex_N424), .Q(mul_ex_Z_19_)
         );
  DLH_X2 mul_ex_Z_reg_18_ ( .G(mul_ex_n26), .D(mul_ex_N425), .Q(mul_ex_Z_18_)
         );
  DLH_X2 mul_ex_Z_reg_17_ ( .G(mul_ex_n26), .D(mul_ex_N426), .Q(mul_ex_Z_17_)
         );
  DLH_X2 mul_ex_Z_reg_16_ ( .G(mul_ex_n26), .D(mul_ex_N427), .Q(mul_ex_Z_16_)
         );
  DLH_X2 mul_ex_Z_reg_15_ ( .G(mul_ex_n26), .D(mul_ex_N428), .Q(mul_ex_Z_15_)
         );
  DLH_X2 mul_ex_Z_reg_14_ ( .G(mul_ex_n26), .D(mul_ex_N429), .Q(mul_ex_Z_14_)
         );
  DLH_X2 mul_ex_Z_reg_13_ ( .G(mul_ex_n26), .D(mul_ex_N430), .Q(mul_ex_Z_13_)
         );
  DLH_X2 mul_ex_Z_reg_12_ ( .G(mul_ex_n26), .D(mul_ex_N431), .Q(mul_ex_Z_12_)
         );
  DLH_X2 mul_ex_Z_reg_11_ ( .G(mul_ex_n26), .D(mul_ex_N432), .Q(mul_ex_Z_11_)
         );
  DLH_X2 mul_ex_Z_reg_10_ ( .G(mul_ex_n25), .D(mul_ex_N433), .Q(mul_ex_Z_10_)
         );
  DLH_X2 mul_ex_Z_reg_9_ ( .G(mul_ex_n25), .D(mul_ex_N434), .Q(mul_ex_Z_9_) );
  DLH_X2 mul_ex_Z_reg_8_ ( .G(mul_ex_n25), .D(mul_ex_N435), .Q(mul_ex_Z_8_) );
  DLH_X2 mul_ex_Z_reg_7_ ( .G(mul_ex_n25), .D(mul_ex_N436), .Q(mul_ex_Z_7_) );
  DLH_X2 mul_ex_Z_reg_6_ ( .G(mul_ex_n25), .D(mul_ex_N437), .Q(mul_ex_Z_6_) );
  DLH_X2 mul_ex_Z_reg_5_ ( .G(mul_ex_n25), .D(mul_ex_N438), .Q(mul_ex_Z_5_) );
  DLH_X2 mul_ex_Z_reg_4_ ( .G(mul_ex_n25), .D(mul_ex_N439), .Q(mul_ex_Z_4_) );
  DLH_X2 mul_ex_Z_reg_3_ ( .G(mul_ex_n25), .D(mul_ex_N440), .Q(mul_ex_Z_3_) );
  DLH_X2 mul_ex_Z_reg_2_ ( .G(mul_ex_n25), .D(mul_ex_N441), .Q(mul_ex_Z_2_) );
  DLH_X2 mul_ex_Z_reg_1_ ( .G(mul_ex_n25), .D(mul_ex_N442), .Q(mul_ex_Z_1_) );
  DLH_X2 mul_ex_Z_reg_0_ ( .G(mul_ex_n25), .D(mul_ex_N443), .Q(mul_ex_Z_0_) );
  DLH_X2 mul_ex_L_reg_31_ ( .G(mul_ex_n30), .D(mul_ex_N379), .Q(mul_ex_L_31_)
         );
  DLH_X2 mul_ex_L_reg_30_ ( .G(mul_ex_n30), .D(mul_ex_N380), .Q(mul_ex_L_30_)
         );
  DLH_X2 mul_ex_L_reg_29_ ( .G(mul_ex_n30), .D(mul_ex_N381), .Q(mul_ex_L_29_)
         );
  DLH_X2 mul_ex_L_reg_28_ ( .G(mul_ex_n30), .D(mul_ex_N382), .Q(mul_ex_L_28_)
         );
  DLH_X2 mul_ex_L_reg_27_ ( .G(mul_ex_n30), .D(mul_ex_N383), .Q(mul_ex_L_27_)
         );
  DLH_X2 mul_ex_L_reg_26_ ( .G(mul_ex_n30), .D(mul_ex_N384), .Q(mul_ex_L_26_)
         );
  DLH_X2 mul_ex_L_reg_25_ ( .G(mul_ex_n30), .D(mul_ex_N385), .Q(mul_ex_L_25_)
         );
  DLH_X2 mul_ex_L_reg_24_ ( .G(mul_ex_n30), .D(mul_ex_N386), .Q(mul_ex_L_24_)
         );
  DLH_X2 mul_ex_L_reg_23_ ( .G(mul_ex_n30), .D(mul_ex_N387), .Q(mul_ex_L_23_)
         );
  DLH_X2 mul_ex_L_reg_22_ ( .G(mul_ex_n30), .D(mul_ex_N388), .Q(mul_ex_L_22_)
         );
  DLH_X2 mul_ex_L_reg_21_ ( .G(mul_ex_n29), .D(mul_ex_N389), .Q(mul_ex_L_21_)
         );
  DLH_X2 mul_ex_L_reg_20_ ( .G(mul_ex_n29), .D(mul_ex_N390), .Q(mul_ex_L_20_)
         );
  DLH_X2 mul_ex_L_reg_19_ ( .G(mul_ex_n29), .D(mul_ex_N391), .Q(mul_ex_L_19_)
         );
  DLH_X2 mul_ex_L_reg_18_ ( .G(mul_ex_n29), .D(mul_ex_N392), .Q(mul_ex_L_18_)
         );
  DLH_X2 mul_ex_L_reg_17_ ( .G(mul_ex_n29), .D(mul_ex_N393), .Q(mul_ex_L_17_)
         );
  DLH_X2 mul_ex_L_reg_16_ ( .G(mul_ex_n29), .D(mul_ex_N394), .Q(mul_ex_L_16_)
         );
  DLH_X2 mul_ex_L_reg_15_ ( .G(mul_ex_n29), .D(mul_ex_N395), .Q(mul_ex_L_15_)
         );
  DLH_X2 mul_ex_L_reg_14_ ( .G(mul_ex_n29), .D(mul_ex_N396), .Q(mul_ex_L_14_)
         );
  DLH_X2 mul_ex_L_reg_13_ ( .G(mul_ex_n29), .D(mul_ex_N397), .Q(mul_ex_L_13_)
         );
  DLH_X2 mul_ex_L_reg_12_ ( .G(mul_ex_n29), .D(mul_ex_N398), .Q(mul_ex_L_12_)
         );
  DLH_X2 mul_ex_L_reg_11_ ( .G(mul_ex_n29), .D(mul_ex_N399), .Q(mul_ex_L_11_)
         );
  DLH_X2 mul_ex_L_reg_10_ ( .G(mul_ex_n28), .D(mul_ex_N400), .Q(mul_ex_L_10_)
         );
  DLH_X2 mul_ex_L_reg_9_ ( .G(mul_ex_n28), .D(mul_ex_N401), .Q(mul_ex_L_9_) );
  DLH_X2 mul_ex_L_reg_8_ ( .G(mul_ex_n28), .D(mul_ex_N402), .Q(mul_ex_L_8_) );
  DLH_X2 mul_ex_L_reg_7_ ( .G(mul_ex_n28), .D(mul_ex_N403), .Q(mul_ex_L_7_) );
  DLH_X2 mul_ex_L_reg_6_ ( .G(mul_ex_n28), .D(mul_ex_N404), .Q(mul_ex_L_6_) );
  DLH_X2 mul_ex_L_reg_5_ ( .G(mul_ex_n28), .D(mul_ex_N405), .Q(mul_ex_L_5_) );
  DLH_X2 mul_ex_L_reg_4_ ( .G(mul_ex_n28), .D(mul_ex_N406), .Q(mul_ex_L_4_) );
  DLH_X2 mul_ex_L_reg_3_ ( .G(mul_ex_n28), .D(mul_ex_N407), .Q(mul_ex_L_3_) );
  DLH_X2 mul_ex_L_reg_2_ ( .G(mul_ex_n28), .D(mul_ex_N408), .Q(mul_ex_L_2_) );
  DLH_X2 mul_ex_L_reg_1_ ( .G(mul_ex_n28), .D(mul_ex_N409), .Q(mul_ex_L_1_) );
  DLH_X2 mul_ex_L_reg_0_ ( .G(mul_ex_n28), .D(mul_ex_N410), .Q(mul_ex_L_0_) );
  DLH_X2 mul_ex_P1_reg_31_ ( .G(mul_ex_n32), .D(mul_ex_N88), .Q(mul_ex_P1[31])
         );
  DLH_X2 mul_ex_P1_reg_30_ ( .G(mul_ex_n32), .D(mul_ex_N89), .Q(mul_ex_P1[30])
         );
  DLH_X2 mul_ex_P1_reg_29_ ( .G(mul_ex_n32), .D(mul_ex_N90), .Q(mul_ex_P1[29])
         );
  DLH_X2 mul_ex_P1_reg_28_ ( .G(mul_ex_N43), .D(mul_ex_N91), .Q(mul_ex_P1[28])
         );
  DLH_X2 mul_ex_P1_reg_27_ ( .G(mul_ex_N43), .D(mul_ex_N92), .Q(mul_ex_P1[27])
         );
  DLH_X2 mul_ex_P1_reg_26_ ( .G(mul_ex_N43), .D(mul_ex_N93), .Q(mul_ex_P1[26])
         );
  DLH_X2 mul_ex_P1_reg_25_ ( .G(mul_ex_N43), .D(mul_ex_N94), .Q(mul_ex_P1[25])
         );
  DLH_X2 mul_ex_P1_reg_24_ ( .G(mul_ex_N43), .D(mul_ex_N95), .Q(mul_ex_P1[24])
         );
  DLH_X2 mul_ex_P1_reg_23_ ( .G(mul_ex_N43), .D(mul_ex_N96), .Q(mul_ex_P1[23])
         );
  DLH_X2 mul_ex_P1_reg_22_ ( .G(mul_ex_N43), .D(mul_ex_N97), .Q(mul_ex_P1[22])
         );
  DLH_X2 mul_ex_P1_reg_21_ ( .G(mul_ex_N43), .D(mul_ex_N98), .Q(mul_ex_P1[21])
         );
  DLH_X2 mul_ex_P1_reg_20_ ( .G(mul_ex_N43), .D(mul_ex_N99), .Q(mul_ex_P1[20])
         );
  DLH_X2 mul_ex_P1_reg_19_ ( .G(mul_ex_N43), .D(mul_ex_N100), .Q(mul_ex_P1[19]) );
  DLH_X2 mul_ex_P1_reg_18_ ( .G(mul_ex_N43), .D(mul_ex_N101), .Q(mul_ex_P1[18]) );
  DLH_X2 mul_ex_P1_reg_17_ ( .G(mul_ex_N43), .D(mul_ex_N102), .Q(mul_ex_P1[17]) );
  DLH_X2 mul_ex_P1_reg_16_ ( .G(mul_ex_N43), .D(mul_ex_N103), .Q(mul_ex_P1[16]) );
  DLH_X2 mul_ex_P1_reg_15_ ( .G(mul_ex_N43), .D(mul_ex_N104), .Q(mul_ex_P1[15]) );
  DLH_X2 mul_ex_P_reg_31_ ( .G(mul_ex_n24), .D(mul_ex_N445), .Q(mul_ex_P[31])
         );
  DLH_X2 mul_ex_P_reg_30_ ( .G(mul_ex_n24), .D(mul_ex_N446), .Q(mul_ex_P[30])
         );
  DLH_X2 mul_ex_P_reg_29_ ( .G(mul_ex_n24), .D(mul_ex_N447), .Q(mul_ex_P[29])
         );
  DLH_X2 mul_ex_P_reg_28_ ( .G(mul_ex_n24), .D(mul_ex_N448), .Q(mul_ex_P[28])
         );
  DLH_X2 mul_ex_P_reg_27_ ( .G(mul_ex_n24), .D(mul_ex_N449), .Q(mul_ex_P[27])
         );
  DLH_X2 mul_ex_P_reg_26_ ( .G(mul_ex_n24), .D(mul_ex_N450), .Q(mul_ex_P[26])
         );
  DLH_X2 mul_ex_P_reg_25_ ( .G(mul_ex_n24), .D(mul_ex_N451), .Q(mul_ex_P[25])
         );
  DLH_X2 mul_ex_P_reg_24_ ( .G(mul_ex_n24), .D(mul_ex_N452), .Q(mul_ex_P[24])
         );
  DLH_X2 mul_ex_P_reg_23_ ( .G(mul_ex_n24), .D(mul_ex_N453), .Q(mul_ex_P[23])
         );
  DLH_X2 mul_ex_P_reg_22_ ( .G(mul_ex_n24), .D(mul_ex_N454), .Q(mul_ex_P[22])
         );
  DLH_X2 mul_ex_P_reg_21_ ( .G(mul_ex_n23), .D(mul_ex_N455), .Q(mul_ex_P[21])
         );
  DLH_X2 mul_ex_P_reg_20_ ( .G(mul_ex_n23), .D(mul_ex_N456), .Q(mul_ex_P[20])
         );
  DLH_X2 mul_ex_P_reg_19_ ( .G(mul_ex_n23), .D(mul_ex_N457), .Q(mul_ex_P[19])
         );
  DLH_X2 mul_ex_P_reg_18_ ( .G(mul_ex_n23), .D(mul_ex_N458), .Q(mul_ex_P[18])
         );
  DLH_X2 mul_ex_P_reg_17_ ( .G(mul_ex_n23), .D(mul_ex_N459), .Q(mul_ex_P[17])
         );
  DLH_X2 mul_ex_P_reg_16_ ( .G(mul_ex_n23), .D(mul_ex_N460), .Q(mul_ex_P[16])
         );
  DLH_X2 mul_ex_P_reg_15_ ( .G(mul_ex_n23), .D(mul_ex_N461), .Q(mul_ex_P[15])
         );
  DLH_X2 mul_ex_P_reg_14_ ( .G(mul_ex_n23), .D(mul_ex_N462), .Q(mul_ex_P[14])
         );
  DLH_X2 mul_ex_P_reg_13_ ( .G(mul_ex_n23), .D(mul_ex_N463), .Q(mul_ex_P[13])
         );
  DLH_X2 mul_ex_P_reg_12_ ( .G(mul_ex_n23), .D(mul_ex_N464), .Q(mul_ex_P[12])
         );
  DLH_X2 mul_ex_P_reg_11_ ( .G(mul_ex_n23), .D(mul_ex_N465), .Q(mul_ex_P[11])
         );
  DLH_X2 mul_ex_P_reg_10_ ( .G(mul_ex_n22), .D(mul_ex_N466), .Q(mul_ex_P[10])
         );
  DLH_X2 mul_ex_P_reg_9_ ( .G(mul_ex_n22), .D(mul_ex_N467), .Q(mul_ex_P[9]) );
  DLH_X2 mul_ex_P_reg_8_ ( .G(mul_ex_n22), .D(mul_ex_N468), .Q(mul_ex_P[8]) );
  DLH_X2 mul_ex_P_reg_7_ ( .G(mul_ex_n22), .D(mul_ex_N469), .Q(mul_ex_P[7]) );
  DLH_X2 mul_ex_P_reg_6_ ( .G(mul_ex_n22), .D(mul_ex_N470), .Q(mul_ex_P[6]) );
  DLH_X2 mul_ex_P_reg_5_ ( .G(mul_ex_n22), .D(mul_ex_N471), .Q(mul_ex_P[5]) );
  DLH_X2 mul_ex_P_reg_4_ ( .G(mul_ex_n22), .D(mul_ex_N472), .Q(mul_ex_P[4]) );
  DLH_X2 mul_ex_P_reg_3_ ( .G(mul_ex_n22), .D(mul_ex_N473), .Q(mul_ex_P[3]) );
  DLH_X2 mul_ex_P_reg_2_ ( .G(mul_ex_n22), .D(mul_ex_N474), .Q(mul_ex_P[2]) );
  DLH_X2 mul_ex_P_reg_1_ ( .G(mul_ex_n22), .D(mul_ex_N475), .Q(mul_ex_P[1]) );
  DLH_X2 mul_ex_P_reg_0_ ( .G(mul_ex_n22), .D(mul_ex_N476), .Q(mul_ex_P[0]) );
  DLH_X2 mul_ex_done_reg ( .G(mul_ex_n8), .D(mul_ex_n18), .Q(mul_done) );
  DLH_X2 mul_ex_P2_reg_31_ ( .G(mul_ex_n15), .D(mul_ex_N105), .Q(mul_ex_P2[31]) );
  DLH_X2 mul_ex_P2_reg_30_ ( .G(mul_ex_n15), .D(mul_ex_N106), .Q(mul_ex_P2[30]) );
  DLH_X2 mul_ex_P2_reg_29_ ( .G(mul_ex_n15), .D(mul_ex_N107), .Q(mul_ex_P2[29]) );
  DLH_X2 mul_ex_P2_reg_28_ ( .G(mul_ex_n15), .D(mul_ex_N108), .Q(mul_ex_P2[28]) );
  DLH_X2 mul_ex_P2_reg_27_ ( .G(mul_ex_n15), .D(mul_ex_N109), .Q(mul_ex_P2[27]) );
  DLH_X2 mul_ex_P2_reg_26_ ( .G(mul_ex_n15), .D(mul_ex_N110), .Q(mul_ex_P2[26]) );
  DLH_X2 mul_ex_P2_reg_25_ ( .G(mul_ex_n15), .D(mul_ex_N111), .Q(mul_ex_P2[25]) );
  DLH_X2 mul_ex_P2_reg_24_ ( .G(mul_ex_n15), .D(mul_ex_N112), .Q(mul_ex_P2[24]) );
  DLH_X2 mul_ex_P2_reg_23_ ( .G(mul_ex_n15), .D(mul_ex_N113), .Q(mul_ex_P2[23]) );
  DLH_X2 mul_ex_P2_reg_22_ ( .G(mul_ex_n15), .D(mul_ex_N114), .Q(mul_ex_P2[22]) );
  DLH_X2 mul_ex_P2_reg_21_ ( .G(mul_ex_n15), .D(mul_ex_N115), .Q(mul_ex_P2[21]) );
  DLH_X2 mul_ex_P2_reg_20_ ( .G(mul_ex_n15), .D(mul_ex_N116), .Q(mul_ex_P2[20]) );
  DLH_X2 mul_ex_P2_reg_19_ ( .G(mul_ex_n15), .D(mul_ex_N117), .Q(mul_ex_P2[19]) );
  DLH_X2 mul_ex_P2_reg_18_ ( .G(mul_ex_n15), .D(mul_ex_N118), .Q(mul_ex_P2[18]) );
  DLH_X2 mul_ex_P2_reg_17_ ( .G(mul_ex_n15), .D(mul_ex_N119), .Q(mul_ex_P2[17]) );
  DLH_X2 mul_ex_P2_reg_16_ ( .G(mul_ex_n17), .D(mul_ex_N120), .Q(mul_ex_P2[16]) );
  DLH_X2 mul_ex_P2_reg_15_ ( .G(mul_ex_n17), .D(mul_ex_N121), .Q(mul_ex_P2[15]) );
  DFF_X2 mul_ex_CurrentState_reg_1_ ( .D(mul_ex_N15), .CK(clk), .Q(
        mul_ex_CurrentState_1_) );
  DFF_X2 mul_ex_CurrentState_reg_0_ ( .D(mul_ex_N16), .CK(clk), .Q(
        mul_ex_CurrentState_0_), .QN(mul_ex_n5) );
  DFF_X2 mul_ex_CurrentState_reg_2_ ( .D(mul_ex_N14), .CK(clk), .Q(
        mul_ex_CurrentState_2_), .QN(mul_ex_n4) );
  AND2_X2 mul_ex_U106 ( .A1(mul_ex_N122), .A2(mul_ex_n16), .ZN(mul_ex_N379) );
  AND2_X2 mul_ex_U105 ( .A1(mul_ex_N123), .A2(mul_ex_n16), .ZN(mul_ex_N380) );
  AND2_X2 mul_ex_U104 ( .A1(mul_ex_N124), .A2(mul_ex_n16), .ZN(mul_ex_N381) );
  AND2_X2 mul_ex_U103 ( .A1(mul_ex_N125), .A2(mul_ex_n16), .ZN(mul_ex_N382) );
  AND2_X2 mul_ex_U102 ( .A1(mul_ex_N126), .A2(mul_ex_n16), .ZN(mul_ex_N383) );
  AND2_X2 mul_ex_U101 ( .A1(mul_ex_N127), .A2(mul_ex_n16), .ZN(mul_ex_N384) );
  AND2_X2 mul_ex_U100 ( .A1(mul_ex_N128), .A2(mul_ex_n16), .ZN(mul_ex_N385) );
  AND2_X2 mul_ex_U99 ( .A1(mul_ex_N129), .A2(mul_ex_n16), .ZN(mul_ex_N386) );
  AND2_X2 mul_ex_U98 ( .A1(mul_ex_N130), .A2(mul_ex_n16), .ZN(mul_ex_N387) );
  AND2_X2 mul_ex_U97 ( .A1(mul_ex_N131), .A2(mul_ex_n16), .ZN(mul_ex_N388) );
  AND2_X2 mul_ex_U96 ( .A1(mul_ex_N132), .A2(mul_ex_n16), .ZN(mul_ex_N389) );
  AND2_X2 mul_ex_U95 ( .A1(mul_ex_N133), .A2(mul_ex_n16), .ZN(mul_ex_N390) );
  AND2_X2 mul_ex_U94 ( .A1(mul_ex_N134), .A2(mul_ex_n16), .ZN(mul_ex_N391) );
  AND2_X2 mul_ex_U93 ( .A1(mul_ex_N135), .A2(mul_ex_n16), .ZN(mul_ex_N392) );
  AND2_X2 mul_ex_U92 ( .A1(mul_ex_N136), .A2(mul_ex_n16), .ZN(mul_ex_N393) );
  AND2_X2 mul_ex_U91 ( .A1(mul_ex_N137), .A2(mul_ex_n16), .ZN(mul_ex_N394) );
  AND2_X2 mul_ex_U90 ( .A1(mul_ex_N138), .A2(mul_ex_n16), .ZN(mul_ex_N395) );
  AND2_X2 mul_ex_U89 ( .A1(mul_ex_N139), .A2(mul_ex_n16), .ZN(mul_ex_N396) );
  AND2_X2 mul_ex_U88 ( .A1(mul_ex_N140), .A2(mul_ex_n16), .ZN(mul_ex_N397) );
  AND2_X2 mul_ex_U87 ( .A1(mul_ex_N141), .A2(mul_ex_n16), .ZN(mul_ex_N398) );
  AND2_X2 mul_ex_U86 ( .A1(mul_ex_N142), .A2(mul_ex_n16), .ZN(mul_ex_N399) );
  AND2_X2 mul_ex_U85 ( .A1(mul_ex_N143), .A2(mul_ex_n16), .ZN(mul_ex_N400) );
  AND2_X2 mul_ex_U84 ( .A1(mul_ex_N144), .A2(mul_ex_n17), .ZN(mul_ex_N401) );
  AND2_X2 mul_ex_U83 ( .A1(mul_ex_N145), .A2(mul_ex_n17), .ZN(mul_ex_N402) );
  AND2_X2 mul_ex_U82 ( .A1(mul_ex_N146), .A2(mul_ex_n17), .ZN(mul_ex_N403) );
  AND2_X2 mul_ex_U81 ( .A1(mul_ex_N147), .A2(mul_ex_n17), .ZN(mul_ex_N404) );
  AND2_X2 mul_ex_U80 ( .A1(mul_ex_N148), .A2(mul_ex_n17), .ZN(mul_ex_N405) );
  AND2_X2 mul_ex_U79 ( .A1(mul_ex_N149), .A2(mul_ex_n17), .ZN(mul_ex_N406) );
  AND2_X2 mul_ex_U78 ( .A1(mul_ex_N150), .A2(mul_ex_n17), .ZN(mul_ex_N407) );
  AND2_X2 mul_ex_U77 ( .A1(mul_ex_N151), .A2(mul_ex_n17), .ZN(mul_ex_N408) );
  AND2_X2 mul_ex_U76 ( .A1(mul_ex_N152), .A2(mul_ex_n17), .ZN(mul_ex_N409) );
  AND2_X2 mul_ex_U75 ( .A1(mul_ex_N153), .A2(mul_ex_n17), .ZN(mul_ex_N410) );
  AND2_X2 mul_ex_U73 ( .A1(mul_ex_N218), .A2(mul_ex_n14), .ZN(mul_ex_N412) );
  AND2_X2 mul_ex_U72 ( .A1(mul_ex_N219), .A2(mul_ex_n14), .ZN(mul_ex_N413) );
  AND2_X2 mul_ex_U71 ( .A1(mul_ex_N220), .A2(mul_ex_n14), .ZN(mul_ex_N414) );
  AND2_X2 mul_ex_U70 ( .A1(mul_ex_N221), .A2(mul_ex_n14), .ZN(mul_ex_N415) );
  AND2_X2 mul_ex_U69 ( .A1(mul_ex_N222), .A2(mul_ex_n14), .ZN(mul_ex_N416) );
  AND2_X2 mul_ex_U68 ( .A1(mul_ex_N223), .A2(mul_ex_n14), .ZN(mul_ex_N417) );
  AND2_X2 mul_ex_U67 ( .A1(mul_ex_N224), .A2(mul_ex_n14), .ZN(mul_ex_N418) );
  AND2_X2 mul_ex_U66 ( .A1(mul_ex_N225), .A2(mul_ex_n14), .ZN(mul_ex_N419) );
  AND2_X2 mul_ex_U65 ( .A1(mul_ex_N226), .A2(mul_ex_n14), .ZN(mul_ex_N420) );
  AND2_X2 mul_ex_U64 ( .A1(mul_ex_N227), .A2(mul_ex_n14), .ZN(mul_ex_N421) );
  AND2_X2 mul_ex_U63 ( .A1(mul_ex_N228), .A2(mul_ex_n13), .ZN(mul_ex_N422) );
  AND2_X2 mul_ex_U62 ( .A1(mul_ex_N229), .A2(mul_ex_n13), .ZN(mul_ex_N423) );
  AND2_X2 mul_ex_U61 ( .A1(mul_ex_N230), .A2(mul_ex_n13), .ZN(mul_ex_N424) );
  AND2_X2 mul_ex_U60 ( .A1(mul_ex_N231), .A2(mul_ex_n13), .ZN(mul_ex_N425) );
  AND2_X2 mul_ex_U59 ( .A1(mul_ex_N232), .A2(mul_ex_n13), .ZN(mul_ex_N426) );
  AND2_X2 mul_ex_U58 ( .A1(mul_ex_N233), .A2(mul_ex_n13), .ZN(mul_ex_N427) );
  AND2_X2 mul_ex_U57 ( .A1(mul_ex_N234), .A2(mul_ex_n13), .ZN(mul_ex_N428) );
  AND2_X2 mul_ex_U56 ( .A1(mul_ex_N235), .A2(mul_ex_n13), .ZN(mul_ex_N429) );
  AND2_X2 mul_ex_U55 ( .A1(mul_ex_N236), .A2(mul_ex_n13), .ZN(mul_ex_N430) );
  AND2_X2 mul_ex_U54 ( .A1(mul_ex_N237), .A2(mul_ex_n13), .ZN(mul_ex_N431) );
  AND2_X2 mul_ex_U53 ( .A1(mul_ex_N238), .A2(mul_ex_n13), .ZN(mul_ex_N432) );
  AND2_X2 mul_ex_U52 ( .A1(mul_ex_N239), .A2(mul_ex_n12), .ZN(mul_ex_N433) );
  AND2_X2 mul_ex_U51 ( .A1(mul_ex_N240), .A2(mul_ex_n12), .ZN(mul_ex_N434) );
  AND2_X2 mul_ex_U50 ( .A1(mul_ex_N241), .A2(mul_ex_n12), .ZN(mul_ex_N435) );
  AND2_X2 mul_ex_U49 ( .A1(mul_ex_N242), .A2(mul_ex_n12), .ZN(mul_ex_N436) );
  AND2_X2 mul_ex_U48 ( .A1(mul_ex_N243), .A2(mul_ex_n12), .ZN(mul_ex_N437) );
  AND2_X2 mul_ex_U47 ( .A1(mul_ex_N244), .A2(mul_ex_n12), .ZN(mul_ex_N438) );
  AND2_X2 mul_ex_U46 ( .A1(mul_ex_N245), .A2(mul_ex_n12), .ZN(mul_ex_N439) );
  AND2_X2 mul_ex_U45 ( .A1(mul_ex_N246), .A2(mul_ex_n12), .ZN(mul_ex_N440) );
  AND2_X2 mul_ex_U44 ( .A1(mul_ex_N247), .A2(mul_ex_n12), .ZN(mul_ex_N441) );
  AND2_X2 mul_ex_U43 ( .A1(mul_ex_N248), .A2(mul_ex_n12), .ZN(mul_ex_N442) );
  AND2_X2 mul_ex_U42 ( .A1(mul_ex_N249), .A2(mul_ex_n12), .ZN(mul_ex_N443) );
  AND2_X2 mul_ex_U40 ( .A1(mul_ex_N154), .A2(mul_ex_n11), .ZN(mul_ex_N445) );
  AND2_X2 mul_ex_U39 ( .A1(mul_ex_N155), .A2(mul_ex_n11), .ZN(mul_ex_N446) );
  AND2_X2 mul_ex_U38 ( .A1(mul_ex_N156), .A2(mul_ex_n11), .ZN(mul_ex_N447) );
  AND2_X2 mul_ex_U37 ( .A1(mul_ex_N157), .A2(mul_ex_n11), .ZN(mul_ex_N448) );
  AND2_X2 mul_ex_U36 ( .A1(mul_ex_N158), .A2(mul_ex_n11), .ZN(mul_ex_N449) );
  AND2_X2 mul_ex_U35 ( .A1(mul_ex_N159), .A2(mul_ex_n11), .ZN(mul_ex_N450) );
  AND2_X2 mul_ex_U34 ( .A1(mul_ex_N160), .A2(mul_ex_n11), .ZN(mul_ex_N451) );
  AND2_X2 mul_ex_U33 ( .A1(mul_ex_N161), .A2(mul_ex_n11), .ZN(mul_ex_N452) );
  AND2_X2 mul_ex_U32 ( .A1(mul_ex_N162), .A2(mul_ex_n11), .ZN(mul_ex_N453) );
  AND2_X2 mul_ex_U31 ( .A1(mul_ex_N163), .A2(mul_ex_n11), .ZN(mul_ex_N454) );
  AND2_X2 mul_ex_U30 ( .A1(mul_ex_N164), .A2(mul_ex_n11), .ZN(mul_ex_N455) );
  AND2_X2 mul_ex_U29 ( .A1(mul_ex_N165), .A2(mul_ex_n11), .ZN(mul_ex_N456) );
  AND2_X2 mul_ex_U28 ( .A1(mul_ex_N166), .A2(mul_ex_n11), .ZN(mul_ex_N457) );
  AND2_X2 mul_ex_U27 ( .A1(mul_ex_N167), .A2(mul_ex_n11), .ZN(mul_ex_N458) );
  AND2_X2 mul_ex_U26 ( .A1(mul_ex_N168), .A2(mul_ex_n11), .ZN(mul_ex_N459) );
  AND2_X2 mul_ex_U25 ( .A1(mul_ex_N169), .A2(mul_ex_n11), .ZN(mul_ex_N460) );
  AND2_X2 mul_ex_U24 ( .A1(mul_ex_N170), .A2(mul_ex_n11), .ZN(mul_ex_N461) );
  AND2_X2 mul_ex_U23 ( .A1(mul_ex_N171), .A2(mul_ex_n11), .ZN(mul_ex_N462) );
  AND2_X2 mul_ex_U22 ( .A1(mul_ex_N172), .A2(mul_ex_n11), .ZN(mul_ex_N463) );
  AND2_X2 mul_ex_U21 ( .A1(mul_ex_N173), .A2(mul_ex_n11), .ZN(mul_ex_N464) );
  AND2_X2 mul_ex_U20 ( .A1(mul_ex_N174), .A2(mul_ex_n11), .ZN(mul_ex_N465) );
  AND2_X2 mul_ex_U19 ( .A1(mul_ex_N175), .A2(mul_ex_n11), .ZN(mul_ex_N466) );
  AND2_X2 mul_ex_U18 ( .A1(mul_ex_N176), .A2(mul_ex_n39), .ZN(mul_ex_N467) );
  AND2_X2 mul_ex_U17 ( .A1(mul_ex_N177), .A2(mul_ex_n39), .ZN(mul_ex_N468) );
  AND2_X2 mul_ex_U16 ( .A1(mul_ex_N178), .A2(mul_ex_n39), .ZN(mul_ex_N469) );
  AND2_X2 mul_ex_U15 ( .A1(mul_ex_N179), .A2(mul_ex_n39), .ZN(mul_ex_N470) );
  AND2_X2 mul_ex_U14 ( .A1(mul_ex_N180), .A2(mul_ex_n39), .ZN(mul_ex_N471) );
  AND2_X2 mul_ex_U13 ( .A1(mul_ex_N181), .A2(mul_ex_n39), .ZN(mul_ex_N472) );
  AND2_X2 mul_ex_U12 ( .A1(mul_ex_N182), .A2(mul_ex_n39), .ZN(mul_ex_N473) );
  AND2_X2 mul_ex_U11 ( .A1(mul_ex_N183), .A2(mul_ex_n39), .ZN(mul_ex_N474) );
  AND2_X2 mul_ex_U10 ( .A1(mul_ex_N184), .A2(mul_ex_n39), .ZN(mul_ex_N475) );
  AND2_X2 mul_ex_U9 ( .A1(mul_ex_N185), .A2(mul_ex_n39), .ZN(mul_ex_N476) );
  AND2_X4 mul_ex_add_85_U2 ( .A1(f2_in[31]), .A2(f2_in[15]), .ZN(
        mul_ex_add_85_n2) );
  XOR2_X2 mul_ex_add_85_U1 ( .A(f2_in[31]), .B(f2_in[15]), .Z(mul_ex_N105) );
  FA_X1 mul_ex_add_85_U1_1 ( .A(f2_in[14]), .B(f2_in[30]), .CI(
        mul_ex_add_85_n2), .CO(mul_ex_add_85_carry[2]), .S(mul_ex_N106) );
  FA_X1 mul_ex_add_85_U1_2 ( .A(f2_in[13]), .B(f2_in[29]), .CI(
        mul_ex_add_85_carry[2]), .CO(mul_ex_add_85_carry[3]), .S(mul_ex_N107)
         );
  FA_X1 mul_ex_add_85_U1_3 ( .A(f2_in[12]), .B(f2_in[28]), .CI(
        mul_ex_add_85_carry[3]), .CO(mul_ex_add_85_carry[4]), .S(mul_ex_N108)
         );
  FA_X1 mul_ex_add_85_U1_4 ( .A(f2_in[11]), .B(f2_in[27]), .CI(
        mul_ex_add_85_carry[4]), .CO(mul_ex_add_85_carry[5]), .S(mul_ex_N109)
         );
  FA_X1 mul_ex_add_85_U1_5 ( .A(f2_in[10]), .B(f2_in[26]), .CI(
        mul_ex_add_85_carry[5]), .CO(mul_ex_add_85_carry[6]), .S(mul_ex_N110)
         );
  FA_X1 mul_ex_add_85_U1_6 ( .A(f2_in[9]), .B(f2_in[25]), .CI(
        mul_ex_add_85_carry[6]), .CO(mul_ex_add_85_carry[7]), .S(mul_ex_N111)
         );
  FA_X1 mul_ex_add_85_U1_7 ( .A(f2_in[8]), .B(f2_in[24]), .CI(
        mul_ex_add_85_carry[7]), .CO(mul_ex_add_85_carry[8]), .S(mul_ex_N112)
         );
  FA_X1 mul_ex_add_85_U1_8 ( .A(f2_in[7]), .B(f2_in[23]), .CI(
        mul_ex_add_85_carry[8]), .CO(mul_ex_add_85_carry[9]), .S(mul_ex_N113)
         );
  FA_X1 mul_ex_add_85_U1_9 ( .A(f2_in[6]), .B(f2_in[22]), .CI(
        mul_ex_add_85_carry[9]), .CO(mul_ex_add_85_carry[10]), .S(mul_ex_N114)
         );
  FA_X1 mul_ex_add_85_U1_10 ( .A(f2_in[5]), .B(f2_in[21]), .CI(
        mul_ex_add_85_carry[10]), .CO(mul_ex_add_85_carry[11]), .S(mul_ex_N115) );
  FA_X1 mul_ex_add_85_U1_11 ( .A(f2_in[4]), .B(f2_in[20]), .CI(
        mul_ex_add_85_carry[11]), .CO(mul_ex_add_85_carry[12]), .S(mul_ex_N116) );
  FA_X1 mul_ex_add_85_U1_12 ( .A(f2_in[3]), .B(f2_in[19]), .CI(
        mul_ex_add_85_carry[12]), .CO(mul_ex_add_85_carry[13]), .S(mul_ex_N117) );
  FA_X1 mul_ex_add_85_U1_13 ( .A(f2_in[2]), .B(f2_in[18]), .CI(
        mul_ex_add_85_carry[13]), .CO(mul_ex_add_85_carry[14]), .S(mul_ex_N118) );
  FA_X1 mul_ex_add_85_U1_14 ( .A(f2_in[1]), .B(f2_in[17]), .CI(
        mul_ex_add_85_carry[14]), .CO(mul_ex_add_85_carry[15]), .S(mul_ex_N119) );
  FA_X1 mul_ex_add_85_U1_15 ( .A(f2_in[0]), .B(f2_in[16]), .CI(
        mul_ex_add_85_carry[15]), .CO(mul_ex_N121), .S(mul_ex_N120) );
  AND2_X4 mul_ex_add_77_U2 ( .A1(f1_in[31]), .A2(f1_in[15]), .ZN(
        mul_ex_add_77_n2) );
  XOR2_X2 mul_ex_add_77_U1 ( .A(f1_in[31]), .B(f1_in[15]), .Z(mul_ex_N88) );
  FA_X1 mul_ex_add_77_U1_1 ( .A(f1_in[14]), .B(f1_in[30]), .CI(
        mul_ex_add_77_n2), .CO(mul_ex_add_77_carry[2]), .S(mul_ex_N89) );
  FA_X1 mul_ex_add_77_U1_2 ( .A(f1_in[13]), .B(f1_in[29]), .CI(
        mul_ex_add_77_carry[2]), .CO(mul_ex_add_77_carry[3]), .S(mul_ex_N90)
         );
  FA_X1 mul_ex_add_77_U1_3 ( .A(f1_in[12]), .B(f1_in[28]), .CI(
        mul_ex_add_77_carry[3]), .CO(mul_ex_add_77_carry[4]), .S(mul_ex_N91)
         );
  FA_X1 mul_ex_add_77_U1_4 ( .A(f1_in[11]), .B(f1_in[27]), .CI(
        mul_ex_add_77_carry[4]), .CO(mul_ex_add_77_carry[5]), .S(mul_ex_N92)
         );
  FA_X1 mul_ex_add_77_U1_5 ( .A(f1_in[10]), .B(f1_in[26]), .CI(
        mul_ex_add_77_carry[5]), .CO(mul_ex_add_77_carry[6]), .S(mul_ex_N93)
         );
  FA_X1 mul_ex_add_77_U1_6 ( .A(f1_in[9]), .B(f1_in[25]), .CI(
        mul_ex_add_77_carry[6]), .CO(mul_ex_add_77_carry[7]), .S(mul_ex_N94)
         );
  FA_X1 mul_ex_add_77_U1_7 ( .A(f1_in[8]), .B(f1_in[24]), .CI(
        mul_ex_add_77_carry[7]), .CO(mul_ex_add_77_carry[8]), .S(mul_ex_N95)
         );
  FA_X1 mul_ex_add_77_U1_8 ( .A(f1_in[7]), .B(f1_in[23]), .CI(
        mul_ex_add_77_carry[8]), .CO(mul_ex_add_77_carry[9]), .S(mul_ex_N96)
         );
  FA_X1 mul_ex_add_77_U1_9 ( .A(f1_in[6]), .B(f1_in[22]), .CI(
        mul_ex_add_77_carry[9]), .CO(mul_ex_add_77_carry[10]), .S(mul_ex_N97)
         );
  FA_X1 mul_ex_add_77_U1_10 ( .A(f1_in[5]), .B(f1_in[21]), .CI(
        mul_ex_add_77_carry[10]), .CO(mul_ex_add_77_carry[11]), .S(mul_ex_N98)
         );
  FA_X1 mul_ex_add_77_U1_11 ( .A(f1_in[4]), .B(f1_in[20]), .CI(
        mul_ex_add_77_carry[11]), .CO(mul_ex_add_77_carry[12]), .S(mul_ex_N99)
         );
  FA_X1 mul_ex_add_77_U1_12 ( .A(f1_in[3]), .B(f1_in[19]), .CI(
        mul_ex_add_77_carry[12]), .CO(mul_ex_add_77_carry[13]), .S(mul_ex_N100) );
  FA_X1 mul_ex_add_77_U1_13 ( .A(f1_in[2]), .B(f1_in[18]), .CI(
        mul_ex_add_77_carry[13]), .CO(mul_ex_add_77_carry[14]), .S(mul_ex_N101) );
  FA_X1 mul_ex_add_77_U1_14 ( .A(f1_in[1]), .B(f1_in[17]), .CI(
        mul_ex_add_77_carry[14]), .CO(mul_ex_add_77_carry[15]), .S(mul_ex_N102) );
  FA_X1 mul_ex_add_77_U1_15 ( .A(f1_in[0]), .B(f1_in[16]), .CI(
        mul_ex_add_77_carry[15]), .CO(mul_ex_N104), .S(mul_ex_N103) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U50 ( .A(mul_ex_L_16_), .Z(
        mul_ex_N265) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U49 ( .A(mul_ex_L_17_), .Z(
        mul_ex_N264) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U48 ( .A(mul_ex_L_18_), .Z(
        mul_ex_N263) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U47 ( .A(mul_ex_L_19_), .Z(
        mul_ex_N262) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U46 ( .A(mul_ex_L_20_), .Z(
        mul_ex_N261) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U45 ( .A(mul_ex_L_21_), .Z(
        mul_ex_N260) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U44 ( .A(mul_ex_L_22_), .Z(
        mul_ex_N259) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U43 ( .A(mul_ex_L_23_), .Z(
        mul_ex_N258) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U42 ( .A(mul_ex_L_24_), .Z(
        mul_ex_N257) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U41 ( .A(mul_ex_L_25_), .Z(
        mul_ex_N256) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U40 ( .A(mul_ex_L_26_), .Z(
        mul_ex_N255) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U39 ( .A(mul_ex_L_27_), .Z(
        mul_ex_N254) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U38 ( .A(mul_ex_L_28_), .Z(
        mul_ex_N253) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U37 ( .A(mul_ex_L_29_), .Z(
        mul_ex_N252) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U36 ( .A(mul_ex_L_30_), .Z(
        mul_ex_N251) );
  BUF_X32 mul_ex_add_1_root_add_0_root_add_98_2_U35 ( .A(mul_ex_L_31_), .Z(
        mul_ex_N250) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U34 ( .A(mul_ex_Z_31_), .B(
        mul_ex_L_15_), .Z(mul_ex_N266) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U33 ( .A1(mul_ex_Z_31_), .A2(
        mul_ex_L_15_), .ZN(mul_ex_add_1_root_add_0_root_add_98_2_n33) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U32 ( .A1(mul_ex_Z_0_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_n10), .ZN(mul_ex_N298) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U31 ( .A(mul_ex_Z_0_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_n10), .Z(mul_ex_N297) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U30 ( .A(mul_ex_Z_1_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_n2), .Z(mul_ex_N296) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U29 ( .A(mul_ex_Z_2_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_n11), .Z(mul_ex_N295) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U28 ( .A(mul_ex_Z_3_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_n3), .Z(mul_ex_N294) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U27 ( .A(mul_ex_Z_4_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_n12), .Z(mul_ex_N293) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U26 ( .A(mul_ex_Z_5_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_n4), .Z(mul_ex_N292) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U25 ( .A(mul_ex_Z_6_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_n13), .Z(mul_ex_N291) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U24 ( .A(mul_ex_Z_7_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_n5), .Z(mul_ex_N290) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U23 ( .A(mul_ex_Z_8_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_n14), .Z(mul_ex_N289) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U22 ( .A(mul_ex_Z_9_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_n6), .Z(mul_ex_N288) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U21 ( .A(mul_ex_Z_10_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_n15), .Z(mul_ex_N287) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U20 ( .A(mul_ex_Z_11_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_n7), .Z(mul_ex_N286) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U19 ( .A(mul_ex_Z_12_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_n16), .Z(mul_ex_N285) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U18 ( .A(mul_ex_Z_13_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_n8), .Z(mul_ex_N284) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U17 ( .A1(mul_ex_Z_15_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_carry_32_), .ZN(
        mul_ex_add_1_root_add_0_root_add_98_2_n17) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U16 ( .A1(mul_ex_Z_13_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_n8), .ZN(
        mul_ex_add_1_root_add_0_root_add_98_2_n16) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U15 ( .A1(mul_ex_Z_11_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_n7), .ZN(
        mul_ex_add_1_root_add_0_root_add_98_2_n15) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U14 ( .A1(mul_ex_Z_9_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_n6), .ZN(
        mul_ex_add_1_root_add_0_root_add_98_2_n14) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U13 ( .A1(mul_ex_Z_7_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_n5), .ZN(
        mul_ex_add_1_root_add_0_root_add_98_2_n13) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U12 ( .A1(mul_ex_Z_5_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_n4), .ZN(
        mul_ex_add_1_root_add_0_root_add_98_2_n12) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U11 ( .A1(mul_ex_Z_3_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_n3), .ZN(
        mul_ex_add_1_root_add_0_root_add_98_2_n11) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U10 ( .A1(mul_ex_Z_1_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_n2), .ZN(
        mul_ex_add_1_root_add_0_root_add_98_2_n10) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U9 ( .A(mul_ex_Z_15_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_carry_32_), .Z(mul_ex_N282) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U8 ( .A1(mul_ex_Z_14_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_n17), .ZN(
        mul_ex_add_1_root_add_0_root_add_98_2_n8) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U7 ( .A1(mul_ex_Z_12_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_n16), .ZN(
        mul_ex_add_1_root_add_0_root_add_98_2_n7) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U6 ( .A1(mul_ex_Z_10_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_n15), .ZN(
        mul_ex_add_1_root_add_0_root_add_98_2_n6) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U5 ( .A1(mul_ex_Z_8_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_n14), .ZN(
        mul_ex_add_1_root_add_0_root_add_98_2_n5) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U4 ( .A1(mul_ex_Z_6_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_n13), .ZN(
        mul_ex_add_1_root_add_0_root_add_98_2_n4) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U3 ( .A1(mul_ex_Z_4_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_n12), .ZN(
        mul_ex_add_1_root_add_0_root_add_98_2_n3) );
  AND2_X4 mul_ex_add_1_root_add_0_root_add_98_2_U2 ( .A1(mul_ex_Z_2_), .A2(
        mul_ex_add_1_root_add_0_root_add_98_2_n11), .ZN(
        mul_ex_add_1_root_add_0_root_add_98_2_n2) );
  XOR2_X2 mul_ex_add_1_root_add_0_root_add_98_2_U1 ( .A(mul_ex_Z_14_), .B(
        mul_ex_add_1_root_add_0_root_add_98_2_n17), .Z(mul_ex_N283) );
  FA_X1 mul_ex_add_1_root_add_0_root_add_98_2_U1_17 ( .A(mul_ex_L_14_), .B(
        mul_ex_Z_30_), .CI(mul_ex_add_1_root_add_0_root_add_98_2_n33), .CO(
        mul_ex_add_1_root_add_0_root_add_98_2_carry_18_), .S(mul_ex_N267) );
  FA_X1 mul_ex_add_1_root_add_0_root_add_98_2_U1_18 ( .A(mul_ex_L_13_), .B(
        mul_ex_Z_29_), .CI(mul_ex_add_1_root_add_0_root_add_98_2_carry_18_), 
        .CO(mul_ex_add_1_root_add_0_root_add_98_2_carry_19_), .S(mul_ex_N268)
         );
  FA_X1 mul_ex_add_1_root_add_0_root_add_98_2_U1_19 ( .A(mul_ex_L_12_), .B(
        mul_ex_Z_28_), .CI(mul_ex_add_1_root_add_0_root_add_98_2_carry_19_), 
        .CO(mul_ex_add_1_root_add_0_root_add_98_2_carry_20_), .S(mul_ex_N269)
         );
  FA_X1 mul_ex_add_1_root_add_0_root_add_98_2_U1_20 ( .A(mul_ex_L_11_), .B(
        mul_ex_Z_27_), .CI(mul_ex_add_1_root_add_0_root_add_98_2_carry_20_), 
        .CO(mul_ex_add_1_root_add_0_root_add_98_2_carry_21_), .S(mul_ex_N270)
         );
  FA_X1 mul_ex_add_1_root_add_0_root_add_98_2_U1_21 ( .A(mul_ex_L_10_), .B(
        mul_ex_Z_26_), .CI(mul_ex_add_1_root_add_0_root_add_98_2_carry_21_), 
        .CO(mul_ex_add_1_root_add_0_root_add_98_2_carry_22_), .S(mul_ex_N271)
         );
  FA_X1 mul_ex_add_1_root_add_0_root_add_98_2_U1_22 ( .A(mul_ex_L_9_), .B(
        mul_ex_Z_25_), .CI(mul_ex_add_1_root_add_0_root_add_98_2_carry_22_), 
        .CO(mul_ex_add_1_root_add_0_root_add_98_2_carry_23_), .S(mul_ex_N272)
         );
  FA_X1 mul_ex_add_1_root_add_0_root_add_98_2_U1_23 ( .A(mul_ex_L_8_), .B(
        mul_ex_Z_24_), .CI(mul_ex_add_1_root_add_0_root_add_98_2_carry_23_), 
        .CO(mul_ex_add_1_root_add_0_root_add_98_2_carry_24_), .S(mul_ex_N273)
         );
  FA_X1 mul_ex_add_1_root_add_0_root_add_98_2_U1_24 ( .A(mul_ex_L_7_), .B(
        mul_ex_Z_23_), .CI(mul_ex_add_1_root_add_0_root_add_98_2_carry_24_), 
        .CO(mul_ex_add_1_root_add_0_root_add_98_2_carry_25_), .S(mul_ex_N274)
         );
  FA_X1 mul_ex_add_1_root_add_0_root_add_98_2_U1_25 ( .A(mul_ex_L_6_), .B(
        mul_ex_Z_22_), .CI(mul_ex_add_1_root_add_0_root_add_98_2_carry_25_), 
        .CO(mul_ex_add_1_root_add_0_root_add_98_2_carry_26_), .S(mul_ex_N275)
         );
  FA_X1 mul_ex_add_1_root_add_0_root_add_98_2_U1_26 ( .A(mul_ex_L_5_), .B(
        mul_ex_Z_21_), .CI(mul_ex_add_1_root_add_0_root_add_98_2_carry_26_), 
        .CO(mul_ex_add_1_root_add_0_root_add_98_2_carry_27_), .S(mul_ex_N276)
         );
  FA_X1 mul_ex_add_1_root_add_0_root_add_98_2_U1_27 ( .A(mul_ex_L_4_), .B(
        mul_ex_Z_20_), .CI(mul_ex_add_1_root_add_0_root_add_98_2_carry_27_), 
        .CO(mul_ex_add_1_root_add_0_root_add_98_2_carry_28_), .S(mul_ex_N277)
         );
  FA_X1 mul_ex_add_1_root_add_0_root_add_98_2_U1_28 ( .A(mul_ex_L_3_), .B(
        mul_ex_Z_19_), .CI(mul_ex_add_1_root_add_0_root_add_98_2_carry_28_), 
        .CO(mul_ex_add_1_root_add_0_root_add_98_2_carry_29_), .S(mul_ex_N278)
         );
  FA_X1 mul_ex_add_1_root_add_0_root_add_98_2_U1_29 ( .A(mul_ex_L_2_), .B(
        mul_ex_Z_18_), .CI(mul_ex_add_1_root_add_0_root_add_98_2_carry_29_), 
        .CO(mul_ex_add_1_root_add_0_root_add_98_2_carry_30_), .S(mul_ex_N279)
         );
  FA_X1 mul_ex_add_1_root_add_0_root_add_98_2_U1_30 ( .A(mul_ex_L_1_), .B(
        mul_ex_Z_17_), .CI(mul_ex_add_1_root_add_0_root_add_98_2_carry_30_), 
        .CO(mul_ex_add_1_root_add_0_root_add_98_2_carry_31_), .S(mul_ex_N280)
         );
  FA_X1 mul_ex_add_1_root_add_0_root_add_98_2_U1_31 ( .A(mul_ex_L_0_), .B(
        mul_ex_Z_16_), .CI(mul_ex_add_1_root_add_0_root_add_98_2_carry_31_), 
        .CO(mul_ex_add_1_root_add_0_root_add_98_2_carry_32_), .S(mul_ex_N281)
         );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U63 ( .A(mul_ex_N281), .Z(
        mul_ex_N345) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U62 ( .A(mul_ex_N280), .Z(
        mul_ex_N344) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U61 ( .A(mul_ex_N279), .Z(
        mul_ex_N343) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U60 ( .A(mul_ex_N278), .Z(
        mul_ex_N342) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U59 ( .A(mul_ex_N277), .Z(
        mul_ex_N341) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U58 ( .A(mul_ex_N276), .Z(
        mul_ex_N340) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U57 ( .A(mul_ex_N275), .Z(
        mul_ex_N339) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U56 ( .A(mul_ex_N274), .Z(
        mul_ex_N338) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U55 ( .A(mul_ex_N273), .Z(
        mul_ex_N337) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U54 ( .A(mul_ex_N272), .Z(
        mul_ex_N336) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U53 ( .A(mul_ex_N271), .Z(
        mul_ex_N335) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U52 ( .A(mul_ex_N270), .Z(
        mul_ex_N334) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U51 ( .A(mul_ex_N269), .Z(
        mul_ex_N333) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U50 ( .A(mul_ex_N268), .Z(
        mul_ex_N332) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U49 ( .A(mul_ex_N267), .Z(
        mul_ex_N331) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U48 ( .A(mul_ex_N266), .Z(
        mul_ex_N330) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U47 ( .A(mul_ex_N265), .Z(
        mul_ex_N329) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U46 ( .A(mul_ex_N264), .Z(
        mul_ex_N328) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U45 ( .A(mul_ex_N263), .Z(
        mul_ex_N327) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U44 ( .A(mul_ex_N262), .Z(
        mul_ex_N326) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U43 ( .A(mul_ex_N261), .Z(
        mul_ex_N325) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U42 ( .A(mul_ex_N260), .Z(
        mul_ex_N324) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U41 ( .A(mul_ex_N259), .Z(
        mul_ex_N323) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U40 ( .A(mul_ex_N258), .Z(
        mul_ex_N322) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U39 ( .A(mul_ex_N257), .Z(
        mul_ex_N321) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U38 ( .A(mul_ex_N256), .Z(
        mul_ex_N320) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U37 ( .A(mul_ex_N255), .Z(
        mul_ex_N319) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U36 ( .A(mul_ex_N254), .Z(
        mul_ex_N318) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U35 ( .A(mul_ex_N253), .Z(
        mul_ex_N317) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U34 ( .A(mul_ex_N252), .Z(
        mul_ex_N316) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U33 ( .A(mul_ex_N251), .Z(
        mul_ex_N315) );
  BUF_X32 mul_ex_add_0_root_add_0_root_add_98_2_U32 ( .A(mul_ex_N250), .Z(
        mul_ex_N314) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U31 ( .A(mul_ex_Z_0_), .B(
        mul_ex_add_0_root_add_0_root_add_98_2_n15), .Z(mul_ex_N377) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U30 ( .A(mul_ex_Z_1_), .B(
        mul_ex_add_0_root_add_0_root_add_98_2_n7), .Z(mul_ex_N376) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U29 ( .A(mul_ex_Z_2_), .B(
        mul_ex_add_0_root_add_0_root_add_98_2_n1), .Z(mul_ex_N375) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U28 ( .A(mul_ex_Z_3_), .B(
        mul_ex_add_0_root_add_0_root_add_98_2_n8), .Z(mul_ex_N374) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U27 ( .A(mul_ex_Z_4_), .B(
        mul_ex_add_0_root_add_0_root_add_98_2_n2), .Z(mul_ex_N373) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U26 ( .A(mul_ex_Z_5_), .B(
        mul_ex_add_0_root_add_0_root_add_98_2_n9), .Z(mul_ex_N372) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U25 ( .A(mul_ex_Z_6_), .B(
        mul_ex_add_0_root_add_0_root_add_98_2_n3), .Z(mul_ex_N371) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U24 ( .A(mul_ex_Z_7_), .B(
        mul_ex_add_0_root_add_0_root_add_98_2_n10), .Z(mul_ex_N370) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U23 ( .A(mul_ex_Z_8_), .B(
        mul_ex_add_0_root_add_0_root_add_98_2_n4), .Z(mul_ex_N369) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U22 ( .A(mul_ex_Z_9_), .B(
        mul_ex_add_0_root_add_0_root_add_98_2_n11), .Z(mul_ex_N368) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U21 ( .A(mul_ex_Z_10_), .B(
        mul_ex_add_0_root_add_0_root_add_98_2_n5), .Z(mul_ex_N367) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U20 ( .A(mul_ex_Z_11_), .B(
        mul_ex_add_0_root_add_0_root_add_98_2_n12), .Z(mul_ex_N366) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U19 ( .A(mul_ex_Z_12_), .B(
        mul_ex_add_0_root_add_0_root_add_98_2_n6), .Z(mul_ex_N365) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U18 ( .A(mul_ex_Z_13_), .B(
        mul_ex_add_0_root_add_0_root_add_98_2_n13), .Z(mul_ex_N364) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U17 ( .A(mul_ex_N282), .B(
        mul_ex_Z_31_), .Z(mul_ex_N346) );
  XOR2_X2 mul_ex_add_0_root_add_0_root_add_98_2_U16 ( .A(mul_ex_Z_14_), .B(
        mul_ex_add_0_root_add_0_root_add_98_2_carry_49_), .Z(mul_ex_N363) );
  AND2_X4 mul_ex_add_0_root_add_0_root_add_98_2_U15 ( .A1(mul_ex_Z_1_), .A2(
        mul_ex_add_0_root_add_0_root_add_98_2_n7), .ZN(
        mul_ex_add_0_root_add_0_root_add_98_2_n15) );
  AND2_X4 mul_ex_add_0_root_add_0_root_add_98_2_U14 ( .A1(mul_ex_N282), .A2(
        mul_ex_Z_31_), .ZN(mul_ex_add_0_root_add_0_root_add_98_2_n14) );
  AND2_X4 mul_ex_add_0_root_add_0_root_add_98_2_U13 ( .A1(mul_ex_Z_14_), .A2(
        mul_ex_add_0_root_add_0_root_add_98_2_carry_49_), .ZN(
        mul_ex_add_0_root_add_0_root_add_98_2_n13) );
  AND2_X4 mul_ex_add_0_root_add_0_root_add_98_2_U12 ( .A1(mul_ex_Z_12_), .A2(
        mul_ex_add_0_root_add_0_root_add_98_2_n6), .ZN(
        mul_ex_add_0_root_add_0_root_add_98_2_n12) );
  AND2_X4 mul_ex_add_0_root_add_0_root_add_98_2_U11 ( .A1(mul_ex_Z_10_), .A2(
        mul_ex_add_0_root_add_0_root_add_98_2_n5), .ZN(
        mul_ex_add_0_root_add_0_root_add_98_2_n11) );
  AND2_X4 mul_ex_add_0_root_add_0_root_add_98_2_U10 ( .A1(mul_ex_Z_8_), .A2(
        mul_ex_add_0_root_add_0_root_add_98_2_n4), .ZN(
        mul_ex_add_0_root_add_0_root_add_98_2_n10) );
  AND2_X4 mul_ex_add_0_root_add_0_root_add_98_2_U9 ( .A1(mul_ex_Z_6_), .A2(
        mul_ex_add_0_root_add_0_root_add_98_2_n3), .ZN(
        mul_ex_add_0_root_add_0_root_add_98_2_n9) );
  AND2_X4 mul_ex_add_0_root_add_0_root_add_98_2_U8 ( .A1(mul_ex_Z_4_), .A2(
        mul_ex_add_0_root_add_0_root_add_98_2_n2), .ZN(
        mul_ex_add_0_root_add_0_root_add_98_2_n8) );
  AND2_X4 mul_ex_add_0_root_add_0_root_add_98_2_U7 ( .A1(mul_ex_Z_2_), .A2(
        mul_ex_add_0_root_add_0_root_add_98_2_n1), .ZN(
        mul_ex_add_0_root_add_0_root_add_98_2_n7) );
  AND2_X4 mul_ex_add_0_root_add_0_root_add_98_2_U6 ( .A1(mul_ex_Z_13_), .A2(
        mul_ex_add_0_root_add_0_root_add_98_2_n13), .ZN(
        mul_ex_add_0_root_add_0_root_add_98_2_n6) );
  AND2_X4 mul_ex_add_0_root_add_0_root_add_98_2_U5 ( .A1(mul_ex_Z_11_), .A2(
        mul_ex_add_0_root_add_0_root_add_98_2_n12), .ZN(
        mul_ex_add_0_root_add_0_root_add_98_2_n5) );
  AND2_X4 mul_ex_add_0_root_add_0_root_add_98_2_U4 ( .A1(mul_ex_Z_9_), .A2(
        mul_ex_add_0_root_add_0_root_add_98_2_n11), .ZN(
        mul_ex_add_0_root_add_0_root_add_98_2_n4) );
  AND2_X4 mul_ex_add_0_root_add_0_root_add_98_2_U3 ( .A1(mul_ex_Z_7_), .A2(
        mul_ex_add_0_root_add_0_root_add_98_2_n10), .ZN(
        mul_ex_add_0_root_add_0_root_add_98_2_n3) );
  AND2_X4 mul_ex_add_0_root_add_0_root_add_98_2_U2 ( .A1(mul_ex_Z_5_), .A2(
        mul_ex_add_0_root_add_0_root_add_98_2_n9), .ZN(
        mul_ex_add_0_root_add_0_root_add_98_2_n2) );
  AND2_X4 mul_ex_add_0_root_add_0_root_add_98_2_U1 ( .A1(mul_ex_Z_3_), .A2(
        mul_ex_add_0_root_add_0_root_add_98_2_n8), .ZN(
        mul_ex_add_0_root_add_0_root_add_98_2_n1) );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_33 ( .A(mul_ex_Z_30_), .B(
        mul_ex_N283), .CI(mul_ex_add_0_root_add_0_root_add_98_2_n14), .CO(
        mul_ex_add_0_root_add_0_root_add_98_2_carry_34_), .S(mul_ex_N347) );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_34 ( .A(mul_ex_Z_29_), .B(
        mul_ex_N284), .CI(mul_ex_add_0_root_add_0_root_add_98_2_carry_34_), 
        .CO(mul_ex_add_0_root_add_0_root_add_98_2_carry_35_), .S(mul_ex_N348)
         );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_35 ( .A(mul_ex_Z_28_), .B(
        mul_ex_N285), .CI(mul_ex_add_0_root_add_0_root_add_98_2_carry_35_), 
        .CO(mul_ex_add_0_root_add_0_root_add_98_2_carry_36_), .S(mul_ex_N349)
         );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_36 ( .A(mul_ex_Z_27_), .B(
        mul_ex_N286), .CI(mul_ex_add_0_root_add_0_root_add_98_2_carry_36_), 
        .CO(mul_ex_add_0_root_add_0_root_add_98_2_carry_37_), .S(mul_ex_N350)
         );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_37 ( .A(mul_ex_Z_26_), .B(
        mul_ex_N287), .CI(mul_ex_add_0_root_add_0_root_add_98_2_carry_37_), 
        .CO(mul_ex_add_0_root_add_0_root_add_98_2_carry_38_), .S(mul_ex_N351)
         );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_38 ( .A(mul_ex_Z_25_), .B(
        mul_ex_N288), .CI(mul_ex_add_0_root_add_0_root_add_98_2_carry_38_), 
        .CO(mul_ex_add_0_root_add_0_root_add_98_2_carry_39_), .S(mul_ex_N352)
         );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_39 ( .A(mul_ex_Z_24_), .B(
        mul_ex_N289), .CI(mul_ex_add_0_root_add_0_root_add_98_2_carry_39_), 
        .CO(mul_ex_add_0_root_add_0_root_add_98_2_carry_40_), .S(mul_ex_N353)
         );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_40 ( .A(mul_ex_Z_23_), .B(
        mul_ex_N290), .CI(mul_ex_add_0_root_add_0_root_add_98_2_carry_40_), 
        .CO(mul_ex_add_0_root_add_0_root_add_98_2_carry_41_), .S(mul_ex_N354)
         );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_41 ( .A(mul_ex_Z_22_), .B(
        mul_ex_N291), .CI(mul_ex_add_0_root_add_0_root_add_98_2_carry_41_), 
        .CO(mul_ex_add_0_root_add_0_root_add_98_2_carry_42_), .S(mul_ex_N355)
         );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_42 ( .A(mul_ex_Z_21_), .B(
        mul_ex_N292), .CI(mul_ex_add_0_root_add_0_root_add_98_2_carry_42_), 
        .CO(mul_ex_add_0_root_add_0_root_add_98_2_carry_43_), .S(mul_ex_N356)
         );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_43 ( .A(mul_ex_Z_20_), .B(
        mul_ex_N293), .CI(mul_ex_add_0_root_add_0_root_add_98_2_carry_43_), 
        .CO(mul_ex_add_0_root_add_0_root_add_98_2_carry_44_), .S(mul_ex_N357)
         );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_44 ( .A(mul_ex_Z_19_), .B(
        mul_ex_N294), .CI(mul_ex_add_0_root_add_0_root_add_98_2_carry_44_), 
        .CO(mul_ex_add_0_root_add_0_root_add_98_2_carry_45_), .S(mul_ex_N358)
         );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_45 ( .A(mul_ex_Z_18_), .B(
        mul_ex_N295), .CI(mul_ex_add_0_root_add_0_root_add_98_2_carry_45_), 
        .CO(mul_ex_add_0_root_add_0_root_add_98_2_carry_46_), .S(mul_ex_N359)
         );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_46 ( .A(mul_ex_Z_17_), .B(
        mul_ex_N296), .CI(mul_ex_add_0_root_add_0_root_add_98_2_carry_46_), 
        .CO(mul_ex_add_0_root_add_0_root_add_98_2_carry_47_), .S(mul_ex_N360)
         );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_47 ( .A(mul_ex_Z_16_), .B(
        mul_ex_N297), .CI(mul_ex_add_0_root_add_0_root_add_98_2_carry_47_), 
        .CO(mul_ex_add_0_root_add_0_root_add_98_2_carry_48_), .S(mul_ex_N361)
         );
  FA_X1 mul_ex_add_0_root_add_0_root_add_98_2_U1_48 ( .A(mul_ex_Z_15_), .B(
        mul_ex_N298), .CI(mul_ex_add_0_root_add_0_root_add_98_2_carry_48_), 
        .CO(mul_ex_add_0_root_add_0_root_add_98_2_carry_49_), .S(mul_ex_N362)
         );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U35 ( .A(mul_ex_L_31_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n33) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U34 ( .A(mul_ex_L_30_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n32) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U33 ( .A(mul_ex_L_29_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n31) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U32 ( .A(mul_ex_L_28_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n30) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U31 ( .A(mul_ex_L_27_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n29) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U30 ( .A(mul_ex_L_26_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n28) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U29 ( .A(mul_ex_L_25_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n27) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U28 ( .A(mul_ex_L_24_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n26) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U27 ( .A(mul_ex_L_23_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n25) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U26 ( .A(mul_ex_L_22_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n24) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U25 ( .A(mul_ex_L_21_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n23) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U24 ( .A(mul_ex_L_20_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n22) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U23 ( .A(mul_ex_L_19_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n21) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U22 ( .A(mul_ex_L_18_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n20) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U21 ( .A(mul_ex_L_17_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n19) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U20 ( .A(mul_ex_L_16_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n18) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U19 ( .A(mul_ex_L_15_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n17) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U18 ( .A(mul_ex_L_14_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n16) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U17 ( .A(mul_ex_L_13_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n15) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U16 ( .A(mul_ex_L_12_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n14) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U15 ( .A(mul_ex_L_11_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n13) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U14 ( .A(mul_ex_L_10_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n12) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U13 ( .A(mul_ex_L_9_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n11) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U12 ( .A(mul_ex_L_8_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n10) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U11 ( .A(mul_ex_L_7_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n9) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U10 ( .A(mul_ex_L_6_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n8) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U9 ( .A(mul_ex_L_5_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n7) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U8 ( .A(mul_ex_L_4_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n6) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U7 ( .A(mul_ex_L_3_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n5) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U6 ( .A(mul_ex_L_2_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n4) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U5 ( .A(mul_ex_L_1_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n3) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U4 ( .A(mul_ex_L_0_), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n2) );
  INV_X4 mul_ex_sub_1_root_sub_0_root_sub_94_2_U3 ( .A(mul_ex_P[31]), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n1) );
  XNOR2_X2 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2 ( .A(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n33), .B(mul_ex_P[31]), .ZN(
        mul_ex_N186) );
  NAND2_X2 mul_ex_sub_1_root_sub_0_root_sub_94_2_U1 ( .A1(mul_ex_L_31_), .A2(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n1), .ZN(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[1]) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_1 ( .A(mul_ex_P[30]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n32), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[1]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[2]), .S(mul_ex_N187) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_2 ( .A(mul_ex_P[29]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n31), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[2]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[3]), .S(mul_ex_N188) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_3 ( .A(mul_ex_P[28]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n30), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[3]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[4]), .S(mul_ex_N189) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_4 ( .A(mul_ex_P[27]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n29), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[4]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[5]), .S(mul_ex_N190) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_5 ( .A(mul_ex_P[26]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n28), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[5]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[6]), .S(mul_ex_N191) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_6 ( .A(mul_ex_P[25]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n27), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[6]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[7]), .S(mul_ex_N192) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_7 ( .A(mul_ex_P[24]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n26), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[7]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[8]), .S(mul_ex_N193) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_8 ( .A(mul_ex_P[23]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n25), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[8]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[9]), .S(mul_ex_N194) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_9 ( .A(mul_ex_P[22]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n24), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[9]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[10]), .S(mul_ex_N195) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_10 ( .A(mul_ex_P[21]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n23), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[10]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[11]), .S(mul_ex_N196) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_11 ( .A(mul_ex_P[20]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n22), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[11]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[12]), .S(mul_ex_N197) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_12 ( .A(mul_ex_P[19]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n21), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[12]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[13]), .S(mul_ex_N198) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_13 ( .A(mul_ex_P[18]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n20), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[13]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[14]), .S(mul_ex_N199) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_14 ( .A(mul_ex_P[17]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n19), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[14]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[15]), .S(mul_ex_N200) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_15 ( .A(mul_ex_P[16]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n18), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[15]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[16]), .S(mul_ex_N201) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_16 ( .A(mul_ex_P[15]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n17), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[16]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[17]), .S(mul_ex_N202) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_17 ( .A(mul_ex_P[14]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n16), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[17]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[18]), .S(mul_ex_N203) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_18 ( .A(mul_ex_P[13]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n15), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[18]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[19]), .S(mul_ex_N204) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_19 ( .A(mul_ex_P[12]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n14), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[19]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[20]), .S(mul_ex_N205) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_20 ( .A(mul_ex_P[11]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n13), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[20]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[21]), .S(mul_ex_N206) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_21 ( .A(mul_ex_P[10]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n12), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[21]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[22]), .S(mul_ex_N207) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_22 ( .A(mul_ex_P[9]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n11), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[22]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[23]), .S(mul_ex_N208) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_23 ( .A(mul_ex_P[8]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n10), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[23]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[24]), .S(mul_ex_N209) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_24 ( .A(mul_ex_P[7]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n9), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[24]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[25]), .S(mul_ex_N210) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_25 ( .A(mul_ex_P[6]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n8), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[25]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[26]), .S(mul_ex_N211) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_26 ( .A(mul_ex_P[5]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n7), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[26]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[27]), .S(mul_ex_N212) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_27 ( .A(mul_ex_P[4]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n6), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[27]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[28]), .S(mul_ex_N213) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_28 ( .A(mul_ex_P[3]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n5), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[28]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[29]), .S(mul_ex_N214) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_29 ( .A(mul_ex_P[2]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n4), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[29]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[30]), .S(mul_ex_N215) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_30 ( .A(mul_ex_P[1]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n3), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[30]), .CO(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[31]), .S(mul_ex_N216) );
  FA_X1 mul_ex_sub_1_root_sub_0_root_sub_94_2_U2_31 ( .A(mul_ex_P[0]), .B(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_n2), .CI(
        mul_ex_sub_1_root_sub_0_root_sub_94_2_carry[31]), .S(mul_ex_N217) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U35 ( .A(mul_ex_H[31]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n33) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U34 ( .A(mul_ex_H[30]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n32) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U33 ( .A(mul_ex_H[29]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n31) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U32 ( .A(mul_ex_H[28]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n30) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U31 ( .A(mul_ex_H[27]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n29) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U30 ( .A(mul_ex_H[26]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n28) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U29 ( .A(mul_ex_H[25]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n27) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U28 ( .A(mul_ex_H[24]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n26) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U27 ( .A(mul_ex_H[23]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n25) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U26 ( .A(mul_ex_H[22]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n24) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U25 ( .A(mul_ex_H[21]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n23) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U24 ( .A(mul_ex_H[20]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n22) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U23 ( .A(mul_ex_H[19]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n21) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U22 ( .A(mul_ex_H[18]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n20) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U21 ( .A(mul_ex_H[17]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n19) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U20 ( .A(mul_ex_H[16]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n18) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U19 ( .A(mul_ex_H[15]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n17) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U18 ( .A(mul_ex_H[14]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n16) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U17 ( .A(mul_ex_H[13]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n15) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U16 ( .A(mul_ex_H[12]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n14) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U15 ( .A(mul_ex_H[11]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n13) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U14 ( .A(mul_ex_H[10]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n12) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U13 ( .A(mul_ex_H[9]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n11) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U12 ( .A(mul_ex_H[8]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n10) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U11 ( .A(mul_ex_H[7]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n9) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U10 ( .A(mul_ex_H[6]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n8) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U9 ( .A(mul_ex_H[5]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n7) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U8 ( .A(mul_ex_H[4]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n6) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U7 ( .A(mul_ex_H[3]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n5) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U6 ( .A(mul_ex_H[2]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n4) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U5 ( .A(mul_ex_H[1]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n3) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U4 ( .A(mul_ex_H[0]), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n2) );
  INV_X4 mul_ex_sub_0_root_sub_0_root_sub_94_2_U3 ( .A(mul_ex_N186), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n1) );
  XNOR2_X2 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2 ( .A(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n33), .B(mul_ex_N186), .ZN(
        mul_ex_N218) );
  NAND2_X2 mul_ex_sub_0_root_sub_0_root_sub_94_2_U1 ( .A1(mul_ex_H[31]), .A2(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n1), .ZN(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[1]) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_1 ( .A(mul_ex_N187), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n32), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[1]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[2]), .S(mul_ex_N219) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_2 ( .A(mul_ex_N188), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n31), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[2]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[3]), .S(mul_ex_N220) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_3 ( .A(mul_ex_N189), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n30), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[3]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[4]), .S(mul_ex_N221) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_4 ( .A(mul_ex_N190), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n29), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[4]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[5]), .S(mul_ex_N222) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_5 ( .A(mul_ex_N191), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n28), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[5]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[6]), .S(mul_ex_N223) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_6 ( .A(mul_ex_N192), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n27), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[6]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[7]), .S(mul_ex_N224) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_7 ( .A(mul_ex_N193), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n26), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[7]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[8]), .S(mul_ex_N225) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_8 ( .A(mul_ex_N194), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n25), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[8]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[9]), .S(mul_ex_N226) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_9 ( .A(mul_ex_N195), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n24), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[9]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[10]), .S(mul_ex_N227) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_10 ( .A(mul_ex_N196), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n23), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[10]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[11]), .S(mul_ex_N228) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_11 ( .A(mul_ex_N197), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n22), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[11]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[12]), .S(mul_ex_N229) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_12 ( .A(mul_ex_N198), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n21), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[12]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[13]), .S(mul_ex_N230) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_13 ( .A(mul_ex_N199), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n20), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[13]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[14]), .S(mul_ex_N231) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_14 ( .A(mul_ex_N200), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n19), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[14]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[15]), .S(mul_ex_N232) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_15 ( .A(mul_ex_N201), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n18), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[15]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[16]), .S(mul_ex_N233) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_16 ( .A(mul_ex_N202), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n17), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[16]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[17]), .S(mul_ex_N234) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_17 ( .A(mul_ex_N203), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n16), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[17]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[18]), .S(mul_ex_N235) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_18 ( .A(mul_ex_N204), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n15), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[18]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[19]), .S(mul_ex_N236) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_19 ( .A(mul_ex_N205), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n14), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[19]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[20]), .S(mul_ex_N237) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_20 ( .A(mul_ex_N206), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n13), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[20]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[21]), .S(mul_ex_N238) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_21 ( .A(mul_ex_N207), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n12), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[21]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[22]), .S(mul_ex_N239) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_22 ( .A(mul_ex_N208), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n11), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[22]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[23]), .S(mul_ex_N240) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_23 ( .A(mul_ex_N209), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n10), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[23]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[24]), .S(mul_ex_N241) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_24 ( .A(mul_ex_N210), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n9), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[24]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[25]), .S(mul_ex_N242) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_25 ( .A(mul_ex_N211), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n8), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[25]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[26]), .S(mul_ex_N243) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_26 ( .A(mul_ex_N212), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n7), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[26]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[27]), .S(mul_ex_N244) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_27 ( .A(mul_ex_N213), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n6), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[27]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[28]), .S(mul_ex_N245) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_28 ( .A(mul_ex_N214), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n5), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[28]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[29]), .S(mul_ex_N246) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_29 ( .A(mul_ex_N215), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n4), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[29]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[30]), .S(mul_ex_N247) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_30 ( .A(mul_ex_N216), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n3), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[30]), .CO(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[31]), .S(mul_ex_N248) );
  FA_X1 mul_ex_sub_0_root_sub_0_root_sub_94_2_U2_31 ( .A(mul_ex_N217), .B(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_n2), .CI(
        mul_ex_sub_0_root_sub_0_root_sub_94_2_carry[31]), .S(mul_ex_N249) );
  INV_X4 mul_ex_mult_90_U811 ( .A(mul_ex_mult_90_n299), .ZN(
        mul_ex_mult_90_SUMB_21__9_) );
  XNOR2_X2 mul_ex_mult_90_U810 ( .A(mul_ex_mult_90_CARRYB_20__9_), .B(
        mul_ex_mult_90_SUMB_20__10_), .ZN(mul_ex_mult_90_n299) );
  INV_X4 mul_ex_mult_90_U809 ( .A(mul_ex_mult_90_n298), .ZN(
        mul_ex_mult_90_CARRYB_21__9_) );
  NAND2_X2 mul_ex_mult_90_U808 ( .A1(mul_ex_mult_90_SUMB_20__10_), .A2(
        mul_ex_mult_90_CARRYB_20__9_), .ZN(mul_ex_mult_90_n298) );
  INV_X4 mul_ex_mult_90_U807 ( .A(mul_ex_mult_90_n297), .ZN(mul_ex_N175) );
  XNOR2_X2 mul_ex_mult_90_U806 ( .A(mul_ex_mult_90_CARRYB_20__0_), .B(
        mul_ex_mult_90_SUMB_20__1_), .ZN(mul_ex_mult_90_n297) );
  INV_X4 mul_ex_mult_90_U805 ( .A(mul_ex_mult_90_n296), .ZN(
        mul_ex_mult_90_CARRYB_21__0_) );
  NAND2_X2 mul_ex_mult_90_U804 ( .A1(mul_ex_mult_90_SUMB_20__1_), .A2(
        mul_ex_mult_90_CARRYB_20__0_), .ZN(mul_ex_mult_90_n296) );
  INV_X4 mul_ex_mult_90_U803 ( .A(mul_ex_mult_90_n295), .ZN(
        mul_ex_mult_90_SUMB_21__1_) );
  XNOR2_X2 mul_ex_mult_90_U802 ( .A(mul_ex_mult_90_CARRYB_20__1_), .B(
        mul_ex_mult_90_SUMB_20__2_), .ZN(mul_ex_mult_90_n295) );
  INV_X4 mul_ex_mult_90_U801 ( .A(mul_ex_mult_90_n294), .ZN(
        mul_ex_mult_90_CARRYB_21__1_) );
  NAND2_X2 mul_ex_mult_90_U800 ( .A1(mul_ex_mult_90_SUMB_20__2_), .A2(
        mul_ex_mult_90_CARRYB_20__1_), .ZN(mul_ex_mult_90_n294) );
  INV_X4 mul_ex_mult_90_U799 ( .A(mul_ex_mult_90_n293), .ZN(
        mul_ex_mult_90_SUMB_21__2_) );
  XNOR2_X2 mul_ex_mult_90_U798 ( .A(mul_ex_mult_90_CARRYB_20__2_), .B(
        mul_ex_mult_90_SUMB_20__3_), .ZN(mul_ex_mult_90_n293) );
  INV_X4 mul_ex_mult_90_U797 ( .A(mul_ex_mult_90_n292), .ZN(
        mul_ex_mult_90_CARRYB_21__2_) );
  NAND2_X2 mul_ex_mult_90_U796 ( .A1(mul_ex_mult_90_SUMB_20__3_), .A2(
        mul_ex_mult_90_CARRYB_20__2_), .ZN(mul_ex_mult_90_n292) );
  INV_X4 mul_ex_mult_90_U795 ( .A(mul_ex_mult_90_n291), .ZN(
        mul_ex_mult_90_SUMB_21__3_) );
  XNOR2_X2 mul_ex_mult_90_U794 ( .A(mul_ex_mult_90_CARRYB_20__3_), .B(
        mul_ex_mult_90_SUMB_20__4_), .ZN(mul_ex_mult_90_n291) );
  INV_X4 mul_ex_mult_90_U793 ( .A(mul_ex_mult_90_n290), .ZN(
        mul_ex_mult_90_CARRYB_21__3_) );
  NAND2_X2 mul_ex_mult_90_U792 ( .A1(mul_ex_mult_90_SUMB_20__4_), .A2(
        mul_ex_mult_90_CARRYB_20__3_), .ZN(mul_ex_mult_90_n290) );
  INV_X4 mul_ex_mult_90_U791 ( .A(mul_ex_mult_90_n289), .ZN(
        mul_ex_mult_90_SUMB_21__4_) );
  XNOR2_X2 mul_ex_mult_90_U790 ( .A(mul_ex_mult_90_CARRYB_20__4_), .B(
        mul_ex_mult_90_SUMB_20__5_), .ZN(mul_ex_mult_90_n289) );
  INV_X4 mul_ex_mult_90_U789 ( .A(mul_ex_mult_90_n288), .ZN(
        mul_ex_mult_90_CARRYB_21__4_) );
  NAND2_X2 mul_ex_mult_90_U788 ( .A1(mul_ex_mult_90_SUMB_20__5_), .A2(
        mul_ex_mult_90_CARRYB_20__4_), .ZN(mul_ex_mult_90_n288) );
  INV_X4 mul_ex_mult_90_U787 ( .A(mul_ex_mult_90_n287), .ZN(
        mul_ex_mult_90_SUMB_21__5_) );
  XNOR2_X2 mul_ex_mult_90_U786 ( .A(mul_ex_mult_90_CARRYB_20__5_), .B(
        mul_ex_mult_90_SUMB_20__6_), .ZN(mul_ex_mult_90_n287) );
  INV_X4 mul_ex_mult_90_U785 ( .A(mul_ex_mult_90_n286), .ZN(
        mul_ex_mult_90_CARRYB_21__5_) );
  NAND2_X2 mul_ex_mult_90_U784 ( .A1(mul_ex_mult_90_SUMB_20__6_), .A2(
        mul_ex_mult_90_CARRYB_20__5_), .ZN(mul_ex_mult_90_n286) );
  INV_X4 mul_ex_mult_90_U783 ( .A(mul_ex_mult_90_n285), .ZN(
        mul_ex_mult_90_SUMB_21__6_) );
  XNOR2_X2 mul_ex_mult_90_U782 ( .A(mul_ex_mult_90_CARRYB_20__6_), .B(
        mul_ex_mult_90_SUMB_20__7_), .ZN(mul_ex_mult_90_n285) );
  INV_X4 mul_ex_mult_90_U781 ( .A(mul_ex_mult_90_n284), .ZN(
        mul_ex_mult_90_CARRYB_21__6_) );
  NAND2_X2 mul_ex_mult_90_U780 ( .A1(mul_ex_mult_90_SUMB_20__7_), .A2(
        mul_ex_mult_90_CARRYB_20__6_), .ZN(mul_ex_mult_90_n284) );
  INV_X4 mul_ex_mult_90_U779 ( .A(mul_ex_mult_90_n283), .ZN(
        mul_ex_mult_90_SUMB_21__7_) );
  XNOR2_X2 mul_ex_mult_90_U778 ( .A(mul_ex_mult_90_CARRYB_20__7_), .B(
        mul_ex_mult_90_SUMB_20__8_), .ZN(mul_ex_mult_90_n283) );
  INV_X4 mul_ex_mult_90_U777 ( .A(mul_ex_mult_90_n282), .ZN(
        mul_ex_mult_90_CARRYB_21__7_) );
  NAND2_X2 mul_ex_mult_90_U776 ( .A1(mul_ex_mult_90_SUMB_20__8_), .A2(
        mul_ex_mult_90_CARRYB_20__7_), .ZN(mul_ex_mult_90_n282) );
  INV_X4 mul_ex_mult_90_U775 ( .A(mul_ex_mult_90_n281), .ZN(
        mul_ex_mult_90_SUMB_21__8_) );
  XNOR2_X2 mul_ex_mult_90_U774 ( .A(mul_ex_mult_90_CARRYB_20__8_), .B(
        mul_ex_mult_90_SUMB_20__9_), .ZN(mul_ex_mult_90_n281) );
  INV_X4 mul_ex_mult_90_U773 ( .A(mul_ex_mult_90_n280), .ZN(
        mul_ex_mult_90_CARRYB_21__8_) );
  NAND2_X2 mul_ex_mult_90_U772 ( .A1(mul_ex_mult_90_SUMB_20__9_), .A2(
        mul_ex_mult_90_CARRYB_20__8_), .ZN(mul_ex_mult_90_n280) );
  INV_X4 mul_ex_mult_90_U771 ( .A(mul_ex_mult_90_n279), .ZN(
        mul_ex_mult_90_SUMB_20__9_) );
  XNOR2_X2 mul_ex_mult_90_U770 ( .A(mul_ex_mult_90_CARRYB_19__9_), .B(
        mul_ex_mult_90_SUMB_19__10_), .ZN(mul_ex_mult_90_n279) );
  INV_X4 mul_ex_mult_90_U769 ( .A(mul_ex_mult_90_n278), .ZN(
        mul_ex_mult_90_CARRYB_20__9_) );
  NAND2_X2 mul_ex_mult_90_U768 ( .A1(mul_ex_mult_90_SUMB_19__10_), .A2(
        mul_ex_mult_90_CARRYB_19__9_), .ZN(mul_ex_mult_90_n278) );
  INV_X4 mul_ex_mult_90_U767 ( .A(mul_ex_mult_90_n277), .ZN(mul_ex_N174) );
  XNOR2_X2 mul_ex_mult_90_U766 ( .A(mul_ex_mult_90_CARRYB_19__0_), .B(
        mul_ex_mult_90_SUMB_19__1_), .ZN(mul_ex_mult_90_n277) );
  INV_X4 mul_ex_mult_90_U765 ( .A(mul_ex_mult_90_n276), .ZN(
        mul_ex_mult_90_CARRYB_20__0_) );
  NAND2_X2 mul_ex_mult_90_U764 ( .A1(mul_ex_mult_90_SUMB_19__1_), .A2(
        mul_ex_mult_90_CARRYB_19__0_), .ZN(mul_ex_mult_90_n276) );
  INV_X4 mul_ex_mult_90_U763 ( .A(mul_ex_mult_90_n275), .ZN(
        mul_ex_mult_90_SUMB_20__10_) );
  XNOR2_X2 mul_ex_mult_90_U762 ( .A(mul_ex_mult_90_CARRYB_19__10_), .B(
        mul_ex_mult_90_SUMB_19__11_), .ZN(mul_ex_mult_90_n275) );
  INV_X4 mul_ex_mult_90_U761 ( .A(mul_ex_mult_90_n274), .ZN(
        mul_ex_mult_90_CARRYB_20__10_) );
  NAND2_X2 mul_ex_mult_90_U760 ( .A1(mul_ex_mult_90_SUMB_19__11_), .A2(
        mul_ex_mult_90_CARRYB_19__10_), .ZN(mul_ex_mult_90_n274) );
  INV_X4 mul_ex_mult_90_U759 ( .A(mul_ex_mult_90_n273), .ZN(
        mul_ex_mult_90_SUMB_20__1_) );
  XNOR2_X2 mul_ex_mult_90_U758 ( .A(mul_ex_mult_90_CARRYB_19__1_), .B(
        mul_ex_mult_90_SUMB_19__2_), .ZN(mul_ex_mult_90_n273) );
  INV_X4 mul_ex_mult_90_U757 ( .A(mul_ex_mult_90_n272), .ZN(
        mul_ex_mult_90_CARRYB_20__1_) );
  NAND2_X2 mul_ex_mult_90_U756 ( .A1(mul_ex_mult_90_SUMB_19__2_), .A2(
        mul_ex_mult_90_CARRYB_19__1_), .ZN(mul_ex_mult_90_n272) );
  INV_X4 mul_ex_mult_90_U755 ( .A(mul_ex_mult_90_n271), .ZN(
        mul_ex_mult_90_SUMB_20__2_) );
  XNOR2_X2 mul_ex_mult_90_U754 ( .A(mul_ex_mult_90_CARRYB_19__2_), .B(
        mul_ex_mult_90_SUMB_19__3_), .ZN(mul_ex_mult_90_n271) );
  INV_X4 mul_ex_mult_90_U753 ( .A(mul_ex_mult_90_n270), .ZN(
        mul_ex_mult_90_CARRYB_20__2_) );
  NAND2_X2 mul_ex_mult_90_U752 ( .A1(mul_ex_mult_90_SUMB_19__3_), .A2(
        mul_ex_mult_90_CARRYB_19__2_), .ZN(mul_ex_mult_90_n270) );
  INV_X4 mul_ex_mult_90_U751 ( .A(mul_ex_mult_90_n269), .ZN(
        mul_ex_mult_90_SUMB_20__3_) );
  XNOR2_X2 mul_ex_mult_90_U750 ( .A(mul_ex_mult_90_CARRYB_19__3_), .B(
        mul_ex_mult_90_SUMB_19__4_), .ZN(mul_ex_mult_90_n269) );
  INV_X4 mul_ex_mult_90_U749 ( .A(mul_ex_mult_90_n268), .ZN(
        mul_ex_mult_90_CARRYB_20__3_) );
  NAND2_X2 mul_ex_mult_90_U748 ( .A1(mul_ex_mult_90_SUMB_19__4_), .A2(
        mul_ex_mult_90_CARRYB_19__3_), .ZN(mul_ex_mult_90_n268) );
  INV_X4 mul_ex_mult_90_U747 ( .A(mul_ex_mult_90_n267), .ZN(
        mul_ex_mult_90_SUMB_20__4_) );
  XNOR2_X2 mul_ex_mult_90_U746 ( .A(mul_ex_mult_90_CARRYB_19__4_), .B(
        mul_ex_mult_90_SUMB_19__5_), .ZN(mul_ex_mult_90_n267) );
  INV_X4 mul_ex_mult_90_U745 ( .A(mul_ex_mult_90_n266), .ZN(
        mul_ex_mult_90_CARRYB_20__4_) );
  NAND2_X2 mul_ex_mult_90_U744 ( .A1(mul_ex_mult_90_SUMB_19__5_), .A2(
        mul_ex_mult_90_CARRYB_19__4_), .ZN(mul_ex_mult_90_n266) );
  INV_X4 mul_ex_mult_90_U743 ( .A(mul_ex_mult_90_n265), .ZN(
        mul_ex_mult_90_SUMB_20__5_) );
  XNOR2_X2 mul_ex_mult_90_U742 ( .A(mul_ex_mult_90_CARRYB_19__5_), .B(
        mul_ex_mult_90_SUMB_19__6_), .ZN(mul_ex_mult_90_n265) );
  INV_X4 mul_ex_mult_90_U741 ( .A(mul_ex_mult_90_n264), .ZN(
        mul_ex_mult_90_CARRYB_20__5_) );
  NAND2_X2 mul_ex_mult_90_U740 ( .A1(mul_ex_mult_90_SUMB_19__6_), .A2(
        mul_ex_mult_90_CARRYB_19__5_), .ZN(mul_ex_mult_90_n264) );
  INV_X4 mul_ex_mult_90_U739 ( .A(mul_ex_mult_90_n263), .ZN(
        mul_ex_mult_90_SUMB_20__6_) );
  XNOR2_X2 mul_ex_mult_90_U738 ( .A(mul_ex_mult_90_CARRYB_19__6_), .B(
        mul_ex_mult_90_SUMB_19__7_), .ZN(mul_ex_mult_90_n263) );
  INV_X4 mul_ex_mult_90_U737 ( .A(mul_ex_mult_90_n262), .ZN(
        mul_ex_mult_90_CARRYB_20__6_) );
  NAND2_X2 mul_ex_mult_90_U736 ( .A1(mul_ex_mult_90_SUMB_19__7_), .A2(
        mul_ex_mult_90_CARRYB_19__6_), .ZN(mul_ex_mult_90_n262) );
  INV_X4 mul_ex_mult_90_U735 ( .A(mul_ex_mult_90_n261), .ZN(
        mul_ex_mult_90_SUMB_20__7_) );
  XNOR2_X2 mul_ex_mult_90_U734 ( .A(mul_ex_mult_90_CARRYB_19__7_), .B(
        mul_ex_mult_90_SUMB_19__8_), .ZN(mul_ex_mult_90_n261) );
  INV_X4 mul_ex_mult_90_U733 ( .A(mul_ex_mult_90_n260), .ZN(
        mul_ex_mult_90_CARRYB_20__7_) );
  NAND2_X2 mul_ex_mult_90_U732 ( .A1(mul_ex_mult_90_SUMB_19__8_), .A2(
        mul_ex_mult_90_CARRYB_19__7_), .ZN(mul_ex_mult_90_n260) );
  INV_X4 mul_ex_mult_90_U731 ( .A(mul_ex_mult_90_n259), .ZN(
        mul_ex_mult_90_SUMB_20__8_) );
  XNOR2_X2 mul_ex_mult_90_U730 ( .A(mul_ex_mult_90_CARRYB_19__8_), .B(
        mul_ex_mult_90_SUMB_19__9_), .ZN(mul_ex_mult_90_n259) );
  INV_X4 mul_ex_mult_90_U729 ( .A(mul_ex_mult_90_n258), .ZN(
        mul_ex_mult_90_CARRYB_20__8_) );
  NAND2_X2 mul_ex_mult_90_U728 ( .A1(mul_ex_mult_90_SUMB_19__9_), .A2(
        mul_ex_mult_90_CARRYB_19__8_), .ZN(mul_ex_mult_90_n258) );
  INV_X4 mul_ex_mult_90_U727 ( .A(mul_ex_mult_90_n257), .ZN(
        mul_ex_mult_90_SUMB_19__9_) );
  XNOR2_X2 mul_ex_mult_90_U726 ( .A(mul_ex_mult_90_CARRYB_18__9_), .B(
        mul_ex_mult_90_SUMB_18__10_), .ZN(mul_ex_mult_90_n257) );
  INV_X4 mul_ex_mult_90_U725 ( .A(mul_ex_mult_90_n256), .ZN(
        mul_ex_mult_90_CARRYB_19__9_) );
  NAND2_X2 mul_ex_mult_90_U724 ( .A1(mul_ex_mult_90_SUMB_18__10_), .A2(
        mul_ex_mult_90_CARRYB_18__9_), .ZN(mul_ex_mult_90_n256) );
  INV_X4 mul_ex_mult_90_U723 ( .A(mul_ex_mult_90_n255), .ZN(mul_ex_N173) );
  XNOR2_X2 mul_ex_mult_90_U722 ( .A(mul_ex_mult_90_CARRYB_18__0_), .B(
        mul_ex_mult_90_SUMB_18__1_), .ZN(mul_ex_mult_90_n255) );
  INV_X4 mul_ex_mult_90_U721 ( .A(mul_ex_mult_90_n254), .ZN(
        mul_ex_mult_90_CARRYB_19__0_) );
  NAND2_X2 mul_ex_mult_90_U720 ( .A1(mul_ex_mult_90_SUMB_18__1_), .A2(
        mul_ex_mult_90_CARRYB_18__0_), .ZN(mul_ex_mult_90_n254) );
  INV_X4 mul_ex_mult_90_U719 ( .A(mul_ex_mult_90_n253), .ZN(
        mul_ex_mult_90_SUMB_19__10_) );
  XNOR2_X2 mul_ex_mult_90_U718 ( .A(mul_ex_mult_90_CARRYB_18__10_), .B(
        mul_ex_mult_90_SUMB_18__11_), .ZN(mul_ex_mult_90_n253) );
  INV_X4 mul_ex_mult_90_U717 ( .A(mul_ex_mult_90_n252), .ZN(
        mul_ex_mult_90_CARRYB_19__10_) );
  NAND2_X2 mul_ex_mult_90_U716 ( .A1(mul_ex_mult_90_SUMB_18__11_), .A2(
        mul_ex_mult_90_CARRYB_18__10_), .ZN(mul_ex_mult_90_n252) );
  INV_X4 mul_ex_mult_90_U715 ( .A(mul_ex_mult_90_n251), .ZN(
        mul_ex_mult_90_SUMB_19__11_) );
  XNOR2_X2 mul_ex_mult_90_U714 ( .A(mul_ex_mult_90_CARRYB_18__11_), .B(
        mul_ex_mult_90_SUMB_18__12_), .ZN(mul_ex_mult_90_n251) );
  INV_X4 mul_ex_mult_90_U713 ( .A(mul_ex_mult_90_n250), .ZN(
        mul_ex_mult_90_CARRYB_19__11_) );
  NAND2_X2 mul_ex_mult_90_U712 ( .A1(mul_ex_mult_90_SUMB_18__12_), .A2(
        mul_ex_mult_90_CARRYB_18__11_), .ZN(mul_ex_mult_90_n250) );
  INV_X4 mul_ex_mult_90_U711 ( .A(mul_ex_mult_90_n249), .ZN(
        mul_ex_mult_90_SUMB_19__1_) );
  XNOR2_X2 mul_ex_mult_90_U710 ( .A(mul_ex_mult_90_CARRYB_18__1_), .B(
        mul_ex_mult_90_SUMB_18__2_), .ZN(mul_ex_mult_90_n249) );
  INV_X4 mul_ex_mult_90_U709 ( .A(mul_ex_mult_90_n248), .ZN(
        mul_ex_mult_90_CARRYB_19__1_) );
  NAND2_X2 mul_ex_mult_90_U708 ( .A1(mul_ex_mult_90_SUMB_18__2_), .A2(
        mul_ex_mult_90_CARRYB_18__1_), .ZN(mul_ex_mult_90_n248) );
  INV_X4 mul_ex_mult_90_U707 ( .A(mul_ex_mult_90_n247), .ZN(
        mul_ex_mult_90_SUMB_19__2_) );
  XNOR2_X2 mul_ex_mult_90_U706 ( .A(mul_ex_mult_90_CARRYB_18__2_), .B(
        mul_ex_mult_90_SUMB_18__3_), .ZN(mul_ex_mult_90_n247) );
  INV_X4 mul_ex_mult_90_U705 ( .A(mul_ex_mult_90_n246), .ZN(
        mul_ex_mult_90_CARRYB_19__2_) );
  NAND2_X2 mul_ex_mult_90_U704 ( .A1(mul_ex_mult_90_SUMB_18__3_), .A2(
        mul_ex_mult_90_CARRYB_18__2_), .ZN(mul_ex_mult_90_n246) );
  INV_X4 mul_ex_mult_90_U703 ( .A(mul_ex_mult_90_n245), .ZN(
        mul_ex_mult_90_SUMB_19__3_) );
  XNOR2_X2 mul_ex_mult_90_U702 ( .A(mul_ex_mult_90_CARRYB_18__3_), .B(
        mul_ex_mult_90_SUMB_18__4_), .ZN(mul_ex_mult_90_n245) );
  INV_X4 mul_ex_mult_90_U701 ( .A(mul_ex_mult_90_n244), .ZN(
        mul_ex_mult_90_CARRYB_19__3_) );
  NAND2_X2 mul_ex_mult_90_U700 ( .A1(mul_ex_mult_90_SUMB_18__4_), .A2(
        mul_ex_mult_90_CARRYB_18__3_), .ZN(mul_ex_mult_90_n244) );
  INV_X4 mul_ex_mult_90_U699 ( .A(mul_ex_mult_90_n243), .ZN(
        mul_ex_mult_90_SUMB_19__4_) );
  XNOR2_X2 mul_ex_mult_90_U698 ( .A(mul_ex_mult_90_CARRYB_18__4_), .B(
        mul_ex_mult_90_SUMB_18__5_), .ZN(mul_ex_mult_90_n243) );
  INV_X4 mul_ex_mult_90_U697 ( .A(mul_ex_mult_90_n242), .ZN(
        mul_ex_mult_90_CARRYB_19__4_) );
  NAND2_X2 mul_ex_mult_90_U696 ( .A1(mul_ex_mult_90_SUMB_18__5_), .A2(
        mul_ex_mult_90_CARRYB_18__4_), .ZN(mul_ex_mult_90_n242) );
  INV_X4 mul_ex_mult_90_U695 ( .A(mul_ex_mult_90_n241), .ZN(
        mul_ex_mult_90_SUMB_19__5_) );
  XNOR2_X2 mul_ex_mult_90_U694 ( .A(mul_ex_mult_90_CARRYB_18__5_), .B(
        mul_ex_mult_90_SUMB_18__6_), .ZN(mul_ex_mult_90_n241) );
  INV_X4 mul_ex_mult_90_U693 ( .A(mul_ex_mult_90_n240), .ZN(
        mul_ex_mult_90_CARRYB_19__5_) );
  NAND2_X2 mul_ex_mult_90_U692 ( .A1(mul_ex_mult_90_SUMB_18__6_), .A2(
        mul_ex_mult_90_CARRYB_18__5_), .ZN(mul_ex_mult_90_n240) );
  INV_X4 mul_ex_mult_90_U691 ( .A(mul_ex_mult_90_n239), .ZN(
        mul_ex_mult_90_SUMB_19__6_) );
  XNOR2_X2 mul_ex_mult_90_U690 ( .A(mul_ex_mult_90_CARRYB_18__6_), .B(
        mul_ex_mult_90_SUMB_18__7_), .ZN(mul_ex_mult_90_n239) );
  INV_X4 mul_ex_mult_90_U689 ( .A(mul_ex_mult_90_n238), .ZN(
        mul_ex_mult_90_CARRYB_19__6_) );
  NAND2_X2 mul_ex_mult_90_U688 ( .A1(mul_ex_mult_90_SUMB_18__7_), .A2(
        mul_ex_mult_90_CARRYB_18__6_), .ZN(mul_ex_mult_90_n238) );
  INV_X4 mul_ex_mult_90_U687 ( .A(mul_ex_mult_90_n237), .ZN(
        mul_ex_mult_90_SUMB_19__7_) );
  XNOR2_X2 mul_ex_mult_90_U686 ( .A(mul_ex_mult_90_CARRYB_18__7_), .B(
        mul_ex_mult_90_SUMB_18__8_), .ZN(mul_ex_mult_90_n237) );
  INV_X4 mul_ex_mult_90_U685 ( .A(mul_ex_mult_90_n236), .ZN(
        mul_ex_mult_90_CARRYB_19__7_) );
  NAND2_X2 mul_ex_mult_90_U684 ( .A1(mul_ex_mult_90_SUMB_18__8_), .A2(
        mul_ex_mult_90_CARRYB_18__7_), .ZN(mul_ex_mult_90_n236) );
  INV_X4 mul_ex_mult_90_U683 ( .A(mul_ex_mult_90_n235), .ZN(
        mul_ex_mult_90_SUMB_19__8_) );
  XNOR2_X2 mul_ex_mult_90_U682 ( .A(mul_ex_mult_90_CARRYB_18__8_), .B(
        mul_ex_mult_90_SUMB_18__9_), .ZN(mul_ex_mult_90_n235) );
  INV_X4 mul_ex_mult_90_U681 ( .A(mul_ex_mult_90_n234), .ZN(
        mul_ex_mult_90_CARRYB_19__8_) );
  NAND2_X2 mul_ex_mult_90_U680 ( .A1(mul_ex_mult_90_SUMB_18__9_), .A2(
        mul_ex_mult_90_CARRYB_18__8_), .ZN(mul_ex_mult_90_n234) );
  INV_X4 mul_ex_mult_90_U679 ( .A(mul_ex_mult_90_n233), .ZN(
        mul_ex_mult_90_SUMB_18__9_) );
  XNOR2_X2 mul_ex_mult_90_U678 ( .A(mul_ex_mult_90_CARRYB_17__9_), .B(
        mul_ex_mult_90_SUMB_17__10_), .ZN(mul_ex_mult_90_n233) );
  INV_X4 mul_ex_mult_90_U677 ( .A(mul_ex_mult_90_n232), .ZN(
        mul_ex_mult_90_CARRYB_18__9_) );
  NAND2_X2 mul_ex_mult_90_U676 ( .A1(mul_ex_mult_90_SUMB_17__10_), .A2(
        mul_ex_mult_90_CARRYB_17__9_), .ZN(mul_ex_mult_90_n232) );
  INV_X4 mul_ex_mult_90_U675 ( .A(mul_ex_mult_90_n231), .ZN(mul_ex_N172) );
  XNOR2_X2 mul_ex_mult_90_U674 ( .A(mul_ex_mult_90_CARRYB_17__0_), .B(
        mul_ex_mult_90_SUMB_17__1_), .ZN(mul_ex_mult_90_n231) );
  INV_X4 mul_ex_mult_90_U673 ( .A(mul_ex_mult_90_n230), .ZN(
        mul_ex_mult_90_CARRYB_18__0_) );
  NAND2_X2 mul_ex_mult_90_U672 ( .A1(mul_ex_mult_90_SUMB_17__1_), .A2(
        mul_ex_mult_90_CARRYB_17__0_), .ZN(mul_ex_mult_90_n230) );
  INV_X4 mul_ex_mult_90_U671 ( .A(mul_ex_mult_90_n229), .ZN(
        mul_ex_mult_90_SUMB_18__10_) );
  XNOR2_X2 mul_ex_mult_90_U670 ( .A(mul_ex_mult_90_CARRYB_17__10_), .B(
        mul_ex_mult_90_SUMB_17__11_), .ZN(mul_ex_mult_90_n229) );
  INV_X4 mul_ex_mult_90_U669 ( .A(mul_ex_mult_90_n228), .ZN(
        mul_ex_mult_90_CARRYB_18__10_) );
  NAND2_X2 mul_ex_mult_90_U668 ( .A1(mul_ex_mult_90_SUMB_17__11_), .A2(
        mul_ex_mult_90_CARRYB_17__10_), .ZN(mul_ex_mult_90_n228) );
  INV_X4 mul_ex_mult_90_U667 ( .A(mul_ex_mult_90_n227), .ZN(
        mul_ex_mult_90_SUMB_18__11_) );
  XNOR2_X2 mul_ex_mult_90_U666 ( .A(mul_ex_mult_90_CARRYB_17__11_), .B(
        mul_ex_mult_90_SUMB_17__12_), .ZN(mul_ex_mult_90_n227) );
  INV_X4 mul_ex_mult_90_U665 ( .A(mul_ex_mult_90_n226), .ZN(
        mul_ex_mult_90_CARRYB_18__11_) );
  NAND2_X2 mul_ex_mult_90_U664 ( .A1(mul_ex_mult_90_SUMB_17__12_), .A2(
        mul_ex_mult_90_CARRYB_17__11_), .ZN(mul_ex_mult_90_n226) );
  INV_X4 mul_ex_mult_90_U663 ( .A(mul_ex_mult_90_n225), .ZN(
        mul_ex_mult_90_SUMB_18__12_) );
  XNOR2_X2 mul_ex_mult_90_U662 ( .A(mul_ex_mult_90_CARRYB_17__12_), .B(
        mul_ex_mult_90_SUMB_17__13_), .ZN(mul_ex_mult_90_n225) );
  INV_X4 mul_ex_mult_90_U661 ( .A(mul_ex_mult_90_n224), .ZN(
        mul_ex_mult_90_CARRYB_18__12_) );
  NAND2_X2 mul_ex_mult_90_U660 ( .A1(mul_ex_mult_90_SUMB_17__13_), .A2(
        mul_ex_mult_90_CARRYB_17__12_), .ZN(mul_ex_mult_90_n224) );
  INV_X4 mul_ex_mult_90_U659 ( .A(mul_ex_mult_90_n223), .ZN(
        mul_ex_mult_90_SUMB_18__1_) );
  XNOR2_X2 mul_ex_mult_90_U658 ( .A(mul_ex_mult_90_CARRYB_17__1_), .B(
        mul_ex_mult_90_SUMB_17__2_), .ZN(mul_ex_mult_90_n223) );
  INV_X4 mul_ex_mult_90_U657 ( .A(mul_ex_mult_90_n222), .ZN(
        mul_ex_mult_90_CARRYB_18__1_) );
  NAND2_X2 mul_ex_mult_90_U656 ( .A1(mul_ex_mult_90_SUMB_17__2_), .A2(
        mul_ex_mult_90_CARRYB_17__1_), .ZN(mul_ex_mult_90_n222) );
  INV_X4 mul_ex_mult_90_U655 ( .A(mul_ex_mult_90_n221), .ZN(
        mul_ex_mult_90_SUMB_18__2_) );
  XNOR2_X2 mul_ex_mult_90_U654 ( .A(mul_ex_mult_90_CARRYB_17__2_), .B(
        mul_ex_mult_90_SUMB_17__3_), .ZN(mul_ex_mult_90_n221) );
  INV_X4 mul_ex_mult_90_U653 ( .A(mul_ex_mult_90_n220), .ZN(
        mul_ex_mult_90_CARRYB_18__2_) );
  NAND2_X2 mul_ex_mult_90_U652 ( .A1(mul_ex_mult_90_SUMB_17__3_), .A2(
        mul_ex_mult_90_CARRYB_17__2_), .ZN(mul_ex_mult_90_n220) );
  INV_X4 mul_ex_mult_90_U651 ( .A(mul_ex_mult_90_n219), .ZN(
        mul_ex_mult_90_SUMB_18__3_) );
  XNOR2_X2 mul_ex_mult_90_U650 ( .A(mul_ex_mult_90_CARRYB_17__3_), .B(
        mul_ex_mult_90_SUMB_17__4_), .ZN(mul_ex_mult_90_n219) );
  INV_X4 mul_ex_mult_90_U649 ( .A(mul_ex_mult_90_n218), .ZN(
        mul_ex_mult_90_CARRYB_18__3_) );
  NAND2_X2 mul_ex_mult_90_U648 ( .A1(mul_ex_mult_90_SUMB_17__4_), .A2(
        mul_ex_mult_90_CARRYB_17__3_), .ZN(mul_ex_mult_90_n218) );
  INV_X4 mul_ex_mult_90_U647 ( .A(mul_ex_mult_90_n217), .ZN(
        mul_ex_mult_90_SUMB_18__4_) );
  XNOR2_X2 mul_ex_mult_90_U646 ( .A(mul_ex_mult_90_CARRYB_17__4_), .B(
        mul_ex_mult_90_SUMB_17__5_), .ZN(mul_ex_mult_90_n217) );
  INV_X4 mul_ex_mult_90_U645 ( .A(mul_ex_mult_90_n216), .ZN(
        mul_ex_mult_90_CARRYB_18__4_) );
  NAND2_X2 mul_ex_mult_90_U644 ( .A1(mul_ex_mult_90_SUMB_17__5_), .A2(
        mul_ex_mult_90_CARRYB_17__4_), .ZN(mul_ex_mult_90_n216) );
  INV_X4 mul_ex_mult_90_U643 ( .A(mul_ex_mult_90_n215), .ZN(
        mul_ex_mult_90_SUMB_18__5_) );
  XNOR2_X2 mul_ex_mult_90_U642 ( .A(mul_ex_mult_90_CARRYB_17__5_), .B(
        mul_ex_mult_90_SUMB_17__6_), .ZN(mul_ex_mult_90_n215) );
  INV_X4 mul_ex_mult_90_U641 ( .A(mul_ex_mult_90_n214), .ZN(
        mul_ex_mult_90_CARRYB_18__5_) );
  NAND2_X2 mul_ex_mult_90_U640 ( .A1(mul_ex_mult_90_SUMB_17__6_), .A2(
        mul_ex_mult_90_CARRYB_17__5_), .ZN(mul_ex_mult_90_n214) );
  INV_X4 mul_ex_mult_90_U639 ( .A(mul_ex_mult_90_n213), .ZN(
        mul_ex_mult_90_SUMB_18__6_) );
  XNOR2_X2 mul_ex_mult_90_U638 ( .A(mul_ex_mult_90_CARRYB_17__6_), .B(
        mul_ex_mult_90_SUMB_17__7_), .ZN(mul_ex_mult_90_n213) );
  INV_X4 mul_ex_mult_90_U637 ( .A(mul_ex_mult_90_n212), .ZN(
        mul_ex_mult_90_CARRYB_18__6_) );
  NAND2_X2 mul_ex_mult_90_U636 ( .A1(mul_ex_mult_90_SUMB_17__7_), .A2(
        mul_ex_mult_90_CARRYB_17__6_), .ZN(mul_ex_mult_90_n212) );
  INV_X4 mul_ex_mult_90_U635 ( .A(mul_ex_mult_90_n211), .ZN(
        mul_ex_mult_90_SUMB_18__7_) );
  XNOR2_X2 mul_ex_mult_90_U634 ( .A(mul_ex_mult_90_CARRYB_17__7_), .B(
        mul_ex_mult_90_SUMB_17__8_), .ZN(mul_ex_mult_90_n211) );
  INV_X4 mul_ex_mult_90_U633 ( .A(mul_ex_mult_90_n210), .ZN(
        mul_ex_mult_90_CARRYB_18__7_) );
  NAND2_X2 mul_ex_mult_90_U632 ( .A1(mul_ex_mult_90_SUMB_17__8_), .A2(
        mul_ex_mult_90_CARRYB_17__7_), .ZN(mul_ex_mult_90_n210) );
  INV_X4 mul_ex_mult_90_U631 ( .A(mul_ex_mult_90_n209), .ZN(
        mul_ex_mult_90_SUMB_18__8_) );
  XNOR2_X2 mul_ex_mult_90_U630 ( .A(mul_ex_mult_90_CARRYB_17__8_), .B(
        mul_ex_mult_90_SUMB_17__9_), .ZN(mul_ex_mult_90_n209) );
  INV_X4 mul_ex_mult_90_U629 ( .A(mul_ex_mult_90_n208), .ZN(
        mul_ex_mult_90_CARRYB_18__8_) );
  NAND2_X2 mul_ex_mult_90_U628 ( .A1(mul_ex_mult_90_SUMB_17__9_), .A2(
        mul_ex_mult_90_CARRYB_17__8_), .ZN(mul_ex_mult_90_n208) );
  INV_X4 mul_ex_mult_90_U627 ( .A(mul_ex_mult_90_n207), .ZN(
        mul_ex_mult_90_SUMB_17__9_) );
  XNOR2_X2 mul_ex_mult_90_U626 ( .A(mul_ex_mult_90_CARRYB_16__9_), .B(
        mul_ex_mult_90_SUMB_16__10_), .ZN(mul_ex_mult_90_n207) );
  INV_X4 mul_ex_mult_90_U625 ( .A(mul_ex_mult_90_n206), .ZN(
        mul_ex_mult_90_CARRYB_17__9_) );
  NAND2_X2 mul_ex_mult_90_U624 ( .A1(mul_ex_mult_90_SUMB_16__10_), .A2(
        mul_ex_mult_90_CARRYB_16__9_), .ZN(mul_ex_mult_90_n206) );
  INV_X4 mul_ex_mult_90_U623 ( .A(mul_ex_mult_90_n205), .ZN(mul_ex_N171) );
  XNOR2_X2 mul_ex_mult_90_U622 ( .A(mul_ex_mult_90_CARRYB_16__0_), .B(
        mul_ex_mult_90_SUMB_16__1_), .ZN(mul_ex_mult_90_n205) );
  INV_X4 mul_ex_mult_90_U621 ( .A(mul_ex_mult_90_n204), .ZN(
        mul_ex_mult_90_CARRYB_17__0_) );
  NAND2_X2 mul_ex_mult_90_U620 ( .A1(mul_ex_mult_90_SUMB_16__1_), .A2(
        mul_ex_mult_90_CARRYB_16__0_), .ZN(mul_ex_mult_90_n204) );
  INV_X4 mul_ex_mult_90_U619 ( .A(mul_ex_mult_90_n203), .ZN(
        mul_ex_mult_90_SUMB_17__10_) );
  XNOR2_X2 mul_ex_mult_90_U618 ( .A(mul_ex_mult_90_CARRYB_16__10_), .B(
        mul_ex_mult_90_SUMB_16__11_), .ZN(mul_ex_mult_90_n203) );
  INV_X4 mul_ex_mult_90_U617 ( .A(mul_ex_mult_90_n202), .ZN(
        mul_ex_mult_90_CARRYB_17__10_) );
  NAND2_X2 mul_ex_mult_90_U616 ( .A1(mul_ex_mult_90_SUMB_16__11_), .A2(
        mul_ex_mult_90_CARRYB_16__10_), .ZN(mul_ex_mult_90_n202) );
  INV_X4 mul_ex_mult_90_U615 ( .A(mul_ex_mult_90_n201), .ZN(
        mul_ex_mult_90_SUMB_17__11_) );
  XNOR2_X2 mul_ex_mult_90_U614 ( .A(mul_ex_mult_90_CARRYB_16__11_), .B(
        mul_ex_mult_90_SUMB_16__12_), .ZN(mul_ex_mult_90_n201) );
  INV_X4 mul_ex_mult_90_U613 ( .A(mul_ex_mult_90_n200), .ZN(
        mul_ex_mult_90_CARRYB_17__11_) );
  NAND2_X2 mul_ex_mult_90_U612 ( .A1(mul_ex_mult_90_SUMB_16__12_), .A2(
        mul_ex_mult_90_CARRYB_16__11_), .ZN(mul_ex_mult_90_n200) );
  INV_X4 mul_ex_mult_90_U611 ( .A(mul_ex_mult_90_n199), .ZN(
        mul_ex_mult_90_SUMB_17__12_) );
  XNOR2_X2 mul_ex_mult_90_U610 ( .A(mul_ex_mult_90_CARRYB_16__12_), .B(
        mul_ex_mult_90_SUMB_16__13_), .ZN(mul_ex_mult_90_n199) );
  INV_X4 mul_ex_mult_90_U609 ( .A(mul_ex_mult_90_n198), .ZN(
        mul_ex_mult_90_CARRYB_17__12_) );
  NAND2_X2 mul_ex_mult_90_U608 ( .A1(mul_ex_mult_90_SUMB_16__13_), .A2(
        mul_ex_mult_90_CARRYB_16__12_), .ZN(mul_ex_mult_90_n198) );
  INV_X4 mul_ex_mult_90_U607 ( .A(mul_ex_mult_90_n197), .ZN(
        mul_ex_mult_90_SUMB_17__13_) );
  XNOR2_X2 mul_ex_mult_90_U606 ( .A(mul_ex_mult_90_CARRYB_16__13_), .B(
        mul_ex_mult_90_SUMB_16__14_), .ZN(mul_ex_mult_90_n197) );
  INV_X4 mul_ex_mult_90_U605 ( .A(mul_ex_mult_90_n196), .ZN(
        mul_ex_mult_90_CARRYB_17__13_) );
  NAND2_X2 mul_ex_mult_90_U604 ( .A1(mul_ex_mult_90_SUMB_16__14_), .A2(
        mul_ex_mult_90_CARRYB_16__13_), .ZN(mul_ex_mult_90_n196) );
  INV_X4 mul_ex_mult_90_U603 ( .A(mul_ex_mult_90_n195), .ZN(
        mul_ex_mult_90_SUMB_17__1_) );
  XNOR2_X2 mul_ex_mult_90_U602 ( .A(mul_ex_mult_90_CARRYB_16__1_), .B(
        mul_ex_mult_90_SUMB_16__2_), .ZN(mul_ex_mult_90_n195) );
  INV_X4 mul_ex_mult_90_U601 ( .A(mul_ex_mult_90_n194), .ZN(
        mul_ex_mult_90_CARRYB_17__1_) );
  NAND2_X2 mul_ex_mult_90_U600 ( .A1(mul_ex_mult_90_SUMB_16__2_), .A2(
        mul_ex_mult_90_CARRYB_16__1_), .ZN(mul_ex_mult_90_n194) );
  INV_X4 mul_ex_mult_90_U599 ( .A(mul_ex_mult_90_n193), .ZN(
        mul_ex_mult_90_SUMB_17__2_) );
  XNOR2_X2 mul_ex_mult_90_U598 ( .A(mul_ex_mult_90_CARRYB_16__2_), .B(
        mul_ex_mult_90_SUMB_16__3_), .ZN(mul_ex_mult_90_n193) );
  INV_X4 mul_ex_mult_90_U597 ( .A(mul_ex_mult_90_n192), .ZN(
        mul_ex_mult_90_CARRYB_17__2_) );
  NAND2_X2 mul_ex_mult_90_U596 ( .A1(mul_ex_mult_90_SUMB_16__3_), .A2(
        mul_ex_mult_90_CARRYB_16__2_), .ZN(mul_ex_mult_90_n192) );
  INV_X4 mul_ex_mult_90_U595 ( .A(mul_ex_mult_90_n191), .ZN(
        mul_ex_mult_90_SUMB_17__3_) );
  XNOR2_X2 mul_ex_mult_90_U594 ( .A(mul_ex_mult_90_CARRYB_16__3_), .B(
        mul_ex_mult_90_SUMB_16__4_), .ZN(mul_ex_mult_90_n191) );
  INV_X4 mul_ex_mult_90_U593 ( .A(mul_ex_mult_90_n190), .ZN(
        mul_ex_mult_90_CARRYB_17__3_) );
  NAND2_X2 mul_ex_mult_90_U592 ( .A1(mul_ex_mult_90_SUMB_16__4_), .A2(
        mul_ex_mult_90_CARRYB_16__3_), .ZN(mul_ex_mult_90_n190) );
  INV_X4 mul_ex_mult_90_U591 ( .A(mul_ex_mult_90_n189), .ZN(
        mul_ex_mult_90_SUMB_17__4_) );
  XNOR2_X2 mul_ex_mult_90_U590 ( .A(mul_ex_mult_90_CARRYB_16__4_), .B(
        mul_ex_mult_90_SUMB_16__5_), .ZN(mul_ex_mult_90_n189) );
  INV_X4 mul_ex_mult_90_U589 ( .A(mul_ex_mult_90_n188), .ZN(
        mul_ex_mult_90_CARRYB_17__4_) );
  NAND2_X2 mul_ex_mult_90_U588 ( .A1(mul_ex_mult_90_SUMB_16__5_), .A2(
        mul_ex_mult_90_CARRYB_16__4_), .ZN(mul_ex_mult_90_n188) );
  INV_X4 mul_ex_mult_90_U587 ( .A(mul_ex_mult_90_n187), .ZN(
        mul_ex_mult_90_SUMB_17__5_) );
  XNOR2_X2 mul_ex_mult_90_U586 ( .A(mul_ex_mult_90_CARRYB_16__5_), .B(
        mul_ex_mult_90_SUMB_16__6_), .ZN(mul_ex_mult_90_n187) );
  INV_X4 mul_ex_mult_90_U585 ( .A(mul_ex_mult_90_n186), .ZN(
        mul_ex_mult_90_CARRYB_17__5_) );
  NAND2_X2 mul_ex_mult_90_U584 ( .A1(mul_ex_mult_90_SUMB_16__6_), .A2(
        mul_ex_mult_90_CARRYB_16__5_), .ZN(mul_ex_mult_90_n186) );
  INV_X4 mul_ex_mult_90_U583 ( .A(mul_ex_mult_90_n185), .ZN(
        mul_ex_mult_90_SUMB_17__6_) );
  XNOR2_X2 mul_ex_mult_90_U582 ( .A(mul_ex_mult_90_CARRYB_16__6_), .B(
        mul_ex_mult_90_SUMB_16__7_), .ZN(mul_ex_mult_90_n185) );
  INV_X4 mul_ex_mult_90_U581 ( .A(mul_ex_mult_90_n184), .ZN(
        mul_ex_mult_90_CARRYB_17__6_) );
  NAND2_X2 mul_ex_mult_90_U580 ( .A1(mul_ex_mult_90_SUMB_16__7_), .A2(
        mul_ex_mult_90_CARRYB_16__6_), .ZN(mul_ex_mult_90_n184) );
  INV_X4 mul_ex_mult_90_U579 ( .A(mul_ex_mult_90_n183), .ZN(
        mul_ex_mult_90_SUMB_17__7_) );
  XNOR2_X2 mul_ex_mult_90_U578 ( .A(mul_ex_mult_90_CARRYB_16__7_), .B(
        mul_ex_mult_90_SUMB_16__8_), .ZN(mul_ex_mult_90_n183) );
  INV_X4 mul_ex_mult_90_U577 ( .A(mul_ex_mult_90_n182), .ZN(
        mul_ex_mult_90_CARRYB_17__7_) );
  NAND2_X2 mul_ex_mult_90_U576 ( .A1(mul_ex_mult_90_SUMB_16__8_), .A2(
        mul_ex_mult_90_CARRYB_16__7_), .ZN(mul_ex_mult_90_n182) );
  INV_X4 mul_ex_mult_90_U575 ( .A(mul_ex_mult_90_n181), .ZN(
        mul_ex_mult_90_SUMB_17__8_) );
  XNOR2_X2 mul_ex_mult_90_U574 ( .A(mul_ex_mult_90_CARRYB_16__8_), .B(
        mul_ex_mult_90_SUMB_16__9_), .ZN(mul_ex_mult_90_n181) );
  INV_X4 mul_ex_mult_90_U573 ( .A(mul_ex_mult_90_n180), .ZN(
        mul_ex_mult_90_CARRYB_17__8_) );
  NAND2_X2 mul_ex_mult_90_U572 ( .A1(mul_ex_mult_90_SUMB_16__9_), .A2(
        mul_ex_mult_90_CARRYB_16__8_), .ZN(mul_ex_mult_90_n180) );
  INV_X4 mul_ex_mult_90_U571 ( .A(mul_ex_mult_90_n179), .ZN(mul_ex_N184) );
  XNOR2_X2 mul_ex_mult_90_U570 ( .A(mul_ex_mult_90_CARRYB_29__0_), .B(
        mul_ex_mult_90_SUMB_29__1_), .ZN(mul_ex_mult_90_n179) );
  INV_X4 mul_ex_mult_90_U569 ( .A(mul_ex_mult_90_n178), .ZN(
        mul_ex_mult_90_CARRYB_30__0_) );
  NAND2_X2 mul_ex_mult_90_U568 ( .A1(mul_ex_mult_90_SUMB_29__1_), .A2(
        mul_ex_mult_90_CARRYB_29__0_), .ZN(mul_ex_mult_90_n178) );
  INV_X4 mul_ex_mult_90_U567 ( .A(mul_ex_mult_90_n177), .ZN(mul_ex_N183) );
  XNOR2_X2 mul_ex_mult_90_U566 ( .A(mul_ex_mult_90_CARRYB_28__0_), .B(
        mul_ex_mult_90_SUMB_28__1_), .ZN(mul_ex_mult_90_n177) );
  INV_X4 mul_ex_mult_90_U565 ( .A(mul_ex_mult_90_n176), .ZN(
        mul_ex_mult_90_CARRYB_29__0_) );
  NAND2_X2 mul_ex_mult_90_U564 ( .A1(mul_ex_mult_90_SUMB_28__1_), .A2(
        mul_ex_mult_90_CARRYB_28__0_), .ZN(mul_ex_mult_90_n176) );
  INV_X4 mul_ex_mult_90_U563 ( .A(mul_ex_mult_90_n175), .ZN(
        mul_ex_mult_90_SUMB_29__1_) );
  XNOR2_X2 mul_ex_mult_90_U562 ( .A(mul_ex_mult_90_CARRYB_28__1_), .B(
        mul_ex_mult_90_SUMB_28__2_), .ZN(mul_ex_mult_90_n175) );
  INV_X4 mul_ex_mult_90_U561 ( .A(mul_ex_mult_90_n174), .ZN(
        mul_ex_mult_90_CARRYB_29__1_) );
  NAND2_X2 mul_ex_mult_90_U560 ( .A1(mul_ex_mult_90_SUMB_28__2_), .A2(
        mul_ex_mult_90_CARRYB_28__1_), .ZN(mul_ex_mult_90_n174) );
  INV_X4 mul_ex_mult_90_U559 ( .A(mul_ex_mult_90_n173), .ZN(mul_ex_N182) );
  XNOR2_X2 mul_ex_mult_90_U558 ( .A(mul_ex_mult_90_CARRYB_27__0_), .B(
        mul_ex_mult_90_SUMB_27__1_), .ZN(mul_ex_mult_90_n173) );
  INV_X4 mul_ex_mult_90_U557 ( .A(mul_ex_mult_90_n172), .ZN(
        mul_ex_mult_90_CARRYB_28__0_) );
  NAND2_X2 mul_ex_mult_90_U556 ( .A1(mul_ex_mult_90_SUMB_27__1_), .A2(
        mul_ex_mult_90_CARRYB_27__0_), .ZN(mul_ex_mult_90_n172) );
  INV_X4 mul_ex_mult_90_U555 ( .A(mul_ex_mult_90_n171), .ZN(
        mul_ex_mult_90_SUMB_28__1_) );
  XNOR2_X2 mul_ex_mult_90_U554 ( .A(mul_ex_mult_90_CARRYB_27__1_), .B(
        mul_ex_mult_90_SUMB_27__2_), .ZN(mul_ex_mult_90_n171) );
  INV_X4 mul_ex_mult_90_U553 ( .A(mul_ex_mult_90_n170), .ZN(
        mul_ex_mult_90_CARRYB_28__1_) );
  NAND2_X2 mul_ex_mult_90_U552 ( .A1(mul_ex_mult_90_SUMB_27__2_), .A2(
        mul_ex_mult_90_CARRYB_27__1_), .ZN(mul_ex_mult_90_n170) );
  INV_X4 mul_ex_mult_90_U551 ( .A(mul_ex_mult_90_n169), .ZN(
        mul_ex_mult_90_SUMB_28__2_) );
  XNOR2_X2 mul_ex_mult_90_U550 ( .A(mul_ex_mult_90_CARRYB_27__2_), .B(
        mul_ex_mult_90_SUMB_27__3_), .ZN(mul_ex_mult_90_n169) );
  INV_X4 mul_ex_mult_90_U549 ( .A(mul_ex_mult_90_n168), .ZN(
        mul_ex_mult_90_CARRYB_28__2_) );
  NAND2_X2 mul_ex_mult_90_U548 ( .A1(mul_ex_mult_90_SUMB_27__3_), .A2(
        mul_ex_mult_90_CARRYB_27__2_), .ZN(mul_ex_mult_90_n168) );
  INV_X4 mul_ex_mult_90_U547 ( .A(mul_ex_mult_90_n167), .ZN(mul_ex_N181) );
  XNOR2_X2 mul_ex_mult_90_U546 ( .A(mul_ex_mult_90_CARRYB_26__0_), .B(
        mul_ex_mult_90_SUMB_26__1_), .ZN(mul_ex_mult_90_n167) );
  INV_X4 mul_ex_mult_90_U545 ( .A(mul_ex_mult_90_n166), .ZN(
        mul_ex_mult_90_CARRYB_27__0_) );
  NAND2_X2 mul_ex_mult_90_U544 ( .A1(mul_ex_mult_90_SUMB_26__1_), .A2(
        mul_ex_mult_90_CARRYB_26__0_), .ZN(mul_ex_mult_90_n166) );
  INV_X4 mul_ex_mult_90_U543 ( .A(mul_ex_mult_90_n165), .ZN(
        mul_ex_mult_90_SUMB_27__1_) );
  XNOR2_X2 mul_ex_mult_90_U542 ( .A(mul_ex_mult_90_CARRYB_26__1_), .B(
        mul_ex_mult_90_SUMB_26__2_), .ZN(mul_ex_mult_90_n165) );
  INV_X4 mul_ex_mult_90_U541 ( .A(mul_ex_mult_90_n164), .ZN(
        mul_ex_mult_90_CARRYB_27__1_) );
  NAND2_X2 mul_ex_mult_90_U540 ( .A1(mul_ex_mult_90_SUMB_26__2_), .A2(
        mul_ex_mult_90_CARRYB_26__1_), .ZN(mul_ex_mult_90_n164) );
  INV_X4 mul_ex_mult_90_U539 ( .A(mul_ex_mult_90_n163), .ZN(
        mul_ex_mult_90_SUMB_27__2_) );
  XNOR2_X2 mul_ex_mult_90_U538 ( .A(mul_ex_mult_90_CARRYB_26__2_), .B(
        mul_ex_mult_90_SUMB_26__3_), .ZN(mul_ex_mult_90_n163) );
  INV_X4 mul_ex_mult_90_U537 ( .A(mul_ex_mult_90_n162), .ZN(
        mul_ex_mult_90_CARRYB_27__2_) );
  NAND2_X2 mul_ex_mult_90_U536 ( .A1(mul_ex_mult_90_SUMB_26__3_), .A2(
        mul_ex_mult_90_CARRYB_26__2_), .ZN(mul_ex_mult_90_n162) );
  INV_X4 mul_ex_mult_90_U535 ( .A(mul_ex_mult_90_n161), .ZN(
        mul_ex_mult_90_SUMB_27__3_) );
  XNOR2_X2 mul_ex_mult_90_U534 ( .A(mul_ex_mult_90_CARRYB_26__3_), .B(
        mul_ex_mult_90_SUMB_26__4_), .ZN(mul_ex_mult_90_n161) );
  INV_X4 mul_ex_mult_90_U533 ( .A(mul_ex_mult_90_n160), .ZN(
        mul_ex_mult_90_CARRYB_27__3_) );
  NAND2_X2 mul_ex_mult_90_U532 ( .A1(mul_ex_mult_90_SUMB_26__4_), .A2(
        mul_ex_mult_90_CARRYB_26__3_), .ZN(mul_ex_mult_90_n160) );
  INV_X4 mul_ex_mult_90_U531 ( .A(mul_ex_mult_90_n159), .ZN(mul_ex_N180) );
  XNOR2_X2 mul_ex_mult_90_U530 ( .A(mul_ex_mult_90_CARRYB_25__0_), .B(
        mul_ex_mult_90_SUMB_25__1_), .ZN(mul_ex_mult_90_n159) );
  INV_X4 mul_ex_mult_90_U529 ( .A(mul_ex_mult_90_n158), .ZN(
        mul_ex_mult_90_CARRYB_26__0_) );
  NAND2_X2 mul_ex_mult_90_U528 ( .A1(mul_ex_mult_90_SUMB_25__1_), .A2(
        mul_ex_mult_90_CARRYB_25__0_), .ZN(mul_ex_mult_90_n158) );
  INV_X4 mul_ex_mult_90_U527 ( .A(mul_ex_mult_90_n157), .ZN(
        mul_ex_mult_90_SUMB_26__1_) );
  XNOR2_X2 mul_ex_mult_90_U526 ( .A(mul_ex_mult_90_CARRYB_25__1_), .B(
        mul_ex_mult_90_SUMB_25__2_), .ZN(mul_ex_mult_90_n157) );
  INV_X4 mul_ex_mult_90_U525 ( .A(mul_ex_mult_90_n156), .ZN(
        mul_ex_mult_90_CARRYB_26__1_) );
  NAND2_X2 mul_ex_mult_90_U524 ( .A1(mul_ex_mult_90_SUMB_25__2_), .A2(
        mul_ex_mult_90_CARRYB_25__1_), .ZN(mul_ex_mult_90_n156) );
  INV_X4 mul_ex_mult_90_U523 ( .A(mul_ex_mult_90_n155), .ZN(
        mul_ex_mult_90_SUMB_26__2_) );
  XNOR2_X2 mul_ex_mult_90_U522 ( .A(mul_ex_mult_90_CARRYB_25__2_), .B(
        mul_ex_mult_90_SUMB_25__3_), .ZN(mul_ex_mult_90_n155) );
  INV_X4 mul_ex_mult_90_U521 ( .A(mul_ex_mult_90_n154), .ZN(
        mul_ex_mult_90_CARRYB_26__2_) );
  NAND2_X2 mul_ex_mult_90_U520 ( .A1(mul_ex_mult_90_SUMB_25__3_), .A2(
        mul_ex_mult_90_CARRYB_25__2_), .ZN(mul_ex_mult_90_n154) );
  INV_X4 mul_ex_mult_90_U519 ( .A(mul_ex_mult_90_n153), .ZN(
        mul_ex_mult_90_SUMB_26__3_) );
  XNOR2_X2 mul_ex_mult_90_U518 ( .A(mul_ex_mult_90_CARRYB_25__3_), .B(
        mul_ex_mult_90_SUMB_25__4_), .ZN(mul_ex_mult_90_n153) );
  INV_X4 mul_ex_mult_90_U517 ( .A(mul_ex_mult_90_n152), .ZN(
        mul_ex_mult_90_CARRYB_26__3_) );
  NAND2_X2 mul_ex_mult_90_U516 ( .A1(mul_ex_mult_90_SUMB_25__4_), .A2(
        mul_ex_mult_90_CARRYB_25__3_), .ZN(mul_ex_mult_90_n152) );
  INV_X4 mul_ex_mult_90_U515 ( .A(mul_ex_mult_90_n151), .ZN(
        mul_ex_mult_90_SUMB_26__4_) );
  XNOR2_X2 mul_ex_mult_90_U514 ( .A(mul_ex_mult_90_CARRYB_25__4_), .B(
        mul_ex_mult_90_SUMB_25__5_), .ZN(mul_ex_mult_90_n151) );
  INV_X4 mul_ex_mult_90_U513 ( .A(mul_ex_mult_90_n150), .ZN(
        mul_ex_mult_90_CARRYB_26__4_) );
  NAND2_X2 mul_ex_mult_90_U512 ( .A1(mul_ex_mult_90_SUMB_25__5_), .A2(
        mul_ex_mult_90_CARRYB_25__4_), .ZN(mul_ex_mult_90_n150) );
  INV_X4 mul_ex_mult_90_U511 ( .A(mul_ex_mult_90_n149), .ZN(mul_ex_N179) );
  XNOR2_X2 mul_ex_mult_90_U510 ( .A(mul_ex_mult_90_CARRYB_24__0_), .B(
        mul_ex_mult_90_SUMB_24__1_), .ZN(mul_ex_mult_90_n149) );
  INV_X4 mul_ex_mult_90_U509 ( .A(mul_ex_mult_90_n148), .ZN(
        mul_ex_mult_90_CARRYB_25__0_) );
  NAND2_X2 mul_ex_mult_90_U508 ( .A1(mul_ex_mult_90_SUMB_24__1_), .A2(
        mul_ex_mult_90_CARRYB_24__0_), .ZN(mul_ex_mult_90_n148) );
  INV_X4 mul_ex_mult_90_U507 ( .A(mul_ex_mult_90_n147), .ZN(
        mul_ex_mult_90_SUMB_25__1_) );
  XNOR2_X2 mul_ex_mult_90_U506 ( .A(mul_ex_mult_90_CARRYB_24__1_), .B(
        mul_ex_mult_90_SUMB_24__2_), .ZN(mul_ex_mult_90_n147) );
  INV_X4 mul_ex_mult_90_U505 ( .A(mul_ex_mult_90_n146), .ZN(
        mul_ex_mult_90_CARRYB_25__1_) );
  NAND2_X2 mul_ex_mult_90_U504 ( .A1(mul_ex_mult_90_SUMB_24__2_), .A2(
        mul_ex_mult_90_CARRYB_24__1_), .ZN(mul_ex_mult_90_n146) );
  INV_X4 mul_ex_mult_90_U503 ( .A(mul_ex_mult_90_n145), .ZN(
        mul_ex_mult_90_SUMB_25__2_) );
  XNOR2_X2 mul_ex_mult_90_U502 ( .A(mul_ex_mult_90_CARRYB_24__2_), .B(
        mul_ex_mult_90_SUMB_24__3_), .ZN(mul_ex_mult_90_n145) );
  INV_X4 mul_ex_mult_90_U501 ( .A(mul_ex_mult_90_n144), .ZN(
        mul_ex_mult_90_CARRYB_25__2_) );
  NAND2_X2 mul_ex_mult_90_U500 ( .A1(mul_ex_mult_90_SUMB_24__3_), .A2(
        mul_ex_mult_90_CARRYB_24__2_), .ZN(mul_ex_mult_90_n144) );
  INV_X4 mul_ex_mult_90_U499 ( .A(mul_ex_mult_90_n143), .ZN(
        mul_ex_mult_90_SUMB_25__3_) );
  XNOR2_X2 mul_ex_mult_90_U498 ( .A(mul_ex_mult_90_CARRYB_24__3_), .B(
        mul_ex_mult_90_SUMB_24__4_), .ZN(mul_ex_mult_90_n143) );
  INV_X4 mul_ex_mult_90_U497 ( .A(mul_ex_mult_90_n142), .ZN(
        mul_ex_mult_90_CARRYB_25__3_) );
  NAND2_X2 mul_ex_mult_90_U205 ( .A1(mul_ex_mult_90_SUMB_24__4_), .A2(
        mul_ex_mult_90_CARRYB_24__3_), .ZN(mul_ex_mult_90_n142) );
  INV_X4 mul_ex_mult_90_U204 ( .A(mul_ex_mult_90_n141), .ZN(
        mul_ex_mult_90_SUMB_25__4_) );
  XNOR2_X2 mul_ex_mult_90_U203 ( .A(mul_ex_mult_90_CARRYB_24__4_), .B(
        mul_ex_mult_90_SUMB_24__5_), .ZN(mul_ex_mult_90_n141) );
  INV_X4 mul_ex_mult_90_U202 ( .A(mul_ex_mult_90_n140), .ZN(
        mul_ex_mult_90_CARRYB_25__4_) );
  NAND2_X2 mul_ex_mult_90_U201 ( .A1(mul_ex_mult_90_SUMB_24__5_), .A2(
        mul_ex_mult_90_CARRYB_24__4_), .ZN(mul_ex_mult_90_n140) );
  INV_X4 mul_ex_mult_90_U200 ( .A(mul_ex_mult_90_n139), .ZN(
        mul_ex_mult_90_SUMB_25__5_) );
  XNOR2_X2 mul_ex_mult_90_U199 ( .A(mul_ex_mult_90_CARRYB_24__5_), .B(
        mul_ex_mult_90_SUMB_24__6_), .ZN(mul_ex_mult_90_n139) );
  INV_X4 mul_ex_mult_90_U198 ( .A(mul_ex_mult_90_n138), .ZN(
        mul_ex_mult_90_CARRYB_25__5_) );
  NAND2_X2 mul_ex_mult_90_U197 ( .A1(mul_ex_mult_90_SUMB_24__6_), .A2(
        mul_ex_mult_90_CARRYB_24__5_), .ZN(mul_ex_mult_90_n138) );
  INV_X4 mul_ex_mult_90_U196 ( .A(mul_ex_mult_90_n137), .ZN(mul_ex_N178) );
  XNOR2_X2 mul_ex_mult_90_U195 ( .A(mul_ex_mult_90_CARRYB_23__0_), .B(
        mul_ex_mult_90_SUMB_23__1_), .ZN(mul_ex_mult_90_n137) );
  INV_X4 mul_ex_mult_90_U194 ( .A(mul_ex_mult_90_n136), .ZN(
        mul_ex_mult_90_CARRYB_24__0_) );
  NAND2_X2 mul_ex_mult_90_U193 ( .A1(mul_ex_mult_90_SUMB_23__1_), .A2(
        mul_ex_mult_90_CARRYB_23__0_), .ZN(mul_ex_mult_90_n136) );
  INV_X4 mul_ex_mult_90_U192 ( .A(mul_ex_mult_90_n135), .ZN(
        mul_ex_mult_90_SUMB_24__1_) );
  XNOR2_X2 mul_ex_mult_90_U191 ( .A(mul_ex_mult_90_CARRYB_23__1_), .B(
        mul_ex_mult_90_SUMB_23__2_), .ZN(mul_ex_mult_90_n135) );
  INV_X4 mul_ex_mult_90_U190 ( .A(mul_ex_mult_90_n134), .ZN(
        mul_ex_mult_90_CARRYB_24__1_) );
  NAND2_X2 mul_ex_mult_90_U189 ( .A1(mul_ex_mult_90_SUMB_23__2_), .A2(
        mul_ex_mult_90_CARRYB_23__1_), .ZN(mul_ex_mult_90_n134) );
  INV_X4 mul_ex_mult_90_U188 ( .A(mul_ex_mult_90_n133), .ZN(
        mul_ex_mult_90_SUMB_24__2_) );
  XNOR2_X2 mul_ex_mult_90_U187 ( .A(mul_ex_mult_90_CARRYB_23__2_), .B(
        mul_ex_mult_90_SUMB_23__3_), .ZN(mul_ex_mult_90_n133) );
  INV_X4 mul_ex_mult_90_U186 ( .A(mul_ex_mult_90_n132), .ZN(
        mul_ex_mult_90_CARRYB_24__2_) );
  NAND2_X2 mul_ex_mult_90_U185 ( .A1(mul_ex_mult_90_SUMB_23__3_), .A2(
        mul_ex_mult_90_CARRYB_23__2_), .ZN(mul_ex_mult_90_n132) );
  INV_X4 mul_ex_mult_90_U184 ( .A(mul_ex_mult_90_n131), .ZN(
        mul_ex_mult_90_SUMB_24__3_) );
  XNOR2_X2 mul_ex_mult_90_U183 ( .A(mul_ex_mult_90_CARRYB_23__3_), .B(
        mul_ex_mult_90_SUMB_23__4_), .ZN(mul_ex_mult_90_n131) );
  INV_X4 mul_ex_mult_90_U182 ( .A(mul_ex_mult_90_n130), .ZN(
        mul_ex_mult_90_CARRYB_24__3_) );
  NAND2_X2 mul_ex_mult_90_U181 ( .A1(mul_ex_mult_90_SUMB_23__4_), .A2(
        mul_ex_mult_90_CARRYB_23__3_), .ZN(mul_ex_mult_90_n130) );
  INV_X4 mul_ex_mult_90_U180 ( .A(mul_ex_mult_90_n129), .ZN(
        mul_ex_mult_90_SUMB_24__4_) );
  XNOR2_X2 mul_ex_mult_90_U179 ( .A(mul_ex_mult_90_CARRYB_23__4_), .B(
        mul_ex_mult_90_SUMB_23__5_), .ZN(mul_ex_mult_90_n129) );
  INV_X4 mul_ex_mult_90_U178 ( .A(mul_ex_mult_90_n128), .ZN(
        mul_ex_mult_90_CARRYB_24__4_) );
  NAND2_X2 mul_ex_mult_90_U177 ( .A1(mul_ex_mult_90_SUMB_23__5_), .A2(
        mul_ex_mult_90_CARRYB_23__4_), .ZN(mul_ex_mult_90_n128) );
  INV_X4 mul_ex_mult_90_U176 ( .A(mul_ex_mult_90_n127), .ZN(
        mul_ex_mult_90_SUMB_24__5_) );
  XNOR2_X2 mul_ex_mult_90_U175 ( .A(mul_ex_mult_90_CARRYB_23__5_), .B(
        mul_ex_mult_90_SUMB_23__6_), .ZN(mul_ex_mult_90_n127) );
  INV_X4 mul_ex_mult_90_U174 ( .A(mul_ex_mult_90_n126), .ZN(
        mul_ex_mult_90_CARRYB_24__5_) );
  NAND2_X2 mul_ex_mult_90_U173 ( .A1(mul_ex_mult_90_SUMB_23__6_), .A2(
        mul_ex_mult_90_CARRYB_23__5_), .ZN(mul_ex_mult_90_n126) );
  INV_X4 mul_ex_mult_90_U172 ( .A(mul_ex_mult_90_n125), .ZN(
        mul_ex_mult_90_SUMB_24__6_) );
  XNOR2_X2 mul_ex_mult_90_U171 ( .A(mul_ex_mult_90_CARRYB_23__6_), .B(
        mul_ex_mult_90_SUMB_23__7_), .ZN(mul_ex_mult_90_n125) );
  INV_X4 mul_ex_mult_90_U170 ( .A(mul_ex_mult_90_n124), .ZN(
        mul_ex_mult_90_CARRYB_24__6_) );
  NAND2_X2 mul_ex_mult_90_U169 ( .A1(mul_ex_mult_90_SUMB_23__7_), .A2(
        mul_ex_mult_90_CARRYB_23__6_), .ZN(mul_ex_mult_90_n124) );
  INV_X4 mul_ex_mult_90_U168 ( .A(mul_ex_mult_90_n123), .ZN(mul_ex_N177) );
  XNOR2_X2 mul_ex_mult_90_U167 ( .A(mul_ex_mult_90_CARRYB_22__0_), .B(
        mul_ex_mult_90_SUMB_22__1_), .ZN(mul_ex_mult_90_n123) );
  INV_X4 mul_ex_mult_90_U166 ( .A(mul_ex_mult_90_n122), .ZN(
        mul_ex_mult_90_CARRYB_23__0_) );
  NAND2_X2 mul_ex_mult_90_U165 ( .A1(mul_ex_mult_90_SUMB_22__1_), .A2(
        mul_ex_mult_90_CARRYB_22__0_), .ZN(mul_ex_mult_90_n122) );
  INV_X4 mul_ex_mult_90_U164 ( .A(mul_ex_mult_90_n121), .ZN(
        mul_ex_mult_90_SUMB_23__1_) );
  XNOR2_X2 mul_ex_mult_90_U163 ( .A(mul_ex_mult_90_CARRYB_22__1_), .B(
        mul_ex_mult_90_SUMB_22__2_), .ZN(mul_ex_mult_90_n121) );
  INV_X4 mul_ex_mult_90_U162 ( .A(mul_ex_mult_90_n120), .ZN(
        mul_ex_mult_90_CARRYB_23__1_) );
  NAND2_X2 mul_ex_mult_90_U161 ( .A1(mul_ex_mult_90_SUMB_22__2_), .A2(
        mul_ex_mult_90_CARRYB_22__1_), .ZN(mul_ex_mult_90_n120) );
  INV_X4 mul_ex_mult_90_U160 ( .A(mul_ex_mult_90_n119), .ZN(
        mul_ex_mult_90_SUMB_23__2_) );
  XNOR2_X2 mul_ex_mult_90_U159 ( .A(mul_ex_mult_90_CARRYB_22__2_), .B(
        mul_ex_mult_90_SUMB_22__3_), .ZN(mul_ex_mult_90_n119) );
  INV_X4 mul_ex_mult_90_U158 ( .A(mul_ex_mult_90_n118), .ZN(
        mul_ex_mult_90_CARRYB_23__2_) );
  NAND2_X2 mul_ex_mult_90_U157 ( .A1(mul_ex_mult_90_SUMB_22__3_), .A2(
        mul_ex_mult_90_CARRYB_22__2_), .ZN(mul_ex_mult_90_n118) );
  INV_X4 mul_ex_mult_90_U156 ( .A(mul_ex_mult_90_n117), .ZN(
        mul_ex_mult_90_SUMB_23__3_) );
  XNOR2_X2 mul_ex_mult_90_U155 ( .A(mul_ex_mult_90_CARRYB_22__3_), .B(
        mul_ex_mult_90_SUMB_22__4_), .ZN(mul_ex_mult_90_n117) );
  INV_X4 mul_ex_mult_90_U154 ( .A(mul_ex_mult_90_n116), .ZN(
        mul_ex_mult_90_CARRYB_23__3_) );
  NAND2_X2 mul_ex_mult_90_U153 ( .A1(mul_ex_mult_90_SUMB_22__4_), .A2(
        mul_ex_mult_90_CARRYB_22__3_), .ZN(mul_ex_mult_90_n116) );
  INV_X4 mul_ex_mult_90_U152 ( .A(mul_ex_mult_90_n115), .ZN(
        mul_ex_mult_90_SUMB_23__4_) );
  XNOR2_X2 mul_ex_mult_90_U151 ( .A(mul_ex_mult_90_CARRYB_22__4_), .B(
        mul_ex_mult_90_SUMB_22__5_), .ZN(mul_ex_mult_90_n115) );
  INV_X4 mul_ex_mult_90_U150 ( .A(mul_ex_mult_90_n114), .ZN(
        mul_ex_mult_90_CARRYB_23__4_) );
  NAND2_X2 mul_ex_mult_90_U149 ( .A1(mul_ex_mult_90_SUMB_22__5_), .A2(
        mul_ex_mult_90_CARRYB_22__4_), .ZN(mul_ex_mult_90_n114) );
  INV_X4 mul_ex_mult_90_U148 ( .A(mul_ex_mult_90_n113), .ZN(
        mul_ex_mult_90_SUMB_23__5_) );
  XNOR2_X2 mul_ex_mult_90_U147 ( .A(mul_ex_mult_90_CARRYB_22__5_), .B(
        mul_ex_mult_90_SUMB_22__6_), .ZN(mul_ex_mult_90_n113) );
  INV_X4 mul_ex_mult_90_U146 ( .A(mul_ex_mult_90_n112), .ZN(
        mul_ex_mult_90_CARRYB_23__5_) );
  NAND2_X2 mul_ex_mult_90_U145 ( .A1(mul_ex_mult_90_SUMB_22__6_), .A2(
        mul_ex_mult_90_CARRYB_22__5_), .ZN(mul_ex_mult_90_n112) );
  INV_X4 mul_ex_mult_90_U144 ( .A(mul_ex_mult_90_n111), .ZN(
        mul_ex_mult_90_SUMB_23__6_) );
  XNOR2_X2 mul_ex_mult_90_U143 ( .A(mul_ex_mult_90_CARRYB_22__6_), .B(
        mul_ex_mult_90_SUMB_22__7_), .ZN(mul_ex_mult_90_n111) );
  INV_X4 mul_ex_mult_90_U142 ( .A(mul_ex_mult_90_n110), .ZN(
        mul_ex_mult_90_CARRYB_23__6_) );
  NAND2_X2 mul_ex_mult_90_U141 ( .A1(mul_ex_mult_90_SUMB_22__7_), .A2(
        mul_ex_mult_90_CARRYB_22__6_), .ZN(mul_ex_mult_90_n110) );
  INV_X4 mul_ex_mult_90_U140 ( .A(mul_ex_mult_90_n109), .ZN(
        mul_ex_mult_90_SUMB_23__7_) );
  XNOR2_X2 mul_ex_mult_90_U139 ( .A(mul_ex_mult_90_CARRYB_22__7_), .B(
        mul_ex_mult_90_SUMB_22__8_), .ZN(mul_ex_mult_90_n109) );
  INV_X4 mul_ex_mult_90_U138 ( .A(mul_ex_mult_90_n108), .ZN(
        mul_ex_mult_90_CARRYB_23__7_) );
  NAND2_X2 mul_ex_mult_90_U137 ( .A1(mul_ex_mult_90_SUMB_22__8_), .A2(
        mul_ex_mult_90_CARRYB_22__7_), .ZN(mul_ex_mult_90_n108) );
  INV_X4 mul_ex_mult_90_U136 ( .A(mul_ex_mult_90_n107), .ZN(mul_ex_N176) );
  XNOR2_X2 mul_ex_mult_90_U135 ( .A(mul_ex_mult_90_CARRYB_21__0_), .B(
        mul_ex_mult_90_SUMB_21__1_), .ZN(mul_ex_mult_90_n107) );
  INV_X4 mul_ex_mult_90_U134 ( .A(mul_ex_mult_90_n106), .ZN(
        mul_ex_mult_90_CARRYB_22__0_) );
  NAND2_X2 mul_ex_mult_90_U133 ( .A1(mul_ex_mult_90_SUMB_21__1_), .A2(
        mul_ex_mult_90_CARRYB_21__0_), .ZN(mul_ex_mult_90_n106) );
  INV_X4 mul_ex_mult_90_U132 ( .A(mul_ex_mult_90_n105), .ZN(
        mul_ex_mult_90_SUMB_22__1_) );
  XNOR2_X2 mul_ex_mult_90_U131 ( .A(mul_ex_mult_90_CARRYB_21__1_), .B(
        mul_ex_mult_90_SUMB_21__2_), .ZN(mul_ex_mult_90_n105) );
  INV_X4 mul_ex_mult_90_U130 ( .A(mul_ex_mult_90_n104), .ZN(
        mul_ex_mult_90_CARRYB_22__1_) );
  NAND2_X2 mul_ex_mult_90_U129 ( .A1(mul_ex_mult_90_SUMB_21__2_), .A2(
        mul_ex_mult_90_CARRYB_21__1_), .ZN(mul_ex_mult_90_n104) );
  INV_X4 mul_ex_mult_90_U128 ( .A(mul_ex_mult_90_n103), .ZN(
        mul_ex_mult_90_SUMB_22__2_) );
  XNOR2_X2 mul_ex_mult_90_U127 ( .A(mul_ex_mult_90_CARRYB_21__2_), .B(
        mul_ex_mult_90_SUMB_21__3_), .ZN(mul_ex_mult_90_n103) );
  INV_X4 mul_ex_mult_90_U126 ( .A(mul_ex_mult_90_n102), .ZN(
        mul_ex_mult_90_CARRYB_22__2_) );
  NAND2_X2 mul_ex_mult_90_U125 ( .A1(mul_ex_mult_90_SUMB_21__3_), .A2(
        mul_ex_mult_90_CARRYB_21__2_), .ZN(mul_ex_mult_90_n102) );
  INV_X4 mul_ex_mult_90_U124 ( .A(mul_ex_mult_90_n101), .ZN(
        mul_ex_mult_90_SUMB_22__3_) );
  XNOR2_X2 mul_ex_mult_90_U123 ( .A(mul_ex_mult_90_CARRYB_21__3_), .B(
        mul_ex_mult_90_SUMB_21__4_), .ZN(mul_ex_mult_90_n101) );
  INV_X4 mul_ex_mult_90_U122 ( .A(mul_ex_mult_90_n100), .ZN(
        mul_ex_mult_90_CARRYB_22__3_) );
  NAND2_X2 mul_ex_mult_90_U121 ( .A1(mul_ex_mult_90_SUMB_21__4_), .A2(
        mul_ex_mult_90_CARRYB_21__3_), .ZN(mul_ex_mult_90_n100) );
  INV_X4 mul_ex_mult_90_U120 ( .A(mul_ex_mult_90_n99), .ZN(
        mul_ex_mult_90_SUMB_22__4_) );
  XNOR2_X2 mul_ex_mult_90_U119 ( .A(mul_ex_mult_90_CARRYB_21__4_), .B(
        mul_ex_mult_90_SUMB_21__5_), .ZN(mul_ex_mult_90_n99) );
  INV_X4 mul_ex_mult_90_U118 ( .A(mul_ex_mult_90_n98), .ZN(
        mul_ex_mult_90_CARRYB_22__4_) );
  NAND2_X2 mul_ex_mult_90_U117 ( .A1(mul_ex_mult_90_SUMB_21__5_), .A2(
        mul_ex_mult_90_CARRYB_21__4_), .ZN(mul_ex_mult_90_n98) );
  INV_X4 mul_ex_mult_90_U116 ( .A(mul_ex_mult_90_n97), .ZN(
        mul_ex_mult_90_SUMB_22__5_) );
  XNOR2_X2 mul_ex_mult_90_U115 ( .A(mul_ex_mult_90_CARRYB_21__5_), .B(
        mul_ex_mult_90_SUMB_21__6_), .ZN(mul_ex_mult_90_n97) );
  INV_X4 mul_ex_mult_90_U114 ( .A(mul_ex_mult_90_n96), .ZN(
        mul_ex_mult_90_CARRYB_22__5_) );
  NAND2_X2 mul_ex_mult_90_U113 ( .A1(mul_ex_mult_90_SUMB_21__6_), .A2(
        mul_ex_mult_90_CARRYB_21__5_), .ZN(mul_ex_mult_90_n96) );
  INV_X4 mul_ex_mult_90_U112 ( .A(mul_ex_mult_90_n95), .ZN(
        mul_ex_mult_90_SUMB_22__6_) );
  XNOR2_X2 mul_ex_mult_90_U111 ( .A(mul_ex_mult_90_CARRYB_21__6_), .B(
        mul_ex_mult_90_SUMB_21__7_), .ZN(mul_ex_mult_90_n95) );
  INV_X4 mul_ex_mult_90_U110 ( .A(mul_ex_mult_90_n94), .ZN(
        mul_ex_mult_90_CARRYB_22__6_) );
  NAND2_X2 mul_ex_mult_90_U109 ( .A1(mul_ex_mult_90_SUMB_21__7_), .A2(
        mul_ex_mult_90_CARRYB_21__6_), .ZN(mul_ex_mult_90_n94) );
  INV_X4 mul_ex_mult_90_U108 ( .A(mul_ex_mult_90_n93), .ZN(
        mul_ex_mult_90_SUMB_22__7_) );
  XNOR2_X2 mul_ex_mult_90_U107 ( .A(mul_ex_mult_90_CARRYB_21__7_), .B(
        mul_ex_mult_90_SUMB_21__8_), .ZN(mul_ex_mult_90_n93) );
  INV_X4 mul_ex_mult_90_U106 ( .A(mul_ex_mult_90_n92), .ZN(
        mul_ex_mult_90_CARRYB_22__7_) );
  NAND2_X2 mul_ex_mult_90_U105 ( .A1(mul_ex_mult_90_SUMB_21__8_), .A2(
        mul_ex_mult_90_CARRYB_21__7_), .ZN(mul_ex_mult_90_n92) );
  INV_X4 mul_ex_mult_90_U104 ( .A(mul_ex_mult_90_n91), .ZN(
        mul_ex_mult_90_SUMB_22__8_) );
  XNOR2_X2 mul_ex_mult_90_U103 ( .A(mul_ex_mult_90_CARRYB_21__8_), .B(
        mul_ex_mult_90_SUMB_21__9_), .ZN(mul_ex_mult_90_n91) );
  INV_X4 mul_ex_mult_90_U102 ( .A(mul_ex_mult_90_n90), .ZN(
        mul_ex_mult_90_CARRYB_22__8_) );
  NAND2_X2 mul_ex_mult_90_U101 ( .A1(mul_ex_mult_90_SUMB_21__9_), .A2(
        mul_ex_mult_90_CARRYB_21__8_), .ZN(mul_ex_mult_90_n90) );
  NOR2_X1 mul_ex_mult_90_U496 ( .A1(mul_ex_mult_90_n54), .A2(
        mul_ex_mult_90_n59), .ZN(mul_ex_N154) );
  NOR2_X1 mul_ex_mult_90_U495 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n89), .ZN(mul_ex_mult_90_ab_0__10_) );
  NOR2_X1 mul_ex_mult_90_U494 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n89), .ZN(mul_ex_mult_90_ab_0__11_) );
  NOR2_X1 mul_ex_mult_90_U493 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n89), .ZN(mul_ex_mult_90_ab_0__12_) );
  NOR2_X1 mul_ex_mult_90_U492 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n89), .ZN(mul_ex_mult_90_ab_0__13_) );
  NOR2_X1 mul_ex_mult_90_U491 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n89), .ZN(mul_ex_mult_90_ab_0__14_) );
  NOR2_X1 mul_ex_mult_90_U490 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n89), .ZN(mul_ex_mult_90_ab_0__15_) );
  NOR2_X1 mul_ex_mult_90_U489 ( .A1(mul_ex_mult_90_n60), .A2(
        mul_ex_mult_90_n89), .ZN(mul_ex_mult_90_ab_0__16_) );
  NOR2_X1 mul_ex_mult_90_U488 ( .A1(mul_ex_mult_90_n53), .A2(
        mul_ex_mult_90_n89), .ZN(mul_ex_mult_90_ab_0__1_) );
  NOR2_X1 mul_ex_mult_90_U487 ( .A1(mul_ex_mult_90_n52), .A2(
        mul_ex_mult_90_n59), .ZN(mul_ex_mult_90_ab_0__2_) );
  NOR2_X1 mul_ex_mult_90_U486 ( .A1(mul_ex_mult_90_n50), .A2(
        mul_ex_mult_90_n59), .ZN(mul_ex_mult_90_ab_0__3_) );
  NOR2_X1 mul_ex_mult_90_U485 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n59), .ZN(mul_ex_mult_90_ab_0__4_) );
  NOR2_X1 mul_ex_mult_90_U484 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n59), .ZN(mul_ex_mult_90_ab_0__5_) );
  NOR2_X1 mul_ex_mult_90_U483 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n59), .ZN(mul_ex_mult_90_ab_0__6_) );
  NOR2_X1 mul_ex_mult_90_U482 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n59), .ZN(mul_ex_mult_90_ab_0__7_) );
  NOR2_X1 mul_ex_mult_90_U481 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n59), .ZN(mul_ex_mult_90_ab_0__8_) );
  NOR2_X1 mul_ex_mult_90_U480 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n59), .ZN(mul_ex_mult_90_ab_0__9_) );
  NOR2_X1 mul_ex_mult_90_U479 ( .A1(mul_ex_mult_90_n54), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__0_) );
  NOR2_X1 mul_ex_mult_90_U478 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__10_) );
  NOR2_X1 mul_ex_mult_90_U477 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__11_) );
  NOR2_X1 mul_ex_mult_90_U476 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__12_) );
  NOR2_X1 mul_ex_mult_90_U475 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__13_) );
  NOR2_X1 mul_ex_mult_90_U474 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__14_) );
  NOR2_X1 mul_ex_mult_90_U473 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__15_) );
  NOR2_X1 mul_ex_mult_90_U472 ( .A1(mul_ex_mult_90_n60), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_SUMB_10__16_) );
  NOR2_X1 mul_ex_mult_90_U471 ( .A1(mul_ex_mult_90_n53), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__1_) );
  NOR2_X1 mul_ex_mult_90_U470 ( .A1(mul_ex_mult_90_n73), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__2_) );
  NOR2_X1 mul_ex_mult_90_U469 ( .A1(mul_ex_mult_90_n50), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__3_) );
  NOR2_X1 mul_ex_mult_90_U468 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__4_) );
  NOR2_X1 mul_ex_mult_90_U467 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__5_) );
  NOR2_X1 mul_ex_mult_90_U466 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__6_) );
  NOR2_X1 mul_ex_mult_90_U465 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__7_) );
  NOR2_X1 mul_ex_mult_90_U464 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__8_) );
  NOR2_X1 mul_ex_mult_90_U463 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n81), .ZN(mul_ex_mult_90_ab_10__9_) );
  NOR2_X1 mul_ex_mult_90_U462 ( .A1(mul_ex_mult_90_n54), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__0_) );
  NOR2_X1 mul_ex_mult_90_U461 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__10_) );
  NOR2_X1 mul_ex_mult_90_U460 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__11_) );
  NOR2_X1 mul_ex_mult_90_U459 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__12_) );
  NOR2_X1 mul_ex_mult_90_U458 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__13_) );
  NOR2_X1 mul_ex_mult_90_U457 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__14_) );
  NOR2_X1 mul_ex_mult_90_U456 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__15_) );
  NOR2_X1 mul_ex_mult_90_U455 ( .A1(mul_ex_mult_90_n60), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_SUMB_11__16_) );
  NOR2_X1 mul_ex_mult_90_U454 ( .A1(mul_ex_mult_90_n53), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__1_) );
  NOR2_X1 mul_ex_mult_90_U453 ( .A1(mul_ex_mult_90_n73), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__2_) );
  NOR2_X1 mul_ex_mult_90_U452 ( .A1(mul_ex_mult_90_n50), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__3_) );
  NOR2_X1 mul_ex_mult_90_U451 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__4_) );
  NOR2_X1 mul_ex_mult_90_U450 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__5_) );
  NOR2_X1 mul_ex_mult_90_U449 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__6_) );
  NOR2_X1 mul_ex_mult_90_U448 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__7_) );
  NOR2_X1 mul_ex_mult_90_U447 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__8_) );
  NOR2_X1 mul_ex_mult_90_U446 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n80), .ZN(mul_ex_mult_90_ab_11__9_) );
  NOR2_X1 mul_ex_mult_90_U445 ( .A1(mul_ex_mult_90_n54), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__0_) );
  NOR2_X1 mul_ex_mult_90_U444 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__10_) );
  NOR2_X1 mul_ex_mult_90_U443 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__11_) );
  NOR2_X1 mul_ex_mult_90_U442 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__12_) );
  NOR2_X1 mul_ex_mult_90_U441 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__13_) );
  NOR2_X1 mul_ex_mult_90_U440 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__14_) );
  NOR2_X1 mul_ex_mult_90_U439 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__15_) );
  NOR2_X1 mul_ex_mult_90_U438 ( .A1(mul_ex_mult_90_n60), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_SUMB_12__16_) );
  NOR2_X1 mul_ex_mult_90_U437 ( .A1(mul_ex_mult_90_n53), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__1_) );
  NOR2_X1 mul_ex_mult_90_U436 ( .A1(mul_ex_mult_90_n73), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__2_) );
  NOR2_X1 mul_ex_mult_90_U435 ( .A1(mul_ex_mult_90_n50), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__3_) );
  NOR2_X1 mul_ex_mult_90_U434 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__4_) );
  NOR2_X1 mul_ex_mult_90_U433 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__5_) );
  NOR2_X1 mul_ex_mult_90_U432 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__6_) );
  NOR2_X1 mul_ex_mult_90_U431 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__7_) );
  NOR2_X1 mul_ex_mult_90_U430 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__8_) );
  NOR2_X1 mul_ex_mult_90_U429 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n79), .ZN(mul_ex_mult_90_ab_12__9_) );
  NOR2_X1 mul_ex_mult_90_U428 ( .A1(mul_ex_mult_90_n54), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__0_) );
  NOR2_X1 mul_ex_mult_90_U427 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__10_) );
  NOR2_X1 mul_ex_mult_90_U426 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__11_) );
  NOR2_X1 mul_ex_mult_90_U425 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__12_) );
  NOR2_X1 mul_ex_mult_90_U424 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__13_) );
  NOR2_X1 mul_ex_mult_90_U423 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__14_) );
  NOR2_X1 mul_ex_mult_90_U422 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__15_) );
  NOR2_X1 mul_ex_mult_90_U421 ( .A1(mul_ex_mult_90_n60), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_SUMB_13__16_) );
  NOR2_X1 mul_ex_mult_90_U420 ( .A1(mul_ex_mult_90_n53), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__1_) );
  NOR2_X1 mul_ex_mult_90_U419 ( .A1(mul_ex_mult_90_n73), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__2_) );
  NOR2_X1 mul_ex_mult_90_U418 ( .A1(mul_ex_mult_90_n50), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__3_) );
  NOR2_X1 mul_ex_mult_90_U417 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__4_) );
  NOR2_X1 mul_ex_mult_90_U416 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__5_) );
  NOR2_X1 mul_ex_mult_90_U415 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__6_) );
  NOR2_X1 mul_ex_mult_90_U414 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__7_) );
  NOR2_X1 mul_ex_mult_90_U413 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__8_) );
  NOR2_X1 mul_ex_mult_90_U412 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n78), .ZN(mul_ex_mult_90_ab_13__9_) );
  NOR2_X1 mul_ex_mult_90_U411 ( .A1(mul_ex_mult_90_n54), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__0_) );
  NOR2_X1 mul_ex_mult_90_U410 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__10_) );
  NOR2_X1 mul_ex_mult_90_U409 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__11_) );
  NOR2_X1 mul_ex_mult_90_U408 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__12_) );
  NOR2_X1 mul_ex_mult_90_U407 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__13_) );
  NOR2_X1 mul_ex_mult_90_U406 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__14_) );
  NOR2_X1 mul_ex_mult_90_U405 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__15_) );
  NOR2_X1 mul_ex_mult_90_U404 ( .A1(mul_ex_mult_90_n60), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_SUMB_14__16_) );
  NOR2_X1 mul_ex_mult_90_U403 ( .A1(mul_ex_mult_90_n53), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__1_) );
  NOR2_X1 mul_ex_mult_90_U402 ( .A1(mul_ex_mult_90_n73), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__2_) );
  NOR2_X1 mul_ex_mult_90_U401 ( .A1(mul_ex_mult_90_n50), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__3_) );
  NOR2_X1 mul_ex_mult_90_U400 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__4_) );
  NOR2_X1 mul_ex_mult_90_U399 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__5_) );
  NOR2_X1 mul_ex_mult_90_U398 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__6_) );
  NOR2_X1 mul_ex_mult_90_U397 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__7_) );
  NOR2_X1 mul_ex_mult_90_U396 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__8_) );
  NOR2_X1 mul_ex_mult_90_U395 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n77), .ZN(mul_ex_mult_90_ab_14__9_) );
  NOR2_X1 mul_ex_mult_90_U394 ( .A1(mul_ex_mult_90_n54), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__0_) );
  NOR2_X1 mul_ex_mult_90_U393 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__10_) );
  NOR2_X1 mul_ex_mult_90_U392 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__11_) );
  NOR2_X1 mul_ex_mult_90_U391 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__12_) );
  NOR2_X1 mul_ex_mult_90_U390 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__13_) );
  NOR2_X1 mul_ex_mult_90_U389 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__14_) );
  NOR2_X1 mul_ex_mult_90_U388 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__15_) );
  NOR2_X1 mul_ex_mult_90_U387 ( .A1(mul_ex_mult_90_n60), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_SUMB_15__16_) );
  NOR2_X1 mul_ex_mult_90_U386 ( .A1(mul_ex_mult_90_n53), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__1_) );
  NOR2_X1 mul_ex_mult_90_U385 ( .A1(mul_ex_mult_90_n73), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__2_) );
  NOR2_X1 mul_ex_mult_90_U384 ( .A1(mul_ex_mult_90_n50), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__3_) );
  NOR2_X1 mul_ex_mult_90_U383 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__4_) );
  NOR2_X1 mul_ex_mult_90_U382 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__5_) );
  NOR2_X1 mul_ex_mult_90_U381 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__6_) );
  NOR2_X1 mul_ex_mult_90_U380 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__7_) );
  NOR2_X1 mul_ex_mult_90_U379 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__8_) );
  NOR2_X1 mul_ex_mult_90_U378 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n76), .ZN(mul_ex_mult_90_ab_15__9_) );
  NOR2_X1 mul_ex_mult_90_U377 ( .A1(mul_ex_mult_90_n54), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__0_) );
  NOR2_X1 mul_ex_mult_90_U376 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__10_) );
  NOR2_X1 mul_ex_mult_90_U375 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__11_) );
  NOR2_X1 mul_ex_mult_90_U374 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__12_) );
  NOR2_X1 mul_ex_mult_90_U373 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__13_) );
  NOR2_X1 mul_ex_mult_90_U372 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__14_) );
  NOR2_X1 mul_ex_mult_90_U371 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__15_) );
  NOR2_X1 mul_ex_mult_90_U370 ( .A1(mul_ex_mult_90_n53), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__1_) );
  NOR2_X1 mul_ex_mult_90_U369 ( .A1(mul_ex_mult_90_n73), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__2_) );
  NOR2_X1 mul_ex_mult_90_U368 ( .A1(mul_ex_mult_90_n50), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__3_) );
  NOR2_X1 mul_ex_mult_90_U367 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__4_) );
  NOR2_X1 mul_ex_mult_90_U366 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__5_) );
  NOR2_X1 mul_ex_mult_90_U365 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__6_) );
  NOR2_X1 mul_ex_mult_90_U364 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__7_) );
  NOR2_X1 mul_ex_mult_90_U363 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__8_) );
  NOR2_X1 mul_ex_mult_90_U362 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n75), .ZN(mul_ex_mult_90_ab_16__9_) );
  NOR2_X1 mul_ex_mult_90_U361 ( .A1(mul_ex_mult_90_n74), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__0_) );
  NOR2_X1 mul_ex_mult_90_U360 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__10_) );
  NOR2_X1 mul_ex_mult_90_U359 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__11_) );
  NOR2_X1 mul_ex_mult_90_U358 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__12_) );
  NOR2_X1 mul_ex_mult_90_U357 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__13_) );
  NOR2_X1 mul_ex_mult_90_U356 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__14_) );
  NOR2_X1 mul_ex_mult_90_U355 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__15_) );
  NOR2_X1 mul_ex_mult_90_U354 ( .A1(mul_ex_mult_90_n60), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__16_) );
  NOR2_X1 mul_ex_mult_90_U353 ( .A1(mul_ex_mult_90_n73), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__2_) );
  NOR2_X1 mul_ex_mult_90_U352 ( .A1(mul_ex_mult_90_n51), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__3_) );
  NOR2_X1 mul_ex_mult_90_U351 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__4_) );
  NOR2_X1 mul_ex_mult_90_U350 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__5_) );
  NOR2_X1 mul_ex_mult_90_U349 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__6_) );
  NOR2_X1 mul_ex_mult_90_U348 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__7_) );
  NOR2_X1 mul_ex_mult_90_U347 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__8_) );
  NOR2_X1 mul_ex_mult_90_U346 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n58), .ZN(mul_ex_mult_90_ab_1__9_) );
  NOR2_X1 mul_ex_mult_90_U345 ( .A1(mul_ex_mult_90_n74), .A2(
        mul_ex_mult_90_n57), .ZN(mul_ex_mult_90_ab_2__0_) );
  NOR2_X1 mul_ex_mult_90_U344 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n88), .ZN(mul_ex_mult_90_ab_2__10_) );
  NOR2_X1 mul_ex_mult_90_U343 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n88), .ZN(mul_ex_mult_90_ab_2__11_) );
  NOR2_X1 mul_ex_mult_90_U342 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n88), .ZN(mul_ex_mult_90_ab_2__12_) );
  NOR2_X1 mul_ex_mult_90_U341 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n88), .ZN(mul_ex_mult_90_ab_2__13_) );
  NOR2_X1 mul_ex_mult_90_U340 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n88), .ZN(mul_ex_mult_90_ab_2__14_) );
  NOR2_X1 mul_ex_mult_90_U339 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n88), .ZN(mul_ex_mult_90_ab_2__15_) );
  NOR2_X1 mul_ex_mult_90_U338 ( .A1(mul_ex_mult_90_n60), .A2(
        mul_ex_mult_90_n88), .ZN(mul_ex_mult_90_SUMB_2__16_) );
  NOR2_X1 mul_ex_mult_90_U337 ( .A1(mul_ex_mult_90_n53), .A2(
        mul_ex_mult_90_n88), .ZN(mul_ex_mult_90_ab_2__1_) );
  NOR2_X1 mul_ex_mult_90_U336 ( .A1(mul_ex_mult_90_n52), .A2(
        mul_ex_mult_90_n57), .ZN(mul_ex_mult_90_ab_2__2_) );
  NOR2_X1 mul_ex_mult_90_U335 ( .A1(mul_ex_mult_90_n51), .A2(
        mul_ex_mult_90_n57), .ZN(mul_ex_mult_90_ab_2__3_) );
  NOR2_X1 mul_ex_mult_90_U334 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n57), .ZN(mul_ex_mult_90_ab_2__4_) );
  NOR2_X1 mul_ex_mult_90_U333 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n57), .ZN(mul_ex_mult_90_ab_2__5_) );
  NOR2_X1 mul_ex_mult_90_U332 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n57), .ZN(mul_ex_mult_90_ab_2__6_) );
  NOR2_X1 mul_ex_mult_90_U331 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n57), .ZN(mul_ex_mult_90_ab_2__7_) );
  NOR2_X1 mul_ex_mult_90_U330 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n57), .ZN(mul_ex_mult_90_ab_2__8_) );
  NOR2_X1 mul_ex_mult_90_U329 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n57), .ZN(mul_ex_mult_90_ab_2__9_) );
  NOR2_X1 mul_ex_mult_90_U328 ( .A1(mul_ex_mult_90_n74), .A2(
        mul_ex_mult_90_n55), .ZN(mul_ex_mult_90_ab_3__0_) );
  NOR2_X1 mul_ex_mult_90_U327 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n55), .ZN(mul_ex_mult_90_ab_3__10_) );
  NOR2_X1 mul_ex_mult_90_U326 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n55), .ZN(mul_ex_mult_90_ab_3__11_) );
  NOR2_X1 mul_ex_mult_90_U325 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n55), .ZN(mul_ex_mult_90_ab_3__12_) );
  NOR2_X1 mul_ex_mult_90_U324 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n55), .ZN(mul_ex_mult_90_ab_3__13_) );
  NOR2_X1 mul_ex_mult_90_U323 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n55), .ZN(mul_ex_mult_90_ab_3__14_) );
  NOR2_X1 mul_ex_mult_90_U322 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n55), .ZN(mul_ex_mult_90_ab_3__15_) );
  NOR2_X1 mul_ex_mult_90_U321 ( .A1(mul_ex_mult_90_n60), .A2(
        mul_ex_mult_90_n55), .ZN(mul_ex_mult_90_SUMB_3__16_) );
  NOR2_X1 mul_ex_mult_90_U320 ( .A1(mul_ex_mult_90_n53), .A2(
        mul_ex_mult_90_n55), .ZN(mul_ex_mult_90_ab_3__1_) );
  NOR2_X1 mul_ex_mult_90_U319 ( .A1(mul_ex_mult_90_n52), .A2(
        mul_ex_mult_90_n56), .ZN(mul_ex_mult_90_ab_3__2_) );
  NOR2_X1 mul_ex_mult_90_U318 ( .A1(mul_ex_mult_90_n51), .A2(
        mul_ex_mult_90_n56), .ZN(mul_ex_mult_90_ab_3__3_) );
  NOR2_X1 mul_ex_mult_90_U317 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n56), .ZN(mul_ex_mult_90_ab_3__4_) );
  NOR2_X1 mul_ex_mult_90_U316 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n56), .ZN(mul_ex_mult_90_ab_3__5_) );
  NOR2_X1 mul_ex_mult_90_U315 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n56), .ZN(mul_ex_mult_90_ab_3__6_) );
  NOR2_X1 mul_ex_mult_90_U314 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n56), .ZN(mul_ex_mult_90_ab_3__7_) );
  NOR2_X1 mul_ex_mult_90_U313 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n56), .ZN(mul_ex_mult_90_ab_3__8_) );
  NOR2_X1 mul_ex_mult_90_U312 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n56), .ZN(mul_ex_mult_90_ab_3__9_) );
  NOR2_X1 mul_ex_mult_90_U311 ( .A1(mul_ex_mult_90_n74), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__0_) );
  NOR2_X1 mul_ex_mult_90_U310 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__10_) );
  NOR2_X1 mul_ex_mult_90_U309 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__11_) );
  NOR2_X1 mul_ex_mult_90_U308 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__12_) );
  NOR2_X1 mul_ex_mult_90_U307 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__13_) );
  NOR2_X1 mul_ex_mult_90_U306 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__14_) );
  NOR2_X1 mul_ex_mult_90_U305 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__15_) );
  NOR2_X1 mul_ex_mult_90_U304 ( .A1(mul_ex_mult_90_n60), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_SUMB_4__16_) );
  NOR2_X1 mul_ex_mult_90_U303 ( .A1(mul_ex_mult_90_n53), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__1_) );
  NOR2_X1 mul_ex_mult_90_U302 ( .A1(mul_ex_mult_90_n52), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__2_) );
  NOR2_X1 mul_ex_mult_90_U301 ( .A1(mul_ex_mult_90_n51), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__3_) );
  NOR2_X1 mul_ex_mult_90_U300 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__4_) );
  NOR2_X1 mul_ex_mult_90_U299 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__5_) );
  NOR2_X1 mul_ex_mult_90_U298 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__6_) );
  NOR2_X1 mul_ex_mult_90_U297 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__7_) );
  NOR2_X1 mul_ex_mult_90_U296 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__8_) );
  NOR2_X1 mul_ex_mult_90_U295 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n87), .ZN(mul_ex_mult_90_ab_4__9_) );
  NOR2_X1 mul_ex_mult_90_U294 ( .A1(mul_ex_mult_90_n74), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__0_) );
  NOR2_X1 mul_ex_mult_90_U293 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__10_) );
  NOR2_X1 mul_ex_mult_90_U292 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__11_) );
  NOR2_X1 mul_ex_mult_90_U291 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__12_) );
  NOR2_X1 mul_ex_mult_90_U290 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__13_) );
  NOR2_X1 mul_ex_mult_90_U289 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__14_) );
  NOR2_X1 mul_ex_mult_90_U288 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__15_) );
  NOR2_X1 mul_ex_mult_90_U287 ( .A1(mul_ex_mult_90_n60), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_SUMB_5__16_) );
  NOR2_X1 mul_ex_mult_90_U286 ( .A1(mul_ex_mult_90_n53), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__1_) );
  NOR2_X1 mul_ex_mult_90_U285 ( .A1(mul_ex_mult_90_n52), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__2_) );
  NOR2_X1 mul_ex_mult_90_U284 ( .A1(mul_ex_mult_90_n51), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__3_) );
  NOR2_X1 mul_ex_mult_90_U283 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__4_) );
  NOR2_X1 mul_ex_mult_90_U282 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__5_) );
  NOR2_X1 mul_ex_mult_90_U281 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__6_) );
  NOR2_X1 mul_ex_mult_90_U280 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__7_) );
  NOR2_X1 mul_ex_mult_90_U279 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__8_) );
  NOR2_X1 mul_ex_mult_90_U278 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n86), .ZN(mul_ex_mult_90_ab_5__9_) );
  NOR2_X1 mul_ex_mult_90_U277 ( .A1(mul_ex_mult_90_n74), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__0_) );
  NOR2_X1 mul_ex_mult_90_U276 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__10_) );
  NOR2_X1 mul_ex_mult_90_U275 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__11_) );
  NOR2_X1 mul_ex_mult_90_U274 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__12_) );
  NOR2_X1 mul_ex_mult_90_U273 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__13_) );
  NOR2_X1 mul_ex_mult_90_U272 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__14_) );
  NOR2_X1 mul_ex_mult_90_U271 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__15_) );
  NOR2_X1 mul_ex_mult_90_U270 ( .A1(mul_ex_mult_90_n60), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_SUMB_6__16_) );
  NOR2_X1 mul_ex_mult_90_U269 ( .A1(mul_ex_mult_90_n53), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__1_) );
  NOR2_X1 mul_ex_mult_90_U268 ( .A1(mul_ex_mult_90_n52), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__2_) );
  NOR2_X1 mul_ex_mult_90_U267 ( .A1(mul_ex_mult_90_n51), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__3_) );
  NOR2_X1 mul_ex_mult_90_U266 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__4_) );
  NOR2_X1 mul_ex_mult_90_U265 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__5_) );
  NOR2_X1 mul_ex_mult_90_U264 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__6_) );
  NOR2_X1 mul_ex_mult_90_U263 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__7_) );
  NOR2_X1 mul_ex_mult_90_U262 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__8_) );
  NOR2_X1 mul_ex_mult_90_U261 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n85), .ZN(mul_ex_mult_90_ab_6__9_) );
  NOR2_X1 mul_ex_mult_90_U260 ( .A1(mul_ex_mult_90_n74), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__0_) );
  NOR2_X1 mul_ex_mult_90_U259 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__10_) );
  NOR2_X1 mul_ex_mult_90_U258 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__11_) );
  NOR2_X1 mul_ex_mult_90_U257 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__12_) );
  NOR2_X1 mul_ex_mult_90_U256 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__13_) );
  NOR2_X1 mul_ex_mult_90_U255 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__14_) );
  NOR2_X1 mul_ex_mult_90_U254 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__15_) );
  NOR2_X1 mul_ex_mult_90_U253 ( .A1(mul_ex_mult_90_n60), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_SUMB_7__16_) );
  NOR2_X1 mul_ex_mult_90_U252 ( .A1(mul_ex_mult_90_n53), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__1_) );
  NOR2_X1 mul_ex_mult_90_U251 ( .A1(mul_ex_mult_90_n52), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__2_) );
  NOR2_X1 mul_ex_mult_90_U250 ( .A1(mul_ex_mult_90_n51), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__3_) );
  NOR2_X1 mul_ex_mult_90_U249 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__4_) );
  NOR2_X1 mul_ex_mult_90_U248 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__5_) );
  NOR2_X1 mul_ex_mult_90_U247 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__6_) );
  NOR2_X1 mul_ex_mult_90_U246 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__7_) );
  NOR2_X1 mul_ex_mult_90_U245 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__8_) );
  NOR2_X1 mul_ex_mult_90_U244 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n84), .ZN(mul_ex_mult_90_ab_7__9_) );
  NOR2_X1 mul_ex_mult_90_U243 ( .A1(mul_ex_mult_90_n74), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__0_) );
  NOR2_X1 mul_ex_mult_90_U242 ( .A1(mul_ex_mult_90_n66), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__10_) );
  NOR2_X1 mul_ex_mult_90_U241 ( .A1(mul_ex_mult_90_n65), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__11_) );
  NOR2_X1 mul_ex_mult_90_U240 ( .A1(mul_ex_mult_90_n64), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__12_) );
  NOR2_X1 mul_ex_mult_90_U239 ( .A1(mul_ex_mult_90_n63), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__13_) );
  NOR2_X1 mul_ex_mult_90_U238 ( .A1(mul_ex_mult_90_n62), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__14_) );
  NOR2_X1 mul_ex_mult_90_U237 ( .A1(mul_ex_mult_90_n61), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__15_) );
  NOR2_X1 mul_ex_mult_90_U236 ( .A1(mul_ex_mult_90_n60), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_SUMB_8__16_) );
  NOR2_X1 mul_ex_mult_90_U235 ( .A1(mul_ex_mult_90_n53), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__1_) );
  NOR2_X1 mul_ex_mult_90_U234 ( .A1(mul_ex_mult_90_n52), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__2_) );
  NOR2_X1 mul_ex_mult_90_U233 ( .A1(mul_ex_mult_90_n51), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__3_) );
  NOR2_X1 mul_ex_mult_90_U232 ( .A1(mul_ex_mult_90_n72), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__4_) );
  NOR2_X1 mul_ex_mult_90_U231 ( .A1(mul_ex_mult_90_n71), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__5_) );
  NOR2_X1 mul_ex_mult_90_U230 ( .A1(mul_ex_mult_90_n70), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__6_) );
  NOR2_X1 mul_ex_mult_90_U229 ( .A1(mul_ex_mult_90_n69), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__7_) );
  NOR2_X1 mul_ex_mult_90_U228 ( .A1(mul_ex_mult_90_n68), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__8_) );
  NOR2_X1 mul_ex_mult_90_U227 ( .A1(mul_ex_mult_90_n67), .A2(
        mul_ex_mult_90_n83), .ZN(mul_ex_mult_90_ab_8__9_) );
  NOR2_X1 mul_ex_mult_90_U226 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n54), .ZN(mul_ex_mult_90_ab_9__0_) );
  NOR2_X1 mul_ex_mult_90_U225 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n66), .ZN(mul_ex_mult_90_ab_9__10_) );
  NOR2_X1 mul_ex_mult_90_U224 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n65), .ZN(mul_ex_mult_90_ab_9__11_) );
  NOR2_X1 mul_ex_mult_90_U223 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n64), .ZN(mul_ex_mult_90_ab_9__12_) );
  NOR2_X1 mul_ex_mult_90_U222 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n63), .ZN(mul_ex_mult_90_ab_9__13_) );
  NOR2_X1 mul_ex_mult_90_U221 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n62), .ZN(mul_ex_mult_90_ab_9__14_) );
  NOR2_X1 mul_ex_mult_90_U220 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n61), .ZN(mul_ex_mult_90_ab_9__15_) );
  NOR2_X1 mul_ex_mult_90_U219 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n60), .ZN(mul_ex_mult_90_SUMB_9__16_) );
  NOR2_X1 mul_ex_mult_90_U218 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n53), .ZN(mul_ex_mult_90_ab_9__1_) );
  NOR2_X1 mul_ex_mult_90_U217 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n52), .ZN(mul_ex_mult_90_ab_9__2_) );
  NOR2_X1 mul_ex_mult_90_U216 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n51), .ZN(mul_ex_mult_90_ab_9__3_) );
  NOR2_X1 mul_ex_mult_90_U215 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n72), .ZN(mul_ex_mult_90_ab_9__4_) );
  NOR2_X1 mul_ex_mult_90_U214 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n71), .ZN(mul_ex_mult_90_ab_9__5_) );
  NOR2_X1 mul_ex_mult_90_U213 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n70), .ZN(mul_ex_mult_90_ab_9__6_) );
  NOR2_X1 mul_ex_mult_90_U212 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n69), .ZN(mul_ex_mult_90_ab_9__7_) );
  NOR2_X1 mul_ex_mult_90_U211 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n68), .ZN(mul_ex_mult_90_ab_9__8_) );
  NOR2_X1 mul_ex_mult_90_U210 ( .A1(mul_ex_mult_90_n82), .A2(
        mul_ex_mult_90_n67), .ZN(mul_ex_mult_90_ab_9__9_) );
  INV_X4 mul_ex_mult_90_U209 ( .A(mul_ex_P1[31]), .ZN(mul_ex_mult_90_n89) );
  INV_X4 mul_ex_mult_90_U208 ( .A(mul_ex_P1[29]), .ZN(mul_ex_mult_90_n88) );
  INV_X4 mul_ex_mult_90_U207 ( .A(mul_ex_P2[31]), .ZN(mul_ex_mult_90_n74) );
  INV_X4 mul_ex_mult_90_U206 ( .A(mul_ex_P2[29]), .ZN(mul_ex_mult_90_n73) );
  INV_X4 mul_ex_mult_90_U100 ( .A(mul_ex_P1[23]), .ZN(mul_ex_mult_90_n83) );
  INV_X4 mul_ex_mult_90_U99 ( .A(mul_ex_P1[24]), .ZN(mul_ex_mult_90_n84) );
  INV_X4 mul_ex_mult_90_U98 ( .A(mul_ex_P1[25]), .ZN(mul_ex_mult_90_n85) );
  INV_X4 mul_ex_mult_90_U97 ( .A(mul_ex_P1[26]), .ZN(mul_ex_mult_90_n86) );
  INV_X4 mul_ex_mult_90_U96 ( .A(mul_ex_P1[27]), .ZN(mul_ex_mult_90_n87) );
  INV_X4 mul_ex_mult_90_U95 ( .A(mul_ex_P2[21]), .ZN(mul_ex_mult_90_n66) );
  INV_X4 mul_ex_mult_90_U94 ( .A(mul_ex_P2[22]), .ZN(mul_ex_mult_90_n67) );
  INV_X4 mul_ex_mult_90_U93 ( .A(mul_ex_P2[23]), .ZN(mul_ex_mult_90_n68) );
  INV_X4 mul_ex_mult_90_U92 ( .A(mul_ex_P2[24]), .ZN(mul_ex_mult_90_n69) );
  INV_X4 mul_ex_mult_90_U91 ( .A(mul_ex_P2[25]), .ZN(mul_ex_mult_90_n70) );
  INV_X4 mul_ex_mult_90_U90 ( .A(mul_ex_P2[26]), .ZN(mul_ex_mult_90_n71) );
  INV_X4 mul_ex_mult_90_U89 ( .A(mul_ex_P2[27]), .ZN(mul_ex_mult_90_n72) );
  INV_X4 mul_ex_mult_90_U88 ( .A(mul_ex_P1[22]), .ZN(mul_ex_mult_90_n82) );
  INV_X4 mul_ex_mult_90_U87 ( .A(mul_ex_P1[15]), .ZN(mul_ex_mult_90_n75) );
  INV_X4 mul_ex_mult_90_U86 ( .A(mul_ex_P2[15]), .ZN(mul_ex_mult_90_n60) );
  INV_X4 mul_ex_mult_90_U85 ( .A(mul_ex_P1[16]), .ZN(mul_ex_mult_90_n76) );
  INV_X4 mul_ex_mult_90_U84 ( .A(mul_ex_P1[17]), .ZN(mul_ex_mult_90_n77) );
  INV_X4 mul_ex_mult_90_U83 ( .A(mul_ex_P1[18]), .ZN(mul_ex_mult_90_n78) );
  INV_X4 mul_ex_mult_90_U82 ( .A(mul_ex_P1[19]), .ZN(mul_ex_mult_90_n79) );
  INV_X4 mul_ex_mult_90_U81 ( .A(mul_ex_P1[20]), .ZN(mul_ex_mult_90_n80) );
  INV_X4 mul_ex_mult_90_U80 ( .A(mul_ex_P1[21]), .ZN(mul_ex_mult_90_n81) );
  INV_X4 mul_ex_mult_90_U79 ( .A(mul_ex_P2[16]), .ZN(mul_ex_mult_90_n61) );
  INV_X4 mul_ex_mult_90_U78 ( .A(mul_ex_P2[17]), .ZN(mul_ex_mult_90_n62) );
  INV_X4 mul_ex_mult_90_U77 ( .A(mul_ex_P2[18]), .ZN(mul_ex_mult_90_n63) );
  INV_X4 mul_ex_mult_90_U76 ( .A(mul_ex_P2[19]), .ZN(mul_ex_mult_90_n64) );
  INV_X4 mul_ex_mult_90_U75 ( .A(mul_ex_P2[20]), .ZN(mul_ex_mult_90_n65) );
  INV_X4 mul_ex_mult_90_U74 ( .A(mul_ex_P1[28]), .ZN(mul_ex_mult_90_n56) );
  INV_X4 mul_ex_mult_90_U73 ( .A(mul_ex_P2[28]), .ZN(mul_ex_mult_90_n51) );
  INV_X4 mul_ex_mult_90_U72 ( .A(mul_ex_P1[28]), .ZN(mul_ex_mult_90_n55) );
  INV_X4 mul_ex_mult_90_U71 ( .A(mul_ex_P1[29]), .ZN(mul_ex_mult_90_n57) );
  INV_X4 mul_ex_mult_90_U70 ( .A(mul_ex_P1[30]), .ZN(mul_ex_mult_90_n58) );
  INV_X4 mul_ex_mult_90_U69 ( .A(mul_ex_P1[31]), .ZN(mul_ex_mult_90_n59) );
  INV_X4 mul_ex_mult_90_U68 ( .A(mul_ex_P2[29]), .ZN(mul_ex_mult_90_n52) );
  INV_X4 mul_ex_mult_90_U67 ( .A(mul_ex_P2[30]), .ZN(mul_ex_mult_90_n53) );
  INV_X4 mul_ex_mult_90_U66 ( .A(mul_ex_P2[31]), .ZN(mul_ex_mult_90_n54) );
  INV_X4 mul_ex_mult_90_U65 ( .A(mul_ex_P2[28]), .ZN(mul_ex_mult_90_n50) );
  AND2_X2 mul_ex_mult_90_U64 ( .A1(mul_ex_P2[30]), .A2(mul_ex_P1[30]), .ZN(
        mul_ex_mult_90_ab_1__1_) );
  XOR2_X2 mul_ex_mult_90_U63 ( .A(mul_ex_mult_90_ab_1__0_), .B(
        mul_ex_mult_90_ab_0__1_), .Z(mul_ex_N155) );
  XOR2_X2 mul_ex_mult_90_U62 ( .A(mul_ex_mult_90_ab_1__1_), .B(
        mul_ex_mult_90_ab_0__2_), .Z(mul_ex_mult_90_n48) );
  XOR2_X2 mul_ex_mult_90_U61 ( .A(mul_ex_mult_90_ab_1__2_), .B(
        mul_ex_mult_90_ab_0__3_), .Z(mul_ex_mult_90_n47) );
  XOR2_X2 mul_ex_mult_90_U60 ( .A(mul_ex_mult_90_ab_1__3_), .B(
        mul_ex_mult_90_ab_0__4_), .Z(mul_ex_mult_90_n46) );
  XOR2_X2 mul_ex_mult_90_U59 ( .A(mul_ex_mult_90_ab_1__4_), .B(
        mul_ex_mult_90_ab_0__5_), .Z(mul_ex_mult_90_n45) );
  XOR2_X2 mul_ex_mult_90_U58 ( .A(mul_ex_mult_90_ab_1__5_), .B(
        mul_ex_mult_90_ab_0__6_), .Z(mul_ex_mult_90_n44) );
  XOR2_X2 mul_ex_mult_90_U57 ( .A(mul_ex_mult_90_ab_1__6_), .B(
        mul_ex_mult_90_ab_0__7_), .Z(mul_ex_mult_90_n43) );
  XOR2_X2 mul_ex_mult_90_U56 ( .A(mul_ex_mult_90_ab_1__7_), .B(
        mul_ex_mult_90_ab_0__8_), .Z(mul_ex_mult_90_n42) );
  XOR2_X2 mul_ex_mult_90_U55 ( .A(mul_ex_mult_90_ab_1__8_), .B(
        mul_ex_mult_90_ab_0__9_), .Z(mul_ex_mult_90_n41) );
  XOR2_X2 mul_ex_mult_90_U54 ( .A(mul_ex_mult_90_ab_1__9_), .B(
        mul_ex_mult_90_ab_0__10_), .Z(mul_ex_mult_90_n40) );
  XOR2_X2 mul_ex_mult_90_U53 ( .A(mul_ex_mult_90_ab_1__10_), .B(
        mul_ex_mult_90_ab_0__11_), .Z(mul_ex_mult_90_n39) );
  XOR2_X2 mul_ex_mult_90_U52 ( .A(mul_ex_mult_90_ab_1__11_), .B(
        mul_ex_mult_90_ab_0__12_), .Z(mul_ex_mult_90_n38) );
  XOR2_X2 mul_ex_mult_90_U51 ( .A(mul_ex_mult_90_ab_1__12_), .B(
        mul_ex_mult_90_ab_0__13_), .Z(mul_ex_mult_90_n37) );
  XOR2_X2 mul_ex_mult_90_U50 ( .A(mul_ex_mult_90_ab_1__13_), .B(
        mul_ex_mult_90_ab_0__14_), .Z(mul_ex_mult_90_n36) );
  XOR2_X2 mul_ex_mult_90_U49 ( .A(mul_ex_mult_90_ab_1__14_), .B(
        mul_ex_mult_90_ab_0__15_), .Z(mul_ex_mult_90_n35) );
  XOR2_X2 mul_ex_mult_90_U48 ( .A(mul_ex_mult_90_ab_1__15_), .B(
        mul_ex_mult_90_ab_0__16_), .Z(mul_ex_mult_90_n34) );
  AND2_X4 mul_ex_mult_90_U47 ( .A1(mul_ex_mult_90_ab_0__1_), .A2(
        mul_ex_mult_90_ab_1__0_), .ZN(mul_ex_mult_90_n33) );
  AND2_X4 mul_ex_mult_90_U46 ( .A1(mul_ex_mult_90_ab_0__2_), .A2(
        mul_ex_mult_90_ab_1__1_), .ZN(mul_ex_mult_90_n32) );
  AND2_X4 mul_ex_mult_90_U45 ( .A1(mul_ex_mult_90_ab_0__3_), .A2(
        mul_ex_mult_90_ab_1__2_), .ZN(mul_ex_mult_90_n31) );
  AND2_X4 mul_ex_mult_90_U44 ( .A1(mul_ex_mult_90_ab_0__4_), .A2(
        mul_ex_mult_90_ab_1__3_), .ZN(mul_ex_mult_90_n30) );
  AND2_X4 mul_ex_mult_90_U43 ( .A1(mul_ex_mult_90_ab_0__5_), .A2(
        mul_ex_mult_90_ab_1__4_), .ZN(mul_ex_mult_90_n29) );
  AND2_X4 mul_ex_mult_90_U42 ( .A1(mul_ex_mult_90_ab_0__6_), .A2(
        mul_ex_mult_90_ab_1__5_), .ZN(mul_ex_mult_90_n28) );
  AND2_X4 mul_ex_mult_90_U41 ( .A1(mul_ex_mult_90_ab_0__7_), .A2(
        mul_ex_mult_90_ab_1__6_), .ZN(mul_ex_mult_90_n27) );
  AND2_X4 mul_ex_mult_90_U40 ( .A1(mul_ex_mult_90_ab_0__8_), .A2(
        mul_ex_mult_90_ab_1__7_), .ZN(mul_ex_mult_90_n26) );
  AND2_X4 mul_ex_mult_90_U39 ( .A1(mul_ex_mult_90_ab_0__9_), .A2(
        mul_ex_mult_90_ab_1__8_), .ZN(mul_ex_mult_90_n25) );
  AND2_X4 mul_ex_mult_90_U38 ( .A1(mul_ex_mult_90_ab_0__10_), .A2(
        mul_ex_mult_90_ab_1__9_), .ZN(mul_ex_mult_90_n24) );
  AND2_X4 mul_ex_mult_90_U37 ( .A1(mul_ex_mult_90_ab_0__11_), .A2(
        mul_ex_mult_90_ab_1__10_), .ZN(mul_ex_mult_90_n23) );
  AND2_X4 mul_ex_mult_90_U36 ( .A1(mul_ex_mult_90_ab_0__12_), .A2(
        mul_ex_mult_90_ab_1__11_), .ZN(mul_ex_mult_90_n22) );
  AND2_X4 mul_ex_mult_90_U35 ( .A1(mul_ex_mult_90_ab_0__13_), .A2(
        mul_ex_mult_90_ab_1__12_), .ZN(mul_ex_mult_90_n21) );
  AND2_X4 mul_ex_mult_90_U34 ( .A1(mul_ex_mult_90_ab_0__14_), .A2(
        mul_ex_mult_90_ab_1__13_), .ZN(mul_ex_mult_90_n20) );
  AND2_X4 mul_ex_mult_90_U33 ( .A1(mul_ex_mult_90_ab_0__15_), .A2(
        mul_ex_mult_90_ab_1__14_), .ZN(mul_ex_mult_90_n19) );
  AND2_X4 mul_ex_mult_90_U32 ( .A1(mul_ex_mult_90_ab_0__16_), .A2(
        mul_ex_mult_90_ab_1__15_), .ZN(mul_ex_mult_90_n18) );
  INV_X4 mul_ex_mult_90_U31 ( .A(mul_ex_mult_90_n17), .ZN(
        mul_ex_mult_90_SUMB_22__9_) );
  XNOR2_X2 mul_ex_mult_90_U30 ( .A(mul_ex_mult_90_CARRYB_21__9_), .B(
        mul_ex_mult_90_SUMB_21__10_), .ZN(mul_ex_mult_90_n17) );
  INV_X4 mul_ex_mult_90_U29 ( .A(mul_ex_mult_90_n16), .ZN(
        mul_ex_mult_90_SUMB_23__8_) );
  XNOR2_X2 mul_ex_mult_90_U28 ( .A(mul_ex_mult_90_CARRYB_22__8_), .B(
        mul_ex_mult_90_SUMB_22__9_), .ZN(mul_ex_mult_90_n16) );
  INV_X4 mul_ex_mult_90_U27 ( .A(mul_ex_mult_90_n15), .ZN(
        mul_ex_mult_90_SUMB_24__7_) );
  XNOR2_X2 mul_ex_mult_90_U26 ( .A(mul_ex_mult_90_CARRYB_23__7_), .B(
        mul_ex_mult_90_SUMB_23__8_), .ZN(mul_ex_mult_90_n15) );
  INV_X4 mul_ex_mult_90_U25 ( .A(mul_ex_mult_90_n14), .ZN(
        mul_ex_mult_90_SUMB_25__6_) );
  XNOR2_X2 mul_ex_mult_90_U24 ( .A(mul_ex_mult_90_CARRYB_24__6_), .B(
        mul_ex_mult_90_SUMB_24__7_), .ZN(mul_ex_mult_90_n14) );
  INV_X4 mul_ex_mult_90_U23 ( .A(mul_ex_mult_90_n13), .ZN(
        mul_ex_mult_90_SUMB_26__5_) );
  XNOR2_X2 mul_ex_mult_90_U22 ( .A(mul_ex_mult_90_CARRYB_25__5_), .B(
        mul_ex_mult_90_SUMB_25__6_), .ZN(mul_ex_mult_90_n13) );
  INV_X4 mul_ex_mult_90_U21 ( .A(mul_ex_mult_90_n12), .ZN(
        mul_ex_mult_90_SUMB_27__4_) );
  XNOR2_X2 mul_ex_mult_90_U20 ( .A(mul_ex_mult_90_CARRYB_26__4_), .B(
        mul_ex_mult_90_SUMB_26__5_), .ZN(mul_ex_mult_90_n12) );
  INV_X4 mul_ex_mult_90_U19 ( .A(mul_ex_mult_90_n11), .ZN(
        mul_ex_mult_90_SUMB_28__3_) );
  XNOR2_X2 mul_ex_mult_90_U18 ( .A(mul_ex_mult_90_CARRYB_27__3_), .B(
        mul_ex_mult_90_SUMB_27__4_), .ZN(mul_ex_mult_90_n11) );
  INV_X4 mul_ex_mult_90_U17 ( .A(mul_ex_mult_90_n10), .ZN(
        mul_ex_mult_90_SUMB_29__2_) );
  XNOR2_X2 mul_ex_mult_90_U16 ( .A(mul_ex_mult_90_CARRYB_28__2_), .B(
        mul_ex_mult_90_SUMB_28__3_), .ZN(mul_ex_mult_90_n10) );
  INV_X4 mul_ex_mult_90_U15 ( .A(mul_ex_mult_90_n9), .ZN(
        mul_ex_mult_90_SUMB_30__1_) );
  XNOR2_X2 mul_ex_mult_90_U14 ( .A(mul_ex_mult_90_CARRYB_29__1_), .B(
        mul_ex_mult_90_SUMB_29__2_), .ZN(mul_ex_mult_90_n9) );
  INV_X4 mul_ex_mult_90_U13 ( .A(mul_ex_mult_90_n8), .ZN(
        mul_ex_mult_90_SUMB_17__14_) );
  XNOR2_X2 mul_ex_mult_90_U12 ( .A(mul_ex_mult_90_CARRYB_16__14_), .B(
        mul_ex_mult_90_SUMB_16__15_), .ZN(mul_ex_mult_90_n8) );
  INV_X4 mul_ex_mult_90_U11 ( .A(mul_ex_mult_90_n7), .ZN(
        mul_ex_mult_90_SUMB_18__13_) );
  XNOR2_X2 mul_ex_mult_90_U10 ( .A(mul_ex_mult_90_CARRYB_17__13_), .B(
        mul_ex_mult_90_SUMB_17__14_), .ZN(mul_ex_mult_90_n7) );
  INV_X4 mul_ex_mult_90_U9 ( .A(mul_ex_mult_90_n6), .ZN(
        mul_ex_mult_90_SUMB_19__12_) );
  XNOR2_X2 mul_ex_mult_90_U8 ( .A(mul_ex_mult_90_CARRYB_18__12_), .B(
        mul_ex_mult_90_SUMB_18__13_), .ZN(mul_ex_mult_90_n6) );
  INV_X4 mul_ex_mult_90_U7 ( .A(mul_ex_mult_90_n5), .ZN(
        mul_ex_mult_90_SUMB_20__11_) );
  XNOR2_X2 mul_ex_mult_90_U6 ( .A(mul_ex_mult_90_CARRYB_19__11_), .B(
        mul_ex_mult_90_SUMB_19__12_), .ZN(mul_ex_mult_90_n5) );
  INV_X4 mul_ex_mult_90_U5 ( .A(mul_ex_mult_90_n4), .ZN(
        mul_ex_mult_90_SUMB_21__10_) );
  XNOR2_X2 mul_ex_mult_90_U4 ( .A(mul_ex_mult_90_CARRYB_20__10_), .B(
        mul_ex_mult_90_SUMB_20__11_), .ZN(mul_ex_mult_90_n4) );
  INV_X4 mul_ex_mult_90_U3 ( .A(mul_ex_mult_90_n3), .ZN(mul_ex_N185) );
  XNOR2_X2 mul_ex_mult_90_U2 ( .A(mul_ex_mult_90_CARRYB_30__0_), .B(
        mul_ex_mult_90_SUMB_30__1_), .ZN(mul_ex_mult_90_n3) );
  FA_X1 mul_ex_mult_90_S2_2_15 ( .A(mul_ex_mult_90_ab_2__15_), .B(
        mul_ex_mult_90_n18), .CI(mul_ex_mult_90_ab_1__16_), .CO(
        mul_ex_mult_90_CARRYB_2__15_), .S(mul_ex_mult_90_SUMB_2__15_) );
  FA_X1 mul_ex_mult_90_S2_2_14 ( .A(mul_ex_mult_90_ab_2__14_), .B(
        mul_ex_mult_90_n19), .CI(mul_ex_mult_90_n34), .CO(
        mul_ex_mult_90_CARRYB_2__14_), .S(mul_ex_mult_90_SUMB_2__14_) );
  FA_X1 mul_ex_mult_90_S2_2_13 ( .A(mul_ex_mult_90_ab_2__13_), .B(
        mul_ex_mult_90_n20), .CI(mul_ex_mult_90_n35), .CO(
        mul_ex_mult_90_CARRYB_2__13_), .S(mul_ex_mult_90_SUMB_2__13_) );
  FA_X1 mul_ex_mult_90_S2_2_12 ( .A(mul_ex_mult_90_ab_2__12_), .B(
        mul_ex_mult_90_n21), .CI(mul_ex_mult_90_n36), .CO(
        mul_ex_mult_90_CARRYB_2__12_), .S(mul_ex_mult_90_SUMB_2__12_) );
  FA_X1 mul_ex_mult_90_S2_2_11 ( .A(mul_ex_mult_90_ab_2__11_), .B(
        mul_ex_mult_90_n22), .CI(mul_ex_mult_90_n37), .CO(
        mul_ex_mult_90_CARRYB_2__11_), .S(mul_ex_mult_90_SUMB_2__11_) );
  FA_X1 mul_ex_mult_90_S2_2_10 ( .A(mul_ex_mult_90_ab_2__10_), .B(
        mul_ex_mult_90_n23), .CI(mul_ex_mult_90_n38), .CO(
        mul_ex_mult_90_CARRYB_2__10_), .S(mul_ex_mult_90_SUMB_2__10_) );
  FA_X1 mul_ex_mult_90_S2_2_9 ( .A(mul_ex_mult_90_ab_2__9_), .B(
        mul_ex_mult_90_n24), .CI(mul_ex_mult_90_n39), .CO(
        mul_ex_mult_90_CARRYB_2__9_), .S(mul_ex_mult_90_SUMB_2__9_) );
  FA_X1 mul_ex_mult_90_S2_2_8 ( .A(mul_ex_mult_90_ab_2__8_), .B(
        mul_ex_mult_90_n25), .CI(mul_ex_mult_90_n40), .CO(
        mul_ex_mult_90_CARRYB_2__8_), .S(mul_ex_mult_90_SUMB_2__8_) );
  FA_X1 mul_ex_mult_90_S2_2_7 ( .A(mul_ex_mult_90_ab_2__7_), .B(
        mul_ex_mult_90_n26), .CI(mul_ex_mult_90_n41), .CO(
        mul_ex_mult_90_CARRYB_2__7_), .S(mul_ex_mult_90_SUMB_2__7_) );
  FA_X1 mul_ex_mult_90_S2_2_6 ( .A(mul_ex_mult_90_ab_2__6_), .B(
        mul_ex_mult_90_n27), .CI(mul_ex_mult_90_n42), .CO(
        mul_ex_mult_90_CARRYB_2__6_), .S(mul_ex_mult_90_SUMB_2__6_) );
  FA_X1 mul_ex_mult_90_S2_2_5 ( .A(mul_ex_mult_90_ab_2__5_), .B(
        mul_ex_mult_90_n28), .CI(mul_ex_mult_90_n43), .CO(
        mul_ex_mult_90_CARRYB_2__5_), .S(mul_ex_mult_90_SUMB_2__5_) );
  FA_X1 mul_ex_mult_90_S2_2_4 ( .A(mul_ex_mult_90_ab_2__4_), .B(
        mul_ex_mult_90_n29), .CI(mul_ex_mult_90_n44), .CO(
        mul_ex_mult_90_CARRYB_2__4_), .S(mul_ex_mult_90_SUMB_2__4_) );
  FA_X1 mul_ex_mult_90_S2_2_3 ( .A(mul_ex_mult_90_ab_2__3_), .B(
        mul_ex_mult_90_n30), .CI(mul_ex_mult_90_n45), .CO(
        mul_ex_mult_90_CARRYB_2__3_), .S(mul_ex_mult_90_SUMB_2__3_) );
  FA_X1 mul_ex_mult_90_S2_2_2 ( .A(mul_ex_mult_90_ab_2__2_), .B(
        mul_ex_mult_90_n31), .CI(mul_ex_mult_90_n46), .CO(
        mul_ex_mult_90_CARRYB_2__2_), .S(mul_ex_mult_90_SUMB_2__2_) );
  FA_X1 mul_ex_mult_90_S2_2_1 ( .A(mul_ex_mult_90_ab_2__1_), .B(
        mul_ex_mult_90_n32), .CI(mul_ex_mult_90_n47), .CO(
        mul_ex_mult_90_CARRYB_2__1_), .S(mul_ex_mult_90_SUMB_2__1_) );
  FA_X1 mul_ex_mult_90_S1_2_0 ( .A(mul_ex_mult_90_ab_2__0_), .B(
        mul_ex_mult_90_n33), .CI(mul_ex_mult_90_n48), .CO(
        mul_ex_mult_90_CARRYB_2__0_), .S(mul_ex_N156) );
  FA_X1 mul_ex_mult_90_S2_3_15 ( .A(mul_ex_mult_90_ab_3__15_), .B(
        mul_ex_mult_90_CARRYB_2__15_), .CI(mul_ex_mult_90_SUMB_2__16_), .CO(
        mul_ex_mult_90_CARRYB_3__15_), .S(mul_ex_mult_90_SUMB_3__15_) );
  FA_X1 mul_ex_mult_90_S2_3_14 ( .A(mul_ex_mult_90_ab_3__14_), .B(
        mul_ex_mult_90_CARRYB_2__14_), .CI(mul_ex_mult_90_SUMB_2__15_), .CO(
        mul_ex_mult_90_CARRYB_3__14_), .S(mul_ex_mult_90_SUMB_3__14_) );
  FA_X1 mul_ex_mult_90_S2_3_13 ( .A(mul_ex_mult_90_ab_3__13_), .B(
        mul_ex_mult_90_CARRYB_2__13_), .CI(mul_ex_mult_90_SUMB_2__14_), .CO(
        mul_ex_mult_90_CARRYB_3__13_), .S(mul_ex_mult_90_SUMB_3__13_) );
  FA_X1 mul_ex_mult_90_S2_3_12 ( .A(mul_ex_mult_90_ab_3__12_), .B(
        mul_ex_mult_90_CARRYB_2__12_), .CI(mul_ex_mult_90_SUMB_2__13_), .CO(
        mul_ex_mult_90_CARRYB_3__12_), .S(mul_ex_mult_90_SUMB_3__12_) );
  FA_X1 mul_ex_mult_90_S2_3_11 ( .A(mul_ex_mult_90_ab_3__11_), .B(
        mul_ex_mult_90_CARRYB_2__11_), .CI(mul_ex_mult_90_SUMB_2__12_), .CO(
        mul_ex_mult_90_CARRYB_3__11_), .S(mul_ex_mult_90_SUMB_3__11_) );
  FA_X1 mul_ex_mult_90_S2_3_10 ( .A(mul_ex_mult_90_ab_3__10_), .B(
        mul_ex_mult_90_CARRYB_2__10_), .CI(mul_ex_mult_90_SUMB_2__11_), .CO(
        mul_ex_mult_90_CARRYB_3__10_), .S(mul_ex_mult_90_SUMB_3__10_) );
  FA_X1 mul_ex_mult_90_S2_3_9 ( .A(mul_ex_mult_90_ab_3__9_), .B(
        mul_ex_mult_90_CARRYB_2__9_), .CI(mul_ex_mult_90_SUMB_2__10_), .CO(
        mul_ex_mult_90_CARRYB_3__9_), .S(mul_ex_mult_90_SUMB_3__9_) );
  FA_X1 mul_ex_mult_90_S2_3_8 ( .A(mul_ex_mult_90_ab_3__8_), .B(
        mul_ex_mult_90_CARRYB_2__8_), .CI(mul_ex_mult_90_SUMB_2__9_), .CO(
        mul_ex_mult_90_CARRYB_3__8_), .S(mul_ex_mult_90_SUMB_3__8_) );
  FA_X1 mul_ex_mult_90_S2_3_7 ( .A(mul_ex_mult_90_ab_3__7_), .B(
        mul_ex_mult_90_CARRYB_2__7_), .CI(mul_ex_mult_90_SUMB_2__8_), .CO(
        mul_ex_mult_90_CARRYB_3__7_), .S(mul_ex_mult_90_SUMB_3__7_) );
  FA_X1 mul_ex_mult_90_S2_3_6 ( .A(mul_ex_mult_90_ab_3__6_), .B(
        mul_ex_mult_90_CARRYB_2__6_), .CI(mul_ex_mult_90_SUMB_2__7_), .CO(
        mul_ex_mult_90_CARRYB_3__6_), .S(mul_ex_mult_90_SUMB_3__6_) );
  FA_X1 mul_ex_mult_90_S2_3_5 ( .A(mul_ex_mult_90_ab_3__5_), .B(
        mul_ex_mult_90_CARRYB_2__5_), .CI(mul_ex_mult_90_SUMB_2__6_), .CO(
        mul_ex_mult_90_CARRYB_3__5_), .S(mul_ex_mult_90_SUMB_3__5_) );
  FA_X1 mul_ex_mult_90_S2_3_4 ( .A(mul_ex_mult_90_ab_3__4_), .B(
        mul_ex_mult_90_CARRYB_2__4_), .CI(mul_ex_mult_90_SUMB_2__5_), .CO(
        mul_ex_mult_90_CARRYB_3__4_), .S(mul_ex_mult_90_SUMB_3__4_) );
  FA_X1 mul_ex_mult_90_S2_3_3 ( .A(mul_ex_mult_90_ab_3__3_), .B(
        mul_ex_mult_90_CARRYB_2__3_), .CI(mul_ex_mult_90_SUMB_2__4_), .CO(
        mul_ex_mult_90_CARRYB_3__3_), .S(mul_ex_mult_90_SUMB_3__3_) );
  FA_X1 mul_ex_mult_90_S2_3_2 ( .A(mul_ex_mult_90_ab_3__2_), .B(
        mul_ex_mult_90_CARRYB_2__2_), .CI(mul_ex_mult_90_SUMB_2__3_), .CO(
        mul_ex_mult_90_CARRYB_3__2_), .S(mul_ex_mult_90_SUMB_3__2_) );
  FA_X1 mul_ex_mult_90_S2_3_1 ( .A(mul_ex_mult_90_ab_3__1_), .B(
        mul_ex_mult_90_CARRYB_2__1_), .CI(mul_ex_mult_90_SUMB_2__2_), .CO(
        mul_ex_mult_90_CARRYB_3__1_), .S(mul_ex_mult_90_SUMB_3__1_) );
  FA_X1 mul_ex_mult_90_S1_3_0 ( .A(mul_ex_mult_90_ab_3__0_), .B(
        mul_ex_mult_90_CARRYB_2__0_), .CI(mul_ex_mult_90_SUMB_2__1_), .CO(
        mul_ex_mult_90_CARRYB_3__0_), .S(mul_ex_N157) );
  FA_X1 mul_ex_mult_90_S2_4_15 ( .A(mul_ex_mult_90_ab_4__15_), .B(
        mul_ex_mult_90_CARRYB_3__15_), .CI(mul_ex_mult_90_SUMB_3__16_), .CO(
        mul_ex_mult_90_CARRYB_4__15_), .S(mul_ex_mult_90_SUMB_4__15_) );
  FA_X1 mul_ex_mult_90_S2_4_14 ( .A(mul_ex_mult_90_ab_4__14_), .B(
        mul_ex_mult_90_CARRYB_3__14_), .CI(mul_ex_mult_90_SUMB_3__15_), .CO(
        mul_ex_mult_90_CARRYB_4__14_), .S(mul_ex_mult_90_SUMB_4__14_) );
  FA_X1 mul_ex_mult_90_S2_4_13 ( .A(mul_ex_mult_90_ab_4__13_), .B(
        mul_ex_mult_90_CARRYB_3__13_), .CI(mul_ex_mult_90_SUMB_3__14_), .CO(
        mul_ex_mult_90_CARRYB_4__13_), .S(mul_ex_mult_90_SUMB_4__13_) );
  FA_X1 mul_ex_mult_90_S2_4_12 ( .A(mul_ex_mult_90_ab_4__12_), .B(
        mul_ex_mult_90_CARRYB_3__12_), .CI(mul_ex_mult_90_SUMB_3__13_), .CO(
        mul_ex_mult_90_CARRYB_4__12_), .S(mul_ex_mult_90_SUMB_4__12_) );
  FA_X1 mul_ex_mult_90_S2_4_11 ( .A(mul_ex_mult_90_ab_4__11_), .B(
        mul_ex_mult_90_CARRYB_3__11_), .CI(mul_ex_mult_90_SUMB_3__12_), .CO(
        mul_ex_mult_90_CARRYB_4__11_), .S(mul_ex_mult_90_SUMB_4__11_) );
  FA_X1 mul_ex_mult_90_S2_4_10 ( .A(mul_ex_mult_90_ab_4__10_), .B(
        mul_ex_mult_90_CARRYB_3__10_), .CI(mul_ex_mult_90_SUMB_3__11_), .CO(
        mul_ex_mult_90_CARRYB_4__10_), .S(mul_ex_mult_90_SUMB_4__10_) );
  FA_X1 mul_ex_mult_90_S2_4_9 ( .A(mul_ex_mult_90_ab_4__9_), .B(
        mul_ex_mult_90_CARRYB_3__9_), .CI(mul_ex_mult_90_SUMB_3__10_), .CO(
        mul_ex_mult_90_CARRYB_4__9_), .S(mul_ex_mult_90_SUMB_4__9_) );
  FA_X1 mul_ex_mult_90_S2_4_8 ( .A(mul_ex_mult_90_ab_4__8_), .B(
        mul_ex_mult_90_CARRYB_3__8_), .CI(mul_ex_mult_90_SUMB_3__9_), .CO(
        mul_ex_mult_90_CARRYB_4__8_), .S(mul_ex_mult_90_SUMB_4__8_) );
  FA_X1 mul_ex_mult_90_S2_4_7 ( .A(mul_ex_mult_90_ab_4__7_), .B(
        mul_ex_mult_90_CARRYB_3__7_), .CI(mul_ex_mult_90_SUMB_3__8_), .CO(
        mul_ex_mult_90_CARRYB_4__7_), .S(mul_ex_mult_90_SUMB_4__7_) );
  FA_X1 mul_ex_mult_90_S2_4_6 ( .A(mul_ex_mult_90_ab_4__6_), .B(
        mul_ex_mult_90_CARRYB_3__6_), .CI(mul_ex_mult_90_SUMB_3__7_), .CO(
        mul_ex_mult_90_CARRYB_4__6_), .S(mul_ex_mult_90_SUMB_4__6_) );
  FA_X1 mul_ex_mult_90_S2_4_5 ( .A(mul_ex_mult_90_ab_4__5_), .B(
        mul_ex_mult_90_CARRYB_3__5_), .CI(mul_ex_mult_90_SUMB_3__6_), .CO(
        mul_ex_mult_90_CARRYB_4__5_), .S(mul_ex_mult_90_SUMB_4__5_) );
  FA_X1 mul_ex_mult_90_S2_4_4 ( .A(mul_ex_mult_90_ab_4__4_), .B(
        mul_ex_mult_90_CARRYB_3__4_), .CI(mul_ex_mult_90_SUMB_3__5_), .CO(
        mul_ex_mult_90_CARRYB_4__4_), .S(mul_ex_mult_90_SUMB_4__4_) );
  FA_X1 mul_ex_mult_90_S2_4_3 ( .A(mul_ex_mult_90_ab_4__3_), .B(
        mul_ex_mult_90_CARRYB_3__3_), .CI(mul_ex_mult_90_SUMB_3__4_), .CO(
        mul_ex_mult_90_CARRYB_4__3_), .S(mul_ex_mult_90_SUMB_4__3_) );
  FA_X1 mul_ex_mult_90_S2_4_2 ( .A(mul_ex_mult_90_ab_4__2_), .B(
        mul_ex_mult_90_CARRYB_3__2_), .CI(mul_ex_mult_90_SUMB_3__3_), .CO(
        mul_ex_mult_90_CARRYB_4__2_), .S(mul_ex_mult_90_SUMB_4__2_) );
  FA_X1 mul_ex_mult_90_S2_4_1 ( .A(mul_ex_mult_90_ab_4__1_), .B(
        mul_ex_mult_90_CARRYB_3__1_), .CI(mul_ex_mult_90_SUMB_3__2_), .CO(
        mul_ex_mult_90_CARRYB_4__1_), .S(mul_ex_mult_90_SUMB_4__1_) );
  FA_X1 mul_ex_mult_90_S1_4_0 ( .A(mul_ex_mult_90_ab_4__0_), .B(
        mul_ex_mult_90_CARRYB_3__0_), .CI(mul_ex_mult_90_SUMB_3__1_), .CO(
        mul_ex_mult_90_CARRYB_4__0_), .S(mul_ex_N158) );
  FA_X1 mul_ex_mult_90_S2_5_15 ( .A(mul_ex_mult_90_ab_5__15_), .B(
        mul_ex_mult_90_CARRYB_4__15_), .CI(mul_ex_mult_90_SUMB_4__16_), .CO(
        mul_ex_mult_90_CARRYB_5__15_), .S(mul_ex_mult_90_SUMB_5__15_) );
  FA_X1 mul_ex_mult_90_S2_5_14 ( .A(mul_ex_mult_90_ab_5__14_), .B(
        mul_ex_mult_90_CARRYB_4__14_), .CI(mul_ex_mult_90_SUMB_4__15_), .CO(
        mul_ex_mult_90_CARRYB_5__14_), .S(mul_ex_mult_90_SUMB_5__14_) );
  FA_X1 mul_ex_mult_90_S2_5_13 ( .A(mul_ex_mult_90_ab_5__13_), .B(
        mul_ex_mult_90_CARRYB_4__13_), .CI(mul_ex_mult_90_SUMB_4__14_), .CO(
        mul_ex_mult_90_CARRYB_5__13_), .S(mul_ex_mult_90_SUMB_5__13_) );
  FA_X1 mul_ex_mult_90_S2_5_12 ( .A(mul_ex_mult_90_ab_5__12_), .B(
        mul_ex_mult_90_CARRYB_4__12_), .CI(mul_ex_mult_90_SUMB_4__13_), .CO(
        mul_ex_mult_90_CARRYB_5__12_), .S(mul_ex_mult_90_SUMB_5__12_) );
  FA_X1 mul_ex_mult_90_S2_5_11 ( .A(mul_ex_mult_90_ab_5__11_), .B(
        mul_ex_mult_90_CARRYB_4__11_), .CI(mul_ex_mult_90_SUMB_4__12_), .CO(
        mul_ex_mult_90_CARRYB_5__11_), .S(mul_ex_mult_90_SUMB_5__11_) );
  FA_X1 mul_ex_mult_90_S2_5_10 ( .A(mul_ex_mult_90_ab_5__10_), .B(
        mul_ex_mult_90_CARRYB_4__10_), .CI(mul_ex_mult_90_SUMB_4__11_), .CO(
        mul_ex_mult_90_CARRYB_5__10_), .S(mul_ex_mult_90_SUMB_5__10_) );
  FA_X1 mul_ex_mult_90_S2_5_9 ( .A(mul_ex_mult_90_ab_5__9_), .B(
        mul_ex_mult_90_CARRYB_4__9_), .CI(mul_ex_mult_90_SUMB_4__10_), .CO(
        mul_ex_mult_90_CARRYB_5__9_), .S(mul_ex_mult_90_SUMB_5__9_) );
  FA_X1 mul_ex_mult_90_S2_5_8 ( .A(mul_ex_mult_90_ab_5__8_), .B(
        mul_ex_mult_90_CARRYB_4__8_), .CI(mul_ex_mult_90_SUMB_4__9_), .CO(
        mul_ex_mult_90_CARRYB_5__8_), .S(mul_ex_mult_90_SUMB_5__8_) );
  FA_X1 mul_ex_mult_90_S2_5_7 ( .A(mul_ex_mult_90_ab_5__7_), .B(
        mul_ex_mult_90_CARRYB_4__7_), .CI(mul_ex_mult_90_SUMB_4__8_), .CO(
        mul_ex_mult_90_CARRYB_5__7_), .S(mul_ex_mult_90_SUMB_5__7_) );
  FA_X1 mul_ex_mult_90_S2_5_6 ( .A(mul_ex_mult_90_ab_5__6_), .B(
        mul_ex_mult_90_CARRYB_4__6_), .CI(mul_ex_mult_90_SUMB_4__7_), .CO(
        mul_ex_mult_90_CARRYB_5__6_), .S(mul_ex_mult_90_SUMB_5__6_) );
  FA_X1 mul_ex_mult_90_S2_5_5 ( .A(mul_ex_mult_90_ab_5__5_), .B(
        mul_ex_mult_90_CARRYB_4__5_), .CI(mul_ex_mult_90_SUMB_4__6_), .CO(
        mul_ex_mult_90_CARRYB_5__5_), .S(mul_ex_mult_90_SUMB_5__5_) );
  FA_X1 mul_ex_mult_90_S2_5_4 ( .A(mul_ex_mult_90_ab_5__4_), .B(
        mul_ex_mult_90_CARRYB_4__4_), .CI(mul_ex_mult_90_SUMB_4__5_), .CO(
        mul_ex_mult_90_CARRYB_5__4_), .S(mul_ex_mult_90_SUMB_5__4_) );
  FA_X1 mul_ex_mult_90_S2_5_3 ( .A(mul_ex_mult_90_ab_5__3_), .B(
        mul_ex_mult_90_CARRYB_4__3_), .CI(mul_ex_mult_90_SUMB_4__4_), .CO(
        mul_ex_mult_90_CARRYB_5__3_), .S(mul_ex_mult_90_SUMB_5__3_) );
  FA_X1 mul_ex_mult_90_S2_5_2 ( .A(mul_ex_mult_90_ab_5__2_), .B(
        mul_ex_mult_90_CARRYB_4__2_), .CI(mul_ex_mult_90_SUMB_4__3_), .CO(
        mul_ex_mult_90_CARRYB_5__2_), .S(mul_ex_mult_90_SUMB_5__2_) );
  FA_X1 mul_ex_mult_90_S2_5_1 ( .A(mul_ex_mult_90_ab_5__1_), .B(
        mul_ex_mult_90_CARRYB_4__1_), .CI(mul_ex_mult_90_SUMB_4__2_), .CO(
        mul_ex_mult_90_CARRYB_5__1_), .S(mul_ex_mult_90_SUMB_5__1_) );
  FA_X1 mul_ex_mult_90_S1_5_0 ( .A(mul_ex_mult_90_ab_5__0_), .B(
        mul_ex_mult_90_CARRYB_4__0_), .CI(mul_ex_mult_90_SUMB_4__1_), .CO(
        mul_ex_mult_90_CARRYB_5__0_), .S(mul_ex_N159) );
  FA_X1 mul_ex_mult_90_S2_6_15 ( .A(mul_ex_mult_90_ab_6__15_), .B(
        mul_ex_mult_90_CARRYB_5__15_), .CI(mul_ex_mult_90_SUMB_5__16_), .CO(
        mul_ex_mult_90_CARRYB_6__15_), .S(mul_ex_mult_90_SUMB_6__15_) );
  FA_X1 mul_ex_mult_90_S2_6_14 ( .A(mul_ex_mult_90_ab_6__14_), .B(
        mul_ex_mult_90_CARRYB_5__14_), .CI(mul_ex_mult_90_SUMB_5__15_), .CO(
        mul_ex_mult_90_CARRYB_6__14_), .S(mul_ex_mult_90_SUMB_6__14_) );
  FA_X1 mul_ex_mult_90_S2_6_13 ( .A(mul_ex_mult_90_ab_6__13_), .B(
        mul_ex_mult_90_CARRYB_5__13_), .CI(mul_ex_mult_90_SUMB_5__14_), .CO(
        mul_ex_mult_90_CARRYB_6__13_), .S(mul_ex_mult_90_SUMB_6__13_) );
  FA_X1 mul_ex_mult_90_S2_6_12 ( .A(mul_ex_mult_90_ab_6__12_), .B(
        mul_ex_mult_90_CARRYB_5__12_), .CI(mul_ex_mult_90_SUMB_5__13_), .CO(
        mul_ex_mult_90_CARRYB_6__12_), .S(mul_ex_mult_90_SUMB_6__12_) );
  FA_X1 mul_ex_mult_90_S2_6_11 ( .A(mul_ex_mult_90_ab_6__11_), .B(
        mul_ex_mult_90_CARRYB_5__11_), .CI(mul_ex_mult_90_SUMB_5__12_), .CO(
        mul_ex_mult_90_CARRYB_6__11_), .S(mul_ex_mult_90_SUMB_6__11_) );
  FA_X1 mul_ex_mult_90_S2_6_10 ( .A(mul_ex_mult_90_ab_6__10_), .B(
        mul_ex_mult_90_CARRYB_5__10_), .CI(mul_ex_mult_90_SUMB_5__11_), .CO(
        mul_ex_mult_90_CARRYB_6__10_), .S(mul_ex_mult_90_SUMB_6__10_) );
  FA_X1 mul_ex_mult_90_S2_6_9 ( .A(mul_ex_mult_90_ab_6__9_), .B(
        mul_ex_mult_90_CARRYB_5__9_), .CI(mul_ex_mult_90_SUMB_5__10_), .CO(
        mul_ex_mult_90_CARRYB_6__9_), .S(mul_ex_mult_90_SUMB_6__9_) );
  FA_X1 mul_ex_mult_90_S2_6_8 ( .A(mul_ex_mult_90_ab_6__8_), .B(
        mul_ex_mult_90_CARRYB_5__8_), .CI(mul_ex_mult_90_SUMB_5__9_), .CO(
        mul_ex_mult_90_CARRYB_6__8_), .S(mul_ex_mult_90_SUMB_6__8_) );
  FA_X1 mul_ex_mult_90_S2_6_7 ( .A(mul_ex_mult_90_ab_6__7_), .B(
        mul_ex_mult_90_CARRYB_5__7_), .CI(mul_ex_mult_90_SUMB_5__8_), .CO(
        mul_ex_mult_90_CARRYB_6__7_), .S(mul_ex_mult_90_SUMB_6__7_) );
  FA_X1 mul_ex_mult_90_S2_6_6 ( .A(mul_ex_mult_90_ab_6__6_), .B(
        mul_ex_mult_90_CARRYB_5__6_), .CI(mul_ex_mult_90_SUMB_5__7_), .CO(
        mul_ex_mult_90_CARRYB_6__6_), .S(mul_ex_mult_90_SUMB_6__6_) );
  FA_X1 mul_ex_mult_90_S2_6_5 ( .A(mul_ex_mult_90_ab_6__5_), .B(
        mul_ex_mult_90_CARRYB_5__5_), .CI(mul_ex_mult_90_SUMB_5__6_), .CO(
        mul_ex_mult_90_CARRYB_6__5_), .S(mul_ex_mult_90_SUMB_6__5_) );
  FA_X1 mul_ex_mult_90_S2_6_4 ( .A(mul_ex_mult_90_ab_6__4_), .B(
        mul_ex_mult_90_CARRYB_5__4_), .CI(mul_ex_mult_90_SUMB_5__5_), .CO(
        mul_ex_mult_90_CARRYB_6__4_), .S(mul_ex_mult_90_SUMB_6__4_) );
  FA_X1 mul_ex_mult_90_S2_6_3 ( .A(mul_ex_mult_90_ab_6__3_), .B(
        mul_ex_mult_90_CARRYB_5__3_), .CI(mul_ex_mult_90_SUMB_5__4_), .CO(
        mul_ex_mult_90_CARRYB_6__3_), .S(mul_ex_mult_90_SUMB_6__3_) );
  FA_X1 mul_ex_mult_90_S2_6_2 ( .A(mul_ex_mult_90_ab_6__2_), .B(
        mul_ex_mult_90_CARRYB_5__2_), .CI(mul_ex_mult_90_SUMB_5__3_), .CO(
        mul_ex_mult_90_CARRYB_6__2_), .S(mul_ex_mult_90_SUMB_6__2_) );
  FA_X1 mul_ex_mult_90_S2_6_1 ( .A(mul_ex_mult_90_ab_6__1_), .B(
        mul_ex_mult_90_CARRYB_5__1_), .CI(mul_ex_mult_90_SUMB_5__2_), .CO(
        mul_ex_mult_90_CARRYB_6__1_), .S(mul_ex_mult_90_SUMB_6__1_) );
  FA_X1 mul_ex_mult_90_S1_6_0 ( .A(mul_ex_mult_90_ab_6__0_), .B(
        mul_ex_mult_90_CARRYB_5__0_), .CI(mul_ex_mult_90_SUMB_5__1_), .CO(
        mul_ex_mult_90_CARRYB_6__0_), .S(mul_ex_N160) );
  FA_X1 mul_ex_mult_90_S2_7_15 ( .A(mul_ex_mult_90_ab_7__15_), .B(
        mul_ex_mult_90_CARRYB_6__15_), .CI(mul_ex_mult_90_SUMB_6__16_), .CO(
        mul_ex_mult_90_CARRYB_7__15_), .S(mul_ex_mult_90_SUMB_7__15_) );
  FA_X1 mul_ex_mult_90_S2_7_14 ( .A(mul_ex_mult_90_ab_7__14_), .B(
        mul_ex_mult_90_CARRYB_6__14_), .CI(mul_ex_mult_90_SUMB_6__15_), .CO(
        mul_ex_mult_90_CARRYB_7__14_), .S(mul_ex_mult_90_SUMB_7__14_) );
  FA_X1 mul_ex_mult_90_S2_7_13 ( .A(mul_ex_mult_90_ab_7__13_), .B(
        mul_ex_mult_90_CARRYB_6__13_), .CI(mul_ex_mult_90_SUMB_6__14_), .CO(
        mul_ex_mult_90_CARRYB_7__13_), .S(mul_ex_mult_90_SUMB_7__13_) );
  FA_X1 mul_ex_mult_90_S2_7_12 ( .A(mul_ex_mult_90_ab_7__12_), .B(
        mul_ex_mult_90_CARRYB_6__12_), .CI(mul_ex_mult_90_SUMB_6__13_), .CO(
        mul_ex_mult_90_CARRYB_7__12_), .S(mul_ex_mult_90_SUMB_7__12_) );
  FA_X1 mul_ex_mult_90_S2_7_11 ( .A(mul_ex_mult_90_ab_7__11_), .B(
        mul_ex_mult_90_CARRYB_6__11_), .CI(mul_ex_mult_90_SUMB_6__12_), .CO(
        mul_ex_mult_90_CARRYB_7__11_), .S(mul_ex_mult_90_SUMB_7__11_) );
  FA_X1 mul_ex_mult_90_S2_7_10 ( .A(mul_ex_mult_90_ab_7__10_), .B(
        mul_ex_mult_90_CARRYB_6__10_), .CI(mul_ex_mult_90_SUMB_6__11_), .CO(
        mul_ex_mult_90_CARRYB_7__10_), .S(mul_ex_mult_90_SUMB_7__10_) );
  FA_X1 mul_ex_mult_90_S2_7_9 ( .A(mul_ex_mult_90_ab_7__9_), .B(
        mul_ex_mult_90_CARRYB_6__9_), .CI(mul_ex_mult_90_SUMB_6__10_), .CO(
        mul_ex_mult_90_CARRYB_7__9_), .S(mul_ex_mult_90_SUMB_7__9_) );
  FA_X1 mul_ex_mult_90_S2_7_8 ( .A(mul_ex_mult_90_ab_7__8_), .B(
        mul_ex_mult_90_CARRYB_6__8_), .CI(mul_ex_mult_90_SUMB_6__9_), .CO(
        mul_ex_mult_90_CARRYB_7__8_), .S(mul_ex_mult_90_SUMB_7__8_) );
  FA_X1 mul_ex_mult_90_S2_7_7 ( .A(mul_ex_mult_90_ab_7__7_), .B(
        mul_ex_mult_90_CARRYB_6__7_), .CI(mul_ex_mult_90_SUMB_6__8_), .CO(
        mul_ex_mult_90_CARRYB_7__7_), .S(mul_ex_mult_90_SUMB_7__7_) );
  FA_X1 mul_ex_mult_90_S2_7_6 ( .A(mul_ex_mult_90_ab_7__6_), .B(
        mul_ex_mult_90_CARRYB_6__6_), .CI(mul_ex_mult_90_SUMB_6__7_), .CO(
        mul_ex_mult_90_CARRYB_7__6_), .S(mul_ex_mult_90_SUMB_7__6_) );
  FA_X1 mul_ex_mult_90_S2_7_5 ( .A(mul_ex_mult_90_ab_7__5_), .B(
        mul_ex_mult_90_CARRYB_6__5_), .CI(mul_ex_mult_90_SUMB_6__6_), .CO(
        mul_ex_mult_90_CARRYB_7__5_), .S(mul_ex_mult_90_SUMB_7__5_) );
  FA_X1 mul_ex_mult_90_S2_7_4 ( .A(mul_ex_mult_90_ab_7__4_), .B(
        mul_ex_mult_90_CARRYB_6__4_), .CI(mul_ex_mult_90_SUMB_6__5_), .CO(
        mul_ex_mult_90_CARRYB_7__4_), .S(mul_ex_mult_90_SUMB_7__4_) );
  FA_X1 mul_ex_mult_90_S2_7_3 ( .A(mul_ex_mult_90_ab_7__3_), .B(
        mul_ex_mult_90_CARRYB_6__3_), .CI(mul_ex_mult_90_SUMB_6__4_), .CO(
        mul_ex_mult_90_CARRYB_7__3_), .S(mul_ex_mult_90_SUMB_7__3_) );
  FA_X1 mul_ex_mult_90_S2_7_2 ( .A(mul_ex_mult_90_ab_7__2_), .B(
        mul_ex_mult_90_CARRYB_6__2_), .CI(mul_ex_mult_90_SUMB_6__3_), .CO(
        mul_ex_mult_90_CARRYB_7__2_), .S(mul_ex_mult_90_SUMB_7__2_) );
  FA_X1 mul_ex_mult_90_S2_7_1 ( .A(mul_ex_mult_90_ab_7__1_), .B(
        mul_ex_mult_90_CARRYB_6__1_), .CI(mul_ex_mult_90_SUMB_6__2_), .CO(
        mul_ex_mult_90_CARRYB_7__1_), .S(mul_ex_mult_90_SUMB_7__1_) );
  FA_X1 mul_ex_mult_90_S1_7_0 ( .A(mul_ex_mult_90_ab_7__0_), .B(
        mul_ex_mult_90_CARRYB_6__0_), .CI(mul_ex_mult_90_SUMB_6__1_), .CO(
        mul_ex_mult_90_CARRYB_7__0_), .S(mul_ex_N161) );
  FA_X1 mul_ex_mult_90_S2_8_15 ( .A(mul_ex_mult_90_ab_8__15_), .B(
        mul_ex_mult_90_CARRYB_7__15_), .CI(mul_ex_mult_90_SUMB_7__16_), .CO(
        mul_ex_mult_90_CARRYB_8__15_), .S(mul_ex_mult_90_SUMB_8__15_) );
  FA_X1 mul_ex_mult_90_S2_8_14 ( .A(mul_ex_mult_90_ab_8__14_), .B(
        mul_ex_mult_90_CARRYB_7__14_), .CI(mul_ex_mult_90_SUMB_7__15_), .CO(
        mul_ex_mult_90_CARRYB_8__14_), .S(mul_ex_mult_90_SUMB_8__14_) );
  FA_X1 mul_ex_mult_90_S2_8_13 ( .A(mul_ex_mult_90_ab_8__13_), .B(
        mul_ex_mult_90_CARRYB_7__13_), .CI(mul_ex_mult_90_SUMB_7__14_), .CO(
        mul_ex_mult_90_CARRYB_8__13_), .S(mul_ex_mult_90_SUMB_8__13_) );
  FA_X1 mul_ex_mult_90_S2_8_12 ( .A(mul_ex_mult_90_ab_8__12_), .B(
        mul_ex_mult_90_CARRYB_7__12_), .CI(mul_ex_mult_90_SUMB_7__13_), .CO(
        mul_ex_mult_90_CARRYB_8__12_), .S(mul_ex_mult_90_SUMB_8__12_) );
  FA_X1 mul_ex_mult_90_S2_8_11 ( .A(mul_ex_mult_90_ab_8__11_), .B(
        mul_ex_mult_90_CARRYB_7__11_), .CI(mul_ex_mult_90_SUMB_7__12_), .CO(
        mul_ex_mult_90_CARRYB_8__11_), .S(mul_ex_mult_90_SUMB_8__11_) );
  FA_X1 mul_ex_mult_90_S2_8_10 ( .A(mul_ex_mult_90_ab_8__10_), .B(
        mul_ex_mult_90_CARRYB_7__10_), .CI(mul_ex_mult_90_SUMB_7__11_), .CO(
        mul_ex_mult_90_CARRYB_8__10_), .S(mul_ex_mult_90_SUMB_8__10_) );
  FA_X1 mul_ex_mult_90_S2_8_9 ( .A(mul_ex_mult_90_ab_8__9_), .B(
        mul_ex_mult_90_CARRYB_7__9_), .CI(mul_ex_mult_90_SUMB_7__10_), .CO(
        mul_ex_mult_90_CARRYB_8__9_), .S(mul_ex_mult_90_SUMB_8__9_) );
  FA_X1 mul_ex_mult_90_S2_8_8 ( .A(mul_ex_mult_90_ab_8__8_), .B(
        mul_ex_mult_90_CARRYB_7__8_), .CI(mul_ex_mult_90_SUMB_7__9_), .CO(
        mul_ex_mult_90_CARRYB_8__8_), .S(mul_ex_mult_90_SUMB_8__8_) );
  FA_X1 mul_ex_mult_90_S2_8_7 ( .A(mul_ex_mult_90_ab_8__7_), .B(
        mul_ex_mult_90_CARRYB_7__7_), .CI(mul_ex_mult_90_SUMB_7__8_), .CO(
        mul_ex_mult_90_CARRYB_8__7_), .S(mul_ex_mult_90_SUMB_8__7_) );
  FA_X1 mul_ex_mult_90_S2_8_6 ( .A(mul_ex_mult_90_ab_8__6_), .B(
        mul_ex_mult_90_CARRYB_7__6_), .CI(mul_ex_mult_90_SUMB_7__7_), .CO(
        mul_ex_mult_90_CARRYB_8__6_), .S(mul_ex_mult_90_SUMB_8__6_) );
  FA_X1 mul_ex_mult_90_S2_8_5 ( .A(mul_ex_mult_90_ab_8__5_), .B(
        mul_ex_mult_90_CARRYB_7__5_), .CI(mul_ex_mult_90_SUMB_7__6_), .CO(
        mul_ex_mult_90_CARRYB_8__5_), .S(mul_ex_mult_90_SUMB_8__5_) );
  FA_X1 mul_ex_mult_90_S2_8_4 ( .A(mul_ex_mult_90_ab_8__4_), .B(
        mul_ex_mult_90_CARRYB_7__4_), .CI(mul_ex_mult_90_SUMB_7__5_), .CO(
        mul_ex_mult_90_CARRYB_8__4_), .S(mul_ex_mult_90_SUMB_8__4_) );
  FA_X1 mul_ex_mult_90_S2_8_3 ( .A(mul_ex_mult_90_ab_8__3_), .B(
        mul_ex_mult_90_CARRYB_7__3_), .CI(mul_ex_mult_90_SUMB_7__4_), .CO(
        mul_ex_mult_90_CARRYB_8__3_), .S(mul_ex_mult_90_SUMB_8__3_) );
  FA_X1 mul_ex_mult_90_S2_8_2 ( .A(mul_ex_mult_90_ab_8__2_), .B(
        mul_ex_mult_90_CARRYB_7__2_), .CI(mul_ex_mult_90_SUMB_7__3_), .CO(
        mul_ex_mult_90_CARRYB_8__2_), .S(mul_ex_mult_90_SUMB_8__2_) );
  FA_X1 mul_ex_mult_90_S2_8_1 ( .A(mul_ex_mult_90_ab_8__1_), .B(
        mul_ex_mult_90_CARRYB_7__1_), .CI(mul_ex_mult_90_SUMB_7__2_), .CO(
        mul_ex_mult_90_CARRYB_8__1_), .S(mul_ex_mult_90_SUMB_8__1_) );
  FA_X1 mul_ex_mult_90_S1_8_0 ( .A(mul_ex_mult_90_ab_8__0_), .B(
        mul_ex_mult_90_CARRYB_7__0_), .CI(mul_ex_mult_90_SUMB_7__1_), .CO(
        mul_ex_mult_90_CARRYB_8__0_), .S(mul_ex_N162) );
  FA_X1 mul_ex_mult_90_S2_9_15 ( .A(mul_ex_mult_90_ab_9__15_), .B(
        mul_ex_mult_90_CARRYB_8__15_), .CI(mul_ex_mult_90_SUMB_8__16_), .CO(
        mul_ex_mult_90_CARRYB_9__15_), .S(mul_ex_mult_90_SUMB_9__15_) );
  FA_X1 mul_ex_mult_90_S2_9_14 ( .A(mul_ex_mult_90_ab_9__14_), .B(
        mul_ex_mult_90_CARRYB_8__14_), .CI(mul_ex_mult_90_SUMB_8__15_), .CO(
        mul_ex_mult_90_CARRYB_9__14_), .S(mul_ex_mult_90_SUMB_9__14_) );
  FA_X1 mul_ex_mult_90_S2_9_13 ( .A(mul_ex_mult_90_ab_9__13_), .B(
        mul_ex_mult_90_CARRYB_8__13_), .CI(mul_ex_mult_90_SUMB_8__14_), .CO(
        mul_ex_mult_90_CARRYB_9__13_), .S(mul_ex_mult_90_SUMB_9__13_) );
  FA_X1 mul_ex_mult_90_S2_9_12 ( .A(mul_ex_mult_90_ab_9__12_), .B(
        mul_ex_mult_90_CARRYB_8__12_), .CI(mul_ex_mult_90_SUMB_8__13_), .CO(
        mul_ex_mult_90_CARRYB_9__12_), .S(mul_ex_mult_90_SUMB_9__12_) );
  FA_X1 mul_ex_mult_90_S2_9_11 ( .A(mul_ex_mult_90_ab_9__11_), .B(
        mul_ex_mult_90_CARRYB_8__11_), .CI(mul_ex_mult_90_SUMB_8__12_), .CO(
        mul_ex_mult_90_CARRYB_9__11_), .S(mul_ex_mult_90_SUMB_9__11_) );
  FA_X1 mul_ex_mult_90_S2_9_10 ( .A(mul_ex_mult_90_ab_9__10_), .B(
        mul_ex_mult_90_CARRYB_8__10_), .CI(mul_ex_mult_90_SUMB_8__11_), .CO(
        mul_ex_mult_90_CARRYB_9__10_), .S(mul_ex_mult_90_SUMB_9__10_) );
  FA_X1 mul_ex_mult_90_S2_9_9 ( .A(mul_ex_mult_90_ab_9__9_), .B(
        mul_ex_mult_90_CARRYB_8__9_), .CI(mul_ex_mult_90_SUMB_8__10_), .CO(
        mul_ex_mult_90_CARRYB_9__9_), .S(mul_ex_mult_90_SUMB_9__9_) );
  FA_X1 mul_ex_mult_90_S2_9_8 ( .A(mul_ex_mult_90_ab_9__8_), .B(
        mul_ex_mult_90_CARRYB_8__8_), .CI(mul_ex_mult_90_SUMB_8__9_), .CO(
        mul_ex_mult_90_CARRYB_9__8_), .S(mul_ex_mult_90_SUMB_9__8_) );
  FA_X1 mul_ex_mult_90_S2_9_7 ( .A(mul_ex_mult_90_ab_9__7_), .B(
        mul_ex_mult_90_CARRYB_8__7_), .CI(mul_ex_mult_90_SUMB_8__8_), .CO(
        mul_ex_mult_90_CARRYB_9__7_), .S(mul_ex_mult_90_SUMB_9__7_) );
  FA_X1 mul_ex_mult_90_S2_9_6 ( .A(mul_ex_mult_90_ab_9__6_), .B(
        mul_ex_mult_90_CARRYB_8__6_), .CI(mul_ex_mult_90_SUMB_8__7_), .CO(
        mul_ex_mult_90_CARRYB_9__6_), .S(mul_ex_mult_90_SUMB_9__6_) );
  FA_X1 mul_ex_mult_90_S2_9_5 ( .A(mul_ex_mult_90_ab_9__5_), .B(
        mul_ex_mult_90_CARRYB_8__5_), .CI(mul_ex_mult_90_SUMB_8__6_), .CO(
        mul_ex_mult_90_CARRYB_9__5_), .S(mul_ex_mult_90_SUMB_9__5_) );
  FA_X1 mul_ex_mult_90_S2_9_4 ( .A(mul_ex_mult_90_ab_9__4_), .B(
        mul_ex_mult_90_CARRYB_8__4_), .CI(mul_ex_mult_90_SUMB_8__5_), .CO(
        mul_ex_mult_90_CARRYB_9__4_), .S(mul_ex_mult_90_SUMB_9__4_) );
  FA_X1 mul_ex_mult_90_S2_9_3 ( .A(mul_ex_mult_90_ab_9__3_), .B(
        mul_ex_mult_90_CARRYB_8__3_), .CI(mul_ex_mult_90_SUMB_8__4_), .CO(
        mul_ex_mult_90_CARRYB_9__3_), .S(mul_ex_mult_90_SUMB_9__3_) );
  FA_X1 mul_ex_mult_90_S2_9_2 ( .A(mul_ex_mult_90_ab_9__2_), .B(
        mul_ex_mult_90_CARRYB_8__2_), .CI(mul_ex_mult_90_SUMB_8__3_), .CO(
        mul_ex_mult_90_CARRYB_9__2_), .S(mul_ex_mult_90_SUMB_9__2_) );
  FA_X1 mul_ex_mult_90_S2_9_1 ( .A(mul_ex_mult_90_ab_9__1_), .B(
        mul_ex_mult_90_CARRYB_8__1_), .CI(mul_ex_mult_90_SUMB_8__2_), .CO(
        mul_ex_mult_90_CARRYB_9__1_), .S(mul_ex_mult_90_SUMB_9__1_) );
  FA_X1 mul_ex_mult_90_S1_9_0 ( .A(mul_ex_mult_90_ab_9__0_), .B(
        mul_ex_mult_90_CARRYB_8__0_), .CI(mul_ex_mult_90_SUMB_8__1_), .CO(
        mul_ex_mult_90_CARRYB_9__0_), .S(mul_ex_N163) );
  FA_X1 mul_ex_mult_90_S2_10_15 ( .A(mul_ex_mult_90_ab_10__15_), .B(
        mul_ex_mult_90_CARRYB_9__15_), .CI(mul_ex_mult_90_SUMB_9__16_), .CO(
        mul_ex_mult_90_CARRYB_10__15_), .S(mul_ex_mult_90_SUMB_10__15_) );
  FA_X1 mul_ex_mult_90_S2_10_14 ( .A(mul_ex_mult_90_ab_10__14_), .B(
        mul_ex_mult_90_CARRYB_9__14_), .CI(mul_ex_mult_90_SUMB_9__15_), .CO(
        mul_ex_mult_90_CARRYB_10__14_), .S(mul_ex_mult_90_SUMB_10__14_) );
  FA_X1 mul_ex_mult_90_S2_10_13 ( .A(mul_ex_mult_90_ab_10__13_), .B(
        mul_ex_mult_90_CARRYB_9__13_), .CI(mul_ex_mult_90_SUMB_9__14_), .CO(
        mul_ex_mult_90_CARRYB_10__13_), .S(mul_ex_mult_90_SUMB_10__13_) );
  FA_X1 mul_ex_mult_90_S2_10_12 ( .A(mul_ex_mult_90_ab_10__12_), .B(
        mul_ex_mult_90_CARRYB_9__12_), .CI(mul_ex_mult_90_SUMB_9__13_), .CO(
        mul_ex_mult_90_CARRYB_10__12_), .S(mul_ex_mult_90_SUMB_10__12_) );
  FA_X1 mul_ex_mult_90_S2_10_11 ( .A(mul_ex_mult_90_ab_10__11_), .B(
        mul_ex_mult_90_CARRYB_9__11_), .CI(mul_ex_mult_90_SUMB_9__12_), .CO(
        mul_ex_mult_90_CARRYB_10__11_), .S(mul_ex_mult_90_SUMB_10__11_) );
  FA_X1 mul_ex_mult_90_S2_10_10 ( .A(mul_ex_mult_90_ab_10__10_), .B(
        mul_ex_mult_90_CARRYB_9__10_), .CI(mul_ex_mult_90_SUMB_9__11_), .CO(
        mul_ex_mult_90_CARRYB_10__10_), .S(mul_ex_mult_90_SUMB_10__10_) );
  FA_X1 mul_ex_mult_90_S2_10_9 ( .A(mul_ex_mult_90_ab_10__9_), .B(
        mul_ex_mult_90_CARRYB_9__9_), .CI(mul_ex_mult_90_SUMB_9__10_), .CO(
        mul_ex_mult_90_CARRYB_10__9_), .S(mul_ex_mult_90_SUMB_10__9_) );
  FA_X1 mul_ex_mult_90_S2_10_8 ( .A(mul_ex_mult_90_ab_10__8_), .B(
        mul_ex_mult_90_CARRYB_9__8_), .CI(mul_ex_mult_90_SUMB_9__9_), .CO(
        mul_ex_mult_90_CARRYB_10__8_), .S(mul_ex_mult_90_SUMB_10__8_) );
  FA_X1 mul_ex_mult_90_S2_10_7 ( .A(mul_ex_mult_90_ab_10__7_), .B(
        mul_ex_mult_90_CARRYB_9__7_), .CI(mul_ex_mult_90_SUMB_9__8_), .CO(
        mul_ex_mult_90_CARRYB_10__7_), .S(mul_ex_mult_90_SUMB_10__7_) );
  FA_X1 mul_ex_mult_90_S2_10_6 ( .A(mul_ex_mult_90_ab_10__6_), .B(
        mul_ex_mult_90_CARRYB_9__6_), .CI(mul_ex_mult_90_SUMB_9__7_), .CO(
        mul_ex_mult_90_CARRYB_10__6_), .S(mul_ex_mult_90_SUMB_10__6_) );
  FA_X1 mul_ex_mult_90_S2_10_5 ( .A(mul_ex_mult_90_ab_10__5_), .B(
        mul_ex_mult_90_CARRYB_9__5_), .CI(mul_ex_mult_90_SUMB_9__6_), .CO(
        mul_ex_mult_90_CARRYB_10__5_), .S(mul_ex_mult_90_SUMB_10__5_) );
  FA_X1 mul_ex_mult_90_S2_10_4 ( .A(mul_ex_mult_90_ab_10__4_), .B(
        mul_ex_mult_90_CARRYB_9__4_), .CI(mul_ex_mult_90_SUMB_9__5_), .CO(
        mul_ex_mult_90_CARRYB_10__4_), .S(mul_ex_mult_90_SUMB_10__4_) );
  FA_X1 mul_ex_mult_90_S2_10_3 ( .A(mul_ex_mult_90_ab_10__3_), .B(
        mul_ex_mult_90_CARRYB_9__3_), .CI(mul_ex_mult_90_SUMB_9__4_), .CO(
        mul_ex_mult_90_CARRYB_10__3_), .S(mul_ex_mult_90_SUMB_10__3_) );
  FA_X1 mul_ex_mult_90_S2_10_2 ( .A(mul_ex_mult_90_ab_10__2_), .B(
        mul_ex_mult_90_CARRYB_9__2_), .CI(mul_ex_mult_90_SUMB_9__3_), .CO(
        mul_ex_mult_90_CARRYB_10__2_), .S(mul_ex_mult_90_SUMB_10__2_) );
  FA_X1 mul_ex_mult_90_S2_10_1 ( .A(mul_ex_mult_90_ab_10__1_), .B(
        mul_ex_mult_90_CARRYB_9__1_), .CI(mul_ex_mult_90_SUMB_9__2_), .CO(
        mul_ex_mult_90_CARRYB_10__1_), .S(mul_ex_mult_90_SUMB_10__1_) );
  FA_X1 mul_ex_mult_90_S1_10_0 ( .A(mul_ex_mult_90_ab_10__0_), .B(
        mul_ex_mult_90_CARRYB_9__0_), .CI(mul_ex_mult_90_SUMB_9__1_), .CO(
        mul_ex_mult_90_CARRYB_10__0_), .S(mul_ex_N164) );
  FA_X1 mul_ex_mult_90_S2_11_15 ( .A(mul_ex_mult_90_ab_11__15_), .B(
        mul_ex_mult_90_CARRYB_10__15_), .CI(mul_ex_mult_90_SUMB_10__16_), .CO(
        mul_ex_mult_90_CARRYB_11__15_), .S(mul_ex_mult_90_SUMB_11__15_) );
  FA_X1 mul_ex_mult_90_S2_11_14 ( .A(mul_ex_mult_90_ab_11__14_), .B(
        mul_ex_mult_90_CARRYB_10__14_), .CI(mul_ex_mult_90_SUMB_10__15_), .CO(
        mul_ex_mult_90_CARRYB_11__14_), .S(mul_ex_mult_90_SUMB_11__14_) );
  FA_X1 mul_ex_mult_90_S2_11_13 ( .A(mul_ex_mult_90_ab_11__13_), .B(
        mul_ex_mult_90_CARRYB_10__13_), .CI(mul_ex_mult_90_SUMB_10__14_), .CO(
        mul_ex_mult_90_CARRYB_11__13_), .S(mul_ex_mult_90_SUMB_11__13_) );
  FA_X1 mul_ex_mult_90_S2_11_12 ( .A(mul_ex_mult_90_ab_11__12_), .B(
        mul_ex_mult_90_CARRYB_10__12_), .CI(mul_ex_mult_90_SUMB_10__13_), .CO(
        mul_ex_mult_90_CARRYB_11__12_), .S(mul_ex_mult_90_SUMB_11__12_) );
  FA_X1 mul_ex_mult_90_S2_11_11 ( .A(mul_ex_mult_90_ab_11__11_), .B(
        mul_ex_mult_90_CARRYB_10__11_), .CI(mul_ex_mult_90_SUMB_10__12_), .CO(
        mul_ex_mult_90_CARRYB_11__11_), .S(mul_ex_mult_90_SUMB_11__11_) );
  FA_X1 mul_ex_mult_90_S2_11_10 ( .A(mul_ex_mult_90_ab_11__10_), .B(
        mul_ex_mult_90_CARRYB_10__10_), .CI(mul_ex_mult_90_SUMB_10__11_), .CO(
        mul_ex_mult_90_CARRYB_11__10_), .S(mul_ex_mult_90_SUMB_11__10_) );
  FA_X1 mul_ex_mult_90_S2_11_9 ( .A(mul_ex_mult_90_ab_11__9_), .B(
        mul_ex_mult_90_CARRYB_10__9_), .CI(mul_ex_mult_90_SUMB_10__10_), .CO(
        mul_ex_mult_90_CARRYB_11__9_), .S(mul_ex_mult_90_SUMB_11__9_) );
  FA_X1 mul_ex_mult_90_S2_11_8 ( .A(mul_ex_mult_90_ab_11__8_), .B(
        mul_ex_mult_90_CARRYB_10__8_), .CI(mul_ex_mult_90_SUMB_10__9_), .CO(
        mul_ex_mult_90_CARRYB_11__8_), .S(mul_ex_mult_90_SUMB_11__8_) );
  FA_X1 mul_ex_mult_90_S2_11_7 ( .A(mul_ex_mult_90_ab_11__7_), .B(
        mul_ex_mult_90_CARRYB_10__7_), .CI(mul_ex_mult_90_SUMB_10__8_), .CO(
        mul_ex_mult_90_CARRYB_11__7_), .S(mul_ex_mult_90_SUMB_11__7_) );
  FA_X1 mul_ex_mult_90_S2_11_6 ( .A(mul_ex_mult_90_ab_11__6_), .B(
        mul_ex_mult_90_CARRYB_10__6_), .CI(mul_ex_mult_90_SUMB_10__7_), .CO(
        mul_ex_mult_90_CARRYB_11__6_), .S(mul_ex_mult_90_SUMB_11__6_) );
  FA_X1 mul_ex_mult_90_S2_11_5 ( .A(mul_ex_mult_90_ab_11__5_), .B(
        mul_ex_mult_90_CARRYB_10__5_), .CI(mul_ex_mult_90_SUMB_10__6_), .CO(
        mul_ex_mult_90_CARRYB_11__5_), .S(mul_ex_mult_90_SUMB_11__5_) );
  FA_X1 mul_ex_mult_90_S2_11_4 ( .A(mul_ex_mult_90_ab_11__4_), .B(
        mul_ex_mult_90_CARRYB_10__4_), .CI(mul_ex_mult_90_SUMB_10__5_), .CO(
        mul_ex_mult_90_CARRYB_11__4_), .S(mul_ex_mult_90_SUMB_11__4_) );
  FA_X1 mul_ex_mult_90_S2_11_3 ( .A(mul_ex_mult_90_ab_11__3_), .B(
        mul_ex_mult_90_CARRYB_10__3_), .CI(mul_ex_mult_90_SUMB_10__4_), .CO(
        mul_ex_mult_90_CARRYB_11__3_), .S(mul_ex_mult_90_SUMB_11__3_) );
  FA_X1 mul_ex_mult_90_S2_11_2 ( .A(mul_ex_mult_90_ab_11__2_), .B(
        mul_ex_mult_90_CARRYB_10__2_), .CI(mul_ex_mult_90_SUMB_10__3_), .CO(
        mul_ex_mult_90_CARRYB_11__2_), .S(mul_ex_mult_90_SUMB_11__2_) );
  FA_X1 mul_ex_mult_90_S2_11_1 ( .A(mul_ex_mult_90_ab_11__1_), .B(
        mul_ex_mult_90_CARRYB_10__1_), .CI(mul_ex_mult_90_SUMB_10__2_), .CO(
        mul_ex_mult_90_CARRYB_11__1_), .S(mul_ex_mult_90_SUMB_11__1_) );
  FA_X1 mul_ex_mult_90_S1_11_0 ( .A(mul_ex_mult_90_ab_11__0_), .B(
        mul_ex_mult_90_CARRYB_10__0_), .CI(mul_ex_mult_90_SUMB_10__1_), .CO(
        mul_ex_mult_90_CARRYB_11__0_), .S(mul_ex_N165) );
  FA_X1 mul_ex_mult_90_S2_12_15 ( .A(mul_ex_mult_90_ab_12__15_), .B(
        mul_ex_mult_90_CARRYB_11__15_), .CI(mul_ex_mult_90_SUMB_11__16_), .CO(
        mul_ex_mult_90_CARRYB_12__15_), .S(mul_ex_mult_90_SUMB_12__15_) );
  FA_X1 mul_ex_mult_90_S2_12_14 ( .A(mul_ex_mult_90_ab_12__14_), .B(
        mul_ex_mult_90_CARRYB_11__14_), .CI(mul_ex_mult_90_SUMB_11__15_), .CO(
        mul_ex_mult_90_CARRYB_12__14_), .S(mul_ex_mult_90_SUMB_12__14_) );
  FA_X1 mul_ex_mult_90_S2_12_13 ( .A(mul_ex_mult_90_ab_12__13_), .B(
        mul_ex_mult_90_CARRYB_11__13_), .CI(mul_ex_mult_90_SUMB_11__14_), .CO(
        mul_ex_mult_90_CARRYB_12__13_), .S(mul_ex_mult_90_SUMB_12__13_) );
  FA_X1 mul_ex_mult_90_S2_12_12 ( .A(mul_ex_mult_90_ab_12__12_), .B(
        mul_ex_mult_90_CARRYB_11__12_), .CI(mul_ex_mult_90_SUMB_11__13_), .CO(
        mul_ex_mult_90_CARRYB_12__12_), .S(mul_ex_mult_90_SUMB_12__12_) );
  FA_X1 mul_ex_mult_90_S2_12_11 ( .A(mul_ex_mult_90_ab_12__11_), .B(
        mul_ex_mult_90_CARRYB_11__11_), .CI(mul_ex_mult_90_SUMB_11__12_), .CO(
        mul_ex_mult_90_CARRYB_12__11_), .S(mul_ex_mult_90_SUMB_12__11_) );
  FA_X1 mul_ex_mult_90_S2_12_10 ( .A(mul_ex_mult_90_ab_12__10_), .B(
        mul_ex_mult_90_CARRYB_11__10_), .CI(mul_ex_mult_90_SUMB_11__11_), .CO(
        mul_ex_mult_90_CARRYB_12__10_), .S(mul_ex_mult_90_SUMB_12__10_) );
  FA_X1 mul_ex_mult_90_S2_12_9 ( .A(mul_ex_mult_90_ab_12__9_), .B(
        mul_ex_mult_90_CARRYB_11__9_), .CI(mul_ex_mult_90_SUMB_11__10_), .CO(
        mul_ex_mult_90_CARRYB_12__9_), .S(mul_ex_mult_90_SUMB_12__9_) );
  FA_X1 mul_ex_mult_90_S2_12_8 ( .A(mul_ex_mult_90_ab_12__8_), .B(
        mul_ex_mult_90_CARRYB_11__8_), .CI(mul_ex_mult_90_SUMB_11__9_), .CO(
        mul_ex_mult_90_CARRYB_12__8_), .S(mul_ex_mult_90_SUMB_12__8_) );
  FA_X1 mul_ex_mult_90_S2_12_7 ( .A(mul_ex_mult_90_ab_12__7_), .B(
        mul_ex_mult_90_CARRYB_11__7_), .CI(mul_ex_mult_90_SUMB_11__8_), .CO(
        mul_ex_mult_90_CARRYB_12__7_), .S(mul_ex_mult_90_SUMB_12__7_) );
  FA_X1 mul_ex_mult_90_S2_12_6 ( .A(mul_ex_mult_90_ab_12__6_), .B(
        mul_ex_mult_90_CARRYB_11__6_), .CI(mul_ex_mult_90_SUMB_11__7_), .CO(
        mul_ex_mult_90_CARRYB_12__6_), .S(mul_ex_mult_90_SUMB_12__6_) );
  FA_X1 mul_ex_mult_90_S2_12_5 ( .A(mul_ex_mult_90_ab_12__5_), .B(
        mul_ex_mult_90_CARRYB_11__5_), .CI(mul_ex_mult_90_SUMB_11__6_), .CO(
        mul_ex_mult_90_CARRYB_12__5_), .S(mul_ex_mult_90_SUMB_12__5_) );
  FA_X1 mul_ex_mult_90_S2_12_4 ( .A(mul_ex_mult_90_ab_12__4_), .B(
        mul_ex_mult_90_CARRYB_11__4_), .CI(mul_ex_mult_90_SUMB_11__5_), .CO(
        mul_ex_mult_90_CARRYB_12__4_), .S(mul_ex_mult_90_SUMB_12__4_) );
  FA_X1 mul_ex_mult_90_S2_12_3 ( .A(mul_ex_mult_90_ab_12__3_), .B(
        mul_ex_mult_90_CARRYB_11__3_), .CI(mul_ex_mult_90_SUMB_11__4_), .CO(
        mul_ex_mult_90_CARRYB_12__3_), .S(mul_ex_mult_90_SUMB_12__3_) );
  FA_X1 mul_ex_mult_90_S2_12_2 ( .A(mul_ex_mult_90_ab_12__2_), .B(
        mul_ex_mult_90_CARRYB_11__2_), .CI(mul_ex_mult_90_SUMB_11__3_), .CO(
        mul_ex_mult_90_CARRYB_12__2_), .S(mul_ex_mult_90_SUMB_12__2_) );
  FA_X1 mul_ex_mult_90_S2_12_1 ( .A(mul_ex_mult_90_ab_12__1_), .B(
        mul_ex_mult_90_CARRYB_11__1_), .CI(mul_ex_mult_90_SUMB_11__2_), .CO(
        mul_ex_mult_90_CARRYB_12__1_), .S(mul_ex_mult_90_SUMB_12__1_) );
  FA_X1 mul_ex_mult_90_S1_12_0 ( .A(mul_ex_mult_90_ab_12__0_), .B(
        mul_ex_mult_90_CARRYB_11__0_), .CI(mul_ex_mult_90_SUMB_11__1_), .CO(
        mul_ex_mult_90_CARRYB_12__0_), .S(mul_ex_N166) );
  FA_X1 mul_ex_mult_90_S2_13_15 ( .A(mul_ex_mult_90_ab_13__15_), .B(
        mul_ex_mult_90_CARRYB_12__15_), .CI(mul_ex_mult_90_SUMB_12__16_), .CO(
        mul_ex_mult_90_CARRYB_13__15_), .S(mul_ex_mult_90_SUMB_13__15_) );
  FA_X1 mul_ex_mult_90_S2_13_14 ( .A(mul_ex_mult_90_ab_13__14_), .B(
        mul_ex_mult_90_CARRYB_12__14_), .CI(mul_ex_mult_90_SUMB_12__15_), .CO(
        mul_ex_mult_90_CARRYB_13__14_), .S(mul_ex_mult_90_SUMB_13__14_) );
  FA_X1 mul_ex_mult_90_S2_13_13 ( .A(mul_ex_mult_90_ab_13__13_), .B(
        mul_ex_mult_90_CARRYB_12__13_), .CI(mul_ex_mult_90_SUMB_12__14_), .CO(
        mul_ex_mult_90_CARRYB_13__13_), .S(mul_ex_mult_90_SUMB_13__13_) );
  FA_X1 mul_ex_mult_90_S2_13_12 ( .A(mul_ex_mult_90_ab_13__12_), .B(
        mul_ex_mult_90_CARRYB_12__12_), .CI(mul_ex_mult_90_SUMB_12__13_), .CO(
        mul_ex_mult_90_CARRYB_13__12_), .S(mul_ex_mult_90_SUMB_13__12_) );
  FA_X1 mul_ex_mult_90_S2_13_11 ( .A(mul_ex_mult_90_ab_13__11_), .B(
        mul_ex_mult_90_CARRYB_12__11_), .CI(mul_ex_mult_90_SUMB_12__12_), .CO(
        mul_ex_mult_90_CARRYB_13__11_), .S(mul_ex_mult_90_SUMB_13__11_) );
  FA_X1 mul_ex_mult_90_S2_13_10 ( .A(mul_ex_mult_90_ab_13__10_), .B(
        mul_ex_mult_90_CARRYB_12__10_), .CI(mul_ex_mult_90_SUMB_12__11_), .CO(
        mul_ex_mult_90_CARRYB_13__10_), .S(mul_ex_mult_90_SUMB_13__10_) );
  FA_X1 mul_ex_mult_90_S2_13_9 ( .A(mul_ex_mult_90_ab_13__9_), .B(
        mul_ex_mult_90_CARRYB_12__9_), .CI(mul_ex_mult_90_SUMB_12__10_), .CO(
        mul_ex_mult_90_CARRYB_13__9_), .S(mul_ex_mult_90_SUMB_13__9_) );
  FA_X1 mul_ex_mult_90_S2_13_8 ( .A(mul_ex_mult_90_ab_13__8_), .B(
        mul_ex_mult_90_CARRYB_12__8_), .CI(mul_ex_mult_90_SUMB_12__9_), .CO(
        mul_ex_mult_90_CARRYB_13__8_), .S(mul_ex_mult_90_SUMB_13__8_) );
  FA_X1 mul_ex_mult_90_S2_13_7 ( .A(mul_ex_mult_90_ab_13__7_), .B(
        mul_ex_mult_90_CARRYB_12__7_), .CI(mul_ex_mult_90_SUMB_12__8_), .CO(
        mul_ex_mult_90_CARRYB_13__7_), .S(mul_ex_mult_90_SUMB_13__7_) );
  FA_X1 mul_ex_mult_90_S2_13_6 ( .A(mul_ex_mult_90_ab_13__6_), .B(
        mul_ex_mult_90_CARRYB_12__6_), .CI(mul_ex_mult_90_SUMB_12__7_), .CO(
        mul_ex_mult_90_CARRYB_13__6_), .S(mul_ex_mult_90_SUMB_13__6_) );
  FA_X1 mul_ex_mult_90_S2_13_5 ( .A(mul_ex_mult_90_ab_13__5_), .B(
        mul_ex_mult_90_CARRYB_12__5_), .CI(mul_ex_mult_90_SUMB_12__6_), .CO(
        mul_ex_mult_90_CARRYB_13__5_), .S(mul_ex_mult_90_SUMB_13__5_) );
  FA_X1 mul_ex_mult_90_S2_13_4 ( .A(mul_ex_mult_90_ab_13__4_), .B(
        mul_ex_mult_90_CARRYB_12__4_), .CI(mul_ex_mult_90_SUMB_12__5_), .CO(
        mul_ex_mult_90_CARRYB_13__4_), .S(mul_ex_mult_90_SUMB_13__4_) );
  FA_X1 mul_ex_mult_90_S2_13_3 ( .A(mul_ex_mult_90_ab_13__3_), .B(
        mul_ex_mult_90_CARRYB_12__3_), .CI(mul_ex_mult_90_SUMB_12__4_), .CO(
        mul_ex_mult_90_CARRYB_13__3_), .S(mul_ex_mult_90_SUMB_13__3_) );
  FA_X1 mul_ex_mult_90_S2_13_2 ( .A(mul_ex_mult_90_ab_13__2_), .B(
        mul_ex_mult_90_CARRYB_12__2_), .CI(mul_ex_mult_90_SUMB_12__3_), .CO(
        mul_ex_mult_90_CARRYB_13__2_), .S(mul_ex_mult_90_SUMB_13__2_) );
  FA_X1 mul_ex_mult_90_S2_13_1 ( .A(mul_ex_mult_90_ab_13__1_), .B(
        mul_ex_mult_90_CARRYB_12__1_), .CI(mul_ex_mult_90_SUMB_12__2_), .CO(
        mul_ex_mult_90_CARRYB_13__1_), .S(mul_ex_mult_90_SUMB_13__1_) );
  FA_X1 mul_ex_mult_90_S1_13_0 ( .A(mul_ex_mult_90_ab_13__0_), .B(
        mul_ex_mult_90_CARRYB_12__0_), .CI(mul_ex_mult_90_SUMB_12__1_), .CO(
        mul_ex_mult_90_CARRYB_13__0_), .S(mul_ex_N167) );
  FA_X1 mul_ex_mult_90_S2_14_15 ( .A(mul_ex_mult_90_ab_14__15_), .B(
        mul_ex_mult_90_CARRYB_13__15_), .CI(mul_ex_mult_90_SUMB_13__16_), .CO(
        mul_ex_mult_90_CARRYB_14__15_), .S(mul_ex_mult_90_SUMB_14__15_) );
  FA_X1 mul_ex_mult_90_S2_14_14 ( .A(mul_ex_mult_90_ab_14__14_), .B(
        mul_ex_mult_90_CARRYB_13__14_), .CI(mul_ex_mult_90_SUMB_13__15_), .CO(
        mul_ex_mult_90_CARRYB_14__14_), .S(mul_ex_mult_90_SUMB_14__14_) );
  FA_X1 mul_ex_mult_90_S2_14_13 ( .A(mul_ex_mult_90_ab_14__13_), .B(
        mul_ex_mult_90_CARRYB_13__13_), .CI(mul_ex_mult_90_SUMB_13__14_), .CO(
        mul_ex_mult_90_CARRYB_14__13_), .S(mul_ex_mult_90_SUMB_14__13_) );
  FA_X1 mul_ex_mult_90_S2_14_12 ( .A(mul_ex_mult_90_ab_14__12_), .B(
        mul_ex_mult_90_CARRYB_13__12_), .CI(mul_ex_mult_90_SUMB_13__13_), .CO(
        mul_ex_mult_90_CARRYB_14__12_), .S(mul_ex_mult_90_SUMB_14__12_) );
  FA_X1 mul_ex_mult_90_S2_14_11 ( .A(mul_ex_mult_90_ab_14__11_), .B(
        mul_ex_mult_90_CARRYB_13__11_), .CI(mul_ex_mult_90_SUMB_13__12_), .CO(
        mul_ex_mult_90_CARRYB_14__11_), .S(mul_ex_mult_90_SUMB_14__11_) );
  FA_X1 mul_ex_mult_90_S2_14_10 ( .A(mul_ex_mult_90_ab_14__10_), .B(
        mul_ex_mult_90_CARRYB_13__10_), .CI(mul_ex_mult_90_SUMB_13__11_), .CO(
        mul_ex_mult_90_CARRYB_14__10_), .S(mul_ex_mult_90_SUMB_14__10_) );
  FA_X1 mul_ex_mult_90_S2_14_9 ( .A(mul_ex_mult_90_ab_14__9_), .B(
        mul_ex_mult_90_CARRYB_13__9_), .CI(mul_ex_mult_90_SUMB_13__10_), .CO(
        mul_ex_mult_90_CARRYB_14__9_), .S(mul_ex_mult_90_SUMB_14__9_) );
  FA_X1 mul_ex_mult_90_S2_14_8 ( .A(mul_ex_mult_90_ab_14__8_), .B(
        mul_ex_mult_90_CARRYB_13__8_), .CI(mul_ex_mult_90_SUMB_13__9_), .CO(
        mul_ex_mult_90_CARRYB_14__8_), .S(mul_ex_mult_90_SUMB_14__8_) );
  FA_X1 mul_ex_mult_90_S2_14_7 ( .A(mul_ex_mult_90_ab_14__7_), .B(
        mul_ex_mult_90_CARRYB_13__7_), .CI(mul_ex_mult_90_SUMB_13__8_), .CO(
        mul_ex_mult_90_CARRYB_14__7_), .S(mul_ex_mult_90_SUMB_14__7_) );
  FA_X1 mul_ex_mult_90_S2_14_6 ( .A(mul_ex_mult_90_ab_14__6_), .B(
        mul_ex_mult_90_CARRYB_13__6_), .CI(mul_ex_mult_90_SUMB_13__7_), .CO(
        mul_ex_mult_90_CARRYB_14__6_), .S(mul_ex_mult_90_SUMB_14__6_) );
  FA_X1 mul_ex_mult_90_S2_14_5 ( .A(mul_ex_mult_90_ab_14__5_), .B(
        mul_ex_mult_90_CARRYB_13__5_), .CI(mul_ex_mult_90_SUMB_13__6_), .CO(
        mul_ex_mult_90_CARRYB_14__5_), .S(mul_ex_mult_90_SUMB_14__5_) );
  FA_X1 mul_ex_mult_90_S2_14_4 ( .A(mul_ex_mult_90_ab_14__4_), .B(
        mul_ex_mult_90_CARRYB_13__4_), .CI(mul_ex_mult_90_SUMB_13__5_), .CO(
        mul_ex_mult_90_CARRYB_14__4_), .S(mul_ex_mult_90_SUMB_14__4_) );
  FA_X1 mul_ex_mult_90_S2_14_3 ( .A(mul_ex_mult_90_ab_14__3_), .B(
        mul_ex_mult_90_CARRYB_13__3_), .CI(mul_ex_mult_90_SUMB_13__4_), .CO(
        mul_ex_mult_90_CARRYB_14__3_), .S(mul_ex_mult_90_SUMB_14__3_) );
  FA_X1 mul_ex_mult_90_S2_14_2 ( .A(mul_ex_mult_90_ab_14__2_), .B(
        mul_ex_mult_90_CARRYB_13__2_), .CI(mul_ex_mult_90_SUMB_13__3_), .CO(
        mul_ex_mult_90_CARRYB_14__2_), .S(mul_ex_mult_90_SUMB_14__2_) );
  FA_X1 mul_ex_mult_90_S2_14_1 ( .A(mul_ex_mult_90_ab_14__1_), .B(
        mul_ex_mult_90_CARRYB_13__1_), .CI(mul_ex_mult_90_SUMB_13__2_), .CO(
        mul_ex_mult_90_CARRYB_14__1_), .S(mul_ex_mult_90_SUMB_14__1_) );
  FA_X1 mul_ex_mult_90_S1_14_0 ( .A(mul_ex_mult_90_ab_14__0_), .B(
        mul_ex_mult_90_CARRYB_13__0_), .CI(mul_ex_mult_90_SUMB_13__1_), .CO(
        mul_ex_mult_90_CARRYB_14__0_), .S(mul_ex_N168) );
  FA_X1 mul_ex_mult_90_S2_15_15 ( .A(mul_ex_mult_90_ab_15__15_), .B(
        mul_ex_mult_90_CARRYB_14__15_), .CI(mul_ex_mult_90_SUMB_14__16_), .CO(
        mul_ex_mult_90_CARRYB_15__15_), .S(mul_ex_mult_90_SUMB_15__15_) );
  FA_X1 mul_ex_mult_90_S2_15_14 ( .A(mul_ex_mult_90_ab_15__14_), .B(
        mul_ex_mult_90_CARRYB_14__14_), .CI(mul_ex_mult_90_SUMB_14__15_), .CO(
        mul_ex_mult_90_CARRYB_15__14_), .S(mul_ex_mult_90_SUMB_15__14_) );
  FA_X1 mul_ex_mult_90_S2_15_13 ( .A(mul_ex_mult_90_ab_15__13_), .B(
        mul_ex_mult_90_CARRYB_14__13_), .CI(mul_ex_mult_90_SUMB_14__14_), .CO(
        mul_ex_mult_90_CARRYB_15__13_), .S(mul_ex_mult_90_SUMB_15__13_) );
  FA_X1 mul_ex_mult_90_S2_15_12 ( .A(mul_ex_mult_90_ab_15__12_), .B(
        mul_ex_mult_90_CARRYB_14__12_), .CI(mul_ex_mult_90_SUMB_14__13_), .CO(
        mul_ex_mult_90_CARRYB_15__12_), .S(mul_ex_mult_90_SUMB_15__12_) );
  FA_X1 mul_ex_mult_90_S2_15_11 ( .A(mul_ex_mult_90_ab_15__11_), .B(
        mul_ex_mult_90_CARRYB_14__11_), .CI(mul_ex_mult_90_SUMB_14__12_), .CO(
        mul_ex_mult_90_CARRYB_15__11_), .S(mul_ex_mult_90_SUMB_15__11_) );
  FA_X1 mul_ex_mult_90_S2_15_10 ( .A(mul_ex_mult_90_ab_15__10_), .B(
        mul_ex_mult_90_CARRYB_14__10_), .CI(mul_ex_mult_90_SUMB_14__11_), .CO(
        mul_ex_mult_90_CARRYB_15__10_), .S(mul_ex_mult_90_SUMB_15__10_) );
  FA_X1 mul_ex_mult_90_S2_15_9 ( .A(mul_ex_mult_90_ab_15__9_), .B(
        mul_ex_mult_90_CARRYB_14__9_), .CI(mul_ex_mult_90_SUMB_14__10_), .CO(
        mul_ex_mult_90_CARRYB_15__9_), .S(mul_ex_mult_90_SUMB_15__9_) );
  FA_X1 mul_ex_mult_90_S2_15_8 ( .A(mul_ex_mult_90_ab_15__8_), .B(
        mul_ex_mult_90_CARRYB_14__8_), .CI(mul_ex_mult_90_SUMB_14__9_), .CO(
        mul_ex_mult_90_CARRYB_15__8_), .S(mul_ex_mult_90_SUMB_15__8_) );
  FA_X1 mul_ex_mult_90_S2_15_7 ( .A(mul_ex_mult_90_ab_15__7_), .B(
        mul_ex_mult_90_CARRYB_14__7_), .CI(mul_ex_mult_90_SUMB_14__8_), .CO(
        mul_ex_mult_90_CARRYB_15__7_), .S(mul_ex_mult_90_SUMB_15__7_) );
  FA_X1 mul_ex_mult_90_S2_15_6 ( .A(mul_ex_mult_90_ab_15__6_), .B(
        mul_ex_mult_90_CARRYB_14__6_), .CI(mul_ex_mult_90_SUMB_14__7_), .CO(
        mul_ex_mult_90_CARRYB_15__6_), .S(mul_ex_mult_90_SUMB_15__6_) );
  FA_X1 mul_ex_mult_90_S2_15_5 ( .A(mul_ex_mult_90_ab_15__5_), .B(
        mul_ex_mult_90_CARRYB_14__5_), .CI(mul_ex_mult_90_SUMB_14__6_), .CO(
        mul_ex_mult_90_CARRYB_15__5_), .S(mul_ex_mult_90_SUMB_15__5_) );
  FA_X1 mul_ex_mult_90_S2_15_4 ( .A(mul_ex_mult_90_ab_15__4_), .B(
        mul_ex_mult_90_CARRYB_14__4_), .CI(mul_ex_mult_90_SUMB_14__5_), .CO(
        mul_ex_mult_90_CARRYB_15__4_), .S(mul_ex_mult_90_SUMB_15__4_) );
  FA_X1 mul_ex_mult_90_S2_15_3 ( .A(mul_ex_mult_90_ab_15__3_), .B(
        mul_ex_mult_90_CARRYB_14__3_), .CI(mul_ex_mult_90_SUMB_14__4_), .CO(
        mul_ex_mult_90_CARRYB_15__3_), .S(mul_ex_mult_90_SUMB_15__3_) );
  FA_X1 mul_ex_mult_90_S2_15_2 ( .A(mul_ex_mult_90_ab_15__2_), .B(
        mul_ex_mult_90_CARRYB_14__2_), .CI(mul_ex_mult_90_SUMB_14__3_), .CO(
        mul_ex_mult_90_CARRYB_15__2_), .S(mul_ex_mult_90_SUMB_15__2_) );
  FA_X1 mul_ex_mult_90_S2_15_1 ( .A(mul_ex_mult_90_ab_15__1_), .B(
        mul_ex_mult_90_CARRYB_14__1_), .CI(mul_ex_mult_90_SUMB_14__2_), .CO(
        mul_ex_mult_90_CARRYB_15__1_), .S(mul_ex_mult_90_SUMB_15__1_) );
  FA_X1 mul_ex_mult_90_S1_15_0 ( .A(mul_ex_mult_90_ab_15__0_), .B(
        mul_ex_mult_90_CARRYB_14__0_), .CI(mul_ex_mult_90_SUMB_14__1_), .CO(
        mul_ex_mult_90_CARRYB_15__0_), .S(mul_ex_N169) );
  FA_X1 mul_ex_mult_90_S2_16_15 ( .A(mul_ex_mult_90_ab_16__15_), .B(
        mul_ex_mult_90_CARRYB_15__15_), .CI(mul_ex_mult_90_SUMB_15__16_), .S(
        mul_ex_mult_90_SUMB_16__15_) );
  FA_X1 mul_ex_mult_90_S2_16_14 ( .A(mul_ex_mult_90_ab_16__14_), .B(
        mul_ex_mult_90_CARRYB_15__14_), .CI(mul_ex_mult_90_SUMB_15__15_), .CO(
        mul_ex_mult_90_CARRYB_16__14_), .S(mul_ex_mult_90_SUMB_16__14_) );
  FA_X1 mul_ex_mult_90_S2_16_13 ( .A(mul_ex_mult_90_ab_16__13_), .B(
        mul_ex_mult_90_CARRYB_15__13_), .CI(mul_ex_mult_90_SUMB_15__14_), .CO(
        mul_ex_mult_90_CARRYB_16__13_), .S(mul_ex_mult_90_SUMB_16__13_) );
  FA_X1 mul_ex_mult_90_S2_16_12 ( .A(mul_ex_mult_90_ab_16__12_), .B(
        mul_ex_mult_90_CARRYB_15__12_), .CI(mul_ex_mult_90_SUMB_15__13_), .CO(
        mul_ex_mult_90_CARRYB_16__12_), .S(mul_ex_mult_90_SUMB_16__12_) );
  FA_X1 mul_ex_mult_90_S2_16_11 ( .A(mul_ex_mult_90_ab_16__11_), .B(
        mul_ex_mult_90_CARRYB_15__11_), .CI(mul_ex_mult_90_SUMB_15__12_), .CO(
        mul_ex_mult_90_CARRYB_16__11_), .S(mul_ex_mult_90_SUMB_16__11_) );
  FA_X1 mul_ex_mult_90_S2_16_10 ( .A(mul_ex_mult_90_ab_16__10_), .B(
        mul_ex_mult_90_CARRYB_15__10_), .CI(mul_ex_mult_90_SUMB_15__11_), .CO(
        mul_ex_mult_90_CARRYB_16__10_), .S(mul_ex_mult_90_SUMB_16__10_) );
  FA_X1 mul_ex_mult_90_S2_16_9 ( .A(mul_ex_mult_90_ab_16__9_), .B(
        mul_ex_mult_90_CARRYB_15__9_), .CI(mul_ex_mult_90_SUMB_15__10_), .CO(
        mul_ex_mult_90_CARRYB_16__9_), .S(mul_ex_mult_90_SUMB_16__9_) );
  FA_X1 mul_ex_mult_90_S2_16_8 ( .A(mul_ex_mult_90_ab_16__8_), .B(
        mul_ex_mult_90_CARRYB_15__8_), .CI(mul_ex_mult_90_SUMB_15__9_), .CO(
        mul_ex_mult_90_CARRYB_16__8_), .S(mul_ex_mult_90_SUMB_16__8_) );
  FA_X1 mul_ex_mult_90_S2_16_7 ( .A(mul_ex_mult_90_ab_16__7_), .B(
        mul_ex_mult_90_CARRYB_15__7_), .CI(mul_ex_mult_90_SUMB_15__8_), .CO(
        mul_ex_mult_90_CARRYB_16__7_), .S(mul_ex_mult_90_SUMB_16__7_) );
  FA_X1 mul_ex_mult_90_S2_16_6 ( .A(mul_ex_mult_90_ab_16__6_), .B(
        mul_ex_mult_90_CARRYB_15__6_), .CI(mul_ex_mult_90_SUMB_15__7_), .CO(
        mul_ex_mult_90_CARRYB_16__6_), .S(mul_ex_mult_90_SUMB_16__6_) );
  FA_X1 mul_ex_mult_90_S2_16_5 ( .A(mul_ex_mult_90_ab_16__5_), .B(
        mul_ex_mult_90_CARRYB_15__5_), .CI(mul_ex_mult_90_SUMB_15__6_), .CO(
        mul_ex_mult_90_CARRYB_16__5_), .S(mul_ex_mult_90_SUMB_16__5_) );
  FA_X1 mul_ex_mult_90_S2_16_4 ( .A(mul_ex_mult_90_ab_16__4_), .B(
        mul_ex_mult_90_CARRYB_15__4_), .CI(mul_ex_mult_90_SUMB_15__5_), .CO(
        mul_ex_mult_90_CARRYB_16__4_), .S(mul_ex_mult_90_SUMB_16__4_) );
  FA_X1 mul_ex_mult_90_S2_16_3 ( .A(mul_ex_mult_90_ab_16__3_), .B(
        mul_ex_mult_90_CARRYB_15__3_), .CI(mul_ex_mult_90_SUMB_15__4_), .CO(
        mul_ex_mult_90_CARRYB_16__3_), .S(mul_ex_mult_90_SUMB_16__3_) );
  FA_X1 mul_ex_mult_90_S2_16_2 ( .A(mul_ex_mult_90_ab_16__2_), .B(
        mul_ex_mult_90_CARRYB_15__2_), .CI(mul_ex_mult_90_SUMB_15__3_), .CO(
        mul_ex_mult_90_CARRYB_16__2_), .S(mul_ex_mult_90_SUMB_16__2_) );
  FA_X1 mul_ex_mult_90_S2_16_1 ( .A(mul_ex_mult_90_ab_16__1_), .B(
        mul_ex_mult_90_CARRYB_15__1_), .CI(mul_ex_mult_90_SUMB_15__2_), .CO(
        mul_ex_mult_90_CARRYB_16__1_), .S(mul_ex_mult_90_SUMB_16__1_) );
  FA_X1 mul_ex_mult_90_S1_16_0 ( .A(mul_ex_mult_90_ab_16__0_), .B(
        mul_ex_mult_90_CARRYB_15__0_), .CI(mul_ex_mult_90_SUMB_15__1_), .CO(
        mul_ex_mult_90_CARRYB_16__0_), .S(mul_ex_N170) );
  NOR2_X1 mul_ex_mult_76_U350 ( .A1(mul_ex_mult_76_n94), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_N56) );
  NOR2_X1 mul_ex_mult_76_U349 ( .A1(mul_ex_mult_76_n84), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_mult_76_ab_0__10_) );
  NOR2_X1 mul_ex_mult_76_U348 ( .A1(mul_ex_mult_76_n83), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_mult_76_ab_0__11_) );
  NOR2_X1 mul_ex_mult_76_U347 ( .A1(mul_ex_mult_76_n82), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_mult_76_ab_0__12_) );
  NOR2_X1 mul_ex_mult_76_U346 ( .A1(mul_ex_mult_76_n81), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_mult_76_ab_0__13_) );
  NOR2_X1 mul_ex_mult_76_U345 ( .A1(mul_ex_mult_76_n80), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_mult_76_ab_0__14_) );
  NOR2_X1 mul_ex_mult_76_U344 ( .A1(mul_ex_mult_76_n79), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_mult_76_ab_0__15_) );
  NOR2_X1 mul_ex_mult_76_U343 ( .A1(mul_ex_mult_76_n93), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_mult_76_ab_0__1_) );
  NOR2_X1 mul_ex_mult_76_U342 ( .A1(mul_ex_mult_76_n92), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_mult_76_ab_0__2_) );
  NOR2_X1 mul_ex_mult_76_U341 ( .A1(mul_ex_mult_76_n91), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_mult_76_ab_0__3_) );
  NOR2_X1 mul_ex_mult_76_U340 ( .A1(mul_ex_mult_76_n90), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_mult_76_ab_0__4_) );
  NOR2_X1 mul_ex_mult_76_U339 ( .A1(mul_ex_mult_76_n89), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_mult_76_ab_0__5_) );
  NOR2_X1 mul_ex_mult_76_U338 ( .A1(mul_ex_mult_76_n88), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_mult_76_ab_0__6_) );
  NOR2_X1 mul_ex_mult_76_U337 ( .A1(mul_ex_mult_76_n87), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_mult_76_ab_0__7_) );
  NOR2_X1 mul_ex_mult_76_U336 ( .A1(mul_ex_mult_76_n86), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_mult_76_ab_0__8_) );
  NOR2_X1 mul_ex_mult_76_U335 ( .A1(mul_ex_mult_76_n85), .A2(
        mul_ex_mult_76_n78), .ZN(mul_ex_mult_76_ab_0__9_) );
  NOR2_X1 mul_ex_mult_76_U334 ( .A1(mul_ex_mult_76_n94), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__0_) );
  NOR2_X1 mul_ex_mult_76_U333 ( .A1(mul_ex_mult_76_n84), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__10_) );
  NOR2_X1 mul_ex_mult_76_U332 ( .A1(mul_ex_mult_76_n83), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__11_) );
  NOR2_X1 mul_ex_mult_76_U331 ( .A1(mul_ex_mult_76_n82), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__12_) );
  NOR2_X1 mul_ex_mult_76_U330 ( .A1(mul_ex_mult_76_n81), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__13_) );
  NOR2_X1 mul_ex_mult_76_U329 ( .A1(mul_ex_mult_76_n80), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__14_) );
  NOR2_X1 mul_ex_mult_76_U328 ( .A1(mul_ex_mult_76_n79), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__15_) );
  NOR2_X1 mul_ex_mult_76_U327 ( .A1(mul_ex_mult_76_n93), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__1_) );
  NOR2_X1 mul_ex_mult_76_U326 ( .A1(mul_ex_mult_76_n92), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__2_) );
  NOR2_X1 mul_ex_mult_76_U325 ( .A1(mul_ex_mult_76_n91), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__3_) );
  NOR2_X1 mul_ex_mult_76_U324 ( .A1(mul_ex_mult_76_n90), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__4_) );
  NOR2_X1 mul_ex_mult_76_U323 ( .A1(mul_ex_mult_76_n89), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__5_) );
  NOR2_X1 mul_ex_mult_76_U322 ( .A1(mul_ex_mult_76_n88), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__6_) );
  NOR2_X1 mul_ex_mult_76_U321 ( .A1(mul_ex_mult_76_n87), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__7_) );
  NOR2_X1 mul_ex_mult_76_U320 ( .A1(mul_ex_mult_76_n86), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__8_) );
  NOR2_X1 mul_ex_mult_76_U319 ( .A1(mul_ex_mult_76_n85), .A2(
        mul_ex_mult_76_n68), .ZN(mul_ex_mult_76_ab_10__9_) );
  NOR2_X1 mul_ex_mult_76_U318 ( .A1(mul_ex_mult_76_n94), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__0_) );
  NOR2_X1 mul_ex_mult_76_U317 ( .A1(mul_ex_mult_76_n84), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__10_) );
  NOR2_X1 mul_ex_mult_76_U316 ( .A1(mul_ex_mult_76_n83), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__11_) );
  NOR2_X1 mul_ex_mult_76_U315 ( .A1(mul_ex_mult_76_n82), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__12_) );
  NOR2_X1 mul_ex_mult_76_U314 ( .A1(mul_ex_mult_76_n81), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__13_) );
  NOR2_X1 mul_ex_mult_76_U313 ( .A1(mul_ex_mult_76_n80), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__14_) );
  NOR2_X1 mul_ex_mult_76_U312 ( .A1(mul_ex_mult_76_n79), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__15_) );
  NOR2_X1 mul_ex_mult_76_U311 ( .A1(mul_ex_mult_76_n93), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__1_) );
  NOR2_X1 mul_ex_mult_76_U310 ( .A1(mul_ex_mult_76_n92), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__2_) );
  NOR2_X1 mul_ex_mult_76_U309 ( .A1(mul_ex_mult_76_n91), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__3_) );
  NOR2_X1 mul_ex_mult_76_U308 ( .A1(mul_ex_mult_76_n90), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__4_) );
  NOR2_X1 mul_ex_mult_76_U307 ( .A1(mul_ex_mult_76_n89), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__5_) );
  NOR2_X1 mul_ex_mult_76_U306 ( .A1(mul_ex_mult_76_n88), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__6_) );
  NOR2_X1 mul_ex_mult_76_U305 ( .A1(mul_ex_mult_76_n87), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__7_) );
  NOR2_X1 mul_ex_mult_76_U304 ( .A1(mul_ex_mult_76_n86), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__8_) );
  NOR2_X1 mul_ex_mult_76_U303 ( .A1(mul_ex_mult_76_n85), .A2(
        mul_ex_mult_76_n67), .ZN(mul_ex_mult_76_ab_11__9_) );
  NOR2_X1 mul_ex_mult_76_U302 ( .A1(mul_ex_mult_76_n94), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__0_) );
  NOR2_X1 mul_ex_mult_76_U301 ( .A1(mul_ex_mult_76_n84), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__10_) );
  NOR2_X1 mul_ex_mult_76_U300 ( .A1(mul_ex_mult_76_n83), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__11_) );
  NOR2_X1 mul_ex_mult_76_U299 ( .A1(mul_ex_mult_76_n82), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__12_) );
  NOR2_X1 mul_ex_mult_76_U298 ( .A1(mul_ex_mult_76_n81), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__13_) );
  NOR2_X1 mul_ex_mult_76_U297 ( .A1(mul_ex_mult_76_n80), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__14_) );
  NOR2_X1 mul_ex_mult_76_U296 ( .A1(mul_ex_mult_76_n79), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__15_) );
  NOR2_X1 mul_ex_mult_76_U295 ( .A1(mul_ex_mult_76_n93), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__1_) );
  NOR2_X1 mul_ex_mult_76_U294 ( .A1(mul_ex_mult_76_n92), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__2_) );
  NOR2_X1 mul_ex_mult_76_U293 ( .A1(mul_ex_mult_76_n91), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__3_) );
  NOR2_X1 mul_ex_mult_76_U292 ( .A1(mul_ex_mult_76_n90), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__4_) );
  NOR2_X1 mul_ex_mult_76_U291 ( .A1(mul_ex_mult_76_n89), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__5_) );
  NOR2_X1 mul_ex_mult_76_U290 ( .A1(mul_ex_mult_76_n88), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__6_) );
  NOR2_X1 mul_ex_mult_76_U289 ( .A1(mul_ex_mult_76_n87), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__7_) );
  NOR2_X1 mul_ex_mult_76_U288 ( .A1(mul_ex_mult_76_n86), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__8_) );
  NOR2_X1 mul_ex_mult_76_U287 ( .A1(mul_ex_mult_76_n85), .A2(
        mul_ex_mult_76_n66), .ZN(mul_ex_mult_76_ab_12__9_) );
  NOR2_X1 mul_ex_mult_76_U286 ( .A1(mul_ex_mult_76_n94), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__0_) );
  NOR2_X1 mul_ex_mult_76_U285 ( .A1(mul_ex_mult_76_n84), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__10_) );
  NOR2_X1 mul_ex_mult_76_U284 ( .A1(mul_ex_mult_76_n83), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__11_) );
  NOR2_X1 mul_ex_mult_76_U283 ( .A1(mul_ex_mult_76_n82), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__12_) );
  NOR2_X1 mul_ex_mult_76_U282 ( .A1(mul_ex_mult_76_n81), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__13_) );
  NOR2_X1 mul_ex_mult_76_U281 ( .A1(mul_ex_mult_76_n80), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__14_) );
  NOR2_X1 mul_ex_mult_76_U280 ( .A1(mul_ex_mult_76_n79), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__15_) );
  NOR2_X1 mul_ex_mult_76_U279 ( .A1(mul_ex_mult_76_n93), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__1_) );
  NOR2_X1 mul_ex_mult_76_U278 ( .A1(mul_ex_mult_76_n92), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__2_) );
  NOR2_X1 mul_ex_mult_76_U277 ( .A1(mul_ex_mult_76_n91), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__3_) );
  NOR2_X1 mul_ex_mult_76_U276 ( .A1(mul_ex_mult_76_n90), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__4_) );
  NOR2_X1 mul_ex_mult_76_U275 ( .A1(mul_ex_mult_76_n89), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__5_) );
  NOR2_X1 mul_ex_mult_76_U274 ( .A1(mul_ex_mult_76_n88), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__6_) );
  NOR2_X1 mul_ex_mult_76_U273 ( .A1(mul_ex_mult_76_n87), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__7_) );
  NOR2_X1 mul_ex_mult_76_U272 ( .A1(mul_ex_mult_76_n86), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__8_) );
  NOR2_X1 mul_ex_mult_76_U271 ( .A1(mul_ex_mult_76_n85), .A2(
        mul_ex_mult_76_n65), .ZN(mul_ex_mult_76_ab_13__9_) );
  NOR2_X1 mul_ex_mult_76_U270 ( .A1(mul_ex_mult_76_n94), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__0_) );
  NOR2_X1 mul_ex_mult_76_U269 ( .A1(mul_ex_mult_76_n84), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__10_) );
  NOR2_X1 mul_ex_mult_76_U268 ( .A1(mul_ex_mult_76_n83), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__11_) );
  NOR2_X1 mul_ex_mult_76_U267 ( .A1(mul_ex_mult_76_n82), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__12_) );
  NOR2_X1 mul_ex_mult_76_U266 ( .A1(mul_ex_mult_76_n81), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__13_) );
  NOR2_X1 mul_ex_mult_76_U265 ( .A1(mul_ex_mult_76_n80), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__14_) );
  NOR2_X1 mul_ex_mult_76_U264 ( .A1(mul_ex_mult_76_n79), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__15_) );
  NOR2_X1 mul_ex_mult_76_U263 ( .A1(mul_ex_mult_76_n93), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__1_) );
  NOR2_X1 mul_ex_mult_76_U262 ( .A1(mul_ex_mult_76_n92), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__2_) );
  NOR2_X1 mul_ex_mult_76_U261 ( .A1(mul_ex_mult_76_n91), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__3_) );
  NOR2_X1 mul_ex_mult_76_U260 ( .A1(mul_ex_mult_76_n90), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__4_) );
  NOR2_X1 mul_ex_mult_76_U259 ( .A1(mul_ex_mult_76_n89), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__5_) );
  NOR2_X1 mul_ex_mult_76_U258 ( .A1(mul_ex_mult_76_n88), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__6_) );
  NOR2_X1 mul_ex_mult_76_U257 ( .A1(mul_ex_mult_76_n87), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__7_) );
  NOR2_X1 mul_ex_mult_76_U256 ( .A1(mul_ex_mult_76_n86), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__8_) );
  NOR2_X1 mul_ex_mult_76_U255 ( .A1(mul_ex_mult_76_n85), .A2(
        mul_ex_mult_76_n64), .ZN(mul_ex_mult_76_ab_14__9_) );
  NOR2_X1 mul_ex_mult_76_U254 ( .A1(mul_ex_mult_76_n94), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__0_) );
  NOR2_X1 mul_ex_mult_76_U253 ( .A1(mul_ex_mult_76_n84), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__10_) );
  NOR2_X1 mul_ex_mult_76_U252 ( .A1(mul_ex_mult_76_n83), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__11_) );
  NOR2_X1 mul_ex_mult_76_U251 ( .A1(mul_ex_mult_76_n82), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__12_) );
  NOR2_X1 mul_ex_mult_76_U250 ( .A1(mul_ex_mult_76_n81), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__13_) );
  NOR2_X1 mul_ex_mult_76_U249 ( .A1(mul_ex_mult_76_n80), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__14_) );
  NOR2_X1 mul_ex_mult_76_U248 ( .A1(mul_ex_mult_76_n79), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__15_) );
  NOR2_X1 mul_ex_mult_76_U247 ( .A1(mul_ex_mult_76_n93), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__1_) );
  NOR2_X1 mul_ex_mult_76_U246 ( .A1(mul_ex_mult_76_n92), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__2_) );
  NOR2_X1 mul_ex_mult_76_U245 ( .A1(mul_ex_mult_76_n91), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__3_) );
  NOR2_X1 mul_ex_mult_76_U244 ( .A1(mul_ex_mult_76_n90), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__4_) );
  NOR2_X1 mul_ex_mult_76_U243 ( .A1(mul_ex_mult_76_n89), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__5_) );
  NOR2_X1 mul_ex_mult_76_U242 ( .A1(mul_ex_mult_76_n88), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__6_) );
  NOR2_X1 mul_ex_mult_76_U241 ( .A1(mul_ex_mult_76_n87), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__7_) );
  NOR2_X1 mul_ex_mult_76_U240 ( .A1(mul_ex_mult_76_n86), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__8_) );
  NOR2_X1 mul_ex_mult_76_U239 ( .A1(mul_ex_mult_76_n85), .A2(
        mul_ex_mult_76_n63), .ZN(mul_ex_mult_76_ab_15__9_) );
  NOR2_X1 mul_ex_mult_76_U238 ( .A1(mul_ex_mult_76_n94), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__0_) );
  NOR2_X1 mul_ex_mult_76_U237 ( .A1(mul_ex_mult_76_n84), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__10_) );
  NOR2_X1 mul_ex_mult_76_U236 ( .A1(mul_ex_mult_76_n83), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__11_) );
  NOR2_X1 mul_ex_mult_76_U235 ( .A1(mul_ex_mult_76_n82), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__12_) );
  NOR2_X1 mul_ex_mult_76_U234 ( .A1(mul_ex_mult_76_n81), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__13_) );
  NOR2_X1 mul_ex_mult_76_U233 ( .A1(mul_ex_mult_76_n80), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__14_) );
  NOR2_X1 mul_ex_mult_76_U232 ( .A1(mul_ex_mult_76_n79), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__15_) );
  NOR2_X1 mul_ex_mult_76_U231 ( .A1(mul_ex_mult_76_n93), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__1_) );
  NOR2_X1 mul_ex_mult_76_U230 ( .A1(mul_ex_mult_76_n92), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__2_) );
  NOR2_X1 mul_ex_mult_76_U229 ( .A1(mul_ex_mult_76_n91), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__3_) );
  NOR2_X1 mul_ex_mult_76_U228 ( .A1(mul_ex_mult_76_n90), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__4_) );
  NOR2_X1 mul_ex_mult_76_U227 ( .A1(mul_ex_mult_76_n89), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__5_) );
  NOR2_X1 mul_ex_mult_76_U226 ( .A1(mul_ex_mult_76_n88), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__6_) );
  NOR2_X1 mul_ex_mult_76_U225 ( .A1(mul_ex_mult_76_n87), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__7_) );
  NOR2_X1 mul_ex_mult_76_U224 ( .A1(mul_ex_mult_76_n86), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__8_) );
  NOR2_X1 mul_ex_mult_76_U223 ( .A1(mul_ex_mult_76_n85), .A2(
        mul_ex_mult_76_n77), .ZN(mul_ex_mult_76_ab_1__9_) );
  NOR2_X1 mul_ex_mult_76_U222 ( .A1(mul_ex_mult_76_n94), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__0_) );
  NOR2_X1 mul_ex_mult_76_U221 ( .A1(mul_ex_mult_76_n84), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__10_) );
  NOR2_X1 mul_ex_mult_76_U220 ( .A1(mul_ex_mult_76_n83), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__11_) );
  NOR2_X1 mul_ex_mult_76_U219 ( .A1(mul_ex_mult_76_n82), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__12_) );
  NOR2_X1 mul_ex_mult_76_U218 ( .A1(mul_ex_mult_76_n81), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__13_) );
  NOR2_X1 mul_ex_mult_76_U217 ( .A1(mul_ex_mult_76_n80), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__14_) );
  NOR2_X1 mul_ex_mult_76_U216 ( .A1(mul_ex_mult_76_n79), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__15_) );
  NOR2_X1 mul_ex_mult_76_U215 ( .A1(mul_ex_mult_76_n93), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__1_) );
  NOR2_X1 mul_ex_mult_76_U214 ( .A1(mul_ex_mult_76_n92), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__2_) );
  NOR2_X1 mul_ex_mult_76_U213 ( .A1(mul_ex_mult_76_n91), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__3_) );
  NOR2_X1 mul_ex_mult_76_U212 ( .A1(mul_ex_mult_76_n90), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__4_) );
  NOR2_X1 mul_ex_mult_76_U211 ( .A1(mul_ex_mult_76_n89), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__5_) );
  NOR2_X1 mul_ex_mult_76_U210 ( .A1(mul_ex_mult_76_n88), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__6_) );
  NOR2_X1 mul_ex_mult_76_U209 ( .A1(mul_ex_mult_76_n87), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__7_) );
  NOR2_X1 mul_ex_mult_76_U208 ( .A1(mul_ex_mult_76_n86), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__8_) );
  NOR2_X1 mul_ex_mult_76_U207 ( .A1(mul_ex_mult_76_n85), .A2(
        mul_ex_mult_76_n76), .ZN(mul_ex_mult_76_ab_2__9_) );
  NOR2_X1 mul_ex_mult_76_U206 ( .A1(mul_ex_mult_76_n94), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__0_) );
  NOR2_X1 mul_ex_mult_76_U205 ( .A1(mul_ex_mult_76_n84), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__10_) );
  NOR2_X1 mul_ex_mult_76_U204 ( .A1(mul_ex_mult_76_n83), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__11_) );
  NOR2_X1 mul_ex_mult_76_U203 ( .A1(mul_ex_mult_76_n82), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__12_) );
  NOR2_X1 mul_ex_mult_76_U202 ( .A1(mul_ex_mult_76_n81), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__13_) );
  NOR2_X1 mul_ex_mult_76_U201 ( .A1(mul_ex_mult_76_n80), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__14_) );
  NOR2_X1 mul_ex_mult_76_U200 ( .A1(mul_ex_mult_76_n79), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__15_) );
  NOR2_X1 mul_ex_mult_76_U199 ( .A1(mul_ex_mult_76_n93), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__1_) );
  NOR2_X1 mul_ex_mult_76_U198 ( .A1(mul_ex_mult_76_n92), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__2_) );
  NOR2_X1 mul_ex_mult_76_U197 ( .A1(mul_ex_mult_76_n91), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__3_) );
  NOR2_X1 mul_ex_mult_76_U196 ( .A1(mul_ex_mult_76_n90), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__4_) );
  NOR2_X1 mul_ex_mult_76_U195 ( .A1(mul_ex_mult_76_n89), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__5_) );
  NOR2_X1 mul_ex_mult_76_U194 ( .A1(mul_ex_mult_76_n88), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__6_) );
  NOR2_X1 mul_ex_mult_76_U193 ( .A1(mul_ex_mult_76_n87), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__7_) );
  NOR2_X1 mul_ex_mult_76_U192 ( .A1(mul_ex_mult_76_n86), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__8_) );
  NOR2_X1 mul_ex_mult_76_U191 ( .A1(mul_ex_mult_76_n85), .A2(
        mul_ex_mult_76_n75), .ZN(mul_ex_mult_76_ab_3__9_) );
  NOR2_X1 mul_ex_mult_76_U190 ( .A1(mul_ex_mult_76_n94), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__0_) );
  NOR2_X1 mul_ex_mult_76_U189 ( .A1(mul_ex_mult_76_n84), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__10_) );
  NOR2_X1 mul_ex_mult_76_U188 ( .A1(mul_ex_mult_76_n83), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__11_) );
  NOR2_X1 mul_ex_mult_76_U187 ( .A1(mul_ex_mult_76_n82), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__12_) );
  NOR2_X1 mul_ex_mult_76_U186 ( .A1(mul_ex_mult_76_n81), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__13_) );
  NOR2_X1 mul_ex_mult_76_U185 ( .A1(mul_ex_mult_76_n80), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__14_) );
  NOR2_X1 mul_ex_mult_76_U184 ( .A1(mul_ex_mult_76_n79), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__15_) );
  NOR2_X1 mul_ex_mult_76_U183 ( .A1(mul_ex_mult_76_n93), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__1_) );
  NOR2_X1 mul_ex_mult_76_U182 ( .A1(mul_ex_mult_76_n92), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__2_) );
  NOR2_X1 mul_ex_mult_76_U181 ( .A1(mul_ex_mult_76_n91), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__3_) );
  NOR2_X1 mul_ex_mult_76_U180 ( .A1(mul_ex_mult_76_n90), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__4_) );
  NOR2_X1 mul_ex_mult_76_U179 ( .A1(mul_ex_mult_76_n89), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__5_) );
  NOR2_X1 mul_ex_mult_76_U178 ( .A1(mul_ex_mult_76_n88), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__6_) );
  NOR2_X1 mul_ex_mult_76_U177 ( .A1(mul_ex_mult_76_n87), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__7_) );
  NOR2_X1 mul_ex_mult_76_U176 ( .A1(mul_ex_mult_76_n86), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__8_) );
  NOR2_X1 mul_ex_mult_76_U175 ( .A1(mul_ex_mult_76_n85), .A2(
        mul_ex_mult_76_n74), .ZN(mul_ex_mult_76_ab_4__9_) );
  NOR2_X1 mul_ex_mult_76_U174 ( .A1(mul_ex_mult_76_n94), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__0_) );
  NOR2_X1 mul_ex_mult_76_U173 ( .A1(mul_ex_mult_76_n84), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__10_) );
  NOR2_X1 mul_ex_mult_76_U172 ( .A1(mul_ex_mult_76_n83), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__11_) );
  NOR2_X1 mul_ex_mult_76_U171 ( .A1(mul_ex_mult_76_n82), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__12_) );
  NOR2_X1 mul_ex_mult_76_U170 ( .A1(mul_ex_mult_76_n81), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__13_) );
  NOR2_X1 mul_ex_mult_76_U169 ( .A1(mul_ex_mult_76_n80), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__14_) );
  NOR2_X1 mul_ex_mult_76_U168 ( .A1(mul_ex_mult_76_n79), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__15_) );
  NOR2_X1 mul_ex_mult_76_U167 ( .A1(mul_ex_mult_76_n93), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__1_) );
  NOR2_X1 mul_ex_mult_76_U166 ( .A1(mul_ex_mult_76_n92), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__2_) );
  NOR2_X1 mul_ex_mult_76_U165 ( .A1(mul_ex_mult_76_n91), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__3_) );
  NOR2_X1 mul_ex_mult_76_U164 ( .A1(mul_ex_mult_76_n90), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__4_) );
  NOR2_X1 mul_ex_mult_76_U163 ( .A1(mul_ex_mult_76_n89), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__5_) );
  NOR2_X1 mul_ex_mult_76_U162 ( .A1(mul_ex_mult_76_n88), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__6_) );
  NOR2_X1 mul_ex_mult_76_U161 ( .A1(mul_ex_mult_76_n87), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__7_) );
  NOR2_X1 mul_ex_mult_76_U160 ( .A1(mul_ex_mult_76_n86), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__8_) );
  NOR2_X1 mul_ex_mult_76_U159 ( .A1(mul_ex_mult_76_n85), .A2(
        mul_ex_mult_76_n73), .ZN(mul_ex_mult_76_ab_5__9_) );
  NOR2_X1 mul_ex_mult_76_U158 ( .A1(mul_ex_mult_76_n94), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__0_) );
  NOR2_X1 mul_ex_mult_76_U157 ( .A1(mul_ex_mult_76_n84), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__10_) );
  NOR2_X1 mul_ex_mult_76_U156 ( .A1(mul_ex_mult_76_n83), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__11_) );
  NOR2_X1 mul_ex_mult_76_U155 ( .A1(mul_ex_mult_76_n82), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__12_) );
  NOR2_X1 mul_ex_mult_76_U154 ( .A1(mul_ex_mult_76_n81), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__13_) );
  NOR2_X1 mul_ex_mult_76_U153 ( .A1(mul_ex_mult_76_n80), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__14_) );
  NOR2_X1 mul_ex_mult_76_U152 ( .A1(mul_ex_mult_76_n79), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__15_) );
  NOR2_X1 mul_ex_mult_76_U151 ( .A1(mul_ex_mult_76_n93), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__1_) );
  NOR2_X1 mul_ex_mult_76_U150 ( .A1(mul_ex_mult_76_n92), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__2_) );
  NOR2_X1 mul_ex_mult_76_U149 ( .A1(mul_ex_mult_76_n91), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__3_) );
  NOR2_X1 mul_ex_mult_76_U148 ( .A1(mul_ex_mult_76_n90), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__4_) );
  NOR2_X1 mul_ex_mult_76_U147 ( .A1(mul_ex_mult_76_n89), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__5_) );
  NOR2_X1 mul_ex_mult_76_U146 ( .A1(mul_ex_mult_76_n88), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__6_) );
  NOR2_X1 mul_ex_mult_76_U145 ( .A1(mul_ex_mult_76_n87), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__7_) );
  NOR2_X1 mul_ex_mult_76_U144 ( .A1(mul_ex_mult_76_n86), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__8_) );
  NOR2_X1 mul_ex_mult_76_U143 ( .A1(mul_ex_mult_76_n85), .A2(
        mul_ex_mult_76_n72), .ZN(mul_ex_mult_76_ab_6__9_) );
  NOR2_X1 mul_ex_mult_76_U142 ( .A1(mul_ex_mult_76_n94), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__0_) );
  NOR2_X1 mul_ex_mult_76_U141 ( .A1(mul_ex_mult_76_n84), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__10_) );
  NOR2_X1 mul_ex_mult_76_U140 ( .A1(mul_ex_mult_76_n83), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__11_) );
  NOR2_X1 mul_ex_mult_76_U139 ( .A1(mul_ex_mult_76_n82), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__12_) );
  NOR2_X1 mul_ex_mult_76_U138 ( .A1(mul_ex_mult_76_n81), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__13_) );
  NOR2_X1 mul_ex_mult_76_U137 ( .A1(mul_ex_mult_76_n80), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__14_) );
  NOR2_X1 mul_ex_mult_76_U136 ( .A1(mul_ex_mult_76_n79), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__15_) );
  NOR2_X1 mul_ex_mult_76_U135 ( .A1(mul_ex_mult_76_n93), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__1_) );
  NOR2_X1 mul_ex_mult_76_U134 ( .A1(mul_ex_mult_76_n92), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__2_) );
  NOR2_X1 mul_ex_mult_76_U133 ( .A1(mul_ex_mult_76_n91), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__3_) );
  NOR2_X1 mul_ex_mult_76_U132 ( .A1(mul_ex_mult_76_n90), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__4_) );
  NOR2_X1 mul_ex_mult_76_U131 ( .A1(mul_ex_mult_76_n89), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__5_) );
  NOR2_X1 mul_ex_mult_76_U130 ( .A1(mul_ex_mult_76_n88), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__6_) );
  NOR2_X1 mul_ex_mult_76_U129 ( .A1(mul_ex_mult_76_n87), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__7_) );
  NOR2_X1 mul_ex_mult_76_U128 ( .A1(mul_ex_mult_76_n86), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__8_) );
  NOR2_X1 mul_ex_mult_76_U127 ( .A1(mul_ex_mult_76_n85), .A2(
        mul_ex_mult_76_n71), .ZN(mul_ex_mult_76_ab_7__9_) );
  NOR2_X1 mul_ex_mult_76_U126 ( .A1(mul_ex_mult_76_n94), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__0_) );
  NOR2_X1 mul_ex_mult_76_U125 ( .A1(mul_ex_mult_76_n84), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__10_) );
  NOR2_X1 mul_ex_mult_76_U124 ( .A1(mul_ex_mult_76_n83), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__11_) );
  NOR2_X1 mul_ex_mult_76_U123 ( .A1(mul_ex_mult_76_n82), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__12_) );
  NOR2_X1 mul_ex_mult_76_U122 ( .A1(mul_ex_mult_76_n81), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__13_) );
  NOR2_X1 mul_ex_mult_76_U121 ( .A1(mul_ex_mult_76_n80), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__14_) );
  NOR2_X1 mul_ex_mult_76_U120 ( .A1(mul_ex_mult_76_n79), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__15_) );
  NOR2_X1 mul_ex_mult_76_U119 ( .A1(mul_ex_mult_76_n93), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__1_) );
  NOR2_X1 mul_ex_mult_76_U118 ( .A1(mul_ex_mult_76_n92), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__2_) );
  NOR2_X1 mul_ex_mult_76_U117 ( .A1(mul_ex_mult_76_n91), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__3_) );
  NOR2_X1 mul_ex_mult_76_U116 ( .A1(mul_ex_mult_76_n90), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__4_) );
  NOR2_X1 mul_ex_mult_76_U115 ( .A1(mul_ex_mult_76_n89), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__5_) );
  NOR2_X1 mul_ex_mult_76_U114 ( .A1(mul_ex_mult_76_n88), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__6_) );
  NOR2_X1 mul_ex_mult_76_U113 ( .A1(mul_ex_mult_76_n87), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__7_) );
  NOR2_X1 mul_ex_mult_76_U112 ( .A1(mul_ex_mult_76_n86), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__8_) );
  NOR2_X1 mul_ex_mult_76_U111 ( .A1(mul_ex_mult_76_n85), .A2(
        mul_ex_mult_76_n70), .ZN(mul_ex_mult_76_ab_8__9_) );
  NOR2_X1 mul_ex_mult_76_U110 ( .A1(mul_ex_mult_76_n69), .A2(
        mul_ex_mult_76_n94), .ZN(mul_ex_mult_76_ab_9__0_) );
  NOR2_X1 mul_ex_mult_76_U109 ( .A1(mul_ex_mult_76_n69), .A2(
        mul_ex_mult_76_n84), .ZN(mul_ex_mult_76_ab_9__10_) );
  NOR2_X1 mul_ex_mult_76_U108 ( .A1(mul_ex_mult_76_n69), .A2(
        mul_ex_mult_76_n83), .ZN(mul_ex_mult_76_ab_9__11_) );
  NOR2_X1 mul_ex_mult_76_U107 ( .A1(mul_ex_mult_76_n69), .A2(
        mul_ex_mult_76_n82), .ZN(mul_ex_mult_76_ab_9__12_) );
  NOR2_X1 mul_ex_mult_76_U106 ( .A1(mul_ex_mult_76_n69), .A2(
        mul_ex_mult_76_n81), .ZN(mul_ex_mult_76_ab_9__13_) );
  NOR2_X1 mul_ex_mult_76_U105 ( .A1(mul_ex_mult_76_n69), .A2(
        mul_ex_mult_76_n80), .ZN(mul_ex_mult_76_ab_9__14_) );
  NOR2_X1 mul_ex_mult_76_U104 ( .A1(mul_ex_mult_76_n69), .A2(
        mul_ex_mult_76_n79), .ZN(mul_ex_mult_76_ab_9__15_) );
  NOR2_X1 mul_ex_mult_76_U103 ( .A1(mul_ex_mult_76_n69), .A2(
        mul_ex_mult_76_n93), .ZN(mul_ex_mult_76_ab_9__1_) );
  NOR2_X1 mul_ex_mult_76_U102 ( .A1(mul_ex_mult_76_n69), .A2(
        mul_ex_mult_76_n92), .ZN(mul_ex_mult_76_ab_9__2_) );
  NOR2_X1 mul_ex_mult_76_U101 ( .A1(mul_ex_mult_76_n69), .A2(
        mul_ex_mult_76_n91), .ZN(mul_ex_mult_76_ab_9__3_) );
  NOR2_X1 mul_ex_mult_76_U100 ( .A1(mul_ex_mult_76_n69), .A2(
        mul_ex_mult_76_n90), .ZN(mul_ex_mult_76_ab_9__4_) );
  NOR2_X1 mul_ex_mult_76_U99 ( .A1(mul_ex_mult_76_n69), .A2(mul_ex_mult_76_n89), .ZN(mul_ex_mult_76_ab_9__5_) );
  NOR2_X1 mul_ex_mult_76_U98 ( .A1(mul_ex_mult_76_n69), .A2(mul_ex_mult_76_n88), .ZN(mul_ex_mult_76_ab_9__6_) );
  NOR2_X1 mul_ex_mult_76_U97 ( .A1(mul_ex_mult_76_n69), .A2(mul_ex_mult_76_n87), .ZN(mul_ex_mult_76_ab_9__7_) );
  NOR2_X1 mul_ex_mult_76_U96 ( .A1(mul_ex_mult_76_n69), .A2(mul_ex_mult_76_n86), .ZN(mul_ex_mult_76_ab_9__8_) );
  NOR2_X1 mul_ex_mult_76_U95 ( .A1(mul_ex_mult_76_n69), .A2(mul_ex_mult_76_n85), .ZN(mul_ex_mult_76_ab_9__9_) );
  INV_X4 mul_ex_mult_76_U93 ( .A(f1_in[13]), .ZN(mul_ex_mult_76_n76) );
  INV_X4 mul_ex_mult_76_U92 ( .A(f1_in[0]), .ZN(mul_ex_mult_76_n63) );
  INV_X4 mul_ex_mult_76_U91 ( .A(f1_in[1]), .ZN(mul_ex_mult_76_n64) );
  INV_X4 mul_ex_mult_76_U90 ( .A(f1_in[2]), .ZN(mul_ex_mult_76_n65) );
  INV_X4 mul_ex_mult_76_U89 ( .A(f1_in[3]), .ZN(mul_ex_mult_76_n66) );
  INV_X4 mul_ex_mult_76_U88 ( .A(f1_in[4]), .ZN(mul_ex_mult_76_n67) );
  INV_X4 mul_ex_mult_76_U87 ( .A(f1_in[5]), .ZN(mul_ex_mult_76_n68) );
  INV_X4 mul_ex_mult_76_U86 ( .A(f1_in[7]), .ZN(mul_ex_mult_76_n70) );
  INV_X4 mul_ex_mult_76_U85 ( .A(f1_in[8]), .ZN(mul_ex_mult_76_n71) );
  INV_X4 mul_ex_mult_76_U84 ( .A(f1_in[9]), .ZN(mul_ex_mult_76_n72) );
  INV_X4 mul_ex_mult_76_U83 ( .A(f1_in[10]), .ZN(mul_ex_mult_76_n73) );
  INV_X4 mul_ex_mult_76_U82 ( .A(f1_in[11]), .ZN(mul_ex_mult_76_n74) );
  INV_X4 mul_ex_mult_76_U81 ( .A(f1_in[12]), .ZN(mul_ex_mult_76_n75) );
  INV_X4 mul_ex_mult_76_U80 ( .A(f1_in[14]), .ZN(mul_ex_mult_76_n77) );
  INV_X4 mul_ex_mult_76_U79 ( .A(f1_in[15]), .ZN(mul_ex_mult_76_n78) );
  INV_X4 mul_ex_mult_76_U78 ( .A(f2_in[15]), .ZN(mul_ex_mult_76_n94) );
  INV_X4 mul_ex_mult_76_U77 ( .A(f2_in[0]), .ZN(mul_ex_mult_76_n79) );
  INV_X4 mul_ex_mult_76_U76 ( .A(f2_in[2]), .ZN(mul_ex_mult_76_n81) );
  INV_X4 mul_ex_mult_76_U75 ( .A(f2_in[1]), .ZN(mul_ex_mult_76_n80) );
  INV_X4 mul_ex_mult_76_U74 ( .A(f2_in[4]), .ZN(mul_ex_mult_76_n83) );
  INV_X4 mul_ex_mult_76_U73 ( .A(f2_in[3]), .ZN(mul_ex_mult_76_n82) );
  INV_X4 mul_ex_mult_76_U72 ( .A(f2_in[6]), .ZN(mul_ex_mult_76_n85) );
  INV_X4 mul_ex_mult_76_U71 ( .A(f2_in[5]), .ZN(mul_ex_mult_76_n84) );
  INV_X4 mul_ex_mult_76_U70 ( .A(f2_in[9]), .ZN(mul_ex_mult_76_n88) );
  INV_X4 mul_ex_mult_76_U69 ( .A(f2_in[10]), .ZN(mul_ex_mult_76_n89) );
  INV_X4 mul_ex_mult_76_U68 ( .A(f2_in[11]), .ZN(mul_ex_mult_76_n90) );
  INV_X4 mul_ex_mult_76_U67 ( .A(f2_in[12]), .ZN(mul_ex_mult_76_n91) );
  INV_X4 mul_ex_mult_76_U66 ( .A(f2_in[13]), .ZN(mul_ex_mult_76_n92) );
  INV_X4 mul_ex_mult_76_U65 ( .A(f2_in[14]), .ZN(mul_ex_mult_76_n93) );
  INV_X4 mul_ex_mult_76_U64 ( .A(f2_in[8]), .ZN(mul_ex_mult_76_n87) );
  INV_X4 mul_ex_mult_76_U63 ( .A(f2_in[7]), .ZN(mul_ex_mult_76_n86) );
  INV_X4 mul_ex_mult_76_U62 ( .A(f1_in[6]), .ZN(mul_ex_mult_76_n69) );
  AND2_X4 mul_ex_mult_76_U61 ( .A1(mul_ex_mult_76_CARRYB_15__14_), .A2(
        mul_ex_mult_76_ab_15__15_), .ZN(mul_ex_mult_76_n62) );
  XOR2_X2 mul_ex_mult_76_U60 ( .A(mul_ex_mult_76_CARRYB_15__0_), .B(
        mul_ex_mult_76_SUMB_15__1_), .Z(mul_ex_mult_76_n61) );
  AND2_X4 mul_ex_mult_76_U59 ( .A1(mul_ex_mult_76_CARRYB_15__0_), .A2(
        mul_ex_mult_76_SUMB_15__1_), .ZN(mul_ex_mult_76_n60) );
  AND2_X4 mul_ex_mult_76_U58 ( .A1(mul_ex_mult_76_CARRYB_15__2_), .A2(
        mul_ex_mult_76_SUMB_15__3_), .ZN(mul_ex_mult_76_n59) );
  AND2_X4 mul_ex_mult_76_U57 ( .A1(mul_ex_mult_76_CARRYB_15__4_), .A2(
        mul_ex_mult_76_SUMB_15__5_), .ZN(mul_ex_mult_76_n58) );
  AND2_X4 mul_ex_mult_76_U56 ( .A1(mul_ex_mult_76_CARRYB_15__6_), .A2(
        mul_ex_mult_76_SUMB_15__7_), .ZN(mul_ex_mult_76_n57) );
  AND2_X4 mul_ex_mult_76_U55 ( .A1(mul_ex_mult_76_CARRYB_15__8_), .A2(
        mul_ex_mult_76_SUMB_15__9_), .ZN(mul_ex_mult_76_n56) );
  AND2_X4 mul_ex_mult_76_U54 ( .A1(mul_ex_mult_76_CARRYB_15__10_), .A2(
        mul_ex_mult_76_SUMB_15__11_), .ZN(mul_ex_mult_76_n55) );
  AND2_X4 mul_ex_mult_76_U53 ( .A1(mul_ex_mult_76_CARRYB_15__12_), .A2(
        mul_ex_mult_76_SUMB_15__13_), .ZN(mul_ex_mult_76_n54) );
  AND2_X4 mul_ex_mult_76_U52 ( .A1(mul_ex_mult_76_CARRYB_15__1_), .A2(
        mul_ex_mult_76_SUMB_15__2_), .ZN(mul_ex_mult_76_n53) );
  AND2_X4 mul_ex_mult_76_U51 ( .A1(mul_ex_mult_76_CARRYB_15__3_), .A2(
        mul_ex_mult_76_SUMB_15__4_), .ZN(mul_ex_mult_76_n52) );
  AND2_X4 mul_ex_mult_76_U50 ( .A1(mul_ex_mult_76_CARRYB_15__5_), .A2(
        mul_ex_mult_76_SUMB_15__6_), .ZN(mul_ex_mult_76_n51) );
  AND2_X4 mul_ex_mult_76_U49 ( .A1(mul_ex_mult_76_CARRYB_15__7_), .A2(
        mul_ex_mult_76_SUMB_15__8_), .ZN(mul_ex_mult_76_n50) );
  AND2_X4 mul_ex_mult_76_U48 ( .A1(mul_ex_mult_76_CARRYB_15__9_), .A2(
        mul_ex_mult_76_SUMB_15__10_), .ZN(mul_ex_mult_76_n49) );
  AND2_X4 mul_ex_mult_76_U47 ( .A1(mul_ex_mult_76_CARRYB_15__11_), .A2(
        mul_ex_mult_76_SUMB_15__12_), .ZN(mul_ex_mult_76_n48) );
  AND2_X4 mul_ex_mult_76_U46 ( .A1(mul_ex_mult_76_CARRYB_15__13_), .A2(
        mul_ex_mult_76_SUMB_15__14_), .ZN(mul_ex_mult_76_n47) );
  XOR2_X2 mul_ex_mult_76_U45 ( .A(mul_ex_mult_76_ab_1__0_), .B(
        mul_ex_mult_76_ab_0__1_), .Z(mul_ex_N57) );
  XOR2_X2 mul_ex_mult_76_U44 ( .A(mul_ex_mult_76_ab_1__1_), .B(
        mul_ex_mult_76_ab_0__2_), .Z(mul_ex_mult_76_n45) );
  XOR2_X2 mul_ex_mult_76_U43 ( .A(mul_ex_mult_76_ab_1__2_), .B(
        mul_ex_mult_76_ab_0__3_), .Z(mul_ex_mult_76_n44) );
  XOR2_X2 mul_ex_mult_76_U42 ( .A(mul_ex_mult_76_ab_1__3_), .B(
        mul_ex_mult_76_ab_0__4_), .Z(mul_ex_mult_76_n43) );
  XOR2_X2 mul_ex_mult_76_U41 ( .A(mul_ex_mult_76_ab_1__4_), .B(
        mul_ex_mult_76_ab_0__5_), .Z(mul_ex_mult_76_n42) );
  XOR2_X2 mul_ex_mult_76_U40 ( .A(mul_ex_mult_76_ab_1__5_), .B(
        mul_ex_mult_76_ab_0__6_), .Z(mul_ex_mult_76_n41) );
  XOR2_X2 mul_ex_mult_76_U39 ( .A(mul_ex_mult_76_ab_1__6_), .B(
        mul_ex_mult_76_ab_0__7_), .Z(mul_ex_mult_76_n40) );
  XOR2_X2 mul_ex_mult_76_U38 ( .A(mul_ex_mult_76_ab_1__7_), .B(
        mul_ex_mult_76_ab_0__8_), .Z(mul_ex_mult_76_n39) );
  XOR2_X2 mul_ex_mult_76_U37 ( .A(mul_ex_mult_76_ab_1__8_), .B(
        mul_ex_mult_76_ab_0__9_), .Z(mul_ex_mult_76_n38) );
  XOR2_X2 mul_ex_mult_76_U36 ( .A(mul_ex_mult_76_ab_1__9_), .B(
        mul_ex_mult_76_ab_0__10_), .Z(mul_ex_mult_76_n37) );
  XOR2_X2 mul_ex_mult_76_U35 ( .A(mul_ex_mult_76_ab_1__10_), .B(
        mul_ex_mult_76_ab_0__11_), .Z(mul_ex_mult_76_n36) );
  XOR2_X2 mul_ex_mult_76_U34 ( .A(mul_ex_mult_76_ab_1__11_), .B(
        mul_ex_mult_76_ab_0__12_), .Z(mul_ex_mult_76_n35) );
  XOR2_X2 mul_ex_mult_76_U33 ( .A(mul_ex_mult_76_ab_1__12_), .B(
        mul_ex_mult_76_ab_0__13_), .Z(mul_ex_mult_76_n34) );
  XOR2_X2 mul_ex_mult_76_U32 ( .A(mul_ex_mult_76_ab_1__13_), .B(
        mul_ex_mult_76_ab_0__14_), .Z(mul_ex_mult_76_n33) );
  XOR2_X2 mul_ex_mult_76_U31 ( .A(mul_ex_mult_76_ab_1__14_), .B(
        mul_ex_mult_76_ab_0__15_), .Z(mul_ex_mult_76_n32) );
  AND2_X4 mul_ex_mult_76_U30 ( .A1(mul_ex_mult_76_ab_0__15_), .A2(
        mul_ex_mult_76_ab_1__14_), .ZN(mul_ex_mult_76_n31) );
  XOR2_X2 mul_ex_mult_76_U29 ( .A(mul_ex_mult_76_CARRYB_15__3_), .B(
        mul_ex_mult_76_SUMB_15__4_), .Z(mul_ex_mult_76_n30) );
  XOR2_X2 mul_ex_mult_76_U28 ( .A(mul_ex_mult_76_CARRYB_15__5_), .B(
        mul_ex_mult_76_SUMB_15__6_), .Z(mul_ex_mult_76_n29) );
  XOR2_X2 mul_ex_mult_76_U27 ( .A(mul_ex_mult_76_CARRYB_15__7_), .B(
        mul_ex_mult_76_SUMB_15__8_), .Z(mul_ex_mult_76_n28) );
  XOR2_X2 mul_ex_mult_76_U26 ( .A(mul_ex_mult_76_CARRYB_15__9_), .B(
        mul_ex_mult_76_SUMB_15__10_), .Z(mul_ex_mult_76_n27) );
  XOR2_X2 mul_ex_mult_76_U25 ( .A(mul_ex_mult_76_CARRYB_15__11_), .B(
        mul_ex_mult_76_SUMB_15__12_), .Z(mul_ex_mult_76_n26) );
  XOR2_X2 mul_ex_mult_76_U24 ( .A(mul_ex_mult_76_CARRYB_15__13_), .B(
        mul_ex_mult_76_SUMB_15__14_), .Z(mul_ex_mult_76_n25) );
  XOR2_X2 mul_ex_mult_76_U23 ( .A(mul_ex_mult_76_CARRYB_15__1_), .B(
        mul_ex_mult_76_SUMB_15__2_), .Z(mul_ex_mult_76_n24) );
  XOR2_X2 mul_ex_mult_76_U22 ( .A(mul_ex_mult_76_CARRYB_15__2_), .B(
        mul_ex_mult_76_SUMB_15__3_), .Z(mul_ex_mult_76_n23) );
  XOR2_X2 mul_ex_mult_76_U21 ( .A(mul_ex_mult_76_CARRYB_15__4_), .B(
        mul_ex_mult_76_SUMB_15__5_), .Z(mul_ex_mult_76_n22) );
  XOR2_X2 mul_ex_mult_76_U20 ( .A(mul_ex_mult_76_CARRYB_15__6_), .B(
        mul_ex_mult_76_SUMB_15__7_), .Z(mul_ex_mult_76_n21) );
  XOR2_X2 mul_ex_mult_76_U19 ( .A(mul_ex_mult_76_CARRYB_15__8_), .B(
        mul_ex_mult_76_SUMB_15__9_), .Z(mul_ex_mult_76_n20) );
  XOR2_X2 mul_ex_mult_76_U18 ( .A(mul_ex_mult_76_CARRYB_15__10_), .B(
        mul_ex_mult_76_SUMB_15__11_), .Z(mul_ex_mult_76_n19) );
  XOR2_X2 mul_ex_mult_76_U17 ( .A(mul_ex_mult_76_CARRYB_15__12_), .B(
        mul_ex_mult_76_SUMB_15__13_), .Z(mul_ex_mult_76_n18) );
  XOR2_X2 mul_ex_mult_76_U16 ( .A(mul_ex_mult_76_CARRYB_15__14_), .B(
        mul_ex_mult_76_ab_15__15_), .Z(mul_ex_mult_76_n17) );
  AND2_X4 mul_ex_mult_76_U15 ( .A1(mul_ex_mult_76_ab_0__1_), .A2(
        mul_ex_mult_76_ab_1__0_), .ZN(mul_ex_mult_76_n16) );
  AND2_X4 mul_ex_mult_76_U14 ( .A1(mul_ex_mult_76_ab_0__2_), .A2(
        mul_ex_mult_76_ab_1__1_), .ZN(mul_ex_mult_76_n15) );
  AND2_X4 mul_ex_mult_76_U13 ( .A1(mul_ex_mult_76_ab_0__3_), .A2(
        mul_ex_mult_76_ab_1__2_), .ZN(mul_ex_mult_76_n14) );
  AND2_X4 mul_ex_mult_76_U12 ( .A1(mul_ex_mult_76_ab_0__4_), .A2(
        mul_ex_mult_76_ab_1__3_), .ZN(mul_ex_mult_76_n13) );
  AND2_X4 mul_ex_mult_76_U11 ( .A1(mul_ex_mult_76_ab_0__5_), .A2(
        mul_ex_mult_76_ab_1__4_), .ZN(mul_ex_mult_76_n12) );
  AND2_X4 mul_ex_mult_76_U10 ( .A1(mul_ex_mult_76_ab_0__6_), .A2(
        mul_ex_mult_76_ab_1__5_), .ZN(mul_ex_mult_76_n11) );
  AND2_X4 mul_ex_mult_76_U9 ( .A1(mul_ex_mult_76_ab_0__7_), .A2(
        mul_ex_mult_76_ab_1__6_), .ZN(mul_ex_mult_76_n10) );
  AND2_X4 mul_ex_mult_76_U8 ( .A1(mul_ex_mult_76_ab_0__8_), .A2(
        mul_ex_mult_76_ab_1__7_), .ZN(mul_ex_mult_76_n9) );
  AND2_X4 mul_ex_mult_76_U7 ( .A1(mul_ex_mult_76_ab_0__9_), .A2(
        mul_ex_mult_76_ab_1__8_), .ZN(mul_ex_mult_76_n8) );
  AND2_X4 mul_ex_mult_76_U6 ( .A1(mul_ex_mult_76_ab_0__10_), .A2(
        mul_ex_mult_76_ab_1__9_), .ZN(mul_ex_mult_76_n7) );
  AND2_X4 mul_ex_mult_76_U5 ( .A1(mul_ex_mult_76_ab_0__11_), .A2(
        mul_ex_mult_76_ab_1__10_), .ZN(mul_ex_mult_76_n6) );
  AND2_X4 mul_ex_mult_76_U4 ( .A1(mul_ex_mult_76_ab_0__12_), .A2(
        mul_ex_mult_76_ab_1__11_), .ZN(mul_ex_mult_76_n5) );
  AND2_X4 mul_ex_mult_76_U3 ( .A1(mul_ex_mult_76_ab_0__13_), .A2(
        mul_ex_mult_76_ab_1__12_), .ZN(mul_ex_mult_76_n4) );
  AND2_X4 mul_ex_mult_76_U2 ( .A1(mul_ex_mult_76_ab_0__14_), .A2(
        mul_ex_mult_76_ab_1__13_), .ZN(mul_ex_mult_76_n3) );
  FA_X1 mul_ex_mult_76_S3_2_14 ( .A(mul_ex_mult_76_ab_2__14_), .B(
        mul_ex_mult_76_n31), .CI(mul_ex_mult_76_ab_1__15_), .CO(
        mul_ex_mult_76_CARRYB_2__14_), .S(mul_ex_mult_76_SUMB_2__14_) );
  FA_X1 mul_ex_mult_76_S2_2_13 ( .A(mul_ex_mult_76_ab_2__13_), .B(
        mul_ex_mult_76_n3), .CI(mul_ex_mult_76_n32), .CO(
        mul_ex_mult_76_CARRYB_2__13_), .S(mul_ex_mult_76_SUMB_2__13_) );
  FA_X1 mul_ex_mult_76_S2_2_12 ( .A(mul_ex_mult_76_ab_2__12_), .B(
        mul_ex_mult_76_n4), .CI(mul_ex_mult_76_n33), .CO(
        mul_ex_mult_76_CARRYB_2__12_), .S(mul_ex_mult_76_SUMB_2__12_) );
  FA_X1 mul_ex_mult_76_S2_2_11 ( .A(mul_ex_mult_76_ab_2__11_), .B(
        mul_ex_mult_76_n5), .CI(mul_ex_mult_76_n34), .CO(
        mul_ex_mult_76_CARRYB_2__11_), .S(mul_ex_mult_76_SUMB_2__11_) );
  FA_X1 mul_ex_mult_76_S2_2_10 ( .A(mul_ex_mult_76_ab_2__10_), .B(
        mul_ex_mult_76_n6), .CI(mul_ex_mult_76_n35), .CO(
        mul_ex_mult_76_CARRYB_2__10_), .S(mul_ex_mult_76_SUMB_2__10_) );
  FA_X1 mul_ex_mult_76_S2_2_9 ( .A(mul_ex_mult_76_ab_2__9_), .B(
        mul_ex_mult_76_n7), .CI(mul_ex_mult_76_n36), .CO(
        mul_ex_mult_76_CARRYB_2__9_), .S(mul_ex_mult_76_SUMB_2__9_) );
  FA_X1 mul_ex_mult_76_S2_2_8 ( .A(mul_ex_mult_76_ab_2__8_), .B(
        mul_ex_mult_76_n8), .CI(mul_ex_mult_76_n37), .CO(
        mul_ex_mult_76_CARRYB_2__8_), .S(mul_ex_mult_76_SUMB_2__8_) );
  FA_X1 mul_ex_mult_76_S2_2_7 ( .A(mul_ex_mult_76_ab_2__7_), .B(
        mul_ex_mult_76_n9), .CI(mul_ex_mult_76_n38), .CO(
        mul_ex_mult_76_CARRYB_2__7_), .S(mul_ex_mult_76_SUMB_2__7_) );
  FA_X1 mul_ex_mult_76_S2_2_6 ( .A(mul_ex_mult_76_ab_2__6_), .B(
        mul_ex_mult_76_n10), .CI(mul_ex_mult_76_n39), .CO(
        mul_ex_mult_76_CARRYB_2__6_), .S(mul_ex_mult_76_SUMB_2__6_) );
  FA_X1 mul_ex_mult_76_S2_2_5 ( .A(mul_ex_mult_76_ab_2__5_), .B(
        mul_ex_mult_76_n11), .CI(mul_ex_mult_76_n40), .CO(
        mul_ex_mult_76_CARRYB_2__5_), .S(mul_ex_mult_76_SUMB_2__5_) );
  FA_X1 mul_ex_mult_76_S2_2_4 ( .A(mul_ex_mult_76_ab_2__4_), .B(
        mul_ex_mult_76_n12), .CI(mul_ex_mult_76_n41), .CO(
        mul_ex_mult_76_CARRYB_2__4_), .S(mul_ex_mult_76_SUMB_2__4_) );
  FA_X1 mul_ex_mult_76_S2_2_3 ( .A(mul_ex_mult_76_ab_2__3_), .B(
        mul_ex_mult_76_n13), .CI(mul_ex_mult_76_n42), .CO(
        mul_ex_mult_76_CARRYB_2__3_), .S(mul_ex_mult_76_SUMB_2__3_) );
  FA_X1 mul_ex_mult_76_S2_2_2 ( .A(mul_ex_mult_76_ab_2__2_), .B(
        mul_ex_mult_76_n14), .CI(mul_ex_mult_76_n43), .CO(
        mul_ex_mult_76_CARRYB_2__2_), .S(mul_ex_mult_76_SUMB_2__2_) );
  FA_X1 mul_ex_mult_76_S2_2_1 ( .A(mul_ex_mult_76_ab_2__1_), .B(
        mul_ex_mult_76_n15), .CI(mul_ex_mult_76_n44), .CO(
        mul_ex_mult_76_CARRYB_2__1_), .S(mul_ex_mult_76_SUMB_2__1_) );
  FA_X1 mul_ex_mult_76_S1_2_0 ( .A(mul_ex_mult_76_ab_2__0_), .B(
        mul_ex_mult_76_n16), .CI(mul_ex_mult_76_n45), .CO(
        mul_ex_mult_76_CARRYB_2__0_), .S(mul_ex_mult_76_A1_0_) );
  FA_X1 mul_ex_mult_76_S3_3_14 ( .A(mul_ex_mult_76_ab_3__14_), .B(
        mul_ex_mult_76_CARRYB_2__14_), .CI(mul_ex_mult_76_ab_2__15_), .CO(
        mul_ex_mult_76_CARRYB_3__14_), .S(mul_ex_mult_76_SUMB_3__14_) );
  FA_X1 mul_ex_mult_76_S2_3_13 ( .A(mul_ex_mult_76_ab_3__13_), .B(
        mul_ex_mult_76_CARRYB_2__13_), .CI(mul_ex_mult_76_SUMB_2__14_), .CO(
        mul_ex_mult_76_CARRYB_3__13_), .S(mul_ex_mult_76_SUMB_3__13_) );
  FA_X1 mul_ex_mult_76_S2_3_12 ( .A(mul_ex_mult_76_ab_3__12_), .B(
        mul_ex_mult_76_CARRYB_2__12_), .CI(mul_ex_mult_76_SUMB_2__13_), .CO(
        mul_ex_mult_76_CARRYB_3__12_), .S(mul_ex_mult_76_SUMB_3__12_) );
  FA_X1 mul_ex_mult_76_S2_3_11 ( .A(mul_ex_mult_76_ab_3__11_), .B(
        mul_ex_mult_76_CARRYB_2__11_), .CI(mul_ex_mult_76_SUMB_2__12_), .CO(
        mul_ex_mult_76_CARRYB_3__11_), .S(mul_ex_mult_76_SUMB_3__11_) );
  FA_X1 mul_ex_mult_76_S2_3_10 ( .A(mul_ex_mult_76_ab_3__10_), .B(
        mul_ex_mult_76_CARRYB_2__10_), .CI(mul_ex_mult_76_SUMB_2__11_), .CO(
        mul_ex_mult_76_CARRYB_3__10_), .S(mul_ex_mult_76_SUMB_3__10_) );
  FA_X1 mul_ex_mult_76_S2_3_9 ( .A(mul_ex_mult_76_ab_3__9_), .B(
        mul_ex_mult_76_CARRYB_2__9_), .CI(mul_ex_mult_76_SUMB_2__10_), .CO(
        mul_ex_mult_76_CARRYB_3__9_), .S(mul_ex_mult_76_SUMB_3__9_) );
  FA_X1 mul_ex_mult_76_S2_3_8 ( .A(mul_ex_mult_76_ab_3__8_), .B(
        mul_ex_mult_76_CARRYB_2__8_), .CI(mul_ex_mult_76_SUMB_2__9_), .CO(
        mul_ex_mult_76_CARRYB_3__8_), .S(mul_ex_mult_76_SUMB_3__8_) );
  FA_X1 mul_ex_mult_76_S2_3_7 ( .A(mul_ex_mult_76_ab_3__7_), .B(
        mul_ex_mult_76_CARRYB_2__7_), .CI(mul_ex_mult_76_SUMB_2__8_), .CO(
        mul_ex_mult_76_CARRYB_3__7_), .S(mul_ex_mult_76_SUMB_3__7_) );
  FA_X1 mul_ex_mult_76_S2_3_6 ( .A(mul_ex_mult_76_ab_3__6_), .B(
        mul_ex_mult_76_CARRYB_2__6_), .CI(mul_ex_mult_76_SUMB_2__7_), .CO(
        mul_ex_mult_76_CARRYB_3__6_), .S(mul_ex_mult_76_SUMB_3__6_) );
  FA_X1 mul_ex_mult_76_S2_3_5 ( .A(mul_ex_mult_76_ab_3__5_), .B(
        mul_ex_mult_76_CARRYB_2__5_), .CI(mul_ex_mult_76_SUMB_2__6_), .CO(
        mul_ex_mult_76_CARRYB_3__5_), .S(mul_ex_mult_76_SUMB_3__5_) );
  FA_X1 mul_ex_mult_76_S2_3_4 ( .A(mul_ex_mult_76_ab_3__4_), .B(
        mul_ex_mult_76_CARRYB_2__4_), .CI(mul_ex_mult_76_SUMB_2__5_), .CO(
        mul_ex_mult_76_CARRYB_3__4_), .S(mul_ex_mult_76_SUMB_3__4_) );
  FA_X1 mul_ex_mult_76_S2_3_3 ( .A(mul_ex_mult_76_ab_3__3_), .B(
        mul_ex_mult_76_CARRYB_2__3_), .CI(mul_ex_mult_76_SUMB_2__4_), .CO(
        mul_ex_mult_76_CARRYB_3__3_), .S(mul_ex_mult_76_SUMB_3__3_) );
  FA_X1 mul_ex_mult_76_S2_3_2 ( .A(mul_ex_mult_76_ab_3__2_), .B(
        mul_ex_mult_76_CARRYB_2__2_), .CI(mul_ex_mult_76_SUMB_2__3_), .CO(
        mul_ex_mult_76_CARRYB_3__2_), .S(mul_ex_mult_76_SUMB_3__2_) );
  FA_X1 mul_ex_mult_76_S2_3_1 ( .A(mul_ex_mult_76_ab_3__1_), .B(
        mul_ex_mult_76_CARRYB_2__1_), .CI(mul_ex_mult_76_SUMB_2__2_), .CO(
        mul_ex_mult_76_CARRYB_3__1_), .S(mul_ex_mult_76_SUMB_3__1_) );
  FA_X1 mul_ex_mult_76_S1_3_0 ( .A(mul_ex_mult_76_ab_3__0_), .B(
        mul_ex_mult_76_CARRYB_2__0_), .CI(mul_ex_mult_76_SUMB_2__1_), .CO(
        mul_ex_mult_76_CARRYB_3__0_), .S(mul_ex_mult_76_A1_1_) );
  FA_X1 mul_ex_mult_76_S3_4_14 ( .A(mul_ex_mult_76_ab_4__14_), .B(
        mul_ex_mult_76_CARRYB_3__14_), .CI(mul_ex_mult_76_ab_3__15_), .CO(
        mul_ex_mult_76_CARRYB_4__14_), .S(mul_ex_mult_76_SUMB_4__14_) );
  FA_X1 mul_ex_mult_76_S2_4_13 ( .A(mul_ex_mult_76_ab_4__13_), .B(
        mul_ex_mult_76_CARRYB_3__13_), .CI(mul_ex_mult_76_SUMB_3__14_), .CO(
        mul_ex_mult_76_CARRYB_4__13_), .S(mul_ex_mult_76_SUMB_4__13_) );
  FA_X1 mul_ex_mult_76_S2_4_12 ( .A(mul_ex_mult_76_ab_4__12_), .B(
        mul_ex_mult_76_CARRYB_3__12_), .CI(mul_ex_mult_76_SUMB_3__13_), .CO(
        mul_ex_mult_76_CARRYB_4__12_), .S(mul_ex_mult_76_SUMB_4__12_) );
  FA_X1 mul_ex_mult_76_S2_4_11 ( .A(mul_ex_mult_76_ab_4__11_), .B(
        mul_ex_mult_76_CARRYB_3__11_), .CI(mul_ex_mult_76_SUMB_3__12_), .CO(
        mul_ex_mult_76_CARRYB_4__11_), .S(mul_ex_mult_76_SUMB_4__11_) );
  FA_X1 mul_ex_mult_76_S2_4_10 ( .A(mul_ex_mult_76_ab_4__10_), .B(
        mul_ex_mult_76_CARRYB_3__10_), .CI(mul_ex_mult_76_SUMB_3__11_), .CO(
        mul_ex_mult_76_CARRYB_4__10_), .S(mul_ex_mult_76_SUMB_4__10_) );
  FA_X1 mul_ex_mult_76_S2_4_9 ( .A(mul_ex_mult_76_ab_4__9_), .B(
        mul_ex_mult_76_CARRYB_3__9_), .CI(mul_ex_mult_76_SUMB_3__10_), .CO(
        mul_ex_mult_76_CARRYB_4__9_), .S(mul_ex_mult_76_SUMB_4__9_) );
  FA_X1 mul_ex_mult_76_S2_4_8 ( .A(mul_ex_mult_76_ab_4__8_), .B(
        mul_ex_mult_76_CARRYB_3__8_), .CI(mul_ex_mult_76_SUMB_3__9_), .CO(
        mul_ex_mult_76_CARRYB_4__8_), .S(mul_ex_mult_76_SUMB_4__8_) );
  FA_X1 mul_ex_mult_76_S2_4_7 ( .A(mul_ex_mult_76_ab_4__7_), .B(
        mul_ex_mult_76_CARRYB_3__7_), .CI(mul_ex_mult_76_SUMB_3__8_), .CO(
        mul_ex_mult_76_CARRYB_4__7_), .S(mul_ex_mult_76_SUMB_4__7_) );
  FA_X1 mul_ex_mult_76_S2_4_6 ( .A(mul_ex_mult_76_ab_4__6_), .B(
        mul_ex_mult_76_CARRYB_3__6_), .CI(mul_ex_mult_76_SUMB_3__7_), .CO(
        mul_ex_mult_76_CARRYB_4__6_), .S(mul_ex_mult_76_SUMB_4__6_) );
  FA_X1 mul_ex_mult_76_S2_4_5 ( .A(mul_ex_mult_76_ab_4__5_), .B(
        mul_ex_mult_76_CARRYB_3__5_), .CI(mul_ex_mult_76_SUMB_3__6_), .CO(
        mul_ex_mult_76_CARRYB_4__5_), .S(mul_ex_mult_76_SUMB_4__5_) );
  FA_X1 mul_ex_mult_76_S2_4_4 ( .A(mul_ex_mult_76_ab_4__4_), .B(
        mul_ex_mult_76_CARRYB_3__4_), .CI(mul_ex_mult_76_SUMB_3__5_), .CO(
        mul_ex_mult_76_CARRYB_4__4_), .S(mul_ex_mult_76_SUMB_4__4_) );
  FA_X1 mul_ex_mult_76_S2_4_3 ( .A(mul_ex_mult_76_ab_4__3_), .B(
        mul_ex_mult_76_CARRYB_3__3_), .CI(mul_ex_mult_76_SUMB_3__4_), .CO(
        mul_ex_mult_76_CARRYB_4__3_), .S(mul_ex_mult_76_SUMB_4__3_) );
  FA_X1 mul_ex_mult_76_S2_4_2 ( .A(mul_ex_mult_76_ab_4__2_), .B(
        mul_ex_mult_76_CARRYB_3__2_), .CI(mul_ex_mult_76_SUMB_3__3_), .CO(
        mul_ex_mult_76_CARRYB_4__2_), .S(mul_ex_mult_76_SUMB_4__2_) );
  FA_X1 mul_ex_mult_76_S2_4_1 ( .A(mul_ex_mult_76_ab_4__1_), .B(
        mul_ex_mult_76_CARRYB_3__1_), .CI(mul_ex_mult_76_SUMB_3__2_), .CO(
        mul_ex_mult_76_CARRYB_4__1_), .S(mul_ex_mult_76_SUMB_4__1_) );
  FA_X1 mul_ex_mult_76_S1_4_0 ( .A(mul_ex_mult_76_ab_4__0_), .B(
        mul_ex_mult_76_CARRYB_3__0_), .CI(mul_ex_mult_76_SUMB_3__1_), .CO(
        mul_ex_mult_76_CARRYB_4__0_), .S(mul_ex_mult_76_A1_2_) );
  FA_X1 mul_ex_mult_76_S3_5_14 ( .A(mul_ex_mult_76_ab_5__14_), .B(
        mul_ex_mult_76_CARRYB_4__14_), .CI(mul_ex_mult_76_ab_4__15_), .CO(
        mul_ex_mult_76_CARRYB_5__14_), .S(mul_ex_mult_76_SUMB_5__14_) );
  FA_X1 mul_ex_mult_76_S2_5_13 ( .A(mul_ex_mult_76_ab_5__13_), .B(
        mul_ex_mult_76_CARRYB_4__13_), .CI(mul_ex_mult_76_SUMB_4__14_), .CO(
        mul_ex_mult_76_CARRYB_5__13_), .S(mul_ex_mult_76_SUMB_5__13_) );
  FA_X1 mul_ex_mult_76_S2_5_12 ( .A(mul_ex_mult_76_ab_5__12_), .B(
        mul_ex_mult_76_CARRYB_4__12_), .CI(mul_ex_mult_76_SUMB_4__13_), .CO(
        mul_ex_mult_76_CARRYB_5__12_), .S(mul_ex_mult_76_SUMB_5__12_) );
  FA_X1 mul_ex_mult_76_S2_5_11 ( .A(mul_ex_mult_76_ab_5__11_), .B(
        mul_ex_mult_76_CARRYB_4__11_), .CI(mul_ex_mult_76_SUMB_4__12_), .CO(
        mul_ex_mult_76_CARRYB_5__11_), .S(mul_ex_mult_76_SUMB_5__11_) );
  FA_X1 mul_ex_mult_76_S2_5_10 ( .A(mul_ex_mult_76_ab_5__10_), .B(
        mul_ex_mult_76_CARRYB_4__10_), .CI(mul_ex_mult_76_SUMB_4__11_), .CO(
        mul_ex_mult_76_CARRYB_5__10_), .S(mul_ex_mult_76_SUMB_5__10_) );
  FA_X1 mul_ex_mult_76_S2_5_9 ( .A(mul_ex_mult_76_ab_5__9_), .B(
        mul_ex_mult_76_CARRYB_4__9_), .CI(mul_ex_mult_76_SUMB_4__10_), .CO(
        mul_ex_mult_76_CARRYB_5__9_), .S(mul_ex_mult_76_SUMB_5__9_) );
  FA_X1 mul_ex_mult_76_S2_5_8 ( .A(mul_ex_mult_76_ab_5__8_), .B(
        mul_ex_mult_76_CARRYB_4__8_), .CI(mul_ex_mult_76_SUMB_4__9_), .CO(
        mul_ex_mult_76_CARRYB_5__8_), .S(mul_ex_mult_76_SUMB_5__8_) );
  FA_X1 mul_ex_mult_76_S2_5_7 ( .A(mul_ex_mult_76_ab_5__7_), .B(
        mul_ex_mult_76_CARRYB_4__7_), .CI(mul_ex_mult_76_SUMB_4__8_), .CO(
        mul_ex_mult_76_CARRYB_5__7_), .S(mul_ex_mult_76_SUMB_5__7_) );
  FA_X1 mul_ex_mult_76_S2_5_6 ( .A(mul_ex_mult_76_ab_5__6_), .B(
        mul_ex_mult_76_CARRYB_4__6_), .CI(mul_ex_mult_76_SUMB_4__7_), .CO(
        mul_ex_mult_76_CARRYB_5__6_), .S(mul_ex_mult_76_SUMB_5__6_) );
  FA_X1 mul_ex_mult_76_S2_5_5 ( .A(mul_ex_mult_76_ab_5__5_), .B(
        mul_ex_mult_76_CARRYB_4__5_), .CI(mul_ex_mult_76_SUMB_4__6_), .CO(
        mul_ex_mult_76_CARRYB_5__5_), .S(mul_ex_mult_76_SUMB_5__5_) );
  FA_X1 mul_ex_mult_76_S2_5_4 ( .A(mul_ex_mult_76_ab_5__4_), .B(
        mul_ex_mult_76_CARRYB_4__4_), .CI(mul_ex_mult_76_SUMB_4__5_), .CO(
        mul_ex_mult_76_CARRYB_5__4_), .S(mul_ex_mult_76_SUMB_5__4_) );
  FA_X1 mul_ex_mult_76_S2_5_3 ( .A(mul_ex_mult_76_ab_5__3_), .B(
        mul_ex_mult_76_CARRYB_4__3_), .CI(mul_ex_mult_76_SUMB_4__4_), .CO(
        mul_ex_mult_76_CARRYB_5__3_), .S(mul_ex_mult_76_SUMB_5__3_) );
  FA_X1 mul_ex_mult_76_S2_5_2 ( .A(mul_ex_mult_76_ab_5__2_), .B(
        mul_ex_mult_76_CARRYB_4__2_), .CI(mul_ex_mult_76_SUMB_4__3_), .CO(
        mul_ex_mult_76_CARRYB_5__2_), .S(mul_ex_mult_76_SUMB_5__2_) );
  FA_X1 mul_ex_mult_76_S2_5_1 ( .A(mul_ex_mult_76_ab_5__1_), .B(
        mul_ex_mult_76_CARRYB_4__1_), .CI(mul_ex_mult_76_SUMB_4__2_), .CO(
        mul_ex_mult_76_CARRYB_5__1_), .S(mul_ex_mult_76_SUMB_5__1_) );
  FA_X1 mul_ex_mult_76_S1_5_0 ( .A(mul_ex_mult_76_ab_5__0_), .B(
        mul_ex_mult_76_CARRYB_4__0_), .CI(mul_ex_mult_76_SUMB_4__1_), .CO(
        mul_ex_mult_76_CARRYB_5__0_), .S(mul_ex_mult_76_A1_3_) );
  FA_X1 mul_ex_mult_76_S3_6_14 ( .A(mul_ex_mult_76_ab_6__14_), .B(
        mul_ex_mult_76_CARRYB_5__14_), .CI(mul_ex_mult_76_ab_5__15_), .CO(
        mul_ex_mult_76_CARRYB_6__14_), .S(mul_ex_mult_76_SUMB_6__14_) );
  FA_X1 mul_ex_mult_76_S2_6_13 ( .A(mul_ex_mult_76_ab_6__13_), .B(
        mul_ex_mult_76_CARRYB_5__13_), .CI(mul_ex_mult_76_SUMB_5__14_), .CO(
        mul_ex_mult_76_CARRYB_6__13_), .S(mul_ex_mult_76_SUMB_6__13_) );
  FA_X1 mul_ex_mult_76_S2_6_12 ( .A(mul_ex_mult_76_ab_6__12_), .B(
        mul_ex_mult_76_CARRYB_5__12_), .CI(mul_ex_mult_76_SUMB_5__13_), .CO(
        mul_ex_mult_76_CARRYB_6__12_), .S(mul_ex_mult_76_SUMB_6__12_) );
  FA_X1 mul_ex_mult_76_S2_6_11 ( .A(mul_ex_mult_76_ab_6__11_), .B(
        mul_ex_mult_76_CARRYB_5__11_), .CI(mul_ex_mult_76_SUMB_5__12_), .CO(
        mul_ex_mult_76_CARRYB_6__11_), .S(mul_ex_mult_76_SUMB_6__11_) );
  FA_X1 mul_ex_mult_76_S2_6_10 ( .A(mul_ex_mult_76_ab_6__10_), .B(
        mul_ex_mult_76_CARRYB_5__10_), .CI(mul_ex_mult_76_SUMB_5__11_), .CO(
        mul_ex_mult_76_CARRYB_6__10_), .S(mul_ex_mult_76_SUMB_6__10_) );
  FA_X1 mul_ex_mult_76_S2_6_9 ( .A(mul_ex_mult_76_ab_6__9_), .B(
        mul_ex_mult_76_CARRYB_5__9_), .CI(mul_ex_mult_76_SUMB_5__10_), .CO(
        mul_ex_mult_76_CARRYB_6__9_), .S(mul_ex_mult_76_SUMB_6__9_) );
  FA_X1 mul_ex_mult_76_S2_6_8 ( .A(mul_ex_mult_76_ab_6__8_), .B(
        mul_ex_mult_76_CARRYB_5__8_), .CI(mul_ex_mult_76_SUMB_5__9_), .CO(
        mul_ex_mult_76_CARRYB_6__8_), .S(mul_ex_mult_76_SUMB_6__8_) );
  FA_X1 mul_ex_mult_76_S2_6_7 ( .A(mul_ex_mult_76_ab_6__7_), .B(
        mul_ex_mult_76_CARRYB_5__7_), .CI(mul_ex_mult_76_SUMB_5__8_), .CO(
        mul_ex_mult_76_CARRYB_6__7_), .S(mul_ex_mult_76_SUMB_6__7_) );
  FA_X1 mul_ex_mult_76_S2_6_6 ( .A(mul_ex_mult_76_ab_6__6_), .B(
        mul_ex_mult_76_CARRYB_5__6_), .CI(mul_ex_mult_76_SUMB_5__7_), .CO(
        mul_ex_mult_76_CARRYB_6__6_), .S(mul_ex_mult_76_SUMB_6__6_) );
  FA_X1 mul_ex_mult_76_S2_6_5 ( .A(mul_ex_mult_76_ab_6__5_), .B(
        mul_ex_mult_76_CARRYB_5__5_), .CI(mul_ex_mult_76_SUMB_5__6_), .CO(
        mul_ex_mult_76_CARRYB_6__5_), .S(mul_ex_mult_76_SUMB_6__5_) );
  FA_X1 mul_ex_mult_76_S2_6_4 ( .A(mul_ex_mult_76_ab_6__4_), .B(
        mul_ex_mult_76_CARRYB_5__4_), .CI(mul_ex_mult_76_SUMB_5__5_), .CO(
        mul_ex_mult_76_CARRYB_6__4_), .S(mul_ex_mult_76_SUMB_6__4_) );
  FA_X1 mul_ex_mult_76_S2_6_3 ( .A(mul_ex_mult_76_ab_6__3_), .B(
        mul_ex_mult_76_CARRYB_5__3_), .CI(mul_ex_mult_76_SUMB_5__4_), .CO(
        mul_ex_mult_76_CARRYB_6__3_), .S(mul_ex_mult_76_SUMB_6__3_) );
  FA_X1 mul_ex_mult_76_S2_6_2 ( .A(mul_ex_mult_76_ab_6__2_), .B(
        mul_ex_mult_76_CARRYB_5__2_), .CI(mul_ex_mult_76_SUMB_5__3_), .CO(
        mul_ex_mult_76_CARRYB_6__2_), .S(mul_ex_mult_76_SUMB_6__2_) );
  FA_X1 mul_ex_mult_76_S2_6_1 ( .A(mul_ex_mult_76_ab_6__1_), .B(
        mul_ex_mult_76_CARRYB_5__1_), .CI(mul_ex_mult_76_SUMB_5__2_), .CO(
        mul_ex_mult_76_CARRYB_6__1_), .S(mul_ex_mult_76_SUMB_6__1_) );
  FA_X1 mul_ex_mult_76_S1_6_0 ( .A(mul_ex_mult_76_ab_6__0_), .B(
        mul_ex_mult_76_CARRYB_5__0_), .CI(mul_ex_mult_76_SUMB_5__1_), .CO(
        mul_ex_mult_76_CARRYB_6__0_), .S(mul_ex_mult_76_A1_4_) );
  FA_X1 mul_ex_mult_76_S3_7_14 ( .A(mul_ex_mult_76_ab_7__14_), .B(
        mul_ex_mult_76_CARRYB_6__14_), .CI(mul_ex_mult_76_ab_6__15_), .CO(
        mul_ex_mult_76_CARRYB_7__14_), .S(mul_ex_mult_76_SUMB_7__14_) );
  FA_X1 mul_ex_mult_76_S2_7_13 ( .A(mul_ex_mult_76_ab_7__13_), .B(
        mul_ex_mult_76_CARRYB_6__13_), .CI(mul_ex_mult_76_SUMB_6__14_), .CO(
        mul_ex_mult_76_CARRYB_7__13_), .S(mul_ex_mult_76_SUMB_7__13_) );
  FA_X1 mul_ex_mult_76_S2_7_12 ( .A(mul_ex_mult_76_ab_7__12_), .B(
        mul_ex_mult_76_CARRYB_6__12_), .CI(mul_ex_mult_76_SUMB_6__13_), .CO(
        mul_ex_mult_76_CARRYB_7__12_), .S(mul_ex_mult_76_SUMB_7__12_) );
  FA_X1 mul_ex_mult_76_S2_7_11 ( .A(mul_ex_mult_76_ab_7__11_), .B(
        mul_ex_mult_76_CARRYB_6__11_), .CI(mul_ex_mult_76_SUMB_6__12_), .CO(
        mul_ex_mult_76_CARRYB_7__11_), .S(mul_ex_mult_76_SUMB_7__11_) );
  FA_X1 mul_ex_mult_76_S2_7_10 ( .A(mul_ex_mult_76_ab_7__10_), .B(
        mul_ex_mult_76_CARRYB_6__10_), .CI(mul_ex_mult_76_SUMB_6__11_), .CO(
        mul_ex_mult_76_CARRYB_7__10_), .S(mul_ex_mult_76_SUMB_7__10_) );
  FA_X1 mul_ex_mult_76_S2_7_9 ( .A(mul_ex_mult_76_ab_7__9_), .B(
        mul_ex_mult_76_CARRYB_6__9_), .CI(mul_ex_mult_76_SUMB_6__10_), .CO(
        mul_ex_mult_76_CARRYB_7__9_), .S(mul_ex_mult_76_SUMB_7__9_) );
  FA_X1 mul_ex_mult_76_S2_7_8 ( .A(mul_ex_mult_76_ab_7__8_), .B(
        mul_ex_mult_76_CARRYB_6__8_), .CI(mul_ex_mult_76_SUMB_6__9_), .CO(
        mul_ex_mult_76_CARRYB_7__8_), .S(mul_ex_mult_76_SUMB_7__8_) );
  FA_X1 mul_ex_mult_76_S2_7_7 ( .A(mul_ex_mult_76_ab_7__7_), .B(
        mul_ex_mult_76_CARRYB_6__7_), .CI(mul_ex_mult_76_SUMB_6__8_), .CO(
        mul_ex_mult_76_CARRYB_7__7_), .S(mul_ex_mult_76_SUMB_7__7_) );
  FA_X1 mul_ex_mult_76_S2_7_6 ( .A(mul_ex_mult_76_ab_7__6_), .B(
        mul_ex_mult_76_CARRYB_6__6_), .CI(mul_ex_mult_76_SUMB_6__7_), .CO(
        mul_ex_mult_76_CARRYB_7__6_), .S(mul_ex_mult_76_SUMB_7__6_) );
  FA_X1 mul_ex_mult_76_S2_7_5 ( .A(mul_ex_mult_76_ab_7__5_), .B(
        mul_ex_mult_76_CARRYB_6__5_), .CI(mul_ex_mult_76_SUMB_6__6_), .CO(
        mul_ex_mult_76_CARRYB_7__5_), .S(mul_ex_mult_76_SUMB_7__5_) );
  FA_X1 mul_ex_mult_76_S2_7_4 ( .A(mul_ex_mult_76_ab_7__4_), .B(
        mul_ex_mult_76_CARRYB_6__4_), .CI(mul_ex_mult_76_SUMB_6__5_), .CO(
        mul_ex_mult_76_CARRYB_7__4_), .S(mul_ex_mult_76_SUMB_7__4_) );
  FA_X1 mul_ex_mult_76_S2_7_3 ( .A(mul_ex_mult_76_ab_7__3_), .B(
        mul_ex_mult_76_CARRYB_6__3_), .CI(mul_ex_mult_76_SUMB_6__4_), .CO(
        mul_ex_mult_76_CARRYB_7__3_), .S(mul_ex_mult_76_SUMB_7__3_) );
  FA_X1 mul_ex_mult_76_S2_7_2 ( .A(mul_ex_mult_76_ab_7__2_), .B(
        mul_ex_mult_76_CARRYB_6__2_), .CI(mul_ex_mult_76_SUMB_6__3_), .CO(
        mul_ex_mult_76_CARRYB_7__2_), .S(mul_ex_mult_76_SUMB_7__2_) );
  FA_X1 mul_ex_mult_76_S2_7_1 ( .A(mul_ex_mult_76_ab_7__1_), .B(
        mul_ex_mult_76_CARRYB_6__1_), .CI(mul_ex_mult_76_SUMB_6__2_), .CO(
        mul_ex_mult_76_CARRYB_7__1_), .S(mul_ex_mult_76_SUMB_7__1_) );
  FA_X1 mul_ex_mult_76_S1_7_0 ( .A(mul_ex_mult_76_ab_7__0_), .B(
        mul_ex_mult_76_CARRYB_6__0_), .CI(mul_ex_mult_76_SUMB_6__1_), .CO(
        mul_ex_mult_76_CARRYB_7__0_), .S(mul_ex_mult_76_A1_5_) );
  FA_X1 mul_ex_mult_76_S3_8_14 ( .A(mul_ex_mult_76_ab_8__14_), .B(
        mul_ex_mult_76_CARRYB_7__14_), .CI(mul_ex_mult_76_ab_7__15_), .CO(
        mul_ex_mult_76_CARRYB_8__14_), .S(mul_ex_mult_76_SUMB_8__14_) );
  FA_X1 mul_ex_mult_76_S2_8_13 ( .A(mul_ex_mult_76_ab_8__13_), .B(
        mul_ex_mult_76_CARRYB_7__13_), .CI(mul_ex_mult_76_SUMB_7__14_), .CO(
        mul_ex_mult_76_CARRYB_8__13_), .S(mul_ex_mult_76_SUMB_8__13_) );
  FA_X1 mul_ex_mult_76_S2_8_12 ( .A(mul_ex_mult_76_ab_8__12_), .B(
        mul_ex_mult_76_CARRYB_7__12_), .CI(mul_ex_mult_76_SUMB_7__13_), .CO(
        mul_ex_mult_76_CARRYB_8__12_), .S(mul_ex_mult_76_SUMB_8__12_) );
  FA_X1 mul_ex_mult_76_S2_8_11 ( .A(mul_ex_mult_76_ab_8__11_), .B(
        mul_ex_mult_76_CARRYB_7__11_), .CI(mul_ex_mult_76_SUMB_7__12_), .CO(
        mul_ex_mult_76_CARRYB_8__11_), .S(mul_ex_mult_76_SUMB_8__11_) );
  FA_X1 mul_ex_mult_76_S2_8_10 ( .A(mul_ex_mult_76_ab_8__10_), .B(
        mul_ex_mult_76_CARRYB_7__10_), .CI(mul_ex_mult_76_SUMB_7__11_), .CO(
        mul_ex_mult_76_CARRYB_8__10_), .S(mul_ex_mult_76_SUMB_8__10_) );
  FA_X1 mul_ex_mult_76_S2_8_9 ( .A(mul_ex_mult_76_ab_8__9_), .B(
        mul_ex_mult_76_CARRYB_7__9_), .CI(mul_ex_mult_76_SUMB_7__10_), .CO(
        mul_ex_mult_76_CARRYB_8__9_), .S(mul_ex_mult_76_SUMB_8__9_) );
  FA_X1 mul_ex_mult_76_S2_8_8 ( .A(mul_ex_mult_76_ab_8__8_), .B(
        mul_ex_mult_76_CARRYB_7__8_), .CI(mul_ex_mult_76_SUMB_7__9_), .CO(
        mul_ex_mult_76_CARRYB_8__8_), .S(mul_ex_mult_76_SUMB_8__8_) );
  FA_X1 mul_ex_mult_76_S2_8_7 ( .A(mul_ex_mult_76_ab_8__7_), .B(
        mul_ex_mult_76_CARRYB_7__7_), .CI(mul_ex_mult_76_SUMB_7__8_), .CO(
        mul_ex_mult_76_CARRYB_8__7_), .S(mul_ex_mult_76_SUMB_8__7_) );
  FA_X1 mul_ex_mult_76_S2_8_6 ( .A(mul_ex_mult_76_ab_8__6_), .B(
        mul_ex_mult_76_CARRYB_7__6_), .CI(mul_ex_mult_76_SUMB_7__7_), .CO(
        mul_ex_mult_76_CARRYB_8__6_), .S(mul_ex_mult_76_SUMB_8__6_) );
  FA_X1 mul_ex_mult_76_S2_8_5 ( .A(mul_ex_mult_76_ab_8__5_), .B(
        mul_ex_mult_76_CARRYB_7__5_), .CI(mul_ex_mult_76_SUMB_7__6_), .CO(
        mul_ex_mult_76_CARRYB_8__5_), .S(mul_ex_mult_76_SUMB_8__5_) );
  FA_X1 mul_ex_mult_76_S2_8_4 ( .A(mul_ex_mult_76_ab_8__4_), .B(
        mul_ex_mult_76_CARRYB_7__4_), .CI(mul_ex_mult_76_SUMB_7__5_), .CO(
        mul_ex_mult_76_CARRYB_8__4_), .S(mul_ex_mult_76_SUMB_8__4_) );
  FA_X1 mul_ex_mult_76_S2_8_3 ( .A(mul_ex_mult_76_ab_8__3_), .B(
        mul_ex_mult_76_CARRYB_7__3_), .CI(mul_ex_mult_76_SUMB_7__4_), .CO(
        mul_ex_mult_76_CARRYB_8__3_), .S(mul_ex_mult_76_SUMB_8__3_) );
  FA_X1 mul_ex_mult_76_S2_8_2 ( .A(mul_ex_mult_76_ab_8__2_), .B(
        mul_ex_mult_76_CARRYB_7__2_), .CI(mul_ex_mult_76_SUMB_7__3_), .CO(
        mul_ex_mult_76_CARRYB_8__2_), .S(mul_ex_mult_76_SUMB_8__2_) );
  FA_X1 mul_ex_mult_76_S2_8_1 ( .A(mul_ex_mult_76_ab_8__1_), .B(
        mul_ex_mult_76_CARRYB_7__1_), .CI(mul_ex_mult_76_SUMB_7__2_), .CO(
        mul_ex_mult_76_CARRYB_8__1_), .S(mul_ex_mult_76_SUMB_8__1_) );
  FA_X1 mul_ex_mult_76_S1_8_0 ( .A(mul_ex_mult_76_ab_8__0_), .B(
        mul_ex_mult_76_CARRYB_7__0_), .CI(mul_ex_mult_76_SUMB_7__1_), .CO(
        mul_ex_mult_76_CARRYB_8__0_), .S(mul_ex_mult_76_A1_6_) );
  FA_X1 mul_ex_mult_76_S3_9_14 ( .A(mul_ex_mult_76_ab_9__14_), .B(
        mul_ex_mult_76_CARRYB_8__14_), .CI(mul_ex_mult_76_ab_8__15_), .CO(
        mul_ex_mult_76_CARRYB_9__14_), .S(mul_ex_mult_76_SUMB_9__14_) );
  FA_X1 mul_ex_mult_76_S2_9_13 ( .A(mul_ex_mult_76_ab_9__13_), .B(
        mul_ex_mult_76_CARRYB_8__13_), .CI(mul_ex_mult_76_SUMB_8__14_), .CO(
        mul_ex_mult_76_CARRYB_9__13_), .S(mul_ex_mult_76_SUMB_9__13_) );
  FA_X1 mul_ex_mult_76_S2_9_12 ( .A(mul_ex_mult_76_ab_9__12_), .B(
        mul_ex_mult_76_CARRYB_8__12_), .CI(mul_ex_mult_76_SUMB_8__13_), .CO(
        mul_ex_mult_76_CARRYB_9__12_), .S(mul_ex_mult_76_SUMB_9__12_) );
  FA_X1 mul_ex_mult_76_S2_9_11 ( .A(mul_ex_mult_76_ab_9__11_), .B(
        mul_ex_mult_76_CARRYB_8__11_), .CI(mul_ex_mult_76_SUMB_8__12_), .CO(
        mul_ex_mult_76_CARRYB_9__11_), .S(mul_ex_mult_76_SUMB_9__11_) );
  FA_X1 mul_ex_mult_76_S2_9_10 ( .A(mul_ex_mult_76_ab_9__10_), .B(
        mul_ex_mult_76_CARRYB_8__10_), .CI(mul_ex_mult_76_SUMB_8__11_), .CO(
        mul_ex_mult_76_CARRYB_9__10_), .S(mul_ex_mult_76_SUMB_9__10_) );
  FA_X1 mul_ex_mult_76_S2_9_9 ( .A(mul_ex_mult_76_ab_9__9_), .B(
        mul_ex_mult_76_CARRYB_8__9_), .CI(mul_ex_mult_76_SUMB_8__10_), .CO(
        mul_ex_mult_76_CARRYB_9__9_), .S(mul_ex_mult_76_SUMB_9__9_) );
  FA_X1 mul_ex_mult_76_S2_9_8 ( .A(mul_ex_mult_76_ab_9__8_), .B(
        mul_ex_mult_76_CARRYB_8__8_), .CI(mul_ex_mult_76_SUMB_8__9_), .CO(
        mul_ex_mult_76_CARRYB_9__8_), .S(mul_ex_mult_76_SUMB_9__8_) );
  FA_X1 mul_ex_mult_76_S2_9_7 ( .A(mul_ex_mult_76_ab_9__7_), .B(
        mul_ex_mult_76_CARRYB_8__7_), .CI(mul_ex_mult_76_SUMB_8__8_), .CO(
        mul_ex_mult_76_CARRYB_9__7_), .S(mul_ex_mult_76_SUMB_9__7_) );
  FA_X1 mul_ex_mult_76_S2_9_6 ( .A(mul_ex_mult_76_ab_9__6_), .B(
        mul_ex_mult_76_CARRYB_8__6_), .CI(mul_ex_mult_76_SUMB_8__7_), .CO(
        mul_ex_mult_76_CARRYB_9__6_), .S(mul_ex_mult_76_SUMB_9__6_) );
  FA_X1 mul_ex_mult_76_S2_9_5 ( .A(mul_ex_mult_76_ab_9__5_), .B(
        mul_ex_mult_76_CARRYB_8__5_), .CI(mul_ex_mult_76_SUMB_8__6_), .CO(
        mul_ex_mult_76_CARRYB_9__5_), .S(mul_ex_mult_76_SUMB_9__5_) );
  FA_X1 mul_ex_mult_76_S2_9_4 ( .A(mul_ex_mult_76_ab_9__4_), .B(
        mul_ex_mult_76_CARRYB_8__4_), .CI(mul_ex_mult_76_SUMB_8__5_), .CO(
        mul_ex_mult_76_CARRYB_9__4_), .S(mul_ex_mult_76_SUMB_9__4_) );
  FA_X1 mul_ex_mult_76_S2_9_3 ( .A(mul_ex_mult_76_ab_9__3_), .B(
        mul_ex_mult_76_CARRYB_8__3_), .CI(mul_ex_mult_76_SUMB_8__4_), .CO(
        mul_ex_mult_76_CARRYB_9__3_), .S(mul_ex_mult_76_SUMB_9__3_) );
  FA_X1 mul_ex_mult_76_S2_9_2 ( .A(mul_ex_mult_76_ab_9__2_), .B(
        mul_ex_mult_76_CARRYB_8__2_), .CI(mul_ex_mult_76_SUMB_8__3_), .CO(
        mul_ex_mult_76_CARRYB_9__2_), .S(mul_ex_mult_76_SUMB_9__2_) );
  FA_X1 mul_ex_mult_76_S2_9_1 ( .A(mul_ex_mult_76_ab_9__1_), .B(
        mul_ex_mult_76_CARRYB_8__1_), .CI(mul_ex_mult_76_SUMB_8__2_), .CO(
        mul_ex_mult_76_CARRYB_9__1_), .S(mul_ex_mult_76_SUMB_9__1_) );
  FA_X1 mul_ex_mult_76_S1_9_0 ( .A(mul_ex_mult_76_ab_9__0_), .B(
        mul_ex_mult_76_CARRYB_8__0_), .CI(mul_ex_mult_76_SUMB_8__1_), .CO(
        mul_ex_mult_76_CARRYB_9__0_), .S(mul_ex_mult_76_A1_7_) );
  FA_X1 mul_ex_mult_76_S3_10_14 ( .A(mul_ex_mult_76_ab_10__14_), .B(
        mul_ex_mult_76_CARRYB_9__14_), .CI(mul_ex_mult_76_ab_9__15_), .CO(
        mul_ex_mult_76_CARRYB_10__14_), .S(mul_ex_mult_76_SUMB_10__14_) );
  FA_X1 mul_ex_mult_76_S2_10_13 ( .A(mul_ex_mult_76_ab_10__13_), .B(
        mul_ex_mult_76_CARRYB_9__13_), .CI(mul_ex_mult_76_SUMB_9__14_), .CO(
        mul_ex_mult_76_CARRYB_10__13_), .S(mul_ex_mult_76_SUMB_10__13_) );
  FA_X1 mul_ex_mult_76_S2_10_12 ( .A(mul_ex_mult_76_ab_10__12_), .B(
        mul_ex_mult_76_CARRYB_9__12_), .CI(mul_ex_mult_76_SUMB_9__13_), .CO(
        mul_ex_mult_76_CARRYB_10__12_), .S(mul_ex_mult_76_SUMB_10__12_) );
  FA_X1 mul_ex_mult_76_S2_10_11 ( .A(mul_ex_mult_76_ab_10__11_), .B(
        mul_ex_mult_76_CARRYB_9__11_), .CI(mul_ex_mult_76_SUMB_9__12_), .CO(
        mul_ex_mult_76_CARRYB_10__11_), .S(mul_ex_mult_76_SUMB_10__11_) );
  FA_X1 mul_ex_mult_76_S2_10_10 ( .A(mul_ex_mult_76_ab_10__10_), .B(
        mul_ex_mult_76_CARRYB_9__10_), .CI(mul_ex_mult_76_SUMB_9__11_), .CO(
        mul_ex_mult_76_CARRYB_10__10_), .S(mul_ex_mult_76_SUMB_10__10_) );
  FA_X1 mul_ex_mult_76_S2_10_9 ( .A(mul_ex_mult_76_ab_10__9_), .B(
        mul_ex_mult_76_CARRYB_9__9_), .CI(mul_ex_mult_76_SUMB_9__10_), .CO(
        mul_ex_mult_76_CARRYB_10__9_), .S(mul_ex_mult_76_SUMB_10__9_) );
  FA_X1 mul_ex_mult_76_S2_10_8 ( .A(mul_ex_mult_76_ab_10__8_), .B(
        mul_ex_mult_76_CARRYB_9__8_), .CI(mul_ex_mult_76_SUMB_9__9_), .CO(
        mul_ex_mult_76_CARRYB_10__8_), .S(mul_ex_mult_76_SUMB_10__8_) );
  FA_X1 mul_ex_mult_76_S2_10_7 ( .A(mul_ex_mult_76_ab_10__7_), .B(
        mul_ex_mult_76_CARRYB_9__7_), .CI(mul_ex_mult_76_SUMB_9__8_), .CO(
        mul_ex_mult_76_CARRYB_10__7_), .S(mul_ex_mult_76_SUMB_10__7_) );
  FA_X1 mul_ex_mult_76_S2_10_6 ( .A(mul_ex_mult_76_ab_10__6_), .B(
        mul_ex_mult_76_CARRYB_9__6_), .CI(mul_ex_mult_76_SUMB_9__7_), .CO(
        mul_ex_mult_76_CARRYB_10__6_), .S(mul_ex_mult_76_SUMB_10__6_) );
  FA_X1 mul_ex_mult_76_S2_10_5 ( .A(mul_ex_mult_76_ab_10__5_), .B(
        mul_ex_mult_76_CARRYB_9__5_), .CI(mul_ex_mult_76_SUMB_9__6_), .CO(
        mul_ex_mult_76_CARRYB_10__5_), .S(mul_ex_mult_76_SUMB_10__5_) );
  FA_X1 mul_ex_mult_76_S2_10_4 ( .A(mul_ex_mult_76_ab_10__4_), .B(
        mul_ex_mult_76_CARRYB_9__4_), .CI(mul_ex_mult_76_SUMB_9__5_), .CO(
        mul_ex_mult_76_CARRYB_10__4_), .S(mul_ex_mult_76_SUMB_10__4_) );
  FA_X1 mul_ex_mult_76_S2_10_3 ( .A(mul_ex_mult_76_ab_10__3_), .B(
        mul_ex_mult_76_CARRYB_9__3_), .CI(mul_ex_mult_76_SUMB_9__4_), .CO(
        mul_ex_mult_76_CARRYB_10__3_), .S(mul_ex_mult_76_SUMB_10__3_) );
  FA_X1 mul_ex_mult_76_S2_10_2 ( .A(mul_ex_mult_76_ab_10__2_), .B(
        mul_ex_mult_76_CARRYB_9__2_), .CI(mul_ex_mult_76_SUMB_9__3_), .CO(
        mul_ex_mult_76_CARRYB_10__2_), .S(mul_ex_mult_76_SUMB_10__2_) );
  FA_X1 mul_ex_mult_76_S2_10_1 ( .A(mul_ex_mult_76_ab_10__1_), .B(
        mul_ex_mult_76_CARRYB_9__1_), .CI(mul_ex_mult_76_SUMB_9__2_), .CO(
        mul_ex_mult_76_CARRYB_10__1_), .S(mul_ex_mult_76_SUMB_10__1_) );
  FA_X1 mul_ex_mult_76_S1_10_0 ( .A(mul_ex_mult_76_ab_10__0_), .B(
        mul_ex_mult_76_CARRYB_9__0_), .CI(mul_ex_mult_76_SUMB_9__1_), .CO(
        mul_ex_mult_76_CARRYB_10__0_), .S(mul_ex_mult_76_A1_8_) );
  FA_X1 mul_ex_mult_76_S3_11_14 ( .A(mul_ex_mult_76_ab_11__14_), .B(
        mul_ex_mult_76_CARRYB_10__14_), .CI(mul_ex_mult_76_ab_10__15_), .CO(
        mul_ex_mult_76_CARRYB_11__14_), .S(mul_ex_mult_76_SUMB_11__14_) );
  FA_X1 mul_ex_mult_76_S2_11_13 ( .A(mul_ex_mult_76_ab_11__13_), .B(
        mul_ex_mult_76_CARRYB_10__13_), .CI(mul_ex_mult_76_SUMB_10__14_), .CO(
        mul_ex_mult_76_CARRYB_11__13_), .S(mul_ex_mult_76_SUMB_11__13_) );
  FA_X1 mul_ex_mult_76_S2_11_12 ( .A(mul_ex_mult_76_ab_11__12_), .B(
        mul_ex_mult_76_CARRYB_10__12_), .CI(mul_ex_mult_76_SUMB_10__13_), .CO(
        mul_ex_mult_76_CARRYB_11__12_), .S(mul_ex_mult_76_SUMB_11__12_) );
  FA_X1 mul_ex_mult_76_S2_11_11 ( .A(mul_ex_mult_76_ab_11__11_), .B(
        mul_ex_mult_76_CARRYB_10__11_), .CI(mul_ex_mult_76_SUMB_10__12_), .CO(
        mul_ex_mult_76_CARRYB_11__11_), .S(mul_ex_mult_76_SUMB_11__11_) );
  FA_X1 mul_ex_mult_76_S2_11_10 ( .A(mul_ex_mult_76_ab_11__10_), .B(
        mul_ex_mult_76_CARRYB_10__10_), .CI(mul_ex_mult_76_SUMB_10__11_), .CO(
        mul_ex_mult_76_CARRYB_11__10_), .S(mul_ex_mult_76_SUMB_11__10_) );
  FA_X1 mul_ex_mult_76_S2_11_9 ( .A(mul_ex_mult_76_ab_11__9_), .B(
        mul_ex_mult_76_CARRYB_10__9_), .CI(mul_ex_mult_76_SUMB_10__10_), .CO(
        mul_ex_mult_76_CARRYB_11__9_), .S(mul_ex_mult_76_SUMB_11__9_) );
  FA_X1 mul_ex_mult_76_S2_11_8 ( .A(mul_ex_mult_76_ab_11__8_), .B(
        mul_ex_mult_76_CARRYB_10__8_), .CI(mul_ex_mult_76_SUMB_10__9_), .CO(
        mul_ex_mult_76_CARRYB_11__8_), .S(mul_ex_mult_76_SUMB_11__8_) );
  FA_X1 mul_ex_mult_76_S2_11_7 ( .A(mul_ex_mult_76_ab_11__7_), .B(
        mul_ex_mult_76_CARRYB_10__7_), .CI(mul_ex_mult_76_SUMB_10__8_), .CO(
        mul_ex_mult_76_CARRYB_11__7_), .S(mul_ex_mult_76_SUMB_11__7_) );
  FA_X1 mul_ex_mult_76_S2_11_6 ( .A(mul_ex_mult_76_ab_11__6_), .B(
        mul_ex_mult_76_CARRYB_10__6_), .CI(mul_ex_mult_76_SUMB_10__7_), .CO(
        mul_ex_mult_76_CARRYB_11__6_), .S(mul_ex_mult_76_SUMB_11__6_) );
  FA_X1 mul_ex_mult_76_S2_11_5 ( .A(mul_ex_mult_76_ab_11__5_), .B(
        mul_ex_mult_76_CARRYB_10__5_), .CI(mul_ex_mult_76_SUMB_10__6_), .CO(
        mul_ex_mult_76_CARRYB_11__5_), .S(mul_ex_mult_76_SUMB_11__5_) );
  FA_X1 mul_ex_mult_76_S2_11_4 ( .A(mul_ex_mult_76_ab_11__4_), .B(
        mul_ex_mult_76_CARRYB_10__4_), .CI(mul_ex_mult_76_SUMB_10__5_), .CO(
        mul_ex_mult_76_CARRYB_11__4_), .S(mul_ex_mult_76_SUMB_11__4_) );
  FA_X1 mul_ex_mult_76_S2_11_3 ( .A(mul_ex_mult_76_ab_11__3_), .B(
        mul_ex_mult_76_CARRYB_10__3_), .CI(mul_ex_mult_76_SUMB_10__4_), .CO(
        mul_ex_mult_76_CARRYB_11__3_), .S(mul_ex_mult_76_SUMB_11__3_) );
  FA_X1 mul_ex_mult_76_S2_11_2 ( .A(mul_ex_mult_76_ab_11__2_), .B(
        mul_ex_mult_76_CARRYB_10__2_), .CI(mul_ex_mult_76_SUMB_10__3_), .CO(
        mul_ex_mult_76_CARRYB_11__2_), .S(mul_ex_mult_76_SUMB_11__2_) );
  FA_X1 mul_ex_mult_76_S2_11_1 ( .A(mul_ex_mult_76_ab_11__1_), .B(
        mul_ex_mult_76_CARRYB_10__1_), .CI(mul_ex_mult_76_SUMB_10__2_), .CO(
        mul_ex_mult_76_CARRYB_11__1_), .S(mul_ex_mult_76_SUMB_11__1_) );
  FA_X1 mul_ex_mult_76_S1_11_0 ( .A(mul_ex_mult_76_ab_11__0_), .B(
        mul_ex_mult_76_CARRYB_10__0_), .CI(mul_ex_mult_76_SUMB_10__1_), .CO(
        mul_ex_mult_76_CARRYB_11__0_), .S(mul_ex_mult_76_A1_9_) );
  FA_X1 mul_ex_mult_76_S3_12_14 ( .A(mul_ex_mult_76_ab_12__14_), .B(
        mul_ex_mult_76_CARRYB_11__14_), .CI(mul_ex_mult_76_ab_11__15_), .CO(
        mul_ex_mult_76_CARRYB_12__14_), .S(mul_ex_mult_76_SUMB_12__14_) );
  FA_X1 mul_ex_mult_76_S2_12_13 ( .A(mul_ex_mult_76_ab_12__13_), .B(
        mul_ex_mult_76_CARRYB_11__13_), .CI(mul_ex_mult_76_SUMB_11__14_), .CO(
        mul_ex_mult_76_CARRYB_12__13_), .S(mul_ex_mult_76_SUMB_12__13_) );
  FA_X1 mul_ex_mult_76_S2_12_12 ( .A(mul_ex_mult_76_ab_12__12_), .B(
        mul_ex_mult_76_CARRYB_11__12_), .CI(mul_ex_mult_76_SUMB_11__13_), .CO(
        mul_ex_mult_76_CARRYB_12__12_), .S(mul_ex_mult_76_SUMB_12__12_) );
  FA_X1 mul_ex_mult_76_S2_12_11 ( .A(mul_ex_mult_76_ab_12__11_), .B(
        mul_ex_mult_76_CARRYB_11__11_), .CI(mul_ex_mult_76_SUMB_11__12_), .CO(
        mul_ex_mult_76_CARRYB_12__11_), .S(mul_ex_mult_76_SUMB_12__11_) );
  FA_X1 mul_ex_mult_76_S2_12_10 ( .A(mul_ex_mult_76_ab_12__10_), .B(
        mul_ex_mult_76_CARRYB_11__10_), .CI(mul_ex_mult_76_SUMB_11__11_), .CO(
        mul_ex_mult_76_CARRYB_12__10_), .S(mul_ex_mult_76_SUMB_12__10_) );
  FA_X1 mul_ex_mult_76_S2_12_9 ( .A(mul_ex_mult_76_ab_12__9_), .B(
        mul_ex_mult_76_CARRYB_11__9_), .CI(mul_ex_mult_76_SUMB_11__10_), .CO(
        mul_ex_mult_76_CARRYB_12__9_), .S(mul_ex_mult_76_SUMB_12__9_) );
  FA_X1 mul_ex_mult_76_S2_12_8 ( .A(mul_ex_mult_76_ab_12__8_), .B(
        mul_ex_mult_76_CARRYB_11__8_), .CI(mul_ex_mult_76_SUMB_11__9_), .CO(
        mul_ex_mult_76_CARRYB_12__8_), .S(mul_ex_mult_76_SUMB_12__8_) );
  FA_X1 mul_ex_mult_76_S2_12_7 ( .A(mul_ex_mult_76_ab_12__7_), .B(
        mul_ex_mult_76_CARRYB_11__7_), .CI(mul_ex_mult_76_SUMB_11__8_), .CO(
        mul_ex_mult_76_CARRYB_12__7_), .S(mul_ex_mult_76_SUMB_12__7_) );
  FA_X1 mul_ex_mult_76_S2_12_6 ( .A(mul_ex_mult_76_ab_12__6_), .B(
        mul_ex_mult_76_CARRYB_11__6_), .CI(mul_ex_mult_76_SUMB_11__7_), .CO(
        mul_ex_mult_76_CARRYB_12__6_), .S(mul_ex_mult_76_SUMB_12__6_) );
  FA_X1 mul_ex_mult_76_S2_12_5 ( .A(mul_ex_mult_76_ab_12__5_), .B(
        mul_ex_mult_76_CARRYB_11__5_), .CI(mul_ex_mult_76_SUMB_11__6_), .CO(
        mul_ex_mult_76_CARRYB_12__5_), .S(mul_ex_mult_76_SUMB_12__5_) );
  FA_X1 mul_ex_mult_76_S2_12_4 ( .A(mul_ex_mult_76_ab_12__4_), .B(
        mul_ex_mult_76_CARRYB_11__4_), .CI(mul_ex_mult_76_SUMB_11__5_), .CO(
        mul_ex_mult_76_CARRYB_12__4_), .S(mul_ex_mult_76_SUMB_12__4_) );
  FA_X1 mul_ex_mult_76_S2_12_3 ( .A(mul_ex_mult_76_ab_12__3_), .B(
        mul_ex_mult_76_CARRYB_11__3_), .CI(mul_ex_mult_76_SUMB_11__4_), .CO(
        mul_ex_mult_76_CARRYB_12__3_), .S(mul_ex_mult_76_SUMB_12__3_) );
  FA_X1 mul_ex_mult_76_S2_12_2 ( .A(mul_ex_mult_76_ab_12__2_), .B(
        mul_ex_mult_76_CARRYB_11__2_), .CI(mul_ex_mult_76_SUMB_11__3_), .CO(
        mul_ex_mult_76_CARRYB_12__2_), .S(mul_ex_mult_76_SUMB_12__2_) );
  FA_X1 mul_ex_mult_76_S2_12_1 ( .A(mul_ex_mult_76_ab_12__1_), .B(
        mul_ex_mult_76_CARRYB_11__1_), .CI(mul_ex_mult_76_SUMB_11__2_), .CO(
        mul_ex_mult_76_CARRYB_12__1_), .S(mul_ex_mult_76_SUMB_12__1_) );
  FA_X1 mul_ex_mult_76_S1_12_0 ( .A(mul_ex_mult_76_ab_12__0_), .B(
        mul_ex_mult_76_CARRYB_11__0_), .CI(mul_ex_mult_76_SUMB_11__1_), .CO(
        mul_ex_mult_76_CARRYB_12__0_), .S(mul_ex_mult_76_A1_10_) );
  FA_X1 mul_ex_mult_76_S3_13_14 ( .A(mul_ex_mult_76_ab_13__14_), .B(
        mul_ex_mult_76_CARRYB_12__14_), .CI(mul_ex_mult_76_ab_12__15_), .CO(
        mul_ex_mult_76_CARRYB_13__14_), .S(mul_ex_mult_76_SUMB_13__14_) );
  FA_X1 mul_ex_mult_76_S2_13_13 ( .A(mul_ex_mult_76_ab_13__13_), .B(
        mul_ex_mult_76_CARRYB_12__13_), .CI(mul_ex_mult_76_SUMB_12__14_), .CO(
        mul_ex_mult_76_CARRYB_13__13_), .S(mul_ex_mult_76_SUMB_13__13_) );
  FA_X1 mul_ex_mult_76_S2_13_12 ( .A(mul_ex_mult_76_ab_13__12_), .B(
        mul_ex_mult_76_CARRYB_12__12_), .CI(mul_ex_mult_76_SUMB_12__13_), .CO(
        mul_ex_mult_76_CARRYB_13__12_), .S(mul_ex_mult_76_SUMB_13__12_) );
  FA_X1 mul_ex_mult_76_S2_13_11 ( .A(mul_ex_mult_76_ab_13__11_), .B(
        mul_ex_mult_76_CARRYB_12__11_), .CI(mul_ex_mult_76_SUMB_12__12_), .CO(
        mul_ex_mult_76_CARRYB_13__11_), .S(mul_ex_mult_76_SUMB_13__11_) );
  FA_X1 mul_ex_mult_76_S2_13_10 ( .A(mul_ex_mult_76_ab_13__10_), .B(
        mul_ex_mult_76_CARRYB_12__10_), .CI(mul_ex_mult_76_SUMB_12__11_), .CO(
        mul_ex_mult_76_CARRYB_13__10_), .S(mul_ex_mult_76_SUMB_13__10_) );
  FA_X1 mul_ex_mult_76_S2_13_9 ( .A(mul_ex_mult_76_ab_13__9_), .B(
        mul_ex_mult_76_CARRYB_12__9_), .CI(mul_ex_mult_76_SUMB_12__10_), .CO(
        mul_ex_mult_76_CARRYB_13__9_), .S(mul_ex_mult_76_SUMB_13__9_) );
  FA_X1 mul_ex_mult_76_S2_13_8 ( .A(mul_ex_mult_76_ab_13__8_), .B(
        mul_ex_mult_76_CARRYB_12__8_), .CI(mul_ex_mult_76_SUMB_12__9_), .CO(
        mul_ex_mult_76_CARRYB_13__8_), .S(mul_ex_mult_76_SUMB_13__8_) );
  FA_X1 mul_ex_mult_76_S2_13_7 ( .A(mul_ex_mult_76_ab_13__7_), .B(
        mul_ex_mult_76_CARRYB_12__7_), .CI(mul_ex_mult_76_SUMB_12__8_), .CO(
        mul_ex_mult_76_CARRYB_13__7_), .S(mul_ex_mult_76_SUMB_13__7_) );
  FA_X1 mul_ex_mult_76_S2_13_6 ( .A(mul_ex_mult_76_ab_13__6_), .B(
        mul_ex_mult_76_CARRYB_12__6_), .CI(mul_ex_mult_76_SUMB_12__7_), .CO(
        mul_ex_mult_76_CARRYB_13__6_), .S(mul_ex_mult_76_SUMB_13__6_) );
  FA_X1 mul_ex_mult_76_S2_13_5 ( .A(mul_ex_mult_76_ab_13__5_), .B(
        mul_ex_mult_76_CARRYB_12__5_), .CI(mul_ex_mult_76_SUMB_12__6_), .CO(
        mul_ex_mult_76_CARRYB_13__5_), .S(mul_ex_mult_76_SUMB_13__5_) );
  FA_X1 mul_ex_mult_76_S2_13_4 ( .A(mul_ex_mult_76_ab_13__4_), .B(
        mul_ex_mult_76_CARRYB_12__4_), .CI(mul_ex_mult_76_SUMB_12__5_), .CO(
        mul_ex_mult_76_CARRYB_13__4_), .S(mul_ex_mult_76_SUMB_13__4_) );
  FA_X1 mul_ex_mult_76_S2_13_3 ( .A(mul_ex_mult_76_ab_13__3_), .B(
        mul_ex_mult_76_CARRYB_12__3_), .CI(mul_ex_mult_76_SUMB_12__4_), .CO(
        mul_ex_mult_76_CARRYB_13__3_), .S(mul_ex_mult_76_SUMB_13__3_) );
  FA_X1 mul_ex_mult_76_S2_13_2 ( .A(mul_ex_mult_76_ab_13__2_), .B(
        mul_ex_mult_76_CARRYB_12__2_), .CI(mul_ex_mult_76_SUMB_12__3_), .CO(
        mul_ex_mult_76_CARRYB_13__2_), .S(mul_ex_mult_76_SUMB_13__2_) );
  FA_X1 mul_ex_mult_76_S2_13_1 ( .A(mul_ex_mult_76_ab_13__1_), .B(
        mul_ex_mult_76_CARRYB_12__1_), .CI(mul_ex_mult_76_SUMB_12__2_), .CO(
        mul_ex_mult_76_CARRYB_13__1_), .S(mul_ex_mult_76_SUMB_13__1_) );
  FA_X1 mul_ex_mult_76_S1_13_0 ( .A(mul_ex_mult_76_ab_13__0_), .B(
        mul_ex_mult_76_CARRYB_12__0_), .CI(mul_ex_mult_76_SUMB_12__1_), .CO(
        mul_ex_mult_76_CARRYB_13__0_), .S(mul_ex_mult_76_A1_11_) );
  FA_X1 mul_ex_mult_76_S3_14_14 ( .A(mul_ex_mult_76_ab_14__14_), .B(
        mul_ex_mult_76_CARRYB_13__14_), .CI(mul_ex_mult_76_ab_13__15_), .CO(
        mul_ex_mult_76_CARRYB_14__14_), .S(mul_ex_mult_76_SUMB_14__14_) );
  FA_X1 mul_ex_mult_76_S2_14_13 ( .A(mul_ex_mult_76_ab_14__13_), .B(
        mul_ex_mult_76_CARRYB_13__13_), .CI(mul_ex_mult_76_SUMB_13__14_), .CO(
        mul_ex_mult_76_CARRYB_14__13_), .S(mul_ex_mult_76_SUMB_14__13_) );
  FA_X1 mul_ex_mult_76_S2_14_12 ( .A(mul_ex_mult_76_ab_14__12_), .B(
        mul_ex_mult_76_CARRYB_13__12_), .CI(mul_ex_mult_76_SUMB_13__13_), .CO(
        mul_ex_mult_76_CARRYB_14__12_), .S(mul_ex_mult_76_SUMB_14__12_) );
  FA_X1 mul_ex_mult_76_S2_14_11 ( .A(mul_ex_mult_76_ab_14__11_), .B(
        mul_ex_mult_76_CARRYB_13__11_), .CI(mul_ex_mult_76_SUMB_13__12_), .CO(
        mul_ex_mult_76_CARRYB_14__11_), .S(mul_ex_mult_76_SUMB_14__11_) );
  FA_X1 mul_ex_mult_76_S2_14_10 ( .A(mul_ex_mult_76_ab_14__10_), .B(
        mul_ex_mult_76_CARRYB_13__10_), .CI(mul_ex_mult_76_SUMB_13__11_), .CO(
        mul_ex_mult_76_CARRYB_14__10_), .S(mul_ex_mult_76_SUMB_14__10_) );
  FA_X1 mul_ex_mult_76_S2_14_9 ( .A(mul_ex_mult_76_ab_14__9_), .B(
        mul_ex_mult_76_CARRYB_13__9_), .CI(mul_ex_mult_76_SUMB_13__10_), .CO(
        mul_ex_mult_76_CARRYB_14__9_), .S(mul_ex_mult_76_SUMB_14__9_) );
  FA_X1 mul_ex_mult_76_S2_14_8 ( .A(mul_ex_mult_76_ab_14__8_), .B(
        mul_ex_mult_76_CARRYB_13__8_), .CI(mul_ex_mult_76_SUMB_13__9_), .CO(
        mul_ex_mult_76_CARRYB_14__8_), .S(mul_ex_mult_76_SUMB_14__8_) );
  FA_X1 mul_ex_mult_76_S2_14_7 ( .A(mul_ex_mult_76_ab_14__7_), .B(
        mul_ex_mult_76_CARRYB_13__7_), .CI(mul_ex_mult_76_SUMB_13__8_), .CO(
        mul_ex_mult_76_CARRYB_14__7_), .S(mul_ex_mult_76_SUMB_14__7_) );
  FA_X1 mul_ex_mult_76_S2_14_6 ( .A(mul_ex_mult_76_ab_14__6_), .B(
        mul_ex_mult_76_CARRYB_13__6_), .CI(mul_ex_mult_76_SUMB_13__7_), .CO(
        mul_ex_mult_76_CARRYB_14__6_), .S(mul_ex_mult_76_SUMB_14__6_) );
  FA_X1 mul_ex_mult_76_S2_14_5 ( .A(mul_ex_mult_76_ab_14__5_), .B(
        mul_ex_mult_76_CARRYB_13__5_), .CI(mul_ex_mult_76_SUMB_13__6_), .CO(
        mul_ex_mult_76_CARRYB_14__5_), .S(mul_ex_mult_76_SUMB_14__5_) );
  FA_X1 mul_ex_mult_76_S2_14_4 ( .A(mul_ex_mult_76_ab_14__4_), .B(
        mul_ex_mult_76_CARRYB_13__4_), .CI(mul_ex_mult_76_SUMB_13__5_), .CO(
        mul_ex_mult_76_CARRYB_14__4_), .S(mul_ex_mult_76_SUMB_14__4_) );
  FA_X1 mul_ex_mult_76_S2_14_3 ( .A(mul_ex_mult_76_ab_14__3_), .B(
        mul_ex_mult_76_CARRYB_13__3_), .CI(mul_ex_mult_76_SUMB_13__4_), .CO(
        mul_ex_mult_76_CARRYB_14__3_), .S(mul_ex_mult_76_SUMB_14__3_) );
  FA_X1 mul_ex_mult_76_S2_14_2 ( .A(mul_ex_mult_76_ab_14__2_), .B(
        mul_ex_mult_76_CARRYB_13__2_), .CI(mul_ex_mult_76_SUMB_13__3_), .CO(
        mul_ex_mult_76_CARRYB_14__2_), .S(mul_ex_mult_76_SUMB_14__2_) );
  FA_X1 mul_ex_mult_76_S2_14_1 ( .A(mul_ex_mult_76_ab_14__1_), .B(
        mul_ex_mult_76_CARRYB_13__1_), .CI(mul_ex_mult_76_SUMB_13__2_), .CO(
        mul_ex_mult_76_CARRYB_14__1_), .S(mul_ex_mult_76_SUMB_14__1_) );
  FA_X1 mul_ex_mult_76_S1_14_0 ( .A(mul_ex_mult_76_ab_14__0_), .B(
        mul_ex_mult_76_CARRYB_13__0_), .CI(mul_ex_mult_76_SUMB_13__1_), .CO(
        mul_ex_mult_76_CARRYB_14__0_), .S(mul_ex_mult_76_A1_12_) );
  FA_X1 mul_ex_mult_76_S5_14 ( .A(mul_ex_mult_76_ab_15__14_), .B(
        mul_ex_mult_76_CARRYB_14__14_), .CI(mul_ex_mult_76_ab_14__15_), .CO(
        mul_ex_mult_76_CARRYB_15__14_), .S(mul_ex_mult_76_SUMB_15__14_) );
  FA_X1 mul_ex_mult_76_S4_13 ( .A(mul_ex_mult_76_ab_15__13_), .B(
        mul_ex_mult_76_CARRYB_14__13_), .CI(mul_ex_mult_76_SUMB_14__14_), .CO(
        mul_ex_mult_76_CARRYB_15__13_), .S(mul_ex_mult_76_SUMB_15__13_) );
  FA_X1 mul_ex_mult_76_S4_12 ( .A(mul_ex_mult_76_ab_15__12_), .B(
        mul_ex_mult_76_CARRYB_14__12_), .CI(mul_ex_mult_76_SUMB_14__13_), .CO(
        mul_ex_mult_76_CARRYB_15__12_), .S(mul_ex_mult_76_SUMB_15__12_) );
  FA_X1 mul_ex_mult_76_S4_11 ( .A(mul_ex_mult_76_ab_15__11_), .B(
        mul_ex_mult_76_CARRYB_14__11_), .CI(mul_ex_mult_76_SUMB_14__12_), .CO(
        mul_ex_mult_76_CARRYB_15__11_), .S(mul_ex_mult_76_SUMB_15__11_) );
  FA_X1 mul_ex_mult_76_S4_10 ( .A(mul_ex_mult_76_ab_15__10_), .B(
        mul_ex_mult_76_CARRYB_14__10_), .CI(mul_ex_mult_76_SUMB_14__11_), .CO(
        mul_ex_mult_76_CARRYB_15__10_), .S(mul_ex_mult_76_SUMB_15__10_) );
  FA_X1 mul_ex_mult_76_S4_9 ( .A(mul_ex_mult_76_ab_15__9_), .B(
        mul_ex_mult_76_CARRYB_14__9_), .CI(mul_ex_mult_76_SUMB_14__10_), .CO(
        mul_ex_mult_76_CARRYB_15__9_), .S(mul_ex_mult_76_SUMB_15__9_) );
  FA_X1 mul_ex_mult_76_S4_8 ( .A(mul_ex_mult_76_ab_15__8_), .B(
        mul_ex_mult_76_CARRYB_14__8_), .CI(mul_ex_mult_76_SUMB_14__9_), .CO(
        mul_ex_mult_76_CARRYB_15__8_), .S(mul_ex_mult_76_SUMB_15__8_) );
  FA_X1 mul_ex_mult_76_S4_7 ( .A(mul_ex_mult_76_ab_15__7_), .B(
        mul_ex_mult_76_CARRYB_14__7_), .CI(mul_ex_mult_76_SUMB_14__8_), .CO(
        mul_ex_mult_76_CARRYB_15__7_), .S(mul_ex_mult_76_SUMB_15__7_) );
  FA_X1 mul_ex_mult_76_S4_6 ( .A(mul_ex_mult_76_ab_15__6_), .B(
        mul_ex_mult_76_CARRYB_14__6_), .CI(mul_ex_mult_76_SUMB_14__7_), .CO(
        mul_ex_mult_76_CARRYB_15__6_), .S(mul_ex_mult_76_SUMB_15__6_) );
  FA_X1 mul_ex_mult_76_S4_5 ( .A(mul_ex_mult_76_ab_15__5_), .B(
        mul_ex_mult_76_CARRYB_14__5_), .CI(mul_ex_mult_76_SUMB_14__6_), .CO(
        mul_ex_mult_76_CARRYB_15__5_), .S(mul_ex_mult_76_SUMB_15__5_) );
  FA_X1 mul_ex_mult_76_S4_4 ( .A(mul_ex_mult_76_ab_15__4_), .B(
        mul_ex_mult_76_CARRYB_14__4_), .CI(mul_ex_mult_76_SUMB_14__5_), .CO(
        mul_ex_mult_76_CARRYB_15__4_), .S(mul_ex_mult_76_SUMB_15__4_) );
  FA_X1 mul_ex_mult_76_S4_3 ( .A(mul_ex_mult_76_ab_15__3_), .B(
        mul_ex_mult_76_CARRYB_14__3_), .CI(mul_ex_mult_76_SUMB_14__4_), .CO(
        mul_ex_mult_76_CARRYB_15__3_), .S(mul_ex_mult_76_SUMB_15__3_) );
  FA_X1 mul_ex_mult_76_S4_2 ( .A(mul_ex_mult_76_ab_15__2_), .B(
        mul_ex_mult_76_CARRYB_14__2_), .CI(mul_ex_mult_76_SUMB_14__3_), .CO(
        mul_ex_mult_76_CARRYB_15__2_), .S(mul_ex_mult_76_SUMB_15__2_) );
  FA_X1 mul_ex_mult_76_S4_1 ( .A(mul_ex_mult_76_ab_15__1_), .B(
        mul_ex_mult_76_CARRYB_14__1_), .CI(mul_ex_mult_76_SUMB_14__2_), .CO(
        mul_ex_mult_76_CARRYB_15__1_), .S(mul_ex_mult_76_SUMB_15__1_) );
  FA_X1 mul_ex_mult_76_S4_0 ( .A(mul_ex_mult_76_ab_15__0_), .B(
        mul_ex_mult_76_CARRYB_14__0_), .CI(mul_ex_mult_76_SUMB_14__1_), .CO(
        mul_ex_mult_76_CARRYB_15__0_), .S(mul_ex_mult_76_SUMB_15__0_) );
  BUF_X32 mul_ex_mult_76_FS_1_U100 ( .A(mul_ex_mult_76_n61), .Z(mul_ex_N72) );
  BUF_X32 mul_ex_mult_76_FS_1_U99 ( .A(mul_ex_mult_76_SUMB_15__0_), .Z(
        mul_ex_N71) );
  BUF_X32 mul_ex_mult_76_FS_1_U98 ( .A(mul_ex_mult_76_A1_12_), .Z(mul_ex_N70)
         );
  BUF_X32 mul_ex_mult_76_FS_1_U97 ( .A(mul_ex_mult_76_A1_11_), .Z(mul_ex_N69)
         );
  BUF_X32 mul_ex_mult_76_FS_1_U96 ( .A(mul_ex_mult_76_A1_10_), .Z(mul_ex_N68)
         );
  BUF_X32 mul_ex_mult_76_FS_1_U95 ( .A(mul_ex_mult_76_A1_9_), .Z(mul_ex_N67)
         );
  BUF_X32 mul_ex_mult_76_FS_1_U94 ( .A(mul_ex_mult_76_A1_8_), .Z(mul_ex_N66)
         );
  BUF_X32 mul_ex_mult_76_FS_1_U93 ( .A(mul_ex_mult_76_A1_7_), .Z(mul_ex_N65)
         );
  BUF_X32 mul_ex_mult_76_FS_1_U92 ( .A(mul_ex_mult_76_A1_6_), .Z(mul_ex_N64)
         );
  BUF_X32 mul_ex_mult_76_FS_1_U91 ( .A(mul_ex_mult_76_A1_5_), .Z(mul_ex_N63)
         );
  BUF_X32 mul_ex_mult_76_FS_1_U90 ( .A(mul_ex_mult_76_A1_4_), .Z(mul_ex_N62)
         );
  BUF_X32 mul_ex_mult_76_FS_1_U89 ( .A(mul_ex_mult_76_A1_3_), .Z(mul_ex_N61)
         );
  BUF_X32 mul_ex_mult_76_FS_1_U88 ( .A(mul_ex_mult_76_A1_2_), .Z(mul_ex_N60)
         );
  BUF_X32 mul_ex_mult_76_FS_1_U87 ( .A(mul_ex_mult_76_A1_1_), .Z(mul_ex_N59)
         );
  BUF_X32 mul_ex_mult_76_FS_1_U86 ( .A(mul_ex_mult_76_A1_0_), .Z(mul_ex_N58)
         );
  NAND2_X1 mul_ex_mult_76_FS_1_U85 ( .A1(mul_ex_mult_76_n60), .A2(
        mul_ex_mult_76_n24), .ZN(mul_ex_mult_76_FS_1_n70) );
  AND2_X1 mul_ex_mult_76_FS_1_U84 ( .A1(mul_ex_mult_76_n53), .A2(
        mul_ex_mult_76_n23), .ZN(mul_ex_mult_76_FS_1_n67) );
  NOR2_X1 mul_ex_mult_76_FS_1_U83 ( .A1(mul_ex_mult_76_n53), .A2(
        mul_ex_mult_76_n23), .ZN(mul_ex_mult_76_FS_1_n68) );
  NOR2_X1 mul_ex_mult_76_FS_1_U82 ( .A1(mul_ex_mult_76_FS_1_n67), .A2(
        mul_ex_mult_76_FS_1_n68), .ZN(mul_ex_mult_76_FS_1_n69) );
  XOR2_X1 mul_ex_mult_76_FS_1_U81 ( .A(mul_ex_mult_76_FS_1_n17), .B(
        mul_ex_mult_76_FS_1_n69), .Z(mul_ex_N74) );
  NOR2_X1 mul_ex_mult_76_FS_1_U80 ( .A1(mul_ex_mult_76_n59), .A2(
        mul_ex_mult_76_n30), .ZN(mul_ex_mult_76_FS_1_n63) );
  NAND2_X1 mul_ex_mult_76_FS_1_U79 ( .A1(mul_ex_mult_76_n59), .A2(
        mul_ex_mult_76_n30), .ZN(mul_ex_mult_76_FS_1_n65) );
  NAND2_X1 mul_ex_mult_76_FS_1_U78 ( .A1(mul_ex_mult_76_FS_1_n15), .A2(
        mul_ex_mult_76_FS_1_n65), .ZN(mul_ex_mult_76_FS_1_n66) );
  AOI21_X1 mul_ex_mult_76_FS_1_U77 ( .B1(mul_ex_mult_76_FS_1_n16), .B2(
        mul_ex_mult_76_FS_1_n17), .A(mul_ex_mult_76_FS_1_n67), .ZN(
        mul_ex_mult_76_FS_1_n64) );
  XOR2_X1 mul_ex_mult_76_FS_1_U76 ( .A(mul_ex_mult_76_FS_1_n66), .B(
        mul_ex_mult_76_FS_1_n64), .Z(mul_ex_N75) );
  OAI21_X1 mul_ex_mult_76_FS_1_U75 ( .B1(mul_ex_mult_76_FS_1_n63), .B2(
        mul_ex_mult_76_FS_1_n64), .A(mul_ex_mult_76_FS_1_n65), .ZN(
        mul_ex_mult_76_FS_1_n59) );
  AND2_X1 mul_ex_mult_76_FS_1_U74 ( .A1(mul_ex_mult_76_n52), .A2(
        mul_ex_mult_76_n22), .ZN(mul_ex_mult_76_FS_1_n60) );
  NOR2_X1 mul_ex_mult_76_FS_1_U73 ( .A1(mul_ex_mult_76_n52), .A2(
        mul_ex_mult_76_n22), .ZN(mul_ex_mult_76_FS_1_n61) );
  NOR2_X1 mul_ex_mult_76_FS_1_U72 ( .A1(mul_ex_mult_76_FS_1_n60), .A2(
        mul_ex_mult_76_FS_1_n61), .ZN(mul_ex_mult_76_FS_1_n62) );
  XOR2_X1 mul_ex_mult_76_FS_1_U71 ( .A(mul_ex_mult_76_FS_1_n59), .B(
        mul_ex_mult_76_FS_1_n62), .Z(mul_ex_N76) );
  NOR2_X1 mul_ex_mult_76_FS_1_U70 ( .A1(mul_ex_mult_76_n58), .A2(
        mul_ex_mult_76_n29), .ZN(mul_ex_mult_76_FS_1_n55) );
  NAND2_X1 mul_ex_mult_76_FS_1_U69 ( .A1(mul_ex_mult_76_n58), .A2(
        mul_ex_mult_76_n29), .ZN(mul_ex_mult_76_FS_1_n57) );
  NAND2_X1 mul_ex_mult_76_FS_1_U68 ( .A1(mul_ex_mult_76_FS_1_n13), .A2(
        mul_ex_mult_76_FS_1_n57), .ZN(mul_ex_mult_76_FS_1_n58) );
  AOI21_X1 mul_ex_mult_76_FS_1_U67 ( .B1(mul_ex_mult_76_FS_1_n14), .B2(
        mul_ex_mult_76_FS_1_n59), .A(mul_ex_mult_76_FS_1_n60), .ZN(
        mul_ex_mult_76_FS_1_n56) );
  XOR2_X1 mul_ex_mult_76_FS_1_U66 ( .A(mul_ex_mult_76_FS_1_n58), .B(
        mul_ex_mult_76_FS_1_n56), .Z(mul_ex_N77) );
  OAI21_X1 mul_ex_mult_76_FS_1_U65 ( .B1(mul_ex_mult_76_FS_1_n55), .B2(
        mul_ex_mult_76_FS_1_n56), .A(mul_ex_mult_76_FS_1_n57), .ZN(
        mul_ex_mult_76_FS_1_n51) );
  AND2_X1 mul_ex_mult_76_FS_1_U64 ( .A1(mul_ex_mult_76_n51), .A2(
        mul_ex_mult_76_n21), .ZN(mul_ex_mult_76_FS_1_n52) );
  NOR2_X1 mul_ex_mult_76_FS_1_U63 ( .A1(mul_ex_mult_76_n51), .A2(
        mul_ex_mult_76_n21), .ZN(mul_ex_mult_76_FS_1_n53) );
  NOR2_X1 mul_ex_mult_76_FS_1_U62 ( .A1(mul_ex_mult_76_FS_1_n52), .A2(
        mul_ex_mult_76_FS_1_n53), .ZN(mul_ex_mult_76_FS_1_n54) );
  XOR2_X1 mul_ex_mult_76_FS_1_U61 ( .A(mul_ex_mult_76_FS_1_n51), .B(
        mul_ex_mult_76_FS_1_n54), .Z(mul_ex_N78) );
  NOR2_X1 mul_ex_mult_76_FS_1_U60 ( .A1(mul_ex_mult_76_n57), .A2(
        mul_ex_mult_76_n28), .ZN(mul_ex_mult_76_FS_1_n47) );
  NAND2_X1 mul_ex_mult_76_FS_1_U59 ( .A1(mul_ex_mult_76_n57), .A2(
        mul_ex_mult_76_n28), .ZN(mul_ex_mult_76_FS_1_n49) );
  NAND2_X1 mul_ex_mult_76_FS_1_U58 ( .A1(mul_ex_mult_76_FS_1_n11), .A2(
        mul_ex_mult_76_FS_1_n49), .ZN(mul_ex_mult_76_FS_1_n50) );
  AOI21_X1 mul_ex_mult_76_FS_1_U57 ( .B1(mul_ex_mult_76_FS_1_n12), .B2(
        mul_ex_mult_76_FS_1_n51), .A(mul_ex_mult_76_FS_1_n52), .ZN(
        mul_ex_mult_76_FS_1_n48) );
  XOR2_X1 mul_ex_mult_76_FS_1_U56 ( .A(mul_ex_mult_76_FS_1_n50), .B(
        mul_ex_mult_76_FS_1_n48), .Z(mul_ex_N79) );
  OAI21_X1 mul_ex_mult_76_FS_1_U55 ( .B1(mul_ex_mult_76_FS_1_n47), .B2(
        mul_ex_mult_76_FS_1_n48), .A(mul_ex_mult_76_FS_1_n49), .ZN(
        mul_ex_mult_76_FS_1_n43) );
  AND2_X1 mul_ex_mult_76_FS_1_U54 ( .A1(mul_ex_mult_76_n50), .A2(
        mul_ex_mult_76_n20), .ZN(mul_ex_mult_76_FS_1_n44) );
  NOR2_X1 mul_ex_mult_76_FS_1_U53 ( .A1(mul_ex_mult_76_n50), .A2(
        mul_ex_mult_76_n20), .ZN(mul_ex_mult_76_FS_1_n45) );
  NOR2_X1 mul_ex_mult_76_FS_1_U52 ( .A1(mul_ex_mult_76_FS_1_n44), .A2(
        mul_ex_mult_76_FS_1_n45), .ZN(mul_ex_mult_76_FS_1_n46) );
  XOR2_X1 mul_ex_mult_76_FS_1_U51 ( .A(mul_ex_mult_76_FS_1_n43), .B(
        mul_ex_mult_76_FS_1_n46), .Z(mul_ex_N80) );
  NOR2_X1 mul_ex_mult_76_FS_1_U50 ( .A1(mul_ex_mult_76_n56), .A2(
        mul_ex_mult_76_n27), .ZN(mul_ex_mult_76_FS_1_n39) );
  NAND2_X1 mul_ex_mult_76_FS_1_U49 ( .A1(mul_ex_mult_76_n56), .A2(
        mul_ex_mult_76_n27), .ZN(mul_ex_mult_76_FS_1_n41) );
  NAND2_X1 mul_ex_mult_76_FS_1_U48 ( .A1(mul_ex_mult_76_FS_1_n9), .A2(
        mul_ex_mult_76_FS_1_n41), .ZN(mul_ex_mult_76_FS_1_n42) );
  AOI21_X1 mul_ex_mult_76_FS_1_U47 ( .B1(mul_ex_mult_76_FS_1_n10), .B2(
        mul_ex_mult_76_FS_1_n43), .A(mul_ex_mult_76_FS_1_n44), .ZN(
        mul_ex_mult_76_FS_1_n40) );
  XOR2_X1 mul_ex_mult_76_FS_1_U46 ( .A(mul_ex_mult_76_FS_1_n42), .B(
        mul_ex_mult_76_FS_1_n40), .Z(mul_ex_N81) );
  OAI21_X1 mul_ex_mult_76_FS_1_U45 ( .B1(mul_ex_mult_76_FS_1_n39), .B2(
        mul_ex_mult_76_FS_1_n40), .A(mul_ex_mult_76_FS_1_n41), .ZN(
        mul_ex_mult_76_FS_1_n35) );
  AND2_X1 mul_ex_mult_76_FS_1_U44 ( .A1(mul_ex_mult_76_n49), .A2(
        mul_ex_mult_76_n19), .ZN(mul_ex_mult_76_FS_1_n36) );
  NOR2_X1 mul_ex_mult_76_FS_1_U43 ( .A1(mul_ex_mult_76_n49), .A2(
        mul_ex_mult_76_n19), .ZN(mul_ex_mult_76_FS_1_n37) );
  NOR2_X1 mul_ex_mult_76_FS_1_U42 ( .A1(mul_ex_mult_76_FS_1_n36), .A2(
        mul_ex_mult_76_FS_1_n37), .ZN(mul_ex_mult_76_FS_1_n38) );
  XOR2_X1 mul_ex_mult_76_FS_1_U41 ( .A(mul_ex_mult_76_FS_1_n35), .B(
        mul_ex_mult_76_FS_1_n38), .Z(mul_ex_N82) );
  NOR2_X1 mul_ex_mult_76_FS_1_U40 ( .A1(mul_ex_mult_76_n55), .A2(
        mul_ex_mult_76_n26), .ZN(mul_ex_mult_76_FS_1_n31) );
  NAND2_X1 mul_ex_mult_76_FS_1_U39 ( .A1(mul_ex_mult_76_n55), .A2(
        mul_ex_mult_76_n26), .ZN(mul_ex_mult_76_FS_1_n33) );
  NAND2_X1 mul_ex_mult_76_FS_1_U38 ( .A1(mul_ex_mult_76_FS_1_n7), .A2(
        mul_ex_mult_76_FS_1_n33), .ZN(mul_ex_mult_76_FS_1_n34) );
  AOI21_X1 mul_ex_mult_76_FS_1_U37 ( .B1(mul_ex_mult_76_FS_1_n8), .B2(
        mul_ex_mult_76_FS_1_n35), .A(mul_ex_mult_76_FS_1_n36), .ZN(
        mul_ex_mult_76_FS_1_n32) );
  XOR2_X1 mul_ex_mult_76_FS_1_U36 ( .A(mul_ex_mult_76_FS_1_n34), .B(
        mul_ex_mult_76_FS_1_n32), .Z(mul_ex_N83) );
  OAI21_X1 mul_ex_mult_76_FS_1_U35 ( .B1(mul_ex_mult_76_FS_1_n31), .B2(
        mul_ex_mult_76_FS_1_n32), .A(mul_ex_mult_76_FS_1_n33), .ZN(
        mul_ex_mult_76_FS_1_n27) );
  AND2_X1 mul_ex_mult_76_FS_1_U34 ( .A1(mul_ex_mult_76_n48), .A2(
        mul_ex_mult_76_n18), .ZN(mul_ex_mult_76_FS_1_n28) );
  NOR2_X1 mul_ex_mult_76_FS_1_U33 ( .A1(mul_ex_mult_76_n48), .A2(
        mul_ex_mult_76_n18), .ZN(mul_ex_mult_76_FS_1_n29) );
  NOR2_X1 mul_ex_mult_76_FS_1_U32 ( .A1(mul_ex_mult_76_FS_1_n28), .A2(
        mul_ex_mult_76_FS_1_n29), .ZN(mul_ex_mult_76_FS_1_n30) );
  XOR2_X1 mul_ex_mult_76_FS_1_U31 ( .A(mul_ex_mult_76_FS_1_n27), .B(
        mul_ex_mult_76_FS_1_n30), .Z(mul_ex_N84) );
  NOR2_X1 mul_ex_mult_76_FS_1_U30 ( .A1(mul_ex_mult_76_n54), .A2(
        mul_ex_mult_76_n25), .ZN(mul_ex_mult_76_FS_1_n23) );
  NAND2_X1 mul_ex_mult_76_FS_1_U29 ( .A1(mul_ex_mult_76_n54), .A2(
        mul_ex_mult_76_n25), .ZN(mul_ex_mult_76_FS_1_n25) );
  NAND2_X1 mul_ex_mult_76_FS_1_U28 ( .A1(mul_ex_mult_76_FS_1_n5), .A2(
        mul_ex_mult_76_FS_1_n25), .ZN(mul_ex_mult_76_FS_1_n26) );
  AOI21_X1 mul_ex_mult_76_FS_1_U27 ( .B1(mul_ex_mult_76_FS_1_n6), .B2(
        mul_ex_mult_76_FS_1_n27), .A(mul_ex_mult_76_FS_1_n28), .ZN(
        mul_ex_mult_76_FS_1_n24) );
  XOR2_X1 mul_ex_mult_76_FS_1_U26 ( .A(mul_ex_mult_76_FS_1_n26), .B(
        mul_ex_mult_76_FS_1_n24), .Z(mul_ex_N85) );
  OAI21_X1 mul_ex_mult_76_FS_1_U25 ( .B1(mul_ex_mult_76_FS_1_n23), .B2(
        mul_ex_mult_76_FS_1_n24), .A(mul_ex_mult_76_FS_1_n25), .ZN(
        mul_ex_mult_76_FS_1_n19) );
  AND2_X1 mul_ex_mult_76_FS_1_U24 ( .A1(mul_ex_mult_76_n47), .A2(
        mul_ex_mult_76_n17), .ZN(mul_ex_mult_76_FS_1_n20) );
  NOR2_X1 mul_ex_mult_76_FS_1_U23 ( .A1(mul_ex_mult_76_n47), .A2(
        mul_ex_mult_76_n17), .ZN(mul_ex_mult_76_FS_1_n21) );
  NOR2_X1 mul_ex_mult_76_FS_1_U22 ( .A1(mul_ex_mult_76_FS_1_n20), .A2(
        mul_ex_mult_76_FS_1_n21), .ZN(mul_ex_mult_76_FS_1_n22) );
  XOR2_X1 mul_ex_mult_76_FS_1_U21 ( .A(mul_ex_mult_76_FS_1_n19), .B(
        mul_ex_mult_76_FS_1_n22), .Z(mul_ex_N86) );
  AOI21_X1 mul_ex_mult_76_FS_1_U20 ( .B1(mul_ex_mult_76_FS_1_n19), .B2(
        mul_ex_mult_76_FS_1_n4), .A(mul_ex_mult_76_FS_1_n20), .ZN(
        mul_ex_mult_76_FS_1_n18) );
  XOR2_X1 mul_ex_mult_76_FS_1_U19 ( .A(mul_ex_mult_76_FS_1_n3), .B(
        mul_ex_mult_76_FS_1_n18), .Z(mul_ex_N87) );
  INV_X4 mul_ex_mult_76_FS_1_U18 ( .A(mul_ex_mult_76_FS_1_n70), .ZN(
        mul_ex_mult_76_FS_1_n17) );
  INV_X4 mul_ex_mult_76_FS_1_U17 ( .A(mul_ex_mult_76_FS_1_n68), .ZN(
        mul_ex_mult_76_FS_1_n16) );
  INV_X4 mul_ex_mult_76_FS_1_U16 ( .A(mul_ex_mult_76_FS_1_n63), .ZN(
        mul_ex_mult_76_FS_1_n15) );
  INV_X4 mul_ex_mult_76_FS_1_U15 ( .A(mul_ex_mult_76_FS_1_n61), .ZN(
        mul_ex_mult_76_FS_1_n14) );
  INV_X4 mul_ex_mult_76_FS_1_U14 ( .A(mul_ex_mult_76_FS_1_n55), .ZN(
        mul_ex_mult_76_FS_1_n13) );
  INV_X4 mul_ex_mult_76_FS_1_U13 ( .A(mul_ex_mult_76_FS_1_n53), .ZN(
        mul_ex_mult_76_FS_1_n12) );
  INV_X4 mul_ex_mult_76_FS_1_U12 ( .A(mul_ex_mult_76_FS_1_n47), .ZN(
        mul_ex_mult_76_FS_1_n11) );
  INV_X4 mul_ex_mult_76_FS_1_U11 ( .A(mul_ex_mult_76_FS_1_n45), .ZN(
        mul_ex_mult_76_FS_1_n10) );
  INV_X4 mul_ex_mult_76_FS_1_U10 ( .A(mul_ex_mult_76_FS_1_n39), .ZN(
        mul_ex_mult_76_FS_1_n9) );
  INV_X4 mul_ex_mult_76_FS_1_U9 ( .A(mul_ex_mult_76_FS_1_n37), .ZN(
        mul_ex_mult_76_FS_1_n8) );
  INV_X4 mul_ex_mult_76_FS_1_U8 ( .A(mul_ex_mult_76_FS_1_n31), .ZN(
        mul_ex_mult_76_FS_1_n7) );
  INV_X4 mul_ex_mult_76_FS_1_U7 ( .A(mul_ex_mult_76_FS_1_n29), .ZN(
        mul_ex_mult_76_FS_1_n6) );
  INV_X4 mul_ex_mult_76_FS_1_U6 ( .A(mul_ex_mult_76_FS_1_n23), .ZN(
        mul_ex_mult_76_FS_1_n5) );
  INV_X4 mul_ex_mult_76_FS_1_U5 ( .A(mul_ex_mult_76_FS_1_n21), .ZN(
        mul_ex_mult_76_FS_1_n4) );
  INV_X4 mul_ex_mult_76_FS_1_U4 ( .A(mul_ex_mult_76_n62), .ZN(
        mul_ex_mult_76_FS_1_n3) );
  AND2_X4 mul_ex_mult_76_FS_1_U3 ( .A1(mul_ex_mult_76_FS_1_n1), .A2(
        mul_ex_mult_76_FS_1_n70), .ZN(mul_ex_N73) );
  OR2_X4 mul_ex_mult_76_FS_1_U2 ( .A1(mul_ex_mult_76_n60), .A2(
        mul_ex_mult_76_n24), .ZN(mul_ex_mult_76_FS_1_n1) );
  NOR2_X1 mul_ex_mult_86_U350 ( .A1(mul_ex_mult_86_n94), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_N122) );
  NOR2_X1 mul_ex_mult_86_U349 ( .A1(mul_ex_mult_86_n84), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_mult_86_ab_0__10_) );
  NOR2_X1 mul_ex_mult_86_U348 ( .A1(mul_ex_mult_86_n83), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_mult_86_ab_0__11_) );
  NOR2_X1 mul_ex_mult_86_U347 ( .A1(mul_ex_mult_86_n82), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_mult_86_ab_0__12_) );
  NOR2_X1 mul_ex_mult_86_U346 ( .A1(mul_ex_mult_86_n81), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_mult_86_ab_0__13_) );
  NOR2_X1 mul_ex_mult_86_U345 ( .A1(mul_ex_mult_86_n80), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_mult_86_ab_0__14_) );
  NOR2_X1 mul_ex_mult_86_U344 ( .A1(mul_ex_mult_86_n79), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_mult_86_ab_0__15_) );
  NOR2_X1 mul_ex_mult_86_U343 ( .A1(mul_ex_mult_86_n93), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_mult_86_ab_0__1_) );
  NOR2_X1 mul_ex_mult_86_U342 ( .A1(mul_ex_mult_86_n92), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_mult_86_ab_0__2_) );
  NOR2_X1 mul_ex_mult_86_U341 ( .A1(mul_ex_mult_86_n91), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_mult_86_ab_0__3_) );
  NOR2_X1 mul_ex_mult_86_U340 ( .A1(mul_ex_mult_86_n90), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_mult_86_ab_0__4_) );
  NOR2_X1 mul_ex_mult_86_U339 ( .A1(mul_ex_mult_86_n89), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_mult_86_ab_0__5_) );
  NOR2_X1 mul_ex_mult_86_U338 ( .A1(mul_ex_mult_86_n88), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_mult_86_ab_0__6_) );
  NOR2_X1 mul_ex_mult_86_U337 ( .A1(mul_ex_mult_86_n87), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_mult_86_ab_0__7_) );
  NOR2_X1 mul_ex_mult_86_U336 ( .A1(mul_ex_mult_86_n86), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_mult_86_ab_0__8_) );
  NOR2_X1 mul_ex_mult_86_U335 ( .A1(mul_ex_mult_86_n85), .A2(
        mul_ex_mult_86_n78), .ZN(mul_ex_mult_86_ab_0__9_) );
  NOR2_X1 mul_ex_mult_86_U334 ( .A1(mul_ex_mult_86_n94), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__0_) );
  NOR2_X1 mul_ex_mult_86_U333 ( .A1(mul_ex_mult_86_n84), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__10_) );
  NOR2_X1 mul_ex_mult_86_U332 ( .A1(mul_ex_mult_86_n83), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__11_) );
  NOR2_X1 mul_ex_mult_86_U331 ( .A1(mul_ex_mult_86_n82), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__12_) );
  NOR2_X1 mul_ex_mult_86_U330 ( .A1(mul_ex_mult_86_n81), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__13_) );
  NOR2_X1 mul_ex_mult_86_U329 ( .A1(mul_ex_mult_86_n80), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__14_) );
  NOR2_X1 mul_ex_mult_86_U328 ( .A1(mul_ex_mult_86_n79), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__15_) );
  NOR2_X1 mul_ex_mult_86_U327 ( .A1(mul_ex_mult_86_n93), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__1_) );
  NOR2_X1 mul_ex_mult_86_U326 ( .A1(mul_ex_mult_86_n92), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__2_) );
  NOR2_X1 mul_ex_mult_86_U325 ( .A1(mul_ex_mult_86_n91), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__3_) );
  NOR2_X1 mul_ex_mult_86_U324 ( .A1(mul_ex_mult_86_n90), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__4_) );
  NOR2_X1 mul_ex_mult_86_U323 ( .A1(mul_ex_mult_86_n89), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__5_) );
  NOR2_X1 mul_ex_mult_86_U322 ( .A1(mul_ex_mult_86_n88), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__6_) );
  NOR2_X1 mul_ex_mult_86_U321 ( .A1(mul_ex_mult_86_n87), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__7_) );
  NOR2_X1 mul_ex_mult_86_U320 ( .A1(mul_ex_mult_86_n86), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__8_) );
  NOR2_X1 mul_ex_mult_86_U319 ( .A1(mul_ex_mult_86_n85), .A2(
        mul_ex_mult_86_n68), .ZN(mul_ex_mult_86_ab_10__9_) );
  NOR2_X1 mul_ex_mult_86_U318 ( .A1(mul_ex_mult_86_n94), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__0_) );
  NOR2_X1 mul_ex_mult_86_U317 ( .A1(mul_ex_mult_86_n84), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__10_) );
  NOR2_X1 mul_ex_mult_86_U316 ( .A1(mul_ex_mult_86_n83), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__11_) );
  NOR2_X1 mul_ex_mult_86_U315 ( .A1(mul_ex_mult_86_n82), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__12_) );
  NOR2_X1 mul_ex_mult_86_U314 ( .A1(mul_ex_mult_86_n81), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__13_) );
  NOR2_X1 mul_ex_mult_86_U313 ( .A1(mul_ex_mult_86_n80), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__14_) );
  NOR2_X1 mul_ex_mult_86_U312 ( .A1(mul_ex_mult_86_n79), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__15_) );
  NOR2_X1 mul_ex_mult_86_U311 ( .A1(mul_ex_mult_86_n93), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__1_) );
  NOR2_X1 mul_ex_mult_86_U310 ( .A1(mul_ex_mult_86_n92), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__2_) );
  NOR2_X1 mul_ex_mult_86_U309 ( .A1(mul_ex_mult_86_n91), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__3_) );
  NOR2_X1 mul_ex_mult_86_U308 ( .A1(mul_ex_mult_86_n90), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__4_) );
  NOR2_X1 mul_ex_mult_86_U307 ( .A1(mul_ex_mult_86_n89), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__5_) );
  NOR2_X1 mul_ex_mult_86_U306 ( .A1(mul_ex_mult_86_n88), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__6_) );
  NOR2_X1 mul_ex_mult_86_U305 ( .A1(mul_ex_mult_86_n87), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__7_) );
  NOR2_X1 mul_ex_mult_86_U304 ( .A1(mul_ex_mult_86_n86), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__8_) );
  NOR2_X1 mul_ex_mult_86_U303 ( .A1(mul_ex_mult_86_n85), .A2(
        mul_ex_mult_86_n67), .ZN(mul_ex_mult_86_ab_11__9_) );
  NOR2_X1 mul_ex_mult_86_U302 ( .A1(mul_ex_mult_86_n94), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__0_) );
  NOR2_X1 mul_ex_mult_86_U301 ( .A1(mul_ex_mult_86_n84), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__10_) );
  NOR2_X1 mul_ex_mult_86_U300 ( .A1(mul_ex_mult_86_n83), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__11_) );
  NOR2_X1 mul_ex_mult_86_U299 ( .A1(mul_ex_mult_86_n82), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__12_) );
  NOR2_X1 mul_ex_mult_86_U298 ( .A1(mul_ex_mult_86_n81), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__13_) );
  NOR2_X1 mul_ex_mult_86_U297 ( .A1(mul_ex_mult_86_n80), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__14_) );
  NOR2_X1 mul_ex_mult_86_U296 ( .A1(mul_ex_mult_86_n79), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__15_) );
  NOR2_X1 mul_ex_mult_86_U295 ( .A1(mul_ex_mult_86_n93), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__1_) );
  NOR2_X1 mul_ex_mult_86_U294 ( .A1(mul_ex_mult_86_n92), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__2_) );
  NOR2_X1 mul_ex_mult_86_U293 ( .A1(mul_ex_mult_86_n91), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__3_) );
  NOR2_X1 mul_ex_mult_86_U292 ( .A1(mul_ex_mult_86_n90), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__4_) );
  NOR2_X1 mul_ex_mult_86_U291 ( .A1(mul_ex_mult_86_n89), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__5_) );
  NOR2_X1 mul_ex_mult_86_U290 ( .A1(mul_ex_mult_86_n88), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__6_) );
  NOR2_X1 mul_ex_mult_86_U289 ( .A1(mul_ex_mult_86_n87), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__7_) );
  NOR2_X1 mul_ex_mult_86_U288 ( .A1(mul_ex_mult_86_n86), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__8_) );
  NOR2_X1 mul_ex_mult_86_U287 ( .A1(mul_ex_mult_86_n85), .A2(
        mul_ex_mult_86_n66), .ZN(mul_ex_mult_86_ab_12__9_) );
  NOR2_X1 mul_ex_mult_86_U286 ( .A1(mul_ex_mult_86_n94), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__0_) );
  NOR2_X1 mul_ex_mult_86_U285 ( .A1(mul_ex_mult_86_n84), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__10_) );
  NOR2_X1 mul_ex_mult_86_U284 ( .A1(mul_ex_mult_86_n83), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__11_) );
  NOR2_X1 mul_ex_mult_86_U283 ( .A1(mul_ex_mult_86_n82), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__12_) );
  NOR2_X1 mul_ex_mult_86_U282 ( .A1(mul_ex_mult_86_n81), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__13_) );
  NOR2_X1 mul_ex_mult_86_U281 ( .A1(mul_ex_mult_86_n80), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__14_) );
  NOR2_X1 mul_ex_mult_86_U280 ( .A1(mul_ex_mult_86_n79), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__15_) );
  NOR2_X1 mul_ex_mult_86_U279 ( .A1(mul_ex_mult_86_n93), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__1_) );
  NOR2_X1 mul_ex_mult_86_U278 ( .A1(mul_ex_mult_86_n92), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__2_) );
  NOR2_X1 mul_ex_mult_86_U277 ( .A1(mul_ex_mult_86_n91), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__3_) );
  NOR2_X1 mul_ex_mult_86_U276 ( .A1(mul_ex_mult_86_n90), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__4_) );
  NOR2_X1 mul_ex_mult_86_U275 ( .A1(mul_ex_mult_86_n89), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__5_) );
  NOR2_X1 mul_ex_mult_86_U274 ( .A1(mul_ex_mult_86_n88), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__6_) );
  NOR2_X1 mul_ex_mult_86_U273 ( .A1(mul_ex_mult_86_n87), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__7_) );
  NOR2_X1 mul_ex_mult_86_U272 ( .A1(mul_ex_mult_86_n86), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__8_) );
  NOR2_X1 mul_ex_mult_86_U271 ( .A1(mul_ex_mult_86_n85), .A2(
        mul_ex_mult_86_n65), .ZN(mul_ex_mult_86_ab_13__9_) );
  NOR2_X1 mul_ex_mult_86_U270 ( .A1(mul_ex_mult_86_n94), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__0_) );
  NOR2_X1 mul_ex_mult_86_U269 ( .A1(mul_ex_mult_86_n84), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__10_) );
  NOR2_X1 mul_ex_mult_86_U268 ( .A1(mul_ex_mult_86_n83), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__11_) );
  NOR2_X1 mul_ex_mult_86_U267 ( .A1(mul_ex_mult_86_n82), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__12_) );
  NOR2_X1 mul_ex_mult_86_U266 ( .A1(mul_ex_mult_86_n81), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__13_) );
  NOR2_X1 mul_ex_mult_86_U265 ( .A1(mul_ex_mult_86_n80), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__14_) );
  NOR2_X1 mul_ex_mult_86_U264 ( .A1(mul_ex_mult_86_n79), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__15_) );
  NOR2_X1 mul_ex_mult_86_U263 ( .A1(mul_ex_mult_86_n93), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__1_) );
  NOR2_X1 mul_ex_mult_86_U262 ( .A1(mul_ex_mult_86_n92), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__2_) );
  NOR2_X1 mul_ex_mult_86_U261 ( .A1(mul_ex_mult_86_n91), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__3_) );
  NOR2_X1 mul_ex_mult_86_U260 ( .A1(mul_ex_mult_86_n90), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__4_) );
  NOR2_X1 mul_ex_mult_86_U259 ( .A1(mul_ex_mult_86_n89), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__5_) );
  NOR2_X1 mul_ex_mult_86_U258 ( .A1(mul_ex_mult_86_n88), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__6_) );
  NOR2_X1 mul_ex_mult_86_U257 ( .A1(mul_ex_mult_86_n87), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__7_) );
  NOR2_X1 mul_ex_mult_86_U256 ( .A1(mul_ex_mult_86_n86), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__8_) );
  NOR2_X1 mul_ex_mult_86_U255 ( .A1(mul_ex_mult_86_n85), .A2(
        mul_ex_mult_86_n64), .ZN(mul_ex_mult_86_ab_14__9_) );
  NOR2_X1 mul_ex_mult_86_U254 ( .A1(mul_ex_mult_86_n94), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__0_) );
  NOR2_X1 mul_ex_mult_86_U253 ( .A1(mul_ex_mult_86_n84), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__10_) );
  NOR2_X1 mul_ex_mult_86_U252 ( .A1(mul_ex_mult_86_n83), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__11_) );
  NOR2_X1 mul_ex_mult_86_U251 ( .A1(mul_ex_mult_86_n82), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__12_) );
  NOR2_X1 mul_ex_mult_86_U250 ( .A1(mul_ex_mult_86_n81), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__13_) );
  NOR2_X1 mul_ex_mult_86_U249 ( .A1(mul_ex_mult_86_n80), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__14_) );
  NOR2_X1 mul_ex_mult_86_U248 ( .A1(mul_ex_mult_86_n79), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__15_) );
  NOR2_X1 mul_ex_mult_86_U247 ( .A1(mul_ex_mult_86_n93), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__1_) );
  NOR2_X1 mul_ex_mult_86_U246 ( .A1(mul_ex_mult_86_n92), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__2_) );
  NOR2_X1 mul_ex_mult_86_U245 ( .A1(mul_ex_mult_86_n91), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__3_) );
  NOR2_X1 mul_ex_mult_86_U244 ( .A1(mul_ex_mult_86_n90), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__4_) );
  NOR2_X1 mul_ex_mult_86_U243 ( .A1(mul_ex_mult_86_n89), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__5_) );
  NOR2_X1 mul_ex_mult_86_U242 ( .A1(mul_ex_mult_86_n88), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__6_) );
  NOR2_X1 mul_ex_mult_86_U241 ( .A1(mul_ex_mult_86_n87), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__7_) );
  NOR2_X1 mul_ex_mult_86_U240 ( .A1(mul_ex_mult_86_n86), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__8_) );
  NOR2_X1 mul_ex_mult_86_U239 ( .A1(mul_ex_mult_86_n85), .A2(
        mul_ex_mult_86_n63), .ZN(mul_ex_mult_86_ab_15__9_) );
  NOR2_X1 mul_ex_mult_86_U238 ( .A1(mul_ex_mult_86_n94), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__0_) );
  NOR2_X1 mul_ex_mult_86_U237 ( .A1(mul_ex_mult_86_n84), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__10_) );
  NOR2_X1 mul_ex_mult_86_U236 ( .A1(mul_ex_mult_86_n83), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__11_) );
  NOR2_X1 mul_ex_mult_86_U235 ( .A1(mul_ex_mult_86_n82), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__12_) );
  NOR2_X1 mul_ex_mult_86_U234 ( .A1(mul_ex_mult_86_n81), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__13_) );
  NOR2_X1 mul_ex_mult_86_U233 ( .A1(mul_ex_mult_86_n80), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__14_) );
  NOR2_X1 mul_ex_mult_86_U232 ( .A1(mul_ex_mult_86_n79), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__15_) );
  NOR2_X1 mul_ex_mult_86_U231 ( .A1(mul_ex_mult_86_n93), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__1_) );
  NOR2_X1 mul_ex_mult_86_U230 ( .A1(mul_ex_mult_86_n92), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__2_) );
  NOR2_X1 mul_ex_mult_86_U229 ( .A1(mul_ex_mult_86_n91), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__3_) );
  NOR2_X1 mul_ex_mult_86_U228 ( .A1(mul_ex_mult_86_n90), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__4_) );
  NOR2_X1 mul_ex_mult_86_U227 ( .A1(mul_ex_mult_86_n89), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__5_) );
  NOR2_X1 mul_ex_mult_86_U226 ( .A1(mul_ex_mult_86_n88), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__6_) );
  NOR2_X1 mul_ex_mult_86_U225 ( .A1(mul_ex_mult_86_n87), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__7_) );
  NOR2_X1 mul_ex_mult_86_U224 ( .A1(mul_ex_mult_86_n86), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__8_) );
  NOR2_X1 mul_ex_mult_86_U223 ( .A1(mul_ex_mult_86_n85), .A2(
        mul_ex_mult_86_n77), .ZN(mul_ex_mult_86_ab_1__9_) );
  NOR2_X1 mul_ex_mult_86_U222 ( .A1(mul_ex_mult_86_n94), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__0_) );
  NOR2_X1 mul_ex_mult_86_U221 ( .A1(mul_ex_mult_86_n84), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__10_) );
  NOR2_X1 mul_ex_mult_86_U220 ( .A1(mul_ex_mult_86_n83), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__11_) );
  NOR2_X1 mul_ex_mult_86_U219 ( .A1(mul_ex_mult_86_n82), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__12_) );
  NOR2_X1 mul_ex_mult_86_U218 ( .A1(mul_ex_mult_86_n81), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__13_) );
  NOR2_X1 mul_ex_mult_86_U217 ( .A1(mul_ex_mult_86_n80), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__14_) );
  NOR2_X1 mul_ex_mult_86_U216 ( .A1(mul_ex_mult_86_n79), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__15_) );
  NOR2_X1 mul_ex_mult_86_U215 ( .A1(mul_ex_mult_86_n93), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__1_) );
  NOR2_X1 mul_ex_mult_86_U214 ( .A1(mul_ex_mult_86_n92), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__2_) );
  NOR2_X1 mul_ex_mult_86_U213 ( .A1(mul_ex_mult_86_n91), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__3_) );
  NOR2_X1 mul_ex_mult_86_U212 ( .A1(mul_ex_mult_86_n90), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__4_) );
  NOR2_X1 mul_ex_mult_86_U211 ( .A1(mul_ex_mult_86_n89), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__5_) );
  NOR2_X1 mul_ex_mult_86_U210 ( .A1(mul_ex_mult_86_n88), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__6_) );
  NOR2_X1 mul_ex_mult_86_U209 ( .A1(mul_ex_mult_86_n87), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__7_) );
  NOR2_X1 mul_ex_mult_86_U208 ( .A1(mul_ex_mult_86_n86), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__8_) );
  NOR2_X1 mul_ex_mult_86_U207 ( .A1(mul_ex_mult_86_n85), .A2(
        mul_ex_mult_86_n76), .ZN(mul_ex_mult_86_ab_2__9_) );
  NOR2_X1 mul_ex_mult_86_U206 ( .A1(mul_ex_mult_86_n94), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__0_) );
  NOR2_X1 mul_ex_mult_86_U205 ( .A1(mul_ex_mult_86_n84), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__10_) );
  NOR2_X1 mul_ex_mult_86_U204 ( .A1(mul_ex_mult_86_n83), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__11_) );
  NOR2_X1 mul_ex_mult_86_U203 ( .A1(mul_ex_mult_86_n82), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__12_) );
  NOR2_X1 mul_ex_mult_86_U202 ( .A1(mul_ex_mult_86_n81), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__13_) );
  NOR2_X1 mul_ex_mult_86_U201 ( .A1(mul_ex_mult_86_n80), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__14_) );
  NOR2_X1 mul_ex_mult_86_U200 ( .A1(mul_ex_mult_86_n79), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__15_) );
  NOR2_X1 mul_ex_mult_86_U199 ( .A1(mul_ex_mult_86_n93), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__1_) );
  NOR2_X1 mul_ex_mult_86_U198 ( .A1(mul_ex_mult_86_n92), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__2_) );
  NOR2_X1 mul_ex_mult_86_U197 ( .A1(mul_ex_mult_86_n91), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__3_) );
  NOR2_X1 mul_ex_mult_86_U196 ( .A1(mul_ex_mult_86_n90), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__4_) );
  NOR2_X1 mul_ex_mult_86_U195 ( .A1(mul_ex_mult_86_n89), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__5_) );
  NOR2_X1 mul_ex_mult_86_U194 ( .A1(mul_ex_mult_86_n88), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__6_) );
  NOR2_X1 mul_ex_mult_86_U193 ( .A1(mul_ex_mult_86_n87), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__7_) );
  NOR2_X1 mul_ex_mult_86_U192 ( .A1(mul_ex_mult_86_n86), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__8_) );
  NOR2_X1 mul_ex_mult_86_U191 ( .A1(mul_ex_mult_86_n85), .A2(
        mul_ex_mult_86_n75), .ZN(mul_ex_mult_86_ab_3__9_) );
  NOR2_X1 mul_ex_mult_86_U190 ( .A1(mul_ex_mult_86_n94), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__0_) );
  NOR2_X1 mul_ex_mult_86_U189 ( .A1(mul_ex_mult_86_n84), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__10_) );
  NOR2_X1 mul_ex_mult_86_U188 ( .A1(mul_ex_mult_86_n83), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__11_) );
  NOR2_X1 mul_ex_mult_86_U187 ( .A1(mul_ex_mult_86_n82), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__12_) );
  NOR2_X1 mul_ex_mult_86_U186 ( .A1(mul_ex_mult_86_n81), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__13_) );
  NOR2_X1 mul_ex_mult_86_U185 ( .A1(mul_ex_mult_86_n80), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__14_) );
  NOR2_X1 mul_ex_mult_86_U184 ( .A1(mul_ex_mult_86_n79), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__15_) );
  NOR2_X1 mul_ex_mult_86_U183 ( .A1(mul_ex_mult_86_n93), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__1_) );
  NOR2_X1 mul_ex_mult_86_U182 ( .A1(mul_ex_mult_86_n92), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__2_) );
  NOR2_X1 mul_ex_mult_86_U181 ( .A1(mul_ex_mult_86_n91), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__3_) );
  NOR2_X1 mul_ex_mult_86_U180 ( .A1(mul_ex_mult_86_n90), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__4_) );
  NOR2_X1 mul_ex_mult_86_U179 ( .A1(mul_ex_mult_86_n89), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__5_) );
  NOR2_X1 mul_ex_mult_86_U178 ( .A1(mul_ex_mult_86_n88), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__6_) );
  NOR2_X1 mul_ex_mult_86_U177 ( .A1(mul_ex_mult_86_n87), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__7_) );
  NOR2_X1 mul_ex_mult_86_U176 ( .A1(mul_ex_mult_86_n86), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__8_) );
  NOR2_X1 mul_ex_mult_86_U175 ( .A1(mul_ex_mult_86_n85), .A2(
        mul_ex_mult_86_n74), .ZN(mul_ex_mult_86_ab_4__9_) );
  NOR2_X1 mul_ex_mult_86_U174 ( .A1(mul_ex_mult_86_n94), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__0_) );
  NOR2_X1 mul_ex_mult_86_U173 ( .A1(mul_ex_mult_86_n84), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__10_) );
  NOR2_X1 mul_ex_mult_86_U172 ( .A1(mul_ex_mult_86_n83), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__11_) );
  NOR2_X1 mul_ex_mult_86_U171 ( .A1(mul_ex_mult_86_n82), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__12_) );
  NOR2_X1 mul_ex_mult_86_U170 ( .A1(mul_ex_mult_86_n81), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__13_) );
  NOR2_X1 mul_ex_mult_86_U169 ( .A1(mul_ex_mult_86_n80), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__14_) );
  NOR2_X1 mul_ex_mult_86_U168 ( .A1(mul_ex_mult_86_n79), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__15_) );
  NOR2_X1 mul_ex_mult_86_U167 ( .A1(mul_ex_mult_86_n93), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__1_) );
  NOR2_X1 mul_ex_mult_86_U166 ( .A1(mul_ex_mult_86_n92), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__2_) );
  NOR2_X1 mul_ex_mult_86_U165 ( .A1(mul_ex_mult_86_n91), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__3_) );
  NOR2_X1 mul_ex_mult_86_U164 ( .A1(mul_ex_mult_86_n90), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__4_) );
  NOR2_X1 mul_ex_mult_86_U163 ( .A1(mul_ex_mult_86_n89), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__5_) );
  NOR2_X1 mul_ex_mult_86_U162 ( .A1(mul_ex_mult_86_n88), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__6_) );
  NOR2_X1 mul_ex_mult_86_U161 ( .A1(mul_ex_mult_86_n87), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__7_) );
  NOR2_X1 mul_ex_mult_86_U160 ( .A1(mul_ex_mult_86_n86), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__8_) );
  NOR2_X1 mul_ex_mult_86_U159 ( .A1(mul_ex_mult_86_n85), .A2(
        mul_ex_mult_86_n73), .ZN(mul_ex_mult_86_ab_5__9_) );
  NOR2_X1 mul_ex_mult_86_U158 ( .A1(mul_ex_mult_86_n94), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__0_) );
  NOR2_X1 mul_ex_mult_86_U157 ( .A1(mul_ex_mult_86_n84), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__10_) );
  NOR2_X1 mul_ex_mult_86_U156 ( .A1(mul_ex_mult_86_n83), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__11_) );
  NOR2_X1 mul_ex_mult_86_U155 ( .A1(mul_ex_mult_86_n82), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__12_) );
  NOR2_X1 mul_ex_mult_86_U154 ( .A1(mul_ex_mult_86_n81), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__13_) );
  NOR2_X1 mul_ex_mult_86_U153 ( .A1(mul_ex_mult_86_n80), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__14_) );
  NOR2_X1 mul_ex_mult_86_U152 ( .A1(mul_ex_mult_86_n79), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__15_) );
  NOR2_X1 mul_ex_mult_86_U151 ( .A1(mul_ex_mult_86_n93), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__1_) );
  NOR2_X1 mul_ex_mult_86_U150 ( .A1(mul_ex_mult_86_n92), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__2_) );
  NOR2_X1 mul_ex_mult_86_U149 ( .A1(mul_ex_mult_86_n91), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__3_) );
  NOR2_X1 mul_ex_mult_86_U148 ( .A1(mul_ex_mult_86_n90), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__4_) );
  NOR2_X1 mul_ex_mult_86_U147 ( .A1(mul_ex_mult_86_n89), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__5_) );
  NOR2_X1 mul_ex_mult_86_U146 ( .A1(mul_ex_mult_86_n88), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__6_) );
  NOR2_X1 mul_ex_mult_86_U145 ( .A1(mul_ex_mult_86_n87), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__7_) );
  NOR2_X1 mul_ex_mult_86_U144 ( .A1(mul_ex_mult_86_n86), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__8_) );
  NOR2_X1 mul_ex_mult_86_U143 ( .A1(mul_ex_mult_86_n85), .A2(
        mul_ex_mult_86_n72), .ZN(mul_ex_mult_86_ab_6__9_) );
  NOR2_X1 mul_ex_mult_86_U142 ( .A1(mul_ex_mult_86_n94), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__0_) );
  NOR2_X1 mul_ex_mult_86_U141 ( .A1(mul_ex_mult_86_n84), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__10_) );
  NOR2_X1 mul_ex_mult_86_U140 ( .A1(mul_ex_mult_86_n83), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__11_) );
  NOR2_X1 mul_ex_mult_86_U139 ( .A1(mul_ex_mult_86_n82), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__12_) );
  NOR2_X1 mul_ex_mult_86_U138 ( .A1(mul_ex_mult_86_n81), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__13_) );
  NOR2_X1 mul_ex_mult_86_U137 ( .A1(mul_ex_mult_86_n80), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__14_) );
  NOR2_X1 mul_ex_mult_86_U136 ( .A1(mul_ex_mult_86_n79), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__15_) );
  NOR2_X1 mul_ex_mult_86_U135 ( .A1(mul_ex_mult_86_n93), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__1_) );
  NOR2_X1 mul_ex_mult_86_U134 ( .A1(mul_ex_mult_86_n92), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__2_) );
  NOR2_X1 mul_ex_mult_86_U133 ( .A1(mul_ex_mult_86_n91), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__3_) );
  NOR2_X1 mul_ex_mult_86_U132 ( .A1(mul_ex_mult_86_n90), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__4_) );
  NOR2_X1 mul_ex_mult_86_U131 ( .A1(mul_ex_mult_86_n89), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__5_) );
  NOR2_X1 mul_ex_mult_86_U130 ( .A1(mul_ex_mult_86_n88), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__6_) );
  NOR2_X1 mul_ex_mult_86_U129 ( .A1(mul_ex_mult_86_n87), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__7_) );
  NOR2_X1 mul_ex_mult_86_U128 ( .A1(mul_ex_mult_86_n86), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__8_) );
  NOR2_X1 mul_ex_mult_86_U127 ( .A1(mul_ex_mult_86_n85), .A2(
        mul_ex_mult_86_n71), .ZN(mul_ex_mult_86_ab_7__9_) );
  NOR2_X1 mul_ex_mult_86_U126 ( .A1(mul_ex_mult_86_n94), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__0_) );
  NOR2_X1 mul_ex_mult_86_U125 ( .A1(mul_ex_mult_86_n84), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__10_) );
  NOR2_X1 mul_ex_mult_86_U124 ( .A1(mul_ex_mult_86_n83), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__11_) );
  NOR2_X1 mul_ex_mult_86_U123 ( .A1(mul_ex_mult_86_n82), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__12_) );
  NOR2_X1 mul_ex_mult_86_U122 ( .A1(mul_ex_mult_86_n81), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__13_) );
  NOR2_X1 mul_ex_mult_86_U121 ( .A1(mul_ex_mult_86_n80), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__14_) );
  NOR2_X1 mul_ex_mult_86_U120 ( .A1(mul_ex_mult_86_n79), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__15_) );
  NOR2_X1 mul_ex_mult_86_U119 ( .A1(mul_ex_mult_86_n93), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__1_) );
  NOR2_X1 mul_ex_mult_86_U118 ( .A1(mul_ex_mult_86_n92), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__2_) );
  NOR2_X1 mul_ex_mult_86_U117 ( .A1(mul_ex_mult_86_n91), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__3_) );
  NOR2_X1 mul_ex_mult_86_U116 ( .A1(mul_ex_mult_86_n90), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__4_) );
  NOR2_X1 mul_ex_mult_86_U115 ( .A1(mul_ex_mult_86_n89), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__5_) );
  NOR2_X1 mul_ex_mult_86_U114 ( .A1(mul_ex_mult_86_n88), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__6_) );
  NOR2_X1 mul_ex_mult_86_U113 ( .A1(mul_ex_mult_86_n87), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__7_) );
  NOR2_X1 mul_ex_mult_86_U112 ( .A1(mul_ex_mult_86_n86), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__8_) );
  NOR2_X1 mul_ex_mult_86_U111 ( .A1(mul_ex_mult_86_n85), .A2(
        mul_ex_mult_86_n70), .ZN(mul_ex_mult_86_ab_8__9_) );
  NOR2_X1 mul_ex_mult_86_U110 ( .A1(mul_ex_mult_86_n69), .A2(
        mul_ex_mult_86_n94), .ZN(mul_ex_mult_86_ab_9__0_) );
  NOR2_X1 mul_ex_mult_86_U109 ( .A1(mul_ex_mult_86_n69), .A2(
        mul_ex_mult_86_n84), .ZN(mul_ex_mult_86_ab_9__10_) );
  NOR2_X1 mul_ex_mult_86_U108 ( .A1(mul_ex_mult_86_n69), .A2(
        mul_ex_mult_86_n83), .ZN(mul_ex_mult_86_ab_9__11_) );
  NOR2_X1 mul_ex_mult_86_U107 ( .A1(mul_ex_mult_86_n69), .A2(
        mul_ex_mult_86_n82), .ZN(mul_ex_mult_86_ab_9__12_) );
  NOR2_X1 mul_ex_mult_86_U106 ( .A1(mul_ex_mult_86_n69), .A2(
        mul_ex_mult_86_n81), .ZN(mul_ex_mult_86_ab_9__13_) );
  NOR2_X1 mul_ex_mult_86_U105 ( .A1(mul_ex_mult_86_n69), .A2(
        mul_ex_mult_86_n80), .ZN(mul_ex_mult_86_ab_9__14_) );
  NOR2_X1 mul_ex_mult_86_U104 ( .A1(mul_ex_mult_86_n69), .A2(
        mul_ex_mult_86_n79), .ZN(mul_ex_mult_86_ab_9__15_) );
  NOR2_X1 mul_ex_mult_86_U103 ( .A1(mul_ex_mult_86_n69), .A2(
        mul_ex_mult_86_n93), .ZN(mul_ex_mult_86_ab_9__1_) );
  NOR2_X1 mul_ex_mult_86_U102 ( .A1(mul_ex_mult_86_n69), .A2(
        mul_ex_mult_86_n92), .ZN(mul_ex_mult_86_ab_9__2_) );
  NOR2_X1 mul_ex_mult_86_U101 ( .A1(mul_ex_mult_86_n69), .A2(
        mul_ex_mult_86_n91), .ZN(mul_ex_mult_86_ab_9__3_) );
  NOR2_X1 mul_ex_mult_86_U100 ( .A1(mul_ex_mult_86_n69), .A2(
        mul_ex_mult_86_n90), .ZN(mul_ex_mult_86_ab_9__4_) );
  NOR2_X1 mul_ex_mult_86_U99 ( .A1(mul_ex_mult_86_n69), .A2(mul_ex_mult_86_n89), .ZN(mul_ex_mult_86_ab_9__5_) );
  NOR2_X1 mul_ex_mult_86_U98 ( .A1(mul_ex_mult_86_n69), .A2(mul_ex_mult_86_n88), .ZN(mul_ex_mult_86_ab_9__6_) );
  NOR2_X1 mul_ex_mult_86_U97 ( .A1(mul_ex_mult_86_n69), .A2(mul_ex_mult_86_n87), .ZN(mul_ex_mult_86_ab_9__7_) );
  NOR2_X1 mul_ex_mult_86_U96 ( .A1(mul_ex_mult_86_n69), .A2(mul_ex_mult_86_n86), .ZN(mul_ex_mult_86_ab_9__8_) );
  NOR2_X1 mul_ex_mult_86_U95 ( .A1(mul_ex_mult_86_n69), .A2(mul_ex_mult_86_n85), .ZN(mul_ex_mult_86_ab_9__9_) );
  INV_X4 mul_ex_mult_86_U93 ( .A(f1_in[16]), .ZN(mul_ex_mult_86_n63) );
  INV_X4 mul_ex_mult_86_U92 ( .A(f1_in[17]), .ZN(mul_ex_mult_86_n64) );
  INV_X4 mul_ex_mult_86_U91 ( .A(f1_in[18]), .ZN(mul_ex_mult_86_n65) );
  INV_X4 mul_ex_mult_86_U90 ( .A(f1_in[19]), .ZN(mul_ex_mult_86_n66) );
  INV_X4 mul_ex_mult_86_U89 ( .A(f1_in[20]), .ZN(mul_ex_mult_86_n67) );
  INV_X4 mul_ex_mult_86_U88 ( .A(f1_in[21]), .ZN(mul_ex_mult_86_n68) );
  INV_X4 mul_ex_mult_86_U87 ( .A(f1_in[29]), .ZN(mul_ex_mult_86_n76) );
  INV_X4 mul_ex_mult_86_U86 ( .A(f1_in[23]), .ZN(mul_ex_mult_86_n70) );
  INV_X4 mul_ex_mult_86_U85 ( .A(f1_in[24]), .ZN(mul_ex_mult_86_n71) );
  INV_X4 mul_ex_mult_86_U84 ( .A(f1_in[25]), .ZN(mul_ex_mult_86_n72) );
  INV_X4 mul_ex_mult_86_U83 ( .A(f1_in[26]), .ZN(mul_ex_mult_86_n73) );
  INV_X4 mul_ex_mult_86_U82 ( .A(f1_in[27]), .ZN(mul_ex_mult_86_n74) );
  INV_X4 mul_ex_mult_86_U81 ( .A(f1_in[28]), .ZN(mul_ex_mult_86_n75) );
  INV_X4 mul_ex_mult_86_U80 ( .A(f1_in[30]), .ZN(mul_ex_mult_86_n77) );
  INV_X4 mul_ex_mult_86_U79 ( .A(f1_in[31]), .ZN(mul_ex_mult_86_n78) );
  INV_X4 mul_ex_mult_86_U78 ( .A(f2_in[31]), .ZN(mul_ex_mult_86_n94) );
  INV_X4 mul_ex_mult_86_U77 ( .A(f2_in[16]), .ZN(mul_ex_mult_86_n79) );
  INV_X4 mul_ex_mult_86_U76 ( .A(f2_in[17]), .ZN(mul_ex_mult_86_n80) );
  INV_X4 mul_ex_mult_86_U75 ( .A(f2_in[19]), .ZN(mul_ex_mult_86_n82) );
  INV_X4 mul_ex_mult_86_U74 ( .A(f2_in[18]), .ZN(mul_ex_mult_86_n81) );
  INV_X4 mul_ex_mult_86_U73 ( .A(f2_in[21]), .ZN(mul_ex_mult_86_n84) );
  INV_X4 mul_ex_mult_86_U72 ( .A(f2_in[20]), .ZN(mul_ex_mult_86_n83) );
  INV_X4 mul_ex_mult_86_U71 ( .A(f2_in[23]), .ZN(mul_ex_mult_86_n86) );
  INV_X4 mul_ex_mult_86_U70 ( .A(f2_in[22]), .ZN(mul_ex_mult_86_n85) );
  INV_X4 mul_ex_mult_86_U69 ( .A(f2_in[25]), .ZN(mul_ex_mult_86_n88) );
  INV_X4 mul_ex_mult_86_U68 ( .A(f2_in[26]), .ZN(mul_ex_mult_86_n89) );
  INV_X4 mul_ex_mult_86_U67 ( .A(f2_in[27]), .ZN(mul_ex_mult_86_n90) );
  INV_X4 mul_ex_mult_86_U66 ( .A(f2_in[28]), .ZN(mul_ex_mult_86_n91) );
  INV_X4 mul_ex_mult_86_U65 ( .A(f2_in[29]), .ZN(mul_ex_mult_86_n92) );
  INV_X4 mul_ex_mult_86_U64 ( .A(f2_in[30]), .ZN(mul_ex_mult_86_n93) );
  INV_X4 mul_ex_mult_86_U63 ( .A(f2_in[24]), .ZN(mul_ex_mult_86_n87) );
  INV_X4 mul_ex_mult_86_U62 ( .A(f1_in[22]), .ZN(mul_ex_mult_86_n69) );
  AND2_X4 mul_ex_mult_86_U61 ( .A1(mul_ex_mult_86_CARRYB_15__14_), .A2(
        mul_ex_mult_86_ab_15__15_), .ZN(mul_ex_mult_86_n62) );
  XOR2_X2 mul_ex_mult_86_U60 ( .A(mul_ex_mult_86_CARRYB_15__0_), .B(
        mul_ex_mult_86_SUMB_15__1_), .Z(mul_ex_mult_86_n61) );
  XOR2_X2 mul_ex_mult_86_U59 ( .A(mul_ex_mult_86_ab_1__0_), .B(
        mul_ex_mult_86_ab_0__1_), .Z(mul_ex_N123) );
  AND2_X4 mul_ex_mult_86_U58 ( .A1(mul_ex_mult_86_CARRYB_15__0_), .A2(
        mul_ex_mult_86_SUMB_15__1_), .ZN(mul_ex_mult_86_n59) );
  AND2_X4 mul_ex_mult_86_U57 ( .A1(mul_ex_mult_86_CARRYB_15__2_), .A2(
        mul_ex_mult_86_SUMB_15__3_), .ZN(mul_ex_mult_86_n58) );
  AND2_X4 mul_ex_mult_86_U56 ( .A1(mul_ex_mult_86_CARRYB_15__4_), .A2(
        mul_ex_mult_86_SUMB_15__5_), .ZN(mul_ex_mult_86_n57) );
  AND2_X4 mul_ex_mult_86_U55 ( .A1(mul_ex_mult_86_CARRYB_15__6_), .A2(
        mul_ex_mult_86_SUMB_15__7_), .ZN(mul_ex_mult_86_n56) );
  AND2_X4 mul_ex_mult_86_U54 ( .A1(mul_ex_mult_86_CARRYB_15__8_), .A2(
        mul_ex_mult_86_SUMB_15__9_), .ZN(mul_ex_mult_86_n55) );
  AND2_X4 mul_ex_mult_86_U53 ( .A1(mul_ex_mult_86_CARRYB_15__10_), .A2(
        mul_ex_mult_86_SUMB_15__11_), .ZN(mul_ex_mult_86_n54) );
  AND2_X4 mul_ex_mult_86_U52 ( .A1(mul_ex_mult_86_CARRYB_15__12_), .A2(
        mul_ex_mult_86_SUMB_15__13_), .ZN(mul_ex_mult_86_n53) );
  AND2_X4 mul_ex_mult_86_U51 ( .A1(mul_ex_mult_86_CARRYB_15__1_), .A2(
        mul_ex_mult_86_SUMB_15__2_), .ZN(mul_ex_mult_86_n52) );
  AND2_X4 mul_ex_mult_86_U50 ( .A1(mul_ex_mult_86_CARRYB_15__3_), .A2(
        mul_ex_mult_86_SUMB_15__4_), .ZN(mul_ex_mult_86_n51) );
  AND2_X4 mul_ex_mult_86_U49 ( .A1(mul_ex_mult_86_CARRYB_15__5_), .A2(
        mul_ex_mult_86_SUMB_15__6_), .ZN(mul_ex_mult_86_n50) );
  AND2_X4 mul_ex_mult_86_U48 ( .A1(mul_ex_mult_86_CARRYB_15__7_), .A2(
        mul_ex_mult_86_SUMB_15__8_), .ZN(mul_ex_mult_86_n49) );
  AND2_X4 mul_ex_mult_86_U47 ( .A1(mul_ex_mult_86_CARRYB_15__9_), .A2(
        mul_ex_mult_86_SUMB_15__10_), .ZN(mul_ex_mult_86_n48) );
  AND2_X4 mul_ex_mult_86_U46 ( .A1(mul_ex_mult_86_CARRYB_15__11_), .A2(
        mul_ex_mult_86_SUMB_15__12_), .ZN(mul_ex_mult_86_n47) );
  AND2_X4 mul_ex_mult_86_U45 ( .A1(mul_ex_mult_86_CARRYB_15__13_), .A2(
        mul_ex_mult_86_SUMB_15__14_), .ZN(mul_ex_mult_86_n46) );
  XOR2_X2 mul_ex_mult_86_U44 ( .A(mul_ex_mult_86_ab_1__1_), .B(
        mul_ex_mult_86_ab_0__2_), .Z(mul_ex_mult_86_n45) );
  XOR2_X2 mul_ex_mult_86_U43 ( .A(mul_ex_mult_86_ab_1__2_), .B(
        mul_ex_mult_86_ab_0__3_), .Z(mul_ex_mult_86_n44) );
  XOR2_X2 mul_ex_mult_86_U42 ( .A(mul_ex_mult_86_ab_1__3_), .B(
        mul_ex_mult_86_ab_0__4_), .Z(mul_ex_mult_86_n43) );
  XOR2_X2 mul_ex_mult_86_U41 ( .A(mul_ex_mult_86_ab_1__4_), .B(
        mul_ex_mult_86_ab_0__5_), .Z(mul_ex_mult_86_n42) );
  XOR2_X2 mul_ex_mult_86_U40 ( .A(mul_ex_mult_86_ab_1__5_), .B(
        mul_ex_mult_86_ab_0__6_), .Z(mul_ex_mult_86_n41) );
  XOR2_X2 mul_ex_mult_86_U39 ( .A(mul_ex_mult_86_ab_1__6_), .B(
        mul_ex_mult_86_ab_0__7_), .Z(mul_ex_mult_86_n40) );
  XOR2_X2 mul_ex_mult_86_U38 ( .A(mul_ex_mult_86_ab_1__7_), .B(
        mul_ex_mult_86_ab_0__8_), .Z(mul_ex_mult_86_n39) );
  XOR2_X2 mul_ex_mult_86_U37 ( .A(mul_ex_mult_86_ab_1__8_), .B(
        mul_ex_mult_86_ab_0__9_), .Z(mul_ex_mult_86_n38) );
  XOR2_X2 mul_ex_mult_86_U36 ( .A(mul_ex_mult_86_ab_1__9_), .B(
        mul_ex_mult_86_ab_0__10_), .Z(mul_ex_mult_86_n37) );
  XOR2_X2 mul_ex_mult_86_U35 ( .A(mul_ex_mult_86_ab_1__10_), .B(
        mul_ex_mult_86_ab_0__11_), .Z(mul_ex_mult_86_n36) );
  XOR2_X2 mul_ex_mult_86_U34 ( .A(mul_ex_mult_86_ab_1__11_), .B(
        mul_ex_mult_86_ab_0__12_), .Z(mul_ex_mult_86_n35) );
  XOR2_X2 mul_ex_mult_86_U33 ( .A(mul_ex_mult_86_ab_1__12_), .B(
        mul_ex_mult_86_ab_0__13_), .Z(mul_ex_mult_86_n34) );
  XOR2_X2 mul_ex_mult_86_U32 ( .A(mul_ex_mult_86_ab_1__13_), .B(
        mul_ex_mult_86_ab_0__14_), .Z(mul_ex_mult_86_n33) );
  XOR2_X2 mul_ex_mult_86_U31 ( .A(mul_ex_mult_86_ab_1__14_), .B(
        mul_ex_mult_86_ab_0__15_), .Z(mul_ex_mult_86_n32) );
  AND2_X4 mul_ex_mult_86_U30 ( .A1(mul_ex_mult_86_ab_0__15_), .A2(
        mul_ex_mult_86_ab_1__14_), .ZN(mul_ex_mult_86_n31) );
  XOR2_X2 mul_ex_mult_86_U29 ( .A(mul_ex_mult_86_CARRYB_15__3_), .B(
        mul_ex_mult_86_SUMB_15__4_), .Z(mul_ex_mult_86_n30) );
  XOR2_X2 mul_ex_mult_86_U28 ( .A(mul_ex_mult_86_CARRYB_15__5_), .B(
        mul_ex_mult_86_SUMB_15__6_), .Z(mul_ex_mult_86_n29) );
  XOR2_X2 mul_ex_mult_86_U27 ( .A(mul_ex_mult_86_CARRYB_15__7_), .B(
        mul_ex_mult_86_SUMB_15__8_), .Z(mul_ex_mult_86_n28) );
  XOR2_X2 mul_ex_mult_86_U26 ( .A(mul_ex_mult_86_CARRYB_15__9_), .B(
        mul_ex_mult_86_SUMB_15__10_), .Z(mul_ex_mult_86_n27) );
  XOR2_X2 mul_ex_mult_86_U25 ( .A(mul_ex_mult_86_CARRYB_15__11_), .B(
        mul_ex_mult_86_SUMB_15__12_), .Z(mul_ex_mult_86_n26) );
  XOR2_X2 mul_ex_mult_86_U24 ( .A(mul_ex_mult_86_CARRYB_15__13_), .B(
        mul_ex_mult_86_SUMB_15__14_), .Z(mul_ex_mult_86_n25) );
  XOR2_X2 mul_ex_mult_86_U23 ( .A(mul_ex_mult_86_CARRYB_15__1_), .B(
        mul_ex_mult_86_SUMB_15__2_), .Z(mul_ex_mult_86_n24) );
  XOR2_X2 mul_ex_mult_86_U22 ( .A(mul_ex_mult_86_CARRYB_15__2_), .B(
        mul_ex_mult_86_SUMB_15__3_), .Z(mul_ex_mult_86_n23) );
  XOR2_X2 mul_ex_mult_86_U21 ( .A(mul_ex_mult_86_CARRYB_15__4_), .B(
        mul_ex_mult_86_SUMB_15__5_), .Z(mul_ex_mult_86_n22) );
  XOR2_X2 mul_ex_mult_86_U20 ( .A(mul_ex_mult_86_CARRYB_15__6_), .B(
        mul_ex_mult_86_SUMB_15__7_), .Z(mul_ex_mult_86_n21) );
  XOR2_X2 mul_ex_mult_86_U19 ( .A(mul_ex_mult_86_CARRYB_15__8_), .B(
        mul_ex_mult_86_SUMB_15__9_), .Z(mul_ex_mult_86_n20) );
  XOR2_X2 mul_ex_mult_86_U18 ( .A(mul_ex_mult_86_CARRYB_15__10_), .B(
        mul_ex_mult_86_SUMB_15__11_), .Z(mul_ex_mult_86_n19) );
  XOR2_X2 mul_ex_mult_86_U17 ( .A(mul_ex_mult_86_CARRYB_15__12_), .B(
        mul_ex_mult_86_SUMB_15__13_), .Z(mul_ex_mult_86_n18) );
  XOR2_X2 mul_ex_mult_86_U16 ( .A(mul_ex_mult_86_CARRYB_15__14_), .B(
        mul_ex_mult_86_ab_15__15_), .Z(mul_ex_mult_86_n17) );
  AND2_X4 mul_ex_mult_86_U15 ( .A1(mul_ex_mult_86_ab_0__1_), .A2(
        mul_ex_mult_86_ab_1__0_), .ZN(mul_ex_mult_86_n16) );
  AND2_X4 mul_ex_mult_86_U14 ( .A1(mul_ex_mult_86_ab_0__2_), .A2(
        mul_ex_mult_86_ab_1__1_), .ZN(mul_ex_mult_86_n15) );
  AND2_X4 mul_ex_mult_86_U13 ( .A1(mul_ex_mult_86_ab_0__3_), .A2(
        mul_ex_mult_86_ab_1__2_), .ZN(mul_ex_mult_86_n14) );
  AND2_X4 mul_ex_mult_86_U12 ( .A1(mul_ex_mult_86_ab_0__4_), .A2(
        mul_ex_mult_86_ab_1__3_), .ZN(mul_ex_mult_86_n13) );
  AND2_X4 mul_ex_mult_86_U11 ( .A1(mul_ex_mult_86_ab_0__5_), .A2(
        mul_ex_mult_86_ab_1__4_), .ZN(mul_ex_mult_86_n12) );
  AND2_X4 mul_ex_mult_86_U10 ( .A1(mul_ex_mult_86_ab_0__6_), .A2(
        mul_ex_mult_86_ab_1__5_), .ZN(mul_ex_mult_86_n11) );
  AND2_X4 mul_ex_mult_86_U9 ( .A1(mul_ex_mult_86_ab_0__7_), .A2(
        mul_ex_mult_86_ab_1__6_), .ZN(mul_ex_mult_86_n10) );
  AND2_X4 mul_ex_mult_86_U8 ( .A1(mul_ex_mult_86_ab_0__8_), .A2(
        mul_ex_mult_86_ab_1__7_), .ZN(mul_ex_mult_86_n9) );
  AND2_X4 mul_ex_mult_86_U7 ( .A1(mul_ex_mult_86_ab_0__9_), .A2(
        mul_ex_mult_86_ab_1__8_), .ZN(mul_ex_mult_86_n8) );
  AND2_X4 mul_ex_mult_86_U6 ( .A1(mul_ex_mult_86_ab_0__10_), .A2(
        mul_ex_mult_86_ab_1__9_), .ZN(mul_ex_mult_86_n7) );
  AND2_X4 mul_ex_mult_86_U5 ( .A1(mul_ex_mult_86_ab_0__11_), .A2(
        mul_ex_mult_86_ab_1__10_), .ZN(mul_ex_mult_86_n6) );
  AND2_X4 mul_ex_mult_86_U4 ( .A1(mul_ex_mult_86_ab_0__12_), .A2(
        mul_ex_mult_86_ab_1__11_), .ZN(mul_ex_mult_86_n5) );
  AND2_X4 mul_ex_mult_86_U3 ( .A1(mul_ex_mult_86_ab_0__13_), .A2(
        mul_ex_mult_86_ab_1__12_), .ZN(mul_ex_mult_86_n4) );
  AND2_X4 mul_ex_mult_86_U2 ( .A1(mul_ex_mult_86_ab_0__14_), .A2(
        mul_ex_mult_86_ab_1__13_), .ZN(mul_ex_mult_86_n3) );
  FA_X1 mul_ex_mult_86_S3_2_14 ( .A(mul_ex_mult_86_ab_2__14_), .B(
        mul_ex_mult_86_n31), .CI(mul_ex_mult_86_ab_1__15_), .CO(
        mul_ex_mult_86_CARRYB_2__14_), .S(mul_ex_mult_86_SUMB_2__14_) );
  FA_X1 mul_ex_mult_86_S2_2_13 ( .A(mul_ex_mult_86_ab_2__13_), .B(
        mul_ex_mult_86_n3), .CI(mul_ex_mult_86_n32), .CO(
        mul_ex_mult_86_CARRYB_2__13_), .S(mul_ex_mult_86_SUMB_2__13_) );
  FA_X1 mul_ex_mult_86_S2_2_12 ( .A(mul_ex_mult_86_ab_2__12_), .B(
        mul_ex_mult_86_n4), .CI(mul_ex_mult_86_n33), .CO(
        mul_ex_mult_86_CARRYB_2__12_), .S(mul_ex_mult_86_SUMB_2__12_) );
  FA_X1 mul_ex_mult_86_S2_2_11 ( .A(mul_ex_mult_86_ab_2__11_), .B(
        mul_ex_mult_86_n5), .CI(mul_ex_mult_86_n34), .CO(
        mul_ex_mult_86_CARRYB_2__11_), .S(mul_ex_mult_86_SUMB_2__11_) );
  FA_X1 mul_ex_mult_86_S2_2_10 ( .A(mul_ex_mult_86_ab_2__10_), .B(
        mul_ex_mult_86_n6), .CI(mul_ex_mult_86_n35), .CO(
        mul_ex_mult_86_CARRYB_2__10_), .S(mul_ex_mult_86_SUMB_2__10_) );
  FA_X1 mul_ex_mult_86_S2_2_9 ( .A(mul_ex_mult_86_ab_2__9_), .B(
        mul_ex_mult_86_n7), .CI(mul_ex_mult_86_n36), .CO(
        mul_ex_mult_86_CARRYB_2__9_), .S(mul_ex_mult_86_SUMB_2__9_) );
  FA_X1 mul_ex_mult_86_S2_2_8 ( .A(mul_ex_mult_86_ab_2__8_), .B(
        mul_ex_mult_86_n8), .CI(mul_ex_mult_86_n37), .CO(
        mul_ex_mult_86_CARRYB_2__8_), .S(mul_ex_mult_86_SUMB_2__8_) );
  FA_X1 mul_ex_mult_86_S2_2_7 ( .A(mul_ex_mult_86_ab_2__7_), .B(
        mul_ex_mult_86_n9), .CI(mul_ex_mult_86_n38), .CO(
        mul_ex_mult_86_CARRYB_2__7_), .S(mul_ex_mult_86_SUMB_2__7_) );
  FA_X1 mul_ex_mult_86_S2_2_6 ( .A(mul_ex_mult_86_ab_2__6_), .B(
        mul_ex_mult_86_n10), .CI(mul_ex_mult_86_n39), .CO(
        mul_ex_mult_86_CARRYB_2__6_), .S(mul_ex_mult_86_SUMB_2__6_) );
  FA_X1 mul_ex_mult_86_S2_2_5 ( .A(mul_ex_mult_86_ab_2__5_), .B(
        mul_ex_mult_86_n11), .CI(mul_ex_mult_86_n40), .CO(
        mul_ex_mult_86_CARRYB_2__5_), .S(mul_ex_mult_86_SUMB_2__5_) );
  FA_X1 mul_ex_mult_86_S2_2_4 ( .A(mul_ex_mult_86_ab_2__4_), .B(
        mul_ex_mult_86_n12), .CI(mul_ex_mult_86_n41), .CO(
        mul_ex_mult_86_CARRYB_2__4_), .S(mul_ex_mult_86_SUMB_2__4_) );
  FA_X1 mul_ex_mult_86_S2_2_3 ( .A(mul_ex_mult_86_ab_2__3_), .B(
        mul_ex_mult_86_n13), .CI(mul_ex_mult_86_n42), .CO(
        mul_ex_mult_86_CARRYB_2__3_), .S(mul_ex_mult_86_SUMB_2__3_) );
  FA_X1 mul_ex_mult_86_S2_2_2 ( .A(mul_ex_mult_86_ab_2__2_), .B(
        mul_ex_mult_86_n14), .CI(mul_ex_mult_86_n43), .CO(
        mul_ex_mult_86_CARRYB_2__2_), .S(mul_ex_mult_86_SUMB_2__2_) );
  FA_X1 mul_ex_mult_86_S2_2_1 ( .A(mul_ex_mult_86_ab_2__1_), .B(
        mul_ex_mult_86_n15), .CI(mul_ex_mult_86_n44), .CO(
        mul_ex_mult_86_CARRYB_2__1_), .S(mul_ex_mult_86_SUMB_2__1_) );
  FA_X1 mul_ex_mult_86_S1_2_0 ( .A(mul_ex_mult_86_ab_2__0_), .B(
        mul_ex_mult_86_n16), .CI(mul_ex_mult_86_n45), .CO(
        mul_ex_mult_86_CARRYB_2__0_), .S(mul_ex_mult_86_A1_0_) );
  FA_X1 mul_ex_mult_86_S3_3_14 ( .A(mul_ex_mult_86_ab_3__14_), .B(
        mul_ex_mult_86_CARRYB_2__14_), .CI(mul_ex_mult_86_ab_2__15_), .CO(
        mul_ex_mult_86_CARRYB_3__14_), .S(mul_ex_mult_86_SUMB_3__14_) );
  FA_X1 mul_ex_mult_86_S2_3_13 ( .A(mul_ex_mult_86_ab_3__13_), .B(
        mul_ex_mult_86_CARRYB_2__13_), .CI(mul_ex_mult_86_SUMB_2__14_), .CO(
        mul_ex_mult_86_CARRYB_3__13_), .S(mul_ex_mult_86_SUMB_3__13_) );
  FA_X1 mul_ex_mult_86_S2_3_12 ( .A(mul_ex_mult_86_ab_3__12_), .B(
        mul_ex_mult_86_CARRYB_2__12_), .CI(mul_ex_mult_86_SUMB_2__13_), .CO(
        mul_ex_mult_86_CARRYB_3__12_), .S(mul_ex_mult_86_SUMB_3__12_) );
  FA_X1 mul_ex_mult_86_S2_3_11 ( .A(mul_ex_mult_86_ab_3__11_), .B(
        mul_ex_mult_86_CARRYB_2__11_), .CI(mul_ex_mult_86_SUMB_2__12_), .CO(
        mul_ex_mult_86_CARRYB_3__11_), .S(mul_ex_mult_86_SUMB_3__11_) );
  FA_X1 mul_ex_mult_86_S2_3_10 ( .A(mul_ex_mult_86_ab_3__10_), .B(
        mul_ex_mult_86_CARRYB_2__10_), .CI(mul_ex_mult_86_SUMB_2__11_), .CO(
        mul_ex_mult_86_CARRYB_3__10_), .S(mul_ex_mult_86_SUMB_3__10_) );
  FA_X1 mul_ex_mult_86_S2_3_9 ( .A(mul_ex_mult_86_ab_3__9_), .B(
        mul_ex_mult_86_CARRYB_2__9_), .CI(mul_ex_mult_86_SUMB_2__10_), .CO(
        mul_ex_mult_86_CARRYB_3__9_), .S(mul_ex_mult_86_SUMB_3__9_) );
  FA_X1 mul_ex_mult_86_S2_3_8 ( .A(mul_ex_mult_86_ab_3__8_), .B(
        mul_ex_mult_86_CARRYB_2__8_), .CI(mul_ex_mult_86_SUMB_2__9_), .CO(
        mul_ex_mult_86_CARRYB_3__8_), .S(mul_ex_mult_86_SUMB_3__8_) );
  FA_X1 mul_ex_mult_86_S2_3_7 ( .A(mul_ex_mult_86_ab_3__7_), .B(
        mul_ex_mult_86_CARRYB_2__7_), .CI(mul_ex_mult_86_SUMB_2__8_), .CO(
        mul_ex_mult_86_CARRYB_3__7_), .S(mul_ex_mult_86_SUMB_3__7_) );
  FA_X1 mul_ex_mult_86_S2_3_6 ( .A(mul_ex_mult_86_ab_3__6_), .B(
        mul_ex_mult_86_CARRYB_2__6_), .CI(mul_ex_mult_86_SUMB_2__7_), .CO(
        mul_ex_mult_86_CARRYB_3__6_), .S(mul_ex_mult_86_SUMB_3__6_) );
  FA_X1 mul_ex_mult_86_S2_3_5 ( .A(mul_ex_mult_86_ab_3__5_), .B(
        mul_ex_mult_86_CARRYB_2__5_), .CI(mul_ex_mult_86_SUMB_2__6_), .CO(
        mul_ex_mult_86_CARRYB_3__5_), .S(mul_ex_mult_86_SUMB_3__5_) );
  FA_X1 mul_ex_mult_86_S2_3_4 ( .A(mul_ex_mult_86_ab_3__4_), .B(
        mul_ex_mult_86_CARRYB_2__4_), .CI(mul_ex_mult_86_SUMB_2__5_), .CO(
        mul_ex_mult_86_CARRYB_3__4_), .S(mul_ex_mult_86_SUMB_3__4_) );
  FA_X1 mul_ex_mult_86_S2_3_3 ( .A(mul_ex_mult_86_ab_3__3_), .B(
        mul_ex_mult_86_CARRYB_2__3_), .CI(mul_ex_mult_86_SUMB_2__4_), .CO(
        mul_ex_mult_86_CARRYB_3__3_), .S(mul_ex_mult_86_SUMB_3__3_) );
  FA_X1 mul_ex_mult_86_S2_3_2 ( .A(mul_ex_mult_86_ab_3__2_), .B(
        mul_ex_mult_86_CARRYB_2__2_), .CI(mul_ex_mult_86_SUMB_2__3_), .CO(
        mul_ex_mult_86_CARRYB_3__2_), .S(mul_ex_mult_86_SUMB_3__2_) );
  FA_X1 mul_ex_mult_86_S2_3_1 ( .A(mul_ex_mult_86_ab_3__1_), .B(
        mul_ex_mult_86_CARRYB_2__1_), .CI(mul_ex_mult_86_SUMB_2__2_), .CO(
        mul_ex_mult_86_CARRYB_3__1_), .S(mul_ex_mult_86_SUMB_3__1_) );
  FA_X1 mul_ex_mult_86_S1_3_0 ( .A(mul_ex_mult_86_ab_3__0_), .B(
        mul_ex_mult_86_CARRYB_2__0_), .CI(mul_ex_mult_86_SUMB_2__1_), .CO(
        mul_ex_mult_86_CARRYB_3__0_), .S(mul_ex_mult_86_A1_1_) );
  FA_X1 mul_ex_mult_86_S3_4_14 ( .A(mul_ex_mult_86_ab_4__14_), .B(
        mul_ex_mult_86_CARRYB_3__14_), .CI(mul_ex_mult_86_ab_3__15_), .CO(
        mul_ex_mult_86_CARRYB_4__14_), .S(mul_ex_mult_86_SUMB_4__14_) );
  FA_X1 mul_ex_mult_86_S2_4_13 ( .A(mul_ex_mult_86_ab_4__13_), .B(
        mul_ex_mult_86_CARRYB_3__13_), .CI(mul_ex_mult_86_SUMB_3__14_), .CO(
        mul_ex_mult_86_CARRYB_4__13_), .S(mul_ex_mult_86_SUMB_4__13_) );
  FA_X1 mul_ex_mult_86_S2_4_12 ( .A(mul_ex_mult_86_ab_4__12_), .B(
        mul_ex_mult_86_CARRYB_3__12_), .CI(mul_ex_mult_86_SUMB_3__13_), .CO(
        mul_ex_mult_86_CARRYB_4__12_), .S(mul_ex_mult_86_SUMB_4__12_) );
  FA_X1 mul_ex_mult_86_S2_4_11 ( .A(mul_ex_mult_86_ab_4__11_), .B(
        mul_ex_mult_86_CARRYB_3__11_), .CI(mul_ex_mult_86_SUMB_3__12_), .CO(
        mul_ex_mult_86_CARRYB_4__11_), .S(mul_ex_mult_86_SUMB_4__11_) );
  FA_X1 mul_ex_mult_86_S2_4_10 ( .A(mul_ex_mult_86_ab_4__10_), .B(
        mul_ex_mult_86_CARRYB_3__10_), .CI(mul_ex_mult_86_SUMB_3__11_), .CO(
        mul_ex_mult_86_CARRYB_4__10_), .S(mul_ex_mult_86_SUMB_4__10_) );
  FA_X1 mul_ex_mult_86_S2_4_9 ( .A(mul_ex_mult_86_ab_4__9_), .B(
        mul_ex_mult_86_CARRYB_3__9_), .CI(mul_ex_mult_86_SUMB_3__10_), .CO(
        mul_ex_mult_86_CARRYB_4__9_), .S(mul_ex_mult_86_SUMB_4__9_) );
  FA_X1 mul_ex_mult_86_S2_4_8 ( .A(mul_ex_mult_86_ab_4__8_), .B(
        mul_ex_mult_86_CARRYB_3__8_), .CI(mul_ex_mult_86_SUMB_3__9_), .CO(
        mul_ex_mult_86_CARRYB_4__8_), .S(mul_ex_mult_86_SUMB_4__8_) );
  FA_X1 mul_ex_mult_86_S2_4_7 ( .A(mul_ex_mult_86_ab_4__7_), .B(
        mul_ex_mult_86_CARRYB_3__7_), .CI(mul_ex_mult_86_SUMB_3__8_), .CO(
        mul_ex_mult_86_CARRYB_4__7_), .S(mul_ex_mult_86_SUMB_4__7_) );
  FA_X1 mul_ex_mult_86_S2_4_6 ( .A(mul_ex_mult_86_ab_4__6_), .B(
        mul_ex_mult_86_CARRYB_3__6_), .CI(mul_ex_mult_86_SUMB_3__7_), .CO(
        mul_ex_mult_86_CARRYB_4__6_), .S(mul_ex_mult_86_SUMB_4__6_) );
  FA_X1 mul_ex_mult_86_S2_4_5 ( .A(mul_ex_mult_86_ab_4__5_), .B(
        mul_ex_mult_86_CARRYB_3__5_), .CI(mul_ex_mult_86_SUMB_3__6_), .CO(
        mul_ex_mult_86_CARRYB_4__5_), .S(mul_ex_mult_86_SUMB_4__5_) );
  FA_X1 mul_ex_mult_86_S2_4_4 ( .A(mul_ex_mult_86_ab_4__4_), .B(
        mul_ex_mult_86_CARRYB_3__4_), .CI(mul_ex_mult_86_SUMB_3__5_), .CO(
        mul_ex_mult_86_CARRYB_4__4_), .S(mul_ex_mult_86_SUMB_4__4_) );
  FA_X1 mul_ex_mult_86_S2_4_3 ( .A(mul_ex_mult_86_ab_4__3_), .B(
        mul_ex_mult_86_CARRYB_3__3_), .CI(mul_ex_mult_86_SUMB_3__4_), .CO(
        mul_ex_mult_86_CARRYB_4__3_), .S(mul_ex_mult_86_SUMB_4__3_) );
  FA_X1 mul_ex_mult_86_S2_4_2 ( .A(mul_ex_mult_86_ab_4__2_), .B(
        mul_ex_mult_86_CARRYB_3__2_), .CI(mul_ex_mult_86_SUMB_3__3_), .CO(
        mul_ex_mult_86_CARRYB_4__2_), .S(mul_ex_mult_86_SUMB_4__2_) );
  FA_X1 mul_ex_mult_86_S2_4_1 ( .A(mul_ex_mult_86_ab_4__1_), .B(
        mul_ex_mult_86_CARRYB_3__1_), .CI(mul_ex_mult_86_SUMB_3__2_), .CO(
        mul_ex_mult_86_CARRYB_4__1_), .S(mul_ex_mult_86_SUMB_4__1_) );
  FA_X1 mul_ex_mult_86_S1_4_0 ( .A(mul_ex_mult_86_ab_4__0_), .B(
        mul_ex_mult_86_CARRYB_3__0_), .CI(mul_ex_mult_86_SUMB_3__1_), .CO(
        mul_ex_mult_86_CARRYB_4__0_), .S(mul_ex_mult_86_A1_2_) );
  FA_X1 mul_ex_mult_86_S3_5_14 ( .A(mul_ex_mult_86_ab_5__14_), .B(
        mul_ex_mult_86_CARRYB_4__14_), .CI(mul_ex_mult_86_ab_4__15_), .CO(
        mul_ex_mult_86_CARRYB_5__14_), .S(mul_ex_mult_86_SUMB_5__14_) );
  FA_X1 mul_ex_mult_86_S2_5_13 ( .A(mul_ex_mult_86_ab_5__13_), .B(
        mul_ex_mult_86_CARRYB_4__13_), .CI(mul_ex_mult_86_SUMB_4__14_), .CO(
        mul_ex_mult_86_CARRYB_5__13_), .S(mul_ex_mult_86_SUMB_5__13_) );
  FA_X1 mul_ex_mult_86_S2_5_12 ( .A(mul_ex_mult_86_ab_5__12_), .B(
        mul_ex_mult_86_CARRYB_4__12_), .CI(mul_ex_mult_86_SUMB_4__13_), .CO(
        mul_ex_mult_86_CARRYB_5__12_), .S(mul_ex_mult_86_SUMB_5__12_) );
  FA_X1 mul_ex_mult_86_S2_5_11 ( .A(mul_ex_mult_86_ab_5__11_), .B(
        mul_ex_mult_86_CARRYB_4__11_), .CI(mul_ex_mult_86_SUMB_4__12_), .CO(
        mul_ex_mult_86_CARRYB_5__11_), .S(mul_ex_mult_86_SUMB_5__11_) );
  FA_X1 mul_ex_mult_86_S2_5_10 ( .A(mul_ex_mult_86_ab_5__10_), .B(
        mul_ex_mult_86_CARRYB_4__10_), .CI(mul_ex_mult_86_SUMB_4__11_), .CO(
        mul_ex_mult_86_CARRYB_5__10_), .S(mul_ex_mult_86_SUMB_5__10_) );
  FA_X1 mul_ex_mult_86_S2_5_9 ( .A(mul_ex_mult_86_ab_5__9_), .B(
        mul_ex_mult_86_CARRYB_4__9_), .CI(mul_ex_mult_86_SUMB_4__10_), .CO(
        mul_ex_mult_86_CARRYB_5__9_), .S(mul_ex_mult_86_SUMB_5__9_) );
  FA_X1 mul_ex_mult_86_S2_5_8 ( .A(mul_ex_mult_86_ab_5__8_), .B(
        mul_ex_mult_86_CARRYB_4__8_), .CI(mul_ex_mult_86_SUMB_4__9_), .CO(
        mul_ex_mult_86_CARRYB_5__8_), .S(mul_ex_mult_86_SUMB_5__8_) );
  FA_X1 mul_ex_mult_86_S2_5_7 ( .A(mul_ex_mult_86_ab_5__7_), .B(
        mul_ex_mult_86_CARRYB_4__7_), .CI(mul_ex_mult_86_SUMB_4__8_), .CO(
        mul_ex_mult_86_CARRYB_5__7_), .S(mul_ex_mult_86_SUMB_5__7_) );
  FA_X1 mul_ex_mult_86_S2_5_6 ( .A(mul_ex_mult_86_ab_5__6_), .B(
        mul_ex_mult_86_CARRYB_4__6_), .CI(mul_ex_mult_86_SUMB_4__7_), .CO(
        mul_ex_mult_86_CARRYB_5__6_), .S(mul_ex_mult_86_SUMB_5__6_) );
  FA_X1 mul_ex_mult_86_S2_5_5 ( .A(mul_ex_mult_86_ab_5__5_), .B(
        mul_ex_mult_86_CARRYB_4__5_), .CI(mul_ex_mult_86_SUMB_4__6_), .CO(
        mul_ex_mult_86_CARRYB_5__5_), .S(mul_ex_mult_86_SUMB_5__5_) );
  FA_X1 mul_ex_mult_86_S2_5_4 ( .A(mul_ex_mult_86_ab_5__4_), .B(
        mul_ex_mult_86_CARRYB_4__4_), .CI(mul_ex_mult_86_SUMB_4__5_), .CO(
        mul_ex_mult_86_CARRYB_5__4_), .S(mul_ex_mult_86_SUMB_5__4_) );
  FA_X1 mul_ex_mult_86_S2_5_3 ( .A(mul_ex_mult_86_ab_5__3_), .B(
        mul_ex_mult_86_CARRYB_4__3_), .CI(mul_ex_mult_86_SUMB_4__4_), .CO(
        mul_ex_mult_86_CARRYB_5__3_), .S(mul_ex_mult_86_SUMB_5__3_) );
  FA_X1 mul_ex_mult_86_S2_5_2 ( .A(mul_ex_mult_86_ab_5__2_), .B(
        mul_ex_mult_86_CARRYB_4__2_), .CI(mul_ex_mult_86_SUMB_4__3_), .CO(
        mul_ex_mult_86_CARRYB_5__2_), .S(mul_ex_mult_86_SUMB_5__2_) );
  FA_X1 mul_ex_mult_86_S2_5_1 ( .A(mul_ex_mult_86_ab_5__1_), .B(
        mul_ex_mult_86_CARRYB_4__1_), .CI(mul_ex_mult_86_SUMB_4__2_), .CO(
        mul_ex_mult_86_CARRYB_5__1_), .S(mul_ex_mult_86_SUMB_5__1_) );
  FA_X1 mul_ex_mult_86_S1_5_0 ( .A(mul_ex_mult_86_ab_5__0_), .B(
        mul_ex_mult_86_CARRYB_4__0_), .CI(mul_ex_mult_86_SUMB_4__1_), .CO(
        mul_ex_mult_86_CARRYB_5__0_), .S(mul_ex_mult_86_A1_3_) );
  FA_X1 mul_ex_mult_86_S3_6_14 ( .A(mul_ex_mult_86_ab_6__14_), .B(
        mul_ex_mult_86_CARRYB_5__14_), .CI(mul_ex_mult_86_ab_5__15_), .CO(
        mul_ex_mult_86_CARRYB_6__14_), .S(mul_ex_mult_86_SUMB_6__14_) );
  FA_X1 mul_ex_mult_86_S2_6_13 ( .A(mul_ex_mult_86_ab_6__13_), .B(
        mul_ex_mult_86_CARRYB_5__13_), .CI(mul_ex_mult_86_SUMB_5__14_), .CO(
        mul_ex_mult_86_CARRYB_6__13_), .S(mul_ex_mult_86_SUMB_6__13_) );
  FA_X1 mul_ex_mult_86_S2_6_12 ( .A(mul_ex_mult_86_ab_6__12_), .B(
        mul_ex_mult_86_CARRYB_5__12_), .CI(mul_ex_mult_86_SUMB_5__13_), .CO(
        mul_ex_mult_86_CARRYB_6__12_), .S(mul_ex_mult_86_SUMB_6__12_) );
  FA_X1 mul_ex_mult_86_S2_6_11 ( .A(mul_ex_mult_86_ab_6__11_), .B(
        mul_ex_mult_86_CARRYB_5__11_), .CI(mul_ex_mult_86_SUMB_5__12_), .CO(
        mul_ex_mult_86_CARRYB_6__11_), .S(mul_ex_mult_86_SUMB_6__11_) );
  FA_X1 mul_ex_mult_86_S2_6_10 ( .A(mul_ex_mult_86_ab_6__10_), .B(
        mul_ex_mult_86_CARRYB_5__10_), .CI(mul_ex_mult_86_SUMB_5__11_), .CO(
        mul_ex_mult_86_CARRYB_6__10_), .S(mul_ex_mult_86_SUMB_6__10_) );
  FA_X1 mul_ex_mult_86_S2_6_9 ( .A(mul_ex_mult_86_ab_6__9_), .B(
        mul_ex_mult_86_CARRYB_5__9_), .CI(mul_ex_mult_86_SUMB_5__10_), .CO(
        mul_ex_mult_86_CARRYB_6__9_), .S(mul_ex_mult_86_SUMB_6__9_) );
  FA_X1 mul_ex_mult_86_S2_6_8 ( .A(mul_ex_mult_86_ab_6__8_), .B(
        mul_ex_mult_86_CARRYB_5__8_), .CI(mul_ex_mult_86_SUMB_5__9_), .CO(
        mul_ex_mult_86_CARRYB_6__8_), .S(mul_ex_mult_86_SUMB_6__8_) );
  FA_X1 mul_ex_mult_86_S2_6_7 ( .A(mul_ex_mult_86_ab_6__7_), .B(
        mul_ex_mult_86_CARRYB_5__7_), .CI(mul_ex_mult_86_SUMB_5__8_), .CO(
        mul_ex_mult_86_CARRYB_6__7_), .S(mul_ex_mult_86_SUMB_6__7_) );
  FA_X1 mul_ex_mult_86_S2_6_6 ( .A(mul_ex_mult_86_ab_6__6_), .B(
        mul_ex_mult_86_CARRYB_5__6_), .CI(mul_ex_mult_86_SUMB_5__7_), .CO(
        mul_ex_mult_86_CARRYB_6__6_), .S(mul_ex_mult_86_SUMB_6__6_) );
  FA_X1 mul_ex_mult_86_S2_6_5 ( .A(mul_ex_mult_86_ab_6__5_), .B(
        mul_ex_mult_86_CARRYB_5__5_), .CI(mul_ex_mult_86_SUMB_5__6_), .CO(
        mul_ex_mult_86_CARRYB_6__5_), .S(mul_ex_mult_86_SUMB_6__5_) );
  FA_X1 mul_ex_mult_86_S2_6_4 ( .A(mul_ex_mult_86_ab_6__4_), .B(
        mul_ex_mult_86_CARRYB_5__4_), .CI(mul_ex_mult_86_SUMB_5__5_), .CO(
        mul_ex_mult_86_CARRYB_6__4_), .S(mul_ex_mult_86_SUMB_6__4_) );
  FA_X1 mul_ex_mult_86_S2_6_3 ( .A(mul_ex_mult_86_ab_6__3_), .B(
        mul_ex_mult_86_CARRYB_5__3_), .CI(mul_ex_mult_86_SUMB_5__4_), .CO(
        mul_ex_mult_86_CARRYB_6__3_), .S(mul_ex_mult_86_SUMB_6__3_) );
  FA_X1 mul_ex_mult_86_S2_6_2 ( .A(mul_ex_mult_86_ab_6__2_), .B(
        mul_ex_mult_86_CARRYB_5__2_), .CI(mul_ex_mult_86_SUMB_5__3_), .CO(
        mul_ex_mult_86_CARRYB_6__2_), .S(mul_ex_mult_86_SUMB_6__2_) );
  FA_X1 mul_ex_mult_86_S2_6_1 ( .A(mul_ex_mult_86_ab_6__1_), .B(
        mul_ex_mult_86_CARRYB_5__1_), .CI(mul_ex_mult_86_SUMB_5__2_), .CO(
        mul_ex_mult_86_CARRYB_6__1_), .S(mul_ex_mult_86_SUMB_6__1_) );
  FA_X1 mul_ex_mult_86_S1_6_0 ( .A(mul_ex_mult_86_ab_6__0_), .B(
        mul_ex_mult_86_CARRYB_5__0_), .CI(mul_ex_mult_86_SUMB_5__1_), .CO(
        mul_ex_mult_86_CARRYB_6__0_), .S(mul_ex_mult_86_A1_4_) );
  FA_X1 mul_ex_mult_86_S3_7_14 ( .A(mul_ex_mult_86_ab_7__14_), .B(
        mul_ex_mult_86_CARRYB_6__14_), .CI(mul_ex_mult_86_ab_6__15_), .CO(
        mul_ex_mult_86_CARRYB_7__14_), .S(mul_ex_mult_86_SUMB_7__14_) );
  FA_X1 mul_ex_mult_86_S2_7_13 ( .A(mul_ex_mult_86_ab_7__13_), .B(
        mul_ex_mult_86_CARRYB_6__13_), .CI(mul_ex_mult_86_SUMB_6__14_), .CO(
        mul_ex_mult_86_CARRYB_7__13_), .S(mul_ex_mult_86_SUMB_7__13_) );
  FA_X1 mul_ex_mult_86_S2_7_12 ( .A(mul_ex_mult_86_ab_7__12_), .B(
        mul_ex_mult_86_CARRYB_6__12_), .CI(mul_ex_mult_86_SUMB_6__13_), .CO(
        mul_ex_mult_86_CARRYB_7__12_), .S(mul_ex_mult_86_SUMB_7__12_) );
  FA_X1 mul_ex_mult_86_S2_7_11 ( .A(mul_ex_mult_86_ab_7__11_), .B(
        mul_ex_mult_86_CARRYB_6__11_), .CI(mul_ex_mult_86_SUMB_6__12_), .CO(
        mul_ex_mult_86_CARRYB_7__11_), .S(mul_ex_mult_86_SUMB_7__11_) );
  FA_X1 mul_ex_mult_86_S2_7_10 ( .A(mul_ex_mult_86_ab_7__10_), .B(
        mul_ex_mult_86_CARRYB_6__10_), .CI(mul_ex_mult_86_SUMB_6__11_), .CO(
        mul_ex_mult_86_CARRYB_7__10_), .S(mul_ex_mult_86_SUMB_7__10_) );
  FA_X1 mul_ex_mult_86_S2_7_9 ( .A(mul_ex_mult_86_ab_7__9_), .B(
        mul_ex_mult_86_CARRYB_6__9_), .CI(mul_ex_mult_86_SUMB_6__10_), .CO(
        mul_ex_mult_86_CARRYB_7__9_), .S(mul_ex_mult_86_SUMB_7__9_) );
  FA_X1 mul_ex_mult_86_S2_7_8 ( .A(mul_ex_mult_86_ab_7__8_), .B(
        mul_ex_mult_86_CARRYB_6__8_), .CI(mul_ex_mult_86_SUMB_6__9_), .CO(
        mul_ex_mult_86_CARRYB_7__8_), .S(mul_ex_mult_86_SUMB_7__8_) );
  FA_X1 mul_ex_mult_86_S2_7_7 ( .A(mul_ex_mult_86_ab_7__7_), .B(
        mul_ex_mult_86_CARRYB_6__7_), .CI(mul_ex_mult_86_SUMB_6__8_), .CO(
        mul_ex_mult_86_CARRYB_7__7_), .S(mul_ex_mult_86_SUMB_7__7_) );
  FA_X1 mul_ex_mult_86_S2_7_6 ( .A(mul_ex_mult_86_ab_7__6_), .B(
        mul_ex_mult_86_CARRYB_6__6_), .CI(mul_ex_mult_86_SUMB_6__7_), .CO(
        mul_ex_mult_86_CARRYB_7__6_), .S(mul_ex_mult_86_SUMB_7__6_) );
  FA_X1 mul_ex_mult_86_S2_7_5 ( .A(mul_ex_mult_86_ab_7__5_), .B(
        mul_ex_mult_86_CARRYB_6__5_), .CI(mul_ex_mult_86_SUMB_6__6_), .CO(
        mul_ex_mult_86_CARRYB_7__5_), .S(mul_ex_mult_86_SUMB_7__5_) );
  FA_X1 mul_ex_mult_86_S2_7_4 ( .A(mul_ex_mult_86_ab_7__4_), .B(
        mul_ex_mult_86_CARRYB_6__4_), .CI(mul_ex_mult_86_SUMB_6__5_), .CO(
        mul_ex_mult_86_CARRYB_7__4_), .S(mul_ex_mult_86_SUMB_7__4_) );
  FA_X1 mul_ex_mult_86_S2_7_3 ( .A(mul_ex_mult_86_ab_7__3_), .B(
        mul_ex_mult_86_CARRYB_6__3_), .CI(mul_ex_mult_86_SUMB_6__4_), .CO(
        mul_ex_mult_86_CARRYB_7__3_), .S(mul_ex_mult_86_SUMB_7__3_) );
  FA_X1 mul_ex_mult_86_S2_7_2 ( .A(mul_ex_mult_86_ab_7__2_), .B(
        mul_ex_mult_86_CARRYB_6__2_), .CI(mul_ex_mult_86_SUMB_6__3_), .CO(
        mul_ex_mult_86_CARRYB_7__2_), .S(mul_ex_mult_86_SUMB_7__2_) );
  FA_X1 mul_ex_mult_86_S2_7_1 ( .A(mul_ex_mult_86_ab_7__1_), .B(
        mul_ex_mult_86_CARRYB_6__1_), .CI(mul_ex_mult_86_SUMB_6__2_), .CO(
        mul_ex_mult_86_CARRYB_7__1_), .S(mul_ex_mult_86_SUMB_7__1_) );
  FA_X1 mul_ex_mult_86_S1_7_0 ( .A(mul_ex_mult_86_ab_7__0_), .B(
        mul_ex_mult_86_CARRYB_6__0_), .CI(mul_ex_mult_86_SUMB_6__1_), .CO(
        mul_ex_mult_86_CARRYB_7__0_), .S(mul_ex_mult_86_A1_5_) );
  FA_X1 mul_ex_mult_86_S3_8_14 ( .A(mul_ex_mult_86_ab_8__14_), .B(
        mul_ex_mult_86_CARRYB_7__14_), .CI(mul_ex_mult_86_ab_7__15_), .CO(
        mul_ex_mult_86_CARRYB_8__14_), .S(mul_ex_mult_86_SUMB_8__14_) );
  FA_X1 mul_ex_mult_86_S2_8_13 ( .A(mul_ex_mult_86_ab_8__13_), .B(
        mul_ex_mult_86_CARRYB_7__13_), .CI(mul_ex_mult_86_SUMB_7__14_), .CO(
        mul_ex_mult_86_CARRYB_8__13_), .S(mul_ex_mult_86_SUMB_8__13_) );
  FA_X1 mul_ex_mult_86_S2_8_12 ( .A(mul_ex_mult_86_ab_8__12_), .B(
        mul_ex_mult_86_CARRYB_7__12_), .CI(mul_ex_mult_86_SUMB_7__13_), .CO(
        mul_ex_mult_86_CARRYB_8__12_), .S(mul_ex_mult_86_SUMB_8__12_) );
  FA_X1 mul_ex_mult_86_S2_8_11 ( .A(mul_ex_mult_86_ab_8__11_), .B(
        mul_ex_mult_86_CARRYB_7__11_), .CI(mul_ex_mult_86_SUMB_7__12_), .CO(
        mul_ex_mult_86_CARRYB_8__11_), .S(mul_ex_mult_86_SUMB_8__11_) );
  FA_X1 mul_ex_mult_86_S2_8_10 ( .A(mul_ex_mult_86_ab_8__10_), .B(
        mul_ex_mult_86_CARRYB_7__10_), .CI(mul_ex_mult_86_SUMB_7__11_), .CO(
        mul_ex_mult_86_CARRYB_8__10_), .S(mul_ex_mult_86_SUMB_8__10_) );
  FA_X1 mul_ex_mult_86_S2_8_9 ( .A(mul_ex_mult_86_ab_8__9_), .B(
        mul_ex_mult_86_CARRYB_7__9_), .CI(mul_ex_mult_86_SUMB_7__10_), .CO(
        mul_ex_mult_86_CARRYB_8__9_), .S(mul_ex_mult_86_SUMB_8__9_) );
  FA_X1 mul_ex_mult_86_S2_8_8 ( .A(mul_ex_mult_86_ab_8__8_), .B(
        mul_ex_mult_86_CARRYB_7__8_), .CI(mul_ex_mult_86_SUMB_7__9_), .CO(
        mul_ex_mult_86_CARRYB_8__8_), .S(mul_ex_mult_86_SUMB_8__8_) );
  FA_X1 mul_ex_mult_86_S2_8_7 ( .A(mul_ex_mult_86_ab_8__7_), .B(
        mul_ex_mult_86_CARRYB_7__7_), .CI(mul_ex_mult_86_SUMB_7__8_), .CO(
        mul_ex_mult_86_CARRYB_8__7_), .S(mul_ex_mult_86_SUMB_8__7_) );
  FA_X1 mul_ex_mult_86_S2_8_6 ( .A(mul_ex_mult_86_ab_8__6_), .B(
        mul_ex_mult_86_CARRYB_7__6_), .CI(mul_ex_mult_86_SUMB_7__7_), .CO(
        mul_ex_mult_86_CARRYB_8__6_), .S(mul_ex_mult_86_SUMB_8__6_) );
  FA_X1 mul_ex_mult_86_S2_8_5 ( .A(mul_ex_mult_86_ab_8__5_), .B(
        mul_ex_mult_86_CARRYB_7__5_), .CI(mul_ex_mult_86_SUMB_7__6_), .CO(
        mul_ex_mult_86_CARRYB_8__5_), .S(mul_ex_mult_86_SUMB_8__5_) );
  FA_X1 mul_ex_mult_86_S2_8_4 ( .A(mul_ex_mult_86_ab_8__4_), .B(
        mul_ex_mult_86_CARRYB_7__4_), .CI(mul_ex_mult_86_SUMB_7__5_), .CO(
        mul_ex_mult_86_CARRYB_8__4_), .S(mul_ex_mult_86_SUMB_8__4_) );
  FA_X1 mul_ex_mult_86_S2_8_3 ( .A(mul_ex_mult_86_ab_8__3_), .B(
        mul_ex_mult_86_CARRYB_7__3_), .CI(mul_ex_mult_86_SUMB_7__4_), .CO(
        mul_ex_mult_86_CARRYB_8__3_), .S(mul_ex_mult_86_SUMB_8__3_) );
  FA_X1 mul_ex_mult_86_S2_8_2 ( .A(mul_ex_mult_86_ab_8__2_), .B(
        mul_ex_mult_86_CARRYB_7__2_), .CI(mul_ex_mult_86_SUMB_7__3_), .CO(
        mul_ex_mult_86_CARRYB_8__2_), .S(mul_ex_mult_86_SUMB_8__2_) );
  FA_X1 mul_ex_mult_86_S2_8_1 ( .A(mul_ex_mult_86_ab_8__1_), .B(
        mul_ex_mult_86_CARRYB_7__1_), .CI(mul_ex_mult_86_SUMB_7__2_), .CO(
        mul_ex_mult_86_CARRYB_8__1_), .S(mul_ex_mult_86_SUMB_8__1_) );
  FA_X1 mul_ex_mult_86_S1_8_0 ( .A(mul_ex_mult_86_ab_8__0_), .B(
        mul_ex_mult_86_CARRYB_7__0_), .CI(mul_ex_mult_86_SUMB_7__1_), .CO(
        mul_ex_mult_86_CARRYB_8__0_), .S(mul_ex_mult_86_A1_6_) );
  FA_X1 mul_ex_mult_86_S3_9_14 ( .A(mul_ex_mult_86_ab_9__14_), .B(
        mul_ex_mult_86_CARRYB_8__14_), .CI(mul_ex_mult_86_ab_8__15_), .CO(
        mul_ex_mult_86_CARRYB_9__14_), .S(mul_ex_mult_86_SUMB_9__14_) );
  FA_X1 mul_ex_mult_86_S2_9_13 ( .A(mul_ex_mult_86_ab_9__13_), .B(
        mul_ex_mult_86_CARRYB_8__13_), .CI(mul_ex_mult_86_SUMB_8__14_), .CO(
        mul_ex_mult_86_CARRYB_9__13_), .S(mul_ex_mult_86_SUMB_9__13_) );
  FA_X1 mul_ex_mult_86_S2_9_12 ( .A(mul_ex_mult_86_ab_9__12_), .B(
        mul_ex_mult_86_CARRYB_8__12_), .CI(mul_ex_mult_86_SUMB_8__13_), .CO(
        mul_ex_mult_86_CARRYB_9__12_), .S(mul_ex_mult_86_SUMB_9__12_) );
  FA_X1 mul_ex_mult_86_S2_9_11 ( .A(mul_ex_mult_86_ab_9__11_), .B(
        mul_ex_mult_86_CARRYB_8__11_), .CI(mul_ex_mult_86_SUMB_8__12_), .CO(
        mul_ex_mult_86_CARRYB_9__11_), .S(mul_ex_mult_86_SUMB_9__11_) );
  FA_X1 mul_ex_mult_86_S2_9_10 ( .A(mul_ex_mult_86_ab_9__10_), .B(
        mul_ex_mult_86_CARRYB_8__10_), .CI(mul_ex_mult_86_SUMB_8__11_), .CO(
        mul_ex_mult_86_CARRYB_9__10_), .S(mul_ex_mult_86_SUMB_9__10_) );
  FA_X1 mul_ex_mult_86_S2_9_9 ( .A(mul_ex_mult_86_ab_9__9_), .B(
        mul_ex_mult_86_CARRYB_8__9_), .CI(mul_ex_mult_86_SUMB_8__10_), .CO(
        mul_ex_mult_86_CARRYB_9__9_), .S(mul_ex_mult_86_SUMB_9__9_) );
  FA_X1 mul_ex_mult_86_S2_9_8 ( .A(mul_ex_mult_86_ab_9__8_), .B(
        mul_ex_mult_86_CARRYB_8__8_), .CI(mul_ex_mult_86_SUMB_8__9_), .CO(
        mul_ex_mult_86_CARRYB_9__8_), .S(mul_ex_mult_86_SUMB_9__8_) );
  FA_X1 mul_ex_mult_86_S2_9_7 ( .A(mul_ex_mult_86_ab_9__7_), .B(
        mul_ex_mult_86_CARRYB_8__7_), .CI(mul_ex_mult_86_SUMB_8__8_), .CO(
        mul_ex_mult_86_CARRYB_9__7_), .S(mul_ex_mult_86_SUMB_9__7_) );
  FA_X1 mul_ex_mult_86_S2_9_6 ( .A(mul_ex_mult_86_ab_9__6_), .B(
        mul_ex_mult_86_CARRYB_8__6_), .CI(mul_ex_mult_86_SUMB_8__7_), .CO(
        mul_ex_mult_86_CARRYB_9__6_), .S(mul_ex_mult_86_SUMB_9__6_) );
  FA_X1 mul_ex_mult_86_S2_9_5 ( .A(mul_ex_mult_86_ab_9__5_), .B(
        mul_ex_mult_86_CARRYB_8__5_), .CI(mul_ex_mult_86_SUMB_8__6_), .CO(
        mul_ex_mult_86_CARRYB_9__5_), .S(mul_ex_mult_86_SUMB_9__5_) );
  FA_X1 mul_ex_mult_86_S2_9_4 ( .A(mul_ex_mult_86_ab_9__4_), .B(
        mul_ex_mult_86_CARRYB_8__4_), .CI(mul_ex_mult_86_SUMB_8__5_), .CO(
        mul_ex_mult_86_CARRYB_9__4_), .S(mul_ex_mult_86_SUMB_9__4_) );
  FA_X1 mul_ex_mult_86_S2_9_3 ( .A(mul_ex_mult_86_ab_9__3_), .B(
        mul_ex_mult_86_CARRYB_8__3_), .CI(mul_ex_mult_86_SUMB_8__4_), .CO(
        mul_ex_mult_86_CARRYB_9__3_), .S(mul_ex_mult_86_SUMB_9__3_) );
  FA_X1 mul_ex_mult_86_S2_9_2 ( .A(mul_ex_mult_86_ab_9__2_), .B(
        mul_ex_mult_86_CARRYB_8__2_), .CI(mul_ex_mult_86_SUMB_8__3_), .CO(
        mul_ex_mult_86_CARRYB_9__2_), .S(mul_ex_mult_86_SUMB_9__2_) );
  FA_X1 mul_ex_mult_86_S2_9_1 ( .A(mul_ex_mult_86_ab_9__1_), .B(
        mul_ex_mult_86_CARRYB_8__1_), .CI(mul_ex_mult_86_SUMB_8__2_), .CO(
        mul_ex_mult_86_CARRYB_9__1_), .S(mul_ex_mult_86_SUMB_9__1_) );
  FA_X1 mul_ex_mult_86_S1_9_0 ( .A(mul_ex_mult_86_ab_9__0_), .B(
        mul_ex_mult_86_CARRYB_8__0_), .CI(mul_ex_mult_86_SUMB_8__1_), .CO(
        mul_ex_mult_86_CARRYB_9__0_), .S(mul_ex_mult_86_A1_7_) );
  FA_X1 mul_ex_mult_86_S3_10_14 ( .A(mul_ex_mult_86_ab_10__14_), .B(
        mul_ex_mult_86_CARRYB_9__14_), .CI(mul_ex_mult_86_ab_9__15_), .CO(
        mul_ex_mult_86_CARRYB_10__14_), .S(mul_ex_mult_86_SUMB_10__14_) );
  FA_X1 mul_ex_mult_86_S2_10_13 ( .A(mul_ex_mult_86_ab_10__13_), .B(
        mul_ex_mult_86_CARRYB_9__13_), .CI(mul_ex_mult_86_SUMB_9__14_), .CO(
        mul_ex_mult_86_CARRYB_10__13_), .S(mul_ex_mult_86_SUMB_10__13_) );
  FA_X1 mul_ex_mult_86_S2_10_12 ( .A(mul_ex_mult_86_ab_10__12_), .B(
        mul_ex_mult_86_CARRYB_9__12_), .CI(mul_ex_mult_86_SUMB_9__13_), .CO(
        mul_ex_mult_86_CARRYB_10__12_), .S(mul_ex_mult_86_SUMB_10__12_) );
  FA_X1 mul_ex_mult_86_S2_10_11 ( .A(mul_ex_mult_86_ab_10__11_), .B(
        mul_ex_mult_86_CARRYB_9__11_), .CI(mul_ex_mult_86_SUMB_9__12_), .CO(
        mul_ex_mult_86_CARRYB_10__11_), .S(mul_ex_mult_86_SUMB_10__11_) );
  FA_X1 mul_ex_mult_86_S2_10_10 ( .A(mul_ex_mult_86_ab_10__10_), .B(
        mul_ex_mult_86_CARRYB_9__10_), .CI(mul_ex_mult_86_SUMB_9__11_), .CO(
        mul_ex_mult_86_CARRYB_10__10_), .S(mul_ex_mult_86_SUMB_10__10_) );
  FA_X1 mul_ex_mult_86_S2_10_9 ( .A(mul_ex_mult_86_ab_10__9_), .B(
        mul_ex_mult_86_CARRYB_9__9_), .CI(mul_ex_mult_86_SUMB_9__10_), .CO(
        mul_ex_mult_86_CARRYB_10__9_), .S(mul_ex_mult_86_SUMB_10__9_) );
  FA_X1 mul_ex_mult_86_S2_10_8 ( .A(mul_ex_mult_86_ab_10__8_), .B(
        mul_ex_mult_86_CARRYB_9__8_), .CI(mul_ex_mult_86_SUMB_9__9_), .CO(
        mul_ex_mult_86_CARRYB_10__8_), .S(mul_ex_mult_86_SUMB_10__8_) );
  FA_X1 mul_ex_mult_86_S2_10_7 ( .A(mul_ex_mult_86_ab_10__7_), .B(
        mul_ex_mult_86_CARRYB_9__7_), .CI(mul_ex_mult_86_SUMB_9__8_), .CO(
        mul_ex_mult_86_CARRYB_10__7_), .S(mul_ex_mult_86_SUMB_10__7_) );
  FA_X1 mul_ex_mult_86_S2_10_6 ( .A(mul_ex_mult_86_ab_10__6_), .B(
        mul_ex_mult_86_CARRYB_9__6_), .CI(mul_ex_mult_86_SUMB_9__7_), .CO(
        mul_ex_mult_86_CARRYB_10__6_), .S(mul_ex_mult_86_SUMB_10__6_) );
  FA_X1 mul_ex_mult_86_S2_10_5 ( .A(mul_ex_mult_86_ab_10__5_), .B(
        mul_ex_mult_86_CARRYB_9__5_), .CI(mul_ex_mult_86_SUMB_9__6_), .CO(
        mul_ex_mult_86_CARRYB_10__5_), .S(mul_ex_mult_86_SUMB_10__5_) );
  FA_X1 mul_ex_mult_86_S2_10_4 ( .A(mul_ex_mult_86_ab_10__4_), .B(
        mul_ex_mult_86_CARRYB_9__4_), .CI(mul_ex_mult_86_SUMB_9__5_), .CO(
        mul_ex_mult_86_CARRYB_10__4_), .S(mul_ex_mult_86_SUMB_10__4_) );
  FA_X1 mul_ex_mult_86_S2_10_3 ( .A(mul_ex_mult_86_ab_10__3_), .B(
        mul_ex_mult_86_CARRYB_9__3_), .CI(mul_ex_mult_86_SUMB_9__4_), .CO(
        mul_ex_mult_86_CARRYB_10__3_), .S(mul_ex_mult_86_SUMB_10__3_) );
  FA_X1 mul_ex_mult_86_S2_10_2 ( .A(mul_ex_mult_86_ab_10__2_), .B(
        mul_ex_mult_86_CARRYB_9__2_), .CI(mul_ex_mult_86_SUMB_9__3_), .CO(
        mul_ex_mult_86_CARRYB_10__2_), .S(mul_ex_mult_86_SUMB_10__2_) );
  FA_X1 mul_ex_mult_86_S2_10_1 ( .A(mul_ex_mult_86_ab_10__1_), .B(
        mul_ex_mult_86_CARRYB_9__1_), .CI(mul_ex_mult_86_SUMB_9__2_), .CO(
        mul_ex_mult_86_CARRYB_10__1_), .S(mul_ex_mult_86_SUMB_10__1_) );
  FA_X1 mul_ex_mult_86_S1_10_0 ( .A(mul_ex_mult_86_ab_10__0_), .B(
        mul_ex_mult_86_CARRYB_9__0_), .CI(mul_ex_mult_86_SUMB_9__1_), .CO(
        mul_ex_mult_86_CARRYB_10__0_), .S(mul_ex_mult_86_A1_8_) );
  FA_X1 mul_ex_mult_86_S3_11_14 ( .A(mul_ex_mult_86_ab_11__14_), .B(
        mul_ex_mult_86_CARRYB_10__14_), .CI(mul_ex_mult_86_ab_10__15_), .CO(
        mul_ex_mult_86_CARRYB_11__14_), .S(mul_ex_mult_86_SUMB_11__14_) );
  FA_X1 mul_ex_mult_86_S2_11_13 ( .A(mul_ex_mult_86_ab_11__13_), .B(
        mul_ex_mult_86_CARRYB_10__13_), .CI(mul_ex_mult_86_SUMB_10__14_), .CO(
        mul_ex_mult_86_CARRYB_11__13_), .S(mul_ex_mult_86_SUMB_11__13_) );
  FA_X1 mul_ex_mult_86_S2_11_12 ( .A(mul_ex_mult_86_ab_11__12_), .B(
        mul_ex_mult_86_CARRYB_10__12_), .CI(mul_ex_mult_86_SUMB_10__13_), .CO(
        mul_ex_mult_86_CARRYB_11__12_), .S(mul_ex_mult_86_SUMB_11__12_) );
  FA_X1 mul_ex_mult_86_S2_11_11 ( .A(mul_ex_mult_86_ab_11__11_), .B(
        mul_ex_mult_86_CARRYB_10__11_), .CI(mul_ex_mult_86_SUMB_10__12_), .CO(
        mul_ex_mult_86_CARRYB_11__11_), .S(mul_ex_mult_86_SUMB_11__11_) );
  FA_X1 mul_ex_mult_86_S2_11_10 ( .A(mul_ex_mult_86_ab_11__10_), .B(
        mul_ex_mult_86_CARRYB_10__10_), .CI(mul_ex_mult_86_SUMB_10__11_), .CO(
        mul_ex_mult_86_CARRYB_11__10_), .S(mul_ex_mult_86_SUMB_11__10_) );
  FA_X1 mul_ex_mult_86_S2_11_9 ( .A(mul_ex_mult_86_ab_11__9_), .B(
        mul_ex_mult_86_CARRYB_10__9_), .CI(mul_ex_mult_86_SUMB_10__10_), .CO(
        mul_ex_mult_86_CARRYB_11__9_), .S(mul_ex_mult_86_SUMB_11__9_) );
  FA_X1 mul_ex_mult_86_S2_11_8 ( .A(mul_ex_mult_86_ab_11__8_), .B(
        mul_ex_mult_86_CARRYB_10__8_), .CI(mul_ex_mult_86_SUMB_10__9_), .CO(
        mul_ex_mult_86_CARRYB_11__8_), .S(mul_ex_mult_86_SUMB_11__8_) );
  FA_X1 mul_ex_mult_86_S2_11_7 ( .A(mul_ex_mult_86_ab_11__7_), .B(
        mul_ex_mult_86_CARRYB_10__7_), .CI(mul_ex_mult_86_SUMB_10__8_), .CO(
        mul_ex_mult_86_CARRYB_11__7_), .S(mul_ex_mult_86_SUMB_11__7_) );
  FA_X1 mul_ex_mult_86_S2_11_6 ( .A(mul_ex_mult_86_ab_11__6_), .B(
        mul_ex_mult_86_CARRYB_10__6_), .CI(mul_ex_mult_86_SUMB_10__7_), .CO(
        mul_ex_mult_86_CARRYB_11__6_), .S(mul_ex_mult_86_SUMB_11__6_) );
  FA_X1 mul_ex_mult_86_S2_11_5 ( .A(mul_ex_mult_86_ab_11__5_), .B(
        mul_ex_mult_86_CARRYB_10__5_), .CI(mul_ex_mult_86_SUMB_10__6_), .CO(
        mul_ex_mult_86_CARRYB_11__5_), .S(mul_ex_mult_86_SUMB_11__5_) );
  FA_X1 mul_ex_mult_86_S2_11_4 ( .A(mul_ex_mult_86_ab_11__4_), .B(
        mul_ex_mult_86_CARRYB_10__4_), .CI(mul_ex_mult_86_SUMB_10__5_), .CO(
        mul_ex_mult_86_CARRYB_11__4_), .S(mul_ex_mult_86_SUMB_11__4_) );
  FA_X1 mul_ex_mult_86_S2_11_3 ( .A(mul_ex_mult_86_ab_11__3_), .B(
        mul_ex_mult_86_CARRYB_10__3_), .CI(mul_ex_mult_86_SUMB_10__4_), .CO(
        mul_ex_mult_86_CARRYB_11__3_), .S(mul_ex_mult_86_SUMB_11__3_) );
  FA_X1 mul_ex_mult_86_S2_11_2 ( .A(mul_ex_mult_86_ab_11__2_), .B(
        mul_ex_mult_86_CARRYB_10__2_), .CI(mul_ex_mult_86_SUMB_10__3_), .CO(
        mul_ex_mult_86_CARRYB_11__2_), .S(mul_ex_mult_86_SUMB_11__2_) );
  FA_X1 mul_ex_mult_86_S2_11_1 ( .A(mul_ex_mult_86_ab_11__1_), .B(
        mul_ex_mult_86_CARRYB_10__1_), .CI(mul_ex_mult_86_SUMB_10__2_), .CO(
        mul_ex_mult_86_CARRYB_11__1_), .S(mul_ex_mult_86_SUMB_11__1_) );
  FA_X1 mul_ex_mult_86_S1_11_0 ( .A(mul_ex_mult_86_ab_11__0_), .B(
        mul_ex_mult_86_CARRYB_10__0_), .CI(mul_ex_mult_86_SUMB_10__1_), .CO(
        mul_ex_mult_86_CARRYB_11__0_), .S(mul_ex_mult_86_A1_9_) );
  FA_X1 mul_ex_mult_86_S3_12_14 ( .A(mul_ex_mult_86_ab_12__14_), .B(
        mul_ex_mult_86_CARRYB_11__14_), .CI(mul_ex_mult_86_ab_11__15_), .CO(
        mul_ex_mult_86_CARRYB_12__14_), .S(mul_ex_mult_86_SUMB_12__14_) );
  FA_X1 mul_ex_mult_86_S2_12_13 ( .A(mul_ex_mult_86_ab_12__13_), .B(
        mul_ex_mult_86_CARRYB_11__13_), .CI(mul_ex_mult_86_SUMB_11__14_), .CO(
        mul_ex_mult_86_CARRYB_12__13_), .S(mul_ex_mult_86_SUMB_12__13_) );
  FA_X1 mul_ex_mult_86_S2_12_12 ( .A(mul_ex_mult_86_ab_12__12_), .B(
        mul_ex_mult_86_CARRYB_11__12_), .CI(mul_ex_mult_86_SUMB_11__13_), .CO(
        mul_ex_mult_86_CARRYB_12__12_), .S(mul_ex_mult_86_SUMB_12__12_) );
  FA_X1 mul_ex_mult_86_S2_12_11 ( .A(mul_ex_mult_86_ab_12__11_), .B(
        mul_ex_mult_86_CARRYB_11__11_), .CI(mul_ex_mult_86_SUMB_11__12_), .CO(
        mul_ex_mult_86_CARRYB_12__11_), .S(mul_ex_mult_86_SUMB_12__11_) );
  FA_X1 mul_ex_mult_86_S2_12_10 ( .A(mul_ex_mult_86_ab_12__10_), .B(
        mul_ex_mult_86_CARRYB_11__10_), .CI(mul_ex_mult_86_SUMB_11__11_), .CO(
        mul_ex_mult_86_CARRYB_12__10_), .S(mul_ex_mult_86_SUMB_12__10_) );
  FA_X1 mul_ex_mult_86_S2_12_9 ( .A(mul_ex_mult_86_ab_12__9_), .B(
        mul_ex_mult_86_CARRYB_11__9_), .CI(mul_ex_mult_86_SUMB_11__10_), .CO(
        mul_ex_mult_86_CARRYB_12__9_), .S(mul_ex_mult_86_SUMB_12__9_) );
  FA_X1 mul_ex_mult_86_S2_12_8 ( .A(mul_ex_mult_86_ab_12__8_), .B(
        mul_ex_mult_86_CARRYB_11__8_), .CI(mul_ex_mult_86_SUMB_11__9_), .CO(
        mul_ex_mult_86_CARRYB_12__8_), .S(mul_ex_mult_86_SUMB_12__8_) );
  FA_X1 mul_ex_mult_86_S2_12_7 ( .A(mul_ex_mult_86_ab_12__7_), .B(
        mul_ex_mult_86_CARRYB_11__7_), .CI(mul_ex_mult_86_SUMB_11__8_), .CO(
        mul_ex_mult_86_CARRYB_12__7_), .S(mul_ex_mult_86_SUMB_12__7_) );
  FA_X1 mul_ex_mult_86_S2_12_6 ( .A(mul_ex_mult_86_ab_12__6_), .B(
        mul_ex_mult_86_CARRYB_11__6_), .CI(mul_ex_mult_86_SUMB_11__7_), .CO(
        mul_ex_mult_86_CARRYB_12__6_), .S(mul_ex_mult_86_SUMB_12__6_) );
  FA_X1 mul_ex_mult_86_S2_12_5 ( .A(mul_ex_mult_86_ab_12__5_), .B(
        mul_ex_mult_86_CARRYB_11__5_), .CI(mul_ex_mult_86_SUMB_11__6_), .CO(
        mul_ex_mult_86_CARRYB_12__5_), .S(mul_ex_mult_86_SUMB_12__5_) );
  FA_X1 mul_ex_mult_86_S2_12_4 ( .A(mul_ex_mult_86_ab_12__4_), .B(
        mul_ex_mult_86_CARRYB_11__4_), .CI(mul_ex_mult_86_SUMB_11__5_), .CO(
        mul_ex_mult_86_CARRYB_12__4_), .S(mul_ex_mult_86_SUMB_12__4_) );
  FA_X1 mul_ex_mult_86_S2_12_3 ( .A(mul_ex_mult_86_ab_12__3_), .B(
        mul_ex_mult_86_CARRYB_11__3_), .CI(mul_ex_mult_86_SUMB_11__4_), .CO(
        mul_ex_mult_86_CARRYB_12__3_), .S(mul_ex_mult_86_SUMB_12__3_) );
  FA_X1 mul_ex_mult_86_S2_12_2 ( .A(mul_ex_mult_86_ab_12__2_), .B(
        mul_ex_mult_86_CARRYB_11__2_), .CI(mul_ex_mult_86_SUMB_11__3_), .CO(
        mul_ex_mult_86_CARRYB_12__2_), .S(mul_ex_mult_86_SUMB_12__2_) );
  FA_X1 mul_ex_mult_86_S2_12_1 ( .A(mul_ex_mult_86_ab_12__1_), .B(
        mul_ex_mult_86_CARRYB_11__1_), .CI(mul_ex_mult_86_SUMB_11__2_), .CO(
        mul_ex_mult_86_CARRYB_12__1_), .S(mul_ex_mult_86_SUMB_12__1_) );
  FA_X1 mul_ex_mult_86_S1_12_0 ( .A(mul_ex_mult_86_ab_12__0_), .B(
        mul_ex_mult_86_CARRYB_11__0_), .CI(mul_ex_mult_86_SUMB_11__1_), .CO(
        mul_ex_mult_86_CARRYB_12__0_), .S(mul_ex_mult_86_A1_10_) );
  FA_X1 mul_ex_mult_86_S3_13_14 ( .A(mul_ex_mult_86_ab_13__14_), .B(
        mul_ex_mult_86_CARRYB_12__14_), .CI(mul_ex_mult_86_ab_12__15_), .CO(
        mul_ex_mult_86_CARRYB_13__14_), .S(mul_ex_mult_86_SUMB_13__14_) );
  FA_X1 mul_ex_mult_86_S2_13_13 ( .A(mul_ex_mult_86_ab_13__13_), .B(
        mul_ex_mult_86_CARRYB_12__13_), .CI(mul_ex_mult_86_SUMB_12__14_), .CO(
        mul_ex_mult_86_CARRYB_13__13_), .S(mul_ex_mult_86_SUMB_13__13_) );
  FA_X1 mul_ex_mult_86_S2_13_12 ( .A(mul_ex_mult_86_ab_13__12_), .B(
        mul_ex_mult_86_CARRYB_12__12_), .CI(mul_ex_mult_86_SUMB_12__13_), .CO(
        mul_ex_mult_86_CARRYB_13__12_), .S(mul_ex_mult_86_SUMB_13__12_) );
  FA_X1 mul_ex_mult_86_S2_13_11 ( .A(mul_ex_mult_86_ab_13__11_), .B(
        mul_ex_mult_86_CARRYB_12__11_), .CI(mul_ex_mult_86_SUMB_12__12_), .CO(
        mul_ex_mult_86_CARRYB_13__11_), .S(mul_ex_mult_86_SUMB_13__11_) );
  FA_X1 mul_ex_mult_86_S2_13_10 ( .A(mul_ex_mult_86_ab_13__10_), .B(
        mul_ex_mult_86_CARRYB_12__10_), .CI(mul_ex_mult_86_SUMB_12__11_), .CO(
        mul_ex_mult_86_CARRYB_13__10_), .S(mul_ex_mult_86_SUMB_13__10_) );
  FA_X1 mul_ex_mult_86_S2_13_9 ( .A(mul_ex_mult_86_ab_13__9_), .B(
        mul_ex_mult_86_CARRYB_12__9_), .CI(mul_ex_mult_86_SUMB_12__10_), .CO(
        mul_ex_mult_86_CARRYB_13__9_), .S(mul_ex_mult_86_SUMB_13__9_) );
  FA_X1 mul_ex_mult_86_S2_13_8 ( .A(mul_ex_mult_86_ab_13__8_), .B(
        mul_ex_mult_86_CARRYB_12__8_), .CI(mul_ex_mult_86_SUMB_12__9_), .CO(
        mul_ex_mult_86_CARRYB_13__8_), .S(mul_ex_mult_86_SUMB_13__8_) );
  FA_X1 mul_ex_mult_86_S2_13_7 ( .A(mul_ex_mult_86_ab_13__7_), .B(
        mul_ex_mult_86_CARRYB_12__7_), .CI(mul_ex_mult_86_SUMB_12__8_), .CO(
        mul_ex_mult_86_CARRYB_13__7_), .S(mul_ex_mult_86_SUMB_13__7_) );
  FA_X1 mul_ex_mult_86_S2_13_6 ( .A(mul_ex_mult_86_ab_13__6_), .B(
        mul_ex_mult_86_CARRYB_12__6_), .CI(mul_ex_mult_86_SUMB_12__7_), .CO(
        mul_ex_mult_86_CARRYB_13__6_), .S(mul_ex_mult_86_SUMB_13__6_) );
  FA_X1 mul_ex_mult_86_S2_13_5 ( .A(mul_ex_mult_86_ab_13__5_), .B(
        mul_ex_mult_86_CARRYB_12__5_), .CI(mul_ex_mult_86_SUMB_12__6_), .CO(
        mul_ex_mult_86_CARRYB_13__5_), .S(mul_ex_mult_86_SUMB_13__5_) );
  FA_X1 mul_ex_mult_86_S2_13_4 ( .A(mul_ex_mult_86_ab_13__4_), .B(
        mul_ex_mult_86_CARRYB_12__4_), .CI(mul_ex_mult_86_SUMB_12__5_), .CO(
        mul_ex_mult_86_CARRYB_13__4_), .S(mul_ex_mult_86_SUMB_13__4_) );
  FA_X1 mul_ex_mult_86_S2_13_3 ( .A(mul_ex_mult_86_ab_13__3_), .B(
        mul_ex_mult_86_CARRYB_12__3_), .CI(mul_ex_mult_86_SUMB_12__4_), .CO(
        mul_ex_mult_86_CARRYB_13__3_), .S(mul_ex_mult_86_SUMB_13__3_) );
  FA_X1 mul_ex_mult_86_S2_13_2 ( .A(mul_ex_mult_86_ab_13__2_), .B(
        mul_ex_mult_86_CARRYB_12__2_), .CI(mul_ex_mult_86_SUMB_12__3_), .CO(
        mul_ex_mult_86_CARRYB_13__2_), .S(mul_ex_mult_86_SUMB_13__2_) );
  FA_X1 mul_ex_mult_86_S2_13_1 ( .A(mul_ex_mult_86_ab_13__1_), .B(
        mul_ex_mult_86_CARRYB_12__1_), .CI(mul_ex_mult_86_SUMB_12__2_), .CO(
        mul_ex_mult_86_CARRYB_13__1_), .S(mul_ex_mult_86_SUMB_13__1_) );
  FA_X1 mul_ex_mult_86_S1_13_0 ( .A(mul_ex_mult_86_ab_13__0_), .B(
        mul_ex_mult_86_CARRYB_12__0_), .CI(mul_ex_mult_86_SUMB_12__1_), .CO(
        mul_ex_mult_86_CARRYB_13__0_), .S(mul_ex_mult_86_A1_11_) );
  FA_X1 mul_ex_mult_86_S3_14_14 ( .A(mul_ex_mult_86_ab_14__14_), .B(
        mul_ex_mult_86_CARRYB_13__14_), .CI(mul_ex_mult_86_ab_13__15_), .CO(
        mul_ex_mult_86_CARRYB_14__14_), .S(mul_ex_mult_86_SUMB_14__14_) );
  FA_X1 mul_ex_mult_86_S2_14_13 ( .A(mul_ex_mult_86_ab_14__13_), .B(
        mul_ex_mult_86_CARRYB_13__13_), .CI(mul_ex_mult_86_SUMB_13__14_), .CO(
        mul_ex_mult_86_CARRYB_14__13_), .S(mul_ex_mult_86_SUMB_14__13_) );
  FA_X1 mul_ex_mult_86_S2_14_12 ( .A(mul_ex_mult_86_ab_14__12_), .B(
        mul_ex_mult_86_CARRYB_13__12_), .CI(mul_ex_mult_86_SUMB_13__13_), .CO(
        mul_ex_mult_86_CARRYB_14__12_), .S(mul_ex_mult_86_SUMB_14__12_) );
  FA_X1 mul_ex_mult_86_S2_14_11 ( .A(mul_ex_mult_86_ab_14__11_), .B(
        mul_ex_mult_86_CARRYB_13__11_), .CI(mul_ex_mult_86_SUMB_13__12_), .CO(
        mul_ex_mult_86_CARRYB_14__11_), .S(mul_ex_mult_86_SUMB_14__11_) );
  FA_X1 mul_ex_mult_86_S2_14_10 ( .A(mul_ex_mult_86_ab_14__10_), .B(
        mul_ex_mult_86_CARRYB_13__10_), .CI(mul_ex_mult_86_SUMB_13__11_), .CO(
        mul_ex_mult_86_CARRYB_14__10_), .S(mul_ex_mult_86_SUMB_14__10_) );
  FA_X1 mul_ex_mult_86_S2_14_9 ( .A(mul_ex_mult_86_ab_14__9_), .B(
        mul_ex_mult_86_CARRYB_13__9_), .CI(mul_ex_mult_86_SUMB_13__10_), .CO(
        mul_ex_mult_86_CARRYB_14__9_), .S(mul_ex_mult_86_SUMB_14__9_) );
  FA_X1 mul_ex_mult_86_S2_14_8 ( .A(mul_ex_mult_86_ab_14__8_), .B(
        mul_ex_mult_86_CARRYB_13__8_), .CI(mul_ex_mult_86_SUMB_13__9_), .CO(
        mul_ex_mult_86_CARRYB_14__8_), .S(mul_ex_mult_86_SUMB_14__8_) );
  FA_X1 mul_ex_mult_86_S2_14_7 ( .A(mul_ex_mult_86_ab_14__7_), .B(
        mul_ex_mult_86_CARRYB_13__7_), .CI(mul_ex_mult_86_SUMB_13__8_), .CO(
        mul_ex_mult_86_CARRYB_14__7_), .S(mul_ex_mult_86_SUMB_14__7_) );
  FA_X1 mul_ex_mult_86_S2_14_6 ( .A(mul_ex_mult_86_ab_14__6_), .B(
        mul_ex_mult_86_CARRYB_13__6_), .CI(mul_ex_mult_86_SUMB_13__7_), .CO(
        mul_ex_mult_86_CARRYB_14__6_), .S(mul_ex_mult_86_SUMB_14__6_) );
  FA_X1 mul_ex_mult_86_S2_14_5 ( .A(mul_ex_mult_86_ab_14__5_), .B(
        mul_ex_mult_86_CARRYB_13__5_), .CI(mul_ex_mult_86_SUMB_13__6_), .CO(
        mul_ex_mult_86_CARRYB_14__5_), .S(mul_ex_mult_86_SUMB_14__5_) );
  FA_X1 mul_ex_mult_86_S2_14_4 ( .A(mul_ex_mult_86_ab_14__4_), .B(
        mul_ex_mult_86_CARRYB_13__4_), .CI(mul_ex_mult_86_SUMB_13__5_), .CO(
        mul_ex_mult_86_CARRYB_14__4_), .S(mul_ex_mult_86_SUMB_14__4_) );
  FA_X1 mul_ex_mult_86_S2_14_3 ( .A(mul_ex_mult_86_ab_14__3_), .B(
        mul_ex_mult_86_CARRYB_13__3_), .CI(mul_ex_mult_86_SUMB_13__4_), .CO(
        mul_ex_mult_86_CARRYB_14__3_), .S(mul_ex_mult_86_SUMB_14__3_) );
  FA_X1 mul_ex_mult_86_S2_14_2 ( .A(mul_ex_mult_86_ab_14__2_), .B(
        mul_ex_mult_86_CARRYB_13__2_), .CI(mul_ex_mult_86_SUMB_13__3_), .CO(
        mul_ex_mult_86_CARRYB_14__2_), .S(mul_ex_mult_86_SUMB_14__2_) );
  FA_X1 mul_ex_mult_86_S2_14_1 ( .A(mul_ex_mult_86_ab_14__1_), .B(
        mul_ex_mult_86_CARRYB_13__1_), .CI(mul_ex_mult_86_SUMB_13__2_), .CO(
        mul_ex_mult_86_CARRYB_14__1_), .S(mul_ex_mult_86_SUMB_14__1_) );
  FA_X1 mul_ex_mult_86_S1_14_0 ( .A(mul_ex_mult_86_ab_14__0_), .B(
        mul_ex_mult_86_CARRYB_13__0_), .CI(mul_ex_mult_86_SUMB_13__1_), .CO(
        mul_ex_mult_86_CARRYB_14__0_), .S(mul_ex_mult_86_A1_12_) );
  FA_X1 mul_ex_mult_86_S5_14 ( .A(mul_ex_mult_86_ab_15__14_), .B(
        mul_ex_mult_86_CARRYB_14__14_), .CI(mul_ex_mult_86_ab_14__15_), .CO(
        mul_ex_mult_86_CARRYB_15__14_), .S(mul_ex_mult_86_SUMB_15__14_) );
  FA_X1 mul_ex_mult_86_S4_13 ( .A(mul_ex_mult_86_ab_15__13_), .B(
        mul_ex_mult_86_CARRYB_14__13_), .CI(mul_ex_mult_86_SUMB_14__14_), .CO(
        mul_ex_mult_86_CARRYB_15__13_), .S(mul_ex_mult_86_SUMB_15__13_) );
  FA_X1 mul_ex_mult_86_S4_12 ( .A(mul_ex_mult_86_ab_15__12_), .B(
        mul_ex_mult_86_CARRYB_14__12_), .CI(mul_ex_mult_86_SUMB_14__13_), .CO(
        mul_ex_mult_86_CARRYB_15__12_), .S(mul_ex_mult_86_SUMB_15__12_) );
  FA_X1 mul_ex_mult_86_S4_11 ( .A(mul_ex_mult_86_ab_15__11_), .B(
        mul_ex_mult_86_CARRYB_14__11_), .CI(mul_ex_mult_86_SUMB_14__12_), .CO(
        mul_ex_mult_86_CARRYB_15__11_), .S(mul_ex_mult_86_SUMB_15__11_) );
  FA_X1 mul_ex_mult_86_S4_10 ( .A(mul_ex_mult_86_ab_15__10_), .B(
        mul_ex_mult_86_CARRYB_14__10_), .CI(mul_ex_mult_86_SUMB_14__11_), .CO(
        mul_ex_mult_86_CARRYB_15__10_), .S(mul_ex_mult_86_SUMB_15__10_) );
  FA_X1 mul_ex_mult_86_S4_9 ( .A(mul_ex_mult_86_ab_15__9_), .B(
        mul_ex_mult_86_CARRYB_14__9_), .CI(mul_ex_mult_86_SUMB_14__10_), .CO(
        mul_ex_mult_86_CARRYB_15__9_), .S(mul_ex_mult_86_SUMB_15__9_) );
  FA_X1 mul_ex_mult_86_S4_8 ( .A(mul_ex_mult_86_ab_15__8_), .B(
        mul_ex_mult_86_CARRYB_14__8_), .CI(mul_ex_mult_86_SUMB_14__9_), .CO(
        mul_ex_mult_86_CARRYB_15__8_), .S(mul_ex_mult_86_SUMB_15__8_) );
  FA_X1 mul_ex_mult_86_S4_7 ( .A(mul_ex_mult_86_ab_15__7_), .B(
        mul_ex_mult_86_CARRYB_14__7_), .CI(mul_ex_mult_86_SUMB_14__8_), .CO(
        mul_ex_mult_86_CARRYB_15__7_), .S(mul_ex_mult_86_SUMB_15__7_) );
  FA_X1 mul_ex_mult_86_S4_6 ( .A(mul_ex_mult_86_ab_15__6_), .B(
        mul_ex_mult_86_CARRYB_14__6_), .CI(mul_ex_mult_86_SUMB_14__7_), .CO(
        mul_ex_mult_86_CARRYB_15__6_), .S(mul_ex_mult_86_SUMB_15__6_) );
  FA_X1 mul_ex_mult_86_S4_5 ( .A(mul_ex_mult_86_ab_15__5_), .B(
        mul_ex_mult_86_CARRYB_14__5_), .CI(mul_ex_mult_86_SUMB_14__6_), .CO(
        mul_ex_mult_86_CARRYB_15__5_), .S(mul_ex_mult_86_SUMB_15__5_) );
  FA_X1 mul_ex_mult_86_S4_4 ( .A(mul_ex_mult_86_ab_15__4_), .B(
        mul_ex_mult_86_CARRYB_14__4_), .CI(mul_ex_mult_86_SUMB_14__5_), .CO(
        mul_ex_mult_86_CARRYB_15__4_), .S(mul_ex_mult_86_SUMB_15__4_) );
  FA_X1 mul_ex_mult_86_S4_3 ( .A(mul_ex_mult_86_ab_15__3_), .B(
        mul_ex_mult_86_CARRYB_14__3_), .CI(mul_ex_mult_86_SUMB_14__4_), .CO(
        mul_ex_mult_86_CARRYB_15__3_), .S(mul_ex_mult_86_SUMB_15__3_) );
  FA_X1 mul_ex_mult_86_S4_2 ( .A(mul_ex_mult_86_ab_15__2_), .B(
        mul_ex_mult_86_CARRYB_14__2_), .CI(mul_ex_mult_86_SUMB_14__3_), .CO(
        mul_ex_mult_86_CARRYB_15__2_), .S(mul_ex_mult_86_SUMB_15__2_) );
  FA_X1 mul_ex_mult_86_S4_1 ( .A(mul_ex_mult_86_ab_15__1_), .B(
        mul_ex_mult_86_CARRYB_14__1_), .CI(mul_ex_mult_86_SUMB_14__2_), .CO(
        mul_ex_mult_86_CARRYB_15__1_), .S(mul_ex_mult_86_SUMB_15__1_) );
  FA_X1 mul_ex_mult_86_S4_0 ( .A(mul_ex_mult_86_ab_15__0_), .B(
        mul_ex_mult_86_CARRYB_14__0_), .CI(mul_ex_mult_86_SUMB_14__1_), .CO(
        mul_ex_mult_86_CARRYB_15__0_), .S(mul_ex_mult_86_SUMB_15__0_) );
  BUF_X32 mul_ex_mult_86_FS_1_U100 ( .A(mul_ex_mult_86_n61), .Z(mul_ex_N138)
         );
  BUF_X32 mul_ex_mult_86_FS_1_U99 ( .A(mul_ex_mult_86_SUMB_15__0_), .Z(
        mul_ex_N137) );
  BUF_X32 mul_ex_mult_86_FS_1_U98 ( .A(mul_ex_mult_86_A1_12_), .Z(mul_ex_N136)
         );
  BUF_X32 mul_ex_mult_86_FS_1_U97 ( .A(mul_ex_mult_86_A1_11_), .Z(mul_ex_N135)
         );
  BUF_X32 mul_ex_mult_86_FS_1_U96 ( .A(mul_ex_mult_86_A1_10_), .Z(mul_ex_N134)
         );
  BUF_X4 mul_ex_mult_86_FS_1_U95 ( .A(mul_ex_mult_86_A1_0_), .Z(mul_ex_N124)
         );
  BUF_X4 mul_ex_mult_86_FS_1_U94 ( .A(mul_ex_mult_86_A1_1_), .Z(mul_ex_N125)
         );
  BUF_X4 mul_ex_mult_86_FS_1_U93 ( .A(mul_ex_mult_86_A1_2_), .Z(mul_ex_N126)
         );
  BUF_X4 mul_ex_mult_86_FS_1_U92 ( .A(mul_ex_mult_86_A1_3_), .Z(mul_ex_N127)
         );
  BUF_X4 mul_ex_mult_86_FS_1_U91 ( .A(mul_ex_mult_86_A1_4_), .Z(mul_ex_N128)
         );
  BUF_X4 mul_ex_mult_86_FS_1_U90 ( .A(mul_ex_mult_86_A1_5_), .Z(mul_ex_N129)
         );
  BUF_X4 mul_ex_mult_86_FS_1_U89 ( .A(mul_ex_mult_86_A1_6_), .Z(mul_ex_N130)
         );
  BUF_X4 mul_ex_mult_86_FS_1_U88 ( .A(mul_ex_mult_86_A1_7_), .Z(mul_ex_N131)
         );
  BUF_X4 mul_ex_mult_86_FS_1_U87 ( .A(mul_ex_mult_86_A1_8_), .Z(mul_ex_N132)
         );
  BUF_X4 mul_ex_mult_86_FS_1_U86 ( .A(mul_ex_mult_86_A1_9_), .Z(mul_ex_N133)
         );
  NAND2_X1 mul_ex_mult_86_FS_1_U85 ( .A1(mul_ex_mult_86_n59), .A2(
        mul_ex_mult_86_n24), .ZN(mul_ex_mult_86_FS_1_n70) );
  AND2_X1 mul_ex_mult_86_FS_1_U84 ( .A1(mul_ex_mult_86_n52), .A2(
        mul_ex_mult_86_n23), .ZN(mul_ex_mult_86_FS_1_n67) );
  NOR2_X1 mul_ex_mult_86_FS_1_U83 ( .A1(mul_ex_mult_86_n52), .A2(
        mul_ex_mult_86_n23), .ZN(mul_ex_mult_86_FS_1_n68) );
  NOR2_X1 mul_ex_mult_86_FS_1_U82 ( .A1(mul_ex_mult_86_FS_1_n67), .A2(
        mul_ex_mult_86_FS_1_n68), .ZN(mul_ex_mult_86_FS_1_n69) );
  XOR2_X1 mul_ex_mult_86_FS_1_U81 ( .A(mul_ex_mult_86_FS_1_n17), .B(
        mul_ex_mult_86_FS_1_n69), .Z(mul_ex_N140) );
  NOR2_X1 mul_ex_mult_86_FS_1_U80 ( .A1(mul_ex_mult_86_n58), .A2(
        mul_ex_mult_86_n30), .ZN(mul_ex_mult_86_FS_1_n63) );
  NAND2_X1 mul_ex_mult_86_FS_1_U79 ( .A1(mul_ex_mult_86_n58), .A2(
        mul_ex_mult_86_n30), .ZN(mul_ex_mult_86_FS_1_n65) );
  NAND2_X1 mul_ex_mult_86_FS_1_U78 ( .A1(mul_ex_mult_86_FS_1_n15), .A2(
        mul_ex_mult_86_FS_1_n65), .ZN(mul_ex_mult_86_FS_1_n66) );
  AOI21_X1 mul_ex_mult_86_FS_1_U77 ( .B1(mul_ex_mult_86_FS_1_n16), .B2(
        mul_ex_mult_86_FS_1_n17), .A(mul_ex_mult_86_FS_1_n67), .ZN(
        mul_ex_mult_86_FS_1_n64) );
  XOR2_X1 mul_ex_mult_86_FS_1_U76 ( .A(mul_ex_mult_86_FS_1_n66), .B(
        mul_ex_mult_86_FS_1_n64), .Z(mul_ex_N141) );
  OAI21_X1 mul_ex_mult_86_FS_1_U75 ( .B1(mul_ex_mult_86_FS_1_n63), .B2(
        mul_ex_mult_86_FS_1_n64), .A(mul_ex_mult_86_FS_1_n65), .ZN(
        mul_ex_mult_86_FS_1_n59) );
  AND2_X1 mul_ex_mult_86_FS_1_U74 ( .A1(mul_ex_mult_86_n51), .A2(
        mul_ex_mult_86_n22), .ZN(mul_ex_mult_86_FS_1_n60) );
  NOR2_X1 mul_ex_mult_86_FS_1_U73 ( .A1(mul_ex_mult_86_n51), .A2(
        mul_ex_mult_86_n22), .ZN(mul_ex_mult_86_FS_1_n61) );
  NOR2_X1 mul_ex_mult_86_FS_1_U72 ( .A1(mul_ex_mult_86_FS_1_n60), .A2(
        mul_ex_mult_86_FS_1_n61), .ZN(mul_ex_mult_86_FS_1_n62) );
  XOR2_X1 mul_ex_mult_86_FS_1_U71 ( .A(mul_ex_mult_86_FS_1_n59), .B(
        mul_ex_mult_86_FS_1_n62), .Z(mul_ex_N142) );
  NOR2_X1 mul_ex_mult_86_FS_1_U70 ( .A1(mul_ex_mult_86_n57), .A2(
        mul_ex_mult_86_n29), .ZN(mul_ex_mult_86_FS_1_n55) );
  NAND2_X1 mul_ex_mult_86_FS_1_U69 ( .A1(mul_ex_mult_86_n57), .A2(
        mul_ex_mult_86_n29), .ZN(mul_ex_mult_86_FS_1_n57) );
  NAND2_X1 mul_ex_mult_86_FS_1_U68 ( .A1(mul_ex_mult_86_FS_1_n13), .A2(
        mul_ex_mult_86_FS_1_n57), .ZN(mul_ex_mult_86_FS_1_n58) );
  AOI21_X1 mul_ex_mult_86_FS_1_U67 ( .B1(mul_ex_mult_86_FS_1_n14), .B2(
        mul_ex_mult_86_FS_1_n59), .A(mul_ex_mult_86_FS_1_n60), .ZN(
        mul_ex_mult_86_FS_1_n56) );
  XOR2_X1 mul_ex_mult_86_FS_1_U66 ( .A(mul_ex_mult_86_FS_1_n58), .B(
        mul_ex_mult_86_FS_1_n56), .Z(mul_ex_N143) );
  OAI21_X1 mul_ex_mult_86_FS_1_U65 ( .B1(mul_ex_mult_86_FS_1_n55), .B2(
        mul_ex_mult_86_FS_1_n56), .A(mul_ex_mult_86_FS_1_n57), .ZN(
        mul_ex_mult_86_FS_1_n51) );
  AND2_X1 mul_ex_mult_86_FS_1_U64 ( .A1(mul_ex_mult_86_n50), .A2(
        mul_ex_mult_86_n21), .ZN(mul_ex_mult_86_FS_1_n52) );
  NOR2_X1 mul_ex_mult_86_FS_1_U63 ( .A1(mul_ex_mult_86_n50), .A2(
        mul_ex_mult_86_n21), .ZN(mul_ex_mult_86_FS_1_n53) );
  NOR2_X1 mul_ex_mult_86_FS_1_U62 ( .A1(mul_ex_mult_86_FS_1_n52), .A2(
        mul_ex_mult_86_FS_1_n53), .ZN(mul_ex_mult_86_FS_1_n54) );
  XOR2_X1 mul_ex_mult_86_FS_1_U61 ( .A(mul_ex_mult_86_FS_1_n51), .B(
        mul_ex_mult_86_FS_1_n54), .Z(mul_ex_N144) );
  NOR2_X1 mul_ex_mult_86_FS_1_U60 ( .A1(mul_ex_mult_86_n56), .A2(
        mul_ex_mult_86_n28), .ZN(mul_ex_mult_86_FS_1_n47) );
  NAND2_X1 mul_ex_mult_86_FS_1_U59 ( .A1(mul_ex_mult_86_n56), .A2(
        mul_ex_mult_86_n28), .ZN(mul_ex_mult_86_FS_1_n49) );
  NAND2_X1 mul_ex_mult_86_FS_1_U58 ( .A1(mul_ex_mult_86_FS_1_n11), .A2(
        mul_ex_mult_86_FS_1_n49), .ZN(mul_ex_mult_86_FS_1_n50) );
  AOI21_X1 mul_ex_mult_86_FS_1_U57 ( .B1(mul_ex_mult_86_FS_1_n12), .B2(
        mul_ex_mult_86_FS_1_n51), .A(mul_ex_mult_86_FS_1_n52), .ZN(
        mul_ex_mult_86_FS_1_n48) );
  XOR2_X1 mul_ex_mult_86_FS_1_U56 ( .A(mul_ex_mult_86_FS_1_n50), .B(
        mul_ex_mult_86_FS_1_n48), .Z(mul_ex_N145) );
  OAI21_X1 mul_ex_mult_86_FS_1_U55 ( .B1(mul_ex_mult_86_FS_1_n47), .B2(
        mul_ex_mult_86_FS_1_n48), .A(mul_ex_mult_86_FS_1_n49), .ZN(
        mul_ex_mult_86_FS_1_n43) );
  AND2_X1 mul_ex_mult_86_FS_1_U54 ( .A1(mul_ex_mult_86_n49), .A2(
        mul_ex_mult_86_n20), .ZN(mul_ex_mult_86_FS_1_n44) );
  NOR2_X1 mul_ex_mult_86_FS_1_U53 ( .A1(mul_ex_mult_86_n49), .A2(
        mul_ex_mult_86_n20), .ZN(mul_ex_mult_86_FS_1_n45) );
  NOR2_X1 mul_ex_mult_86_FS_1_U52 ( .A1(mul_ex_mult_86_FS_1_n44), .A2(
        mul_ex_mult_86_FS_1_n45), .ZN(mul_ex_mult_86_FS_1_n46) );
  XOR2_X1 mul_ex_mult_86_FS_1_U51 ( .A(mul_ex_mult_86_FS_1_n43), .B(
        mul_ex_mult_86_FS_1_n46), .Z(mul_ex_N146) );
  NOR2_X1 mul_ex_mult_86_FS_1_U50 ( .A1(mul_ex_mult_86_n55), .A2(
        mul_ex_mult_86_n27), .ZN(mul_ex_mult_86_FS_1_n39) );
  NAND2_X1 mul_ex_mult_86_FS_1_U49 ( .A1(mul_ex_mult_86_n55), .A2(
        mul_ex_mult_86_n27), .ZN(mul_ex_mult_86_FS_1_n41) );
  NAND2_X1 mul_ex_mult_86_FS_1_U48 ( .A1(mul_ex_mult_86_FS_1_n9), .A2(
        mul_ex_mult_86_FS_1_n41), .ZN(mul_ex_mult_86_FS_1_n42) );
  AOI21_X1 mul_ex_mult_86_FS_1_U47 ( .B1(mul_ex_mult_86_FS_1_n10), .B2(
        mul_ex_mult_86_FS_1_n43), .A(mul_ex_mult_86_FS_1_n44), .ZN(
        mul_ex_mult_86_FS_1_n40) );
  XOR2_X1 mul_ex_mult_86_FS_1_U46 ( .A(mul_ex_mult_86_FS_1_n42), .B(
        mul_ex_mult_86_FS_1_n40), .Z(mul_ex_N147) );
  OAI21_X1 mul_ex_mult_86_FS_1_U45 ( .B1(mul_ex_mult_86_FS_1_n39), .B2(
        mul_ex_mult_86_FS_1_n40), .A(mul_ex_mult_86_FS_1_n41), .ZN(
        mul_ex_mult_86_FS_1_n35) );
  AND2_X1 mul_ex_mult_86_FS_1_U44 ( .A1(mul_ex_mult_86_n48), .A2(
        mul_ex_mult_86_n19), .ZN(mul_ex_mult_86_FS_1_n36) );
  NOR2_X1 mul_ex_mult_86_FS_1_U43 ( .A1(mul_ex_mult_86_n48), .A2(
        mul_ex_mult_86_n19), .ZN(mul_ex_mult_86_FS_1_n37) );
  NOR2_X1 mul_ex_mult_86_FS_1_U42 ( .A1(mul_ex_mult_86_FS_1_n36), .A2(
        mul_ex_mult_86_FS_1_n37), .ZN(mul_ex_mult_86_FS_1_n38) );
  XOR2_X1 mul_ex_mult_86_FS_1_U41 ( .A(mul_ex_mult_86_FS_1_n35), .B(
        mul_ex_mult_86_FS_1_n38), .Z(mul_ex_N148) );
  NOR2_X1 mul_ex_mult_86_FS_1_U40 ( .A1(mul_ex_mult_86_n54), .A2(
        mul_ex_mult_86_n26), .ZN(mul_ex_mult_86_FS_1_n31) );
  NAND2_X1 mul_ex_mult_86_FS_1_U39 ( .A1(mul_ex_mult_86_n54), .A2(
        mul_ex_mult_86_n26), .ZN(mul_ex_mult_86_FS_1_n33) );
  NAND2_X1 mul_ex_mult_86_FS_1_U38 ( .A1(mul_ex_mult_86_FS_1_n7), .A2(
        mul_ex_mult_86_FS_1_n33), .ZN(mul_ex_mult_86_FS_1_n34) );
  AOI21_X1 mul_ex_mult_86_FS_1_U37 ( .B1(mul_ex_mult_86_FS_1_n8), .B2(
        mul_ex_mult_86_FS_1_n35), .A(mul_ex_mult_86_FS_1_n36), .ZN(
        mul_ex_mult_86_FS_1_n32) );
  XOR2_X1 mul_ex_mult_86_FS_1_U36 ( .A(mul_ex_mult_86_FS_1_n34), .B(
        mul_ex_mult_86_FS_1_n32), .Z(mul_ex_N149) );
  OAI21_X1 mul_ex_mult_86_FS_1_U35 ( .B1(mul_ex_mult_86_FS_1_n31), .B2(
        mul_ex_mult_86_FS_1_n32), .A(mul_ex_mult_86_FS_1_n33), .ZN(
        mul_ex_mult_86_FS_1_n27) );
  AND2_X1 mul_ex_mult_86_FS_1_U34 ( .A1(mul_ex_mult_86_n47), .A2(
        mul_ex_mult_86_n18), .ZN(mul_ex_mult_86_FS_1_n28) );
  NOR2_X1 mul_ex_mult_86_FS_1_U33 ( .A1(mul_ex_mult_86_n47), .A2(
        mul_ex_mult_86_n18), .ZN(mul_ex_mult_86_FS_1_n29) );
  NOR2_X1 mul_ex_mult_86_FS_1_U32 ( .A1(mul_ex_mult_86_FS_1_n28), .A2(
        mul_ex_mult_86_FS_1_n29), .ZN(mul_ex_mult_86_FS_1_n30) );
  XOR2_X1 mul_ex_mult_86_FS_1_U31 ( .A(mul_ex_mult_86_FS_1_n27), .B(
        mul_ex_mult_86_FS_1_n30), .Z(mul_ex_N150) );
  NOR2_X1 mul_ex_mult_86_FS_1_U30 ( .A1(mul_ex_mult_86_n53), .A2(
        mul_ex_mult_86_n25), .ZN(mul_ex_mult_86_FS_1_n23) );
  NAND2_X1 mul_ex_mult_86_FS_1_U29 ( .A1(mul_ex_mult_86_n53), .A2(
        mul_ex_mult_86_n25), .ZN(mul_ex_mult_86_FS_1_n25) );
  NAND2_X1 mul_ex_mult_86_FS_1_U28 ( .A1(mul_ex_mult_86_FS_1_n5), .A2(
        mul_ex_mult_86_FS_1_n25), .ZN(mul_ex_mult_86_FS_1_n26) );
  AOI21_X1 mul_ex_mult_86_FS_1_U27 ( .B1(mul_ex_mult_86_FS_1_n6), .B2(
        mul_ex_mult_86_FS_1_n27), .A(mul_ex_mult_86_FS_1_n28), .ZN(
        mul_ex_mult_86_FS_1_n24) );
  XOR2_X1 mul_ex_mult_86_FS_1_U26 ( .A(mul_ex_mult_86_FS_1_n26), .B(
        mul_ex_mult_86_FS_1_n24), .Z(mul_ex_N151) );
  OAI21_X1 mul_ex_mult_86_FS_1_U25 ( .B1(mul_ex_mult_86_FS_1_n23), .B2(
        mul_ex_mult_86_FS_1_n24), .A(mul_ex_mult_86_FS_1_n25), .ZN(
        mul_ex_mult_86_FS_1_n19) );
  AND2_X1 mul_ex_mult_86_FS_1_U24 ( .A1(mul_ex_mult_86_n46), .A2(
        mul_ex_mult_86_n17), .ZN(mul_ex_mult_86_FS_1_n20) );
  NOR2_X1 mul_ex_mult_86_FS_1_U23 ( .A1(mul_ex_mult_86_n46), .A2(
        mul_ex_mult_86_n17), .ZN(mul_ex_mult_86_FS_1_n21) );
  NOR2_X1 mul_ex_mult_86_FS_1_U22 ( .A1(mul_ex_mult_86_FS_1_n20), .A2(
        mul_ex_mult_86_FS_1_n21), .ZN(mul_ex_mult_86_FS_1_n22) );
  XOR2_X1 mul_ex_mult_86_FS_1_U21 ( .A(mul_ex_mult_86_FS_1_n19), .B(
        mul_ex_mult_86_FS_1_n22), .Z(mul_ex_N152) );
  AOI21_X1 mul_ex_mult_86_FS_1_U20 ( .B1(mul_ex_mult_86_FS_1_n19), .B2(
        mul_ex_mult_86_FS_1_n4), .A(mul_ex_mult_86_FS_1_n20), .ZN(
        mul_ex_mult_86_FS_1_n18) );
  XOR2_X1 mul_ex_mult_86_FS_1_U19 ( .A(mul_ex_mult_86_FS_1_n3), .B(
        mul_ex_mult_86_FS_1_n18), .Z(mul_ex_N153) );
  INV_X4 mul_ex_mult_86_FS_1_U18 ( .A(mul_ex_mult_86_FS_1_n70), .ZN(
        mul_ex_mult_86_FS_1_n17) );
  INV_X4 mul_ex_mult_86_FS_1_U17 ( .A(mul_ex_mult_86_FS_1_n68), .ZN(
        mul_ex_mult_86_FS_1_n16) );
  INV_X4 mul_ex_mult_86_FS_1_U16 ( .A(mul_ex_mult_86_FS_1_n63), .ZN(
        mul_ex_mult_86_FS_1_n15) );
  INV_X4 mul_ex_mult_86_FS_1_U15 ( .A(mul_ex_mult_86_FS_1_n61), .ZN(
        mul_ex_mult_86_FS_1_n14) );
  INV_X4 mul_ex_mult_86_FS_1_U14 ( .A(mul_ex_mult_86_FS_1_n55), .ZN(
        mul_ex_mult_86_FS_1_n13) );
  INV_X4 mul_ex_mult_86_FS_1_U13 ( .A(mul_ex_mult_86_FS_1_n53), .ZN(
        mul_ex_mult_86_FS_1_n12) );
  INV_X4 mul_ex_mult_86_FS_1_U12 ( .A(mul_ex_mult_86_FS_1_n47), .ZN(
        mul_ex_mult_86_FS_1_n11) );
  INV_X4 mul_ex_mult_86_FS_1_U11 ( .A(mul_ex_mult_86_FS_1_n45), .ZN(
        mul_ex_mult_86_FS_1_n10) );
  INV_X4 mul_ex_mult_86_FS_1_U10 ( .A(mul_ex_mult_86_FS_1_n39), .ZN(
        mul_ex_mult_86_FS_1_n9) );
  INV_X4 mul_ex_mult_86_FS_1_U9 ( .A(mul_ex_mult_86_FS_1_n37), .ZN(
        mul_ex_mult_86_FS_1_n8) );
  INV_X4 mul_ex_mult_86_FS_1_U8 ( .A(mul_ex_mult_86_FS_1_n31), .ZN(
        mul_ex_mult_86_FS_1_n7) );
  INV_X4 mul_ex_mult_86_FS_1_U7 ( .A(mul_ex_mult_86_FS_1_n29), .ZN(
        mul_ex_mult_86_FS_1_n6) );
  INV_X4 mul_ex_mult_86_FS_1_U6 ( .A(mul_ex_mult_86_FS_1_n23), .ZN(
        mul_ex_mult_86_FS_1_n5) );
  INV_X4 mul_ex_mult_86_FS_1_U5 ( .A(mul_ex_mult_86_FS_1_n21), .ZN(
        mul_ex_mult_86_FS_1_n4) );
  INV_X4 mul_ex_mult_86_FS_1_U4 ( .A(mul_ex_mult_86_n62), .ZN(
        mul_ex_mult_86_FS_1_n3) );
  AND2_X4 mul_ex_mult_86_FS_1_U3 ( .A1(mul_ex_mult_86_FS_1_n1), .A2(
        mul_ex_mult_86_FS_1_n70), .ZN(mul_ex_N139) );
  OR2_X4 mul_ex_mult_86_FS_1_U2 ( .A1(mul_ex_mult_86_n59), .A2(
        mul_ex_mult_86_n24), .ZN(mul_ex_mult_86_FS_1_n1) );
  INV_X4 CHOOSE_MULT_OR_INT_U8 ( .A(movi2fp_in), .ZN(CHOOSE_MULT_OR_INT_n1) );
  INV_X4 CHOOSE_MULT_OR_INT_U7 ( .A(movi2fp_in), .ZN(CHOOSE_MULT_OR_INT_n8) );
  INV_X4 CHOOSE_MULT_OR_INT_U6 ( .A(CHOOSE_MULT_OR_INT_n8), .ZN(
        CHOOSE_MULT_OR_INT_n7) );
  INV_X4 CHOOSE_MULT_OR_INT_U5 ( .A(CHOOSE_MULT_OR_INT_n1), .ZN(
        CHOOSE_MULT_OR_INT_n2) );
  INV_X4 CHOOSE_MULT_OR_INT_U4 ( .A(CHOOSE_MULT_OR_INT_n1), .ZN(
        CHOOSE_MULT_OR_INT_n3) );
  INV_X4 CHOOSE_MULT_OR_INT_U3 ( .A(CHOOSE_MULT_OR_INT_n1), .ZN(
        CHOOSE_MULT_OR_INT_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_U2 ( .A(CHOOSE_MULT_OR_INT_n8), .ZN(
        CHOOSE_MULT_OR_INT_n5) );
  INV_X4 CHOOSE_MULT_OR_INT_U1 ( .A(CHOOSE_MULT_OR_INT_n8), .ZN(
        CHOOSE_MULT_OR_INT_n6) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_0__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n2), 
        .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_0__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_0__MUX_U1 ( .A1(mul_result_long[0]), 
        .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_0__MUX_n2), .ZN(fbusW[0]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_1__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n2), 
        .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_1__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_1__MUX_U1 ( .A1(mul_result_long[1]), 
        .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_1__MUX_n2), .ZN(fbusW[1]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_2__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n2), 
        .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_2__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_2__MUX_U1 ( .A1(mul_result_long[2]), 
        .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_2__MUX_n2), .ZN(fbusW[2]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_3__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n2), 
        .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_3__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_3__MUX_U1 ( .A1(mul_result_long[3]), 
        .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_3__MUX_n2), .ZN(fbusW[3]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_4__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n2), 
        .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_4__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_4__MUX_U1 ( .A1(mul_result_long[4]), 
        .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_4__MUX_n2), .ZN(fbusW[4]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_5__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n2), 
        .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_5__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_5__MUX_U1 ( .A1(mul_result_long[5]), 
        .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_5__MUX_n2), .ZN(fbusW[5]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_6__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n2), 
        .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_6__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_6__MUX_U1 ( .A1(mul_result_long[6]), 
        .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_6__MUX_n2), .ZN(fbusW[6]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_7__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n2), 
        .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_7__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_7__MUX_U1 ( .A1(mul_result_long[7]), 
        .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_7__MUX_n2), .ZN(fbusW[7]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_8__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n2), 
        .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_8__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_8__MUX_U1 ( .A1(mul_result_long[8]), 
        .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_8__MUX_n2), .ZN(fbusW[8]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_9__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n2), 
        .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_9__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_9__MUX_U1 ( .A1(mul_result_long[9]), 
        .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_9__MUX_n2), .ZN(fbusW[9]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_10__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n2), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_10__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_10__MUX_U1 ( .A1(mul_result_long[10]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_10__MUX_n2), .ZN(fbusW[10]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_11__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n2), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_11__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_11__MUX_U1 ( .A1(mul_result_long[11]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_11__MUX_n2), .ZN(fbusW[11]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_12__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n3), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_12__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_12__MUX_U1 ( .A1(mul_result_long[12]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_12__MUX_n2), .ZN(fbusW[12]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_13__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n3), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_13__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_13__MUX_U1 ( .A1(mul_result_long[13]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_13__MUX_n2), .ZN(fbusW[13]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_14__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n3), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_14__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_14__MUX_U1 ( .A1(mul_result_long[14]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_14__MUX_n2), .ZN(fbusW[14]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_15__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n3), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_15__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_15__MUX_U1 ( .A1(mul_result_long[15]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_15__MUX_n2), .ZN(fbusW[15]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_16__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n3), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_16__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_16__MUX_U1 ( .A1(mul_result_long[16]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_16__MUX_n2), .ZN(fbusW[16]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_17__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n3), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_17__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_17__MUX_U1 ( .A1(mul_result_long[17]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_17__MUX_n2), .ZN(fbusW[17]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_18__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n3), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_18__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_18__MUX_U1 ( .A1(mul_result_long[18]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_18__MUX_n2), .ZN(fbusW[18]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_19__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n3), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_19__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_19__MUX_U1 ( .A1(mul_result_long[19]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_19__MUX_n2), .ZN(fbusW[19]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_20__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n3), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_20__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_20__MUX_U1 ( .A1(mul_result_long[20]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_20__MUX_n2), .ZN(fbusW[20]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_21__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n3), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_21__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_21__MUX_U1 ( .A1(mul_result_long[21]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_21__MUX_n2), .ZN(fbusW[21]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_22__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n3), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_22__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_22__MUX_U1 ( .A1(mul_result_long[22]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_22__MUX_n2), .ZN(fbusW[22]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_23__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n3), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_23__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_23__MUX_U1 ( .A1(mul_result_long[23]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_23__MUX_n2), .ZN(fbusW[23]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_24__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n4), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_24__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_24__MUX_U1 ( .A1(mul_result_long[24]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_24__MUX_n2), .ZN(fbusW[24]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_25__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n4), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_25__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_25__MUX_U1 ( .A1(mul_result_long[25]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_25__MUX_n2), .ZN(fbusW[25]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_26__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n4), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_26__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_26__MUX_U1 ( .A1(mul_result_long[26]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_26__MUX_n2), .ZN(fbusW[26]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_27__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n4), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_27__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_27__MUX_U1 ( .A1(mul_result_long[27]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_27__MUX_n2), .ZN(fbusW[27]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_28__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n4), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_28__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_28__MUX_U1 ( .A1(mul_result_long[28]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_28__MUX_n2), .ZN(fbusW[28]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_29__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n4), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_29__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_29__MUX_U1 ( .A1(mul_result_long[29]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_29__MUX_n2), .ZN(fbusW[29]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_30__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n4), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_30__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_30__MUX_U1 ( .A1(mul_result_long[30]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_30__MUX_n2), .ZN(fbusW[30]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_31__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n4), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_31__MUX_n2) );
  AND2_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_31__MUX_U1 ( .A1(mul_result_long[31]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_31__MUX_n2), .ZN(fbusW[31]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_32__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_32__MUX_n4), .ZN(fbusW[32]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_32__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n4), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_32__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_32__MUX_U1 ( .A1(
        mul_result_long[32]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_32__MUX_n1), 
        .B1(opA_in[0]), .B2(CHOOSE_MULT_OR_INT_n4), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_32__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_33__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_33__MUX_n4), .ZN(fbusW[33]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_33__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n4), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_33__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_33__MUX_U1 ( .A1(
        mul_result_long[33]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_33__MUX_n1), 
        .B1(opA_in[1]), .B2(CHOOSE_MULT_OR_INT_n4), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_33__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_34__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_34__MUX_n4), .ZN(fbusW[34]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_34__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n4), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_34__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_34__MUX_U1 ( .A1(
        mul_result_long[34]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_34__MUX_n1), 
        .B1(opA_in[2]), .B2(CHOOSE_MULT_OR_INT_n4), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_34__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_35__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_35__MUX_n4), .ZN(fbusW[35]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_35__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n4), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_35__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_35__MUX_U1 ( .A1(
        mul_result_long[35]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_35__MUX_n1), 
        .B1(opA_in[3]), .B2(CHOOSE_MULT_OR_INT_n4), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_35__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_36__MUX_U4 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_36__MUX_n5), .ZN(fbusW[36]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_36__MUX_U3 ( .A(CHOOSE_MULT_OR_INT_n5), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_36__MUX_n2) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_36__MUX_U2 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_36__MUX_n2), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_36__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_36__MUX_U1 ( .A1(
        mul_result_long[36]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_36__MUX_n2), 
        .B1(opA_in[4]), .B2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_36__MUX_n1), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_36__MUX_n5) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_37__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_37__MUX_n4), .ZN(fbusW[37]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_37__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n5), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_37__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_37__MUX_U1 ( .A1(
        mul_result_long[37]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_37__MUX_n1), 
        .B1(opA_in[5]), .B2(CHOOSE_MULT_OR_INT_n5), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_37__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_38__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_38__MUX_n4), .ZN(fbusW[38]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_38__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n5), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_38__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_38__MUX_U1 ( .A1(
        mul_result_long[38]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_38__MUX_n1), 
        .B1(opA_in[6]), .B2(CHOOSE_MULT_OR_INT_n5), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_38__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_39__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_39__MUX_n4), .ZN(fbusW[39]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_39__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n5), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_39__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_39__MUX_U1 ( .A1(
        mul_result_long[39]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_39__MUX_n1), 
        .B1(opA_in[7]), .B2(CHOOSE_MULT_OR_INT_n5), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_39__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_40__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_40__MUX_n4), .ZN(fbusW[40]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_40__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n5), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_40__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_40__MUX_U1 ( .A1(
        mul_result_long[40]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_40__MUX_n1), 
        .B1(opA_in[8]), .B2(CHOOSE_MULT_OR_INT_n5), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_40__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_41__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_41__MUX_n4), .ZN(fbusW[41]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_41__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n5), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_41__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_41__MUX_U1 ( .A1(
        mul_result_long[41]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_41__MUX_n1), 
        .B1(opA_in[9]), .B2(CHOOSE_MULT_OR_INT_n5), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_41__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_42__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_42__MUX_n4), .ZN(fbusW[42]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_42__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n5), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_42__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_42__MUX_U1 ( .A1(
        mul_result_long[42]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_42__MUX_n1), 
        .B1(opA_in[10]), .B2(CHOOSE_MULT_OR_INT_n5), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_42__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_43__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_43__MUX_n4), .ZN(fbusW[43]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_43__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n5), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_43__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_43__MUX_U1 ( .A1(
        mul_result_long[43]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_43__MUX_n1), 
        .B1(opA_in[11]), .B2(CHOOSE_MULT_OR_INT_n5), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_43__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_44__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_44__MUX_n4), .ZN(fbusW[44]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_44__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n5), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_44__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_44__MUX_U1 ( .A1(
        mul_result_long[44]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_44__MUX_n1), 
        .B1(opA_in[12]), .B2(CHOOSE_MULT_OR_INT_n5), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_44__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_45__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_45__MUX_n4), .ZN(fbusW[45]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_45__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n5), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_45__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_45__MUX_U1 ( .A1(
        mul_result_long[45]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_45__MUX_n1), 
        .B1(opA_in[13]), .B2(CHOOSE_MULT_OR_INT_n5), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_45__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_46__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_46__MUX_n4), .ZN(fbusW[46]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_46__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n5), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_46__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_46__MUX_U1 ( .A1(
        mul_result_long[46]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_46__MUX_n1), 
        .B1(opA_in[14]), .B2(CHOOSE_MULT_OR_INT_n5), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_46__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_47__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_47__MUX_n4), .ZN(fbusW[47]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_47__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n5), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_47__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_47__MUX_U1 ( .A1(
        mul_result_long[47]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_47__MUX_n1), 
        .B1(opA_in[15]), .B2(CHOOSE_MULT_OR_INT_n5), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_47__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_48__MUX_U4 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_48__MUX_n5), .ZN(fbusW[48]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_48__MUX_U3 ( .A(CHOOSE_MULT_OR_INT_n6), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_48__MUX_n2) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_48__MUX_U2 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_48__MUX_n2), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_48__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_48__MUX_U1 ( .A1(
        mul_result_long[48]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_48__MUX_n2), 
        .B1(opA_in[16]), .B2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_48__MUX_n1), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_48__MUX_n5) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_49__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_49__MUX_n4), .ZN(fbusW[49]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_49__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n6), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_49__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_49__MUX_U1 ( .A1(
        mul_result_long[49]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_49__MUX_n1), 
        .B1(opA_in[17]), .B2(CHOOSE_MULT_OR_INT_n6), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_49__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_50__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_50__MUX_n4), .ZN(fbusW[50]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_50__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n6), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_50__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_50__MUX_U1 ( .A1(
        mul_result_long[50]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_50__MUX_n1), 
        .B1(opA_in[18]), .B2(CHOOSE_MULT_OR_INT_n6), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_50__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_51__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_51__MUX_n4), .ZN(fbusW[51]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_51__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n6), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_51__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_51__MUX_U1 ( .A1(
        mul_result_long[51]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_51__MUX_n1), 
        .B1(opA_in[19]), .B2(CHOOSE_MULT_OR_INT_n6), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_51__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_52__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_52__MUX_n4), .ZN(fbusW[52]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_52__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n6), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_52__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_52__MUX_U1 ( .A1(
        mul_result_long[52]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_52__MUX_n1), 
        .B1(opA_in[20]), .B2(CHOOSE_MULT_OR_INT_n6), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_52__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_53__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_53__MUX_n4), .ZN(fbusW[53]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_53__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n6), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_53__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_53__MUX_U1 ( .A1(
        mul_result_long[53]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_53__MUX_n1), 
        .B1(opA_in[21]), .B2(CHOOSE_MULT_OR_INT_n6), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_53__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_54__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_54__MUX_n4), .ZN(fbusW[54]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_54__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n6), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_54__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_54__MUX_U1 ( .A1(
        mul_result_long[54]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_54__MUX_n1), 
        .B1(opA_in[22]), .B2(CHOOSE_MULT_OR_INT_n6), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_54__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_55__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_55__MUX_n4), .ZN(fbusW[55]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_55__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n6), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_55__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_55__MUX_U1 ( .A1(
        mul_result_long[55]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_55__MUX_n1), 
        .B1(opA_in[23]), .B2(CHOOSE_MULT_OR_INT_n6), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_55__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_56__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_56__MUX_n4), .ZN(fbusW[56]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_56__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n6), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_56__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_56__MUX_U1 ( .A1(
        mul_result_long[56]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_56__MUX_n1), 
        .B1(opA_in[24]), .B2(CHOOSE_MULT_OR_INT_n6), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_56__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_57__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_57__MUX_n4), .ZN(fbusW[57]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_57__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n6), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_57__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_57__MUX_U1 ( .A1(
        mul_result_long[57]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_57__MUX_n1), 
        .B1(opA_in[25]), .B2(CHOOSE_MULT_OR_INT_n6), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_57__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_58__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_58__MUX_n4), .ZN(fbusW[58]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_58__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n6), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_58__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_58__MUX_U1 ( .A1(
        mul_result_long[58]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_58__MUX_n1), 
        .B1(opA_in[26]), .B2(CHOOSE_MULT_OR_INT_n6), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_58__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_59__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_59__MUX_n4), .ZN(fbusW[59]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_59__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n6), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_59__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_59__MUX_U1 ( .A1(
        mul_result_long[59]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_59__MUX_n1), 
        .B1(opA_in[27]), .B2(CHOOSE_MULT_OR_INT_n6), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_59__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_60__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_60__MUX_n4), .ZN(fbusW[60]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_60__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n7), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_60__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_60__MUX_U1 ( .A1(
        mul_result_long[60]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_60__MUX_n1), 
        .B1(opA_in[28]), .B2(CHOOSE_MULT_OR_INT_n7), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_60__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_61__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_61__MUX_n4), .ZN(fbusW[61]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_61__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n7), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_61__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_61__MUX_U1 ( .A1(
        mul_result_long[61]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_61__MUX_n1), 
        .B1(opA_in[29]), .B2(CHOOSE_MULT_OR_INT_n7), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_61__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_62__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_62__MUX_n4), .ZN(fbusW[62]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_62__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n7), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_62__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_62__MUX_U1 ( .A1(
        mul_result_long[62]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_62__MUX_n1), 
        .B1(opA_in[30]), .B2(CHOOSE_MULT_OR_INT_n7), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_62__MUX_n4) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_63__MUX_U3 ( .A(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_63__MUX_n4), .ZN(fbusW[63]) );
  INV_X4 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_63__MUX_U2 ( .A(CHOOSE_MULT_OR_INT_n7), .ZN(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_63__MUX_n1) );
  AOI22_X2 CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_63__MUX_U1 ( .A1(
        mul_result_long[63]), .A2(CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_63__MUX_n1), 
        .B1(opA_in[31]), .B2(CHOOSE_MULT_OR_INT_n7), .ZN(
        CHOOSE_MULT_OR_INT_MUX2TO1_NBIT_63__MUX_n4) );
  INV_X4 decide_if_leap_U3 ( .A(decide_if_leap_n2), .ZN(leap_out) );
  AOI21_X2 decide_if_leap_U1 ( .B1(decide_if_leap_n3), .B2(branch_in), .A(
        jump_in), .ZN(decide_if_leap_n2) );
  XNOR2_X2 decide_if_leap_U2 ( .A(decide_if_leap_zeroBit), .B(branchZero_in), 
        .ZN(decide_if_leap_n3) );
  NOR2_X2 decide_if_leap_ZERO_A_U1 ( .A1(decide_if_leap_ZERO_A_n1), .A2(
        decide_if_leap_ZERO_A_n2), .ZN(decide_if_leap_zeroBit) );
  NOR4_X2 decide_if_leap_ZERO_A_U11 ( .A1(opA_in[27]), .A2(opA_in[26]), .A3(
        opA_in[25]), .A4(opA_in[24]), .ZN(decide_if_leap_ZERO_A_n7) );
  NOR4_X2 decide_if_leap_ZERO_A_U10 ( .A1(opA_in[30]), .A2(opA_in[2]), .A3(
        opA_in[29]), .A4(opA_in[28]), .ZN(decide_if_leap_ZERO_A_n8) );
  NOR4_X2 decide_if_leap_ZERO_A_U9 ( .A1(opA_in[5]), .A2(opA_in[4]), .A3(
        opA_in[3]), .A4(opA_in[31]), .ZN(decide_if_leap_ZERO_A_n9) );
  NOR4_X2 decide_if_leap_ZERO_A_U8 ( .A1(opA_in[9]), .A2(opA_in[8]), .A3(
        opA_in[7]), .A4(opA_in[6]), .ZN(decide_if_leap_ZERO_A_n10) );
  NAND4_X2 decide_if_leap_ZERO_A_U7 ( .A1(decide_if_leap_ZERO_A_n7), .A2(
        decide_if_leap_ZERO_A_n8), .A3(decide_if_leap_ZERO_A_n9), .A4(
        decide_if_leap_ZERO_A_n10), .ZN(decide_if_leap_ZERO_A_n1) );
  NOR4_X2 decide_if_leap_ZERO_A_U6 ( .A1(opA_in[12]), .A2(opA_in[11]), .A3(
        opA_in[10]), .A4(opA_in[0]), .ZN(decide_if_leap_ZERO_A_n3) );
  NOR4_X2 decide_if_leap_ZERO_A_U5 ( .A1(opA_in[16]), .A2(opA_in[15]), .A3(
        opA_in[14]), .A4(opA_in[13]), .ZN(decide_if_leap_ZERO_A_n4) );
  NOR4_X2 decide_if_leap_ZERO_A_U4 ( .A1(opA_in[1]), .A2(opA_in[19]), .A3(
        opA_in[18]), .A4(opA_in[17]), .ZN(decide_if_leap_ZERO_A_n5) );
  NOR4_X2 decide_if_leap_ZERO_A_U3 ( .A1(opA_in[23]), .A2(opA_in[22]), .A3(
        opA_in[21]), .A4(opA_in[20]), .ZN(decide_if_leap_ZERO_A_n6) );
  NAND4_X2 decide_if_leap_ZERO_A_U2 ( .A1(decide_if_leap_ZERO_A_n3), .A2(
        decide_if_leap_ZERO_A_n4), .A3(decide_if_leap_ZERO_A_n5), .A4(
        decide_if_leap_ZERO_A_n6), .ZN(decide_if_leap_ZERO_A_n2) );
  INV_X32 EXTEND_IMM16_U34 ( .A(EXTEND_IMM16_n18), .ZN(imm16_32[15]) );
  INV_X32 EXTEND_IMM16_U33 ( .A(EXTEND_IMM16_n18), .ZN(imm16_32[14]) );
  INV_X32 EXTEND_IMM16_U32 ( .A(EXTEND_IMM16_n18), .ZN(imm16_32[13]) );
  INV_X32 EXTEND_IMM16_U31 ( .A(EXTEND_IMM16_n18), .ZN(imm16_32[12]) );
  INV_X32 EXTEND_IMM16_U30 ( .A(EXTEND_IMM16_n18), .ZN(imm16_32[11]) );
  INV_X32 EXTEND_IMM16_U29 ( .A(EXTEND_IMM16_n18), .ZN(imm16_32[10]) );
  INV_X32 EXTEND_IMM16_U28 ( .A(EXTEND_IMM16_n18), .ZN(imm16_32[9]) );
  INV_X32 EXTEND_IMM16_U27 ( .A(EXTEND_IMM16_n18), .ZN(imm16_32[8]) );
  INV_X32 EXTEND_IMM16_U26 ( .A(EXTEND_IMM16_n18), .ZN(imm16_32[7]) );
  INV_X32 EXTEND_IMM16_U25 ( .A(EXTEND_IMM16_n18), .ZN(imm16_32[6]) );
  INV_X32 EXTEND_IMM16_U24 ( .A(EXTEND_IMM16_n18), .ZN(imm16_32[5]) );
  INV_X32 EXTEND_IMM16_U23 ( .A(EXTEND_IMM16_n18), .ZN(imm16_32[4]) );
  INV_X32 EXTEND_IMM16_U22 ( .A(EXTEND_IMM16_n18), .ZN(imm16_32[3]) );
  INV_X32 EXTEND_IMM16_U21 ( .A(EXTEND_IMM16_n18), .ZN(imm16_32[2]) );
  INV_X32 EXTEND_IMM16_U20 ( .A(EXTEND_IMM16_n18), .ZN(imm16_32[1]) );
  INV_X32 EXTEND_IMM16_U19 ( .A(imm16_32[0]), .ZN(EXTEND_IMM16_n18) );
  BUF_X32 EXTEND_IMM16_U18 ( .A(offset16_in[0]), .Z(imm16_32[16]) );
  BUF_X32 EXTEND_IMM16_U17 ( .A(offset16_in[1]), .Z(imm16_32[17]) );
  BUF_X32 EXTEND_IMM16_U16 ( .A(offset16_in[2]), .Z(imm16_32[18]) );
  BUF_X32 EXTEND_IMM16_U15 ( .A(offset16_in[3]), .Z(imm16_32[19]) );
  BUF_X32 EXTEND_IMM16_U14 ( .A(offset16_in[4]), .Z(imm16_32[20]) );
  BUF_X32 EXTEND_IMM16_U13 ( .A(offset16_in[5]), .Z(imm16_32[21]) );
  BUF_X32 EXTEND_IMM16_U12 ( .A(offset16_in[6]), .Z(imm16_32[22]) );
  BUF_X32 EXTEND_IMM16_U11 ( .A(offset16_in[7]), .Z(imm16_32[23]) );
  BUF_X32 EXTEND_IMM16_U10 ( .A(offset16_in[8]), .Z(imm16_32[24]) );
  BUF_X32 EXTEND_IMM16_U9 ( .A(offset16_in[9]), .Z(imm16_32[25]) );
  BUF_X32 EXTEND_IMM16_U8 ( .A(offset16_in[10]), .Z(imm16_32[26]) );
  BUF_X32 EXTEND_IMM16_U7 ( .A(offset16_in[11]), .Z(imm16_32[27]) );
  BUF_X32 EXTEND_IMM16_U6 ( .A(offset16_in[12]), .Z(imm16_32[28]) );
  BUF_X32 EXTEND_IMM16_U5 ( .A(offset16_in[13]), .Z(imm16_32[29]) );
  BUF_X32 EXTEND_IMM16_U4 ( .A(offset16_in[14]), .Z(imm16_32[30]) );
  BUF_X32 EXTEND_IMM16_U3 ( .A(offset16_in[15]), .Z(imm16_32[31]) );
  BUF_X32 EXTEND_IMM16_SELECT_EXTEND_U1 ( .A(offset16_in[0]), .Z(imm16_32[0])
         );
  BUF_X32 EXTEND_IMM26_U33 ( .A(imm26_32[0]), .Z(imm26_32[5]) );
  BUF_X32 EXTEND_IMM26_U32 ( .A(imm26_32[0]), .Z(imm26_32[4]) );
  BUF_X32 EXTEND_IMM26_U31 ( .A(imm26_32[0]), .Z(imm26_32[3]) );
  BUF_X32 EXTEND_IMM26_U30 ( .A(imm26_32[0]), .Z(imm26_32[2]) );
  BUF_X32 EXTEND_IMM26_U29 ( .A(imm26_32[0]), .Z(imm26_32[1]) );
  BUF_X32 EXTEND_IMM26_U28 ( .A(offset26_in[0]), .Z(imm26_32[6]) );
  BUF_X32 EXTEND_IMM26_U27 ( .A(offset26_in[1]), .Z(imm26_32[7]) );
  BUF_X32 EXTEND_IMM26_U26 ( .A(offset26_in[2]), .Z(imm26_32[8]) );
  BUF_X32 EXTEND_IMM26_U25 ( .A(offset26_in[3]), .Z(imm26_32[9]) );
  BUF_X32 EXTEND_IMM26_U24 ( .A(offset26_in[4]), .Z(imm26_32[10]) );
  BUF_X32 EXTEND_IMM26_U23 ( .A(offset26_in[5]), .Z(imm26_32[11]) );
  BUF_X32 EXTEND_IMM26_U22 ( .A(offset26_in[6]), .Z(imm26_32[12]) );
  BUF_X32 EXTEND_IMM26_U21 ( .A(offset26_in[7]), .Z(imm26_32[13]) );
  BUF_X32 EXTEND_IMM26_U20 ( .A(offset26_in[8]), .Z(imm26_32[14]) );
  BUF_X32 EXTEND_IMM26_U19 ( .A(offset26_in[9]), .Z(imm26_32[15]) );
  BUF_X32 EXTEND_IMM26_U18 ( .A(offset26_in[10]), .Z(imm26_32[16]) );
  BUF_X32 EXTEND_IMM26_U17 ( .A(offset26_in[11]), .Z(imm26_32[17]) );
  BUF_X32 EXTEND_IMM26_U16 ( .A(offset26_in[12]), .Z(imm26_32[18]) );
  BUF_X32 EXTEND_IMM26_U15 ( .A(offset26_in[13]), .Z(imm26_32[19]) );
  BUF_X32 EXTEND_IMM26_U14 ( .A(offset26_in[14]), .Z(imm26_32[20]) );
  BUF_X32 EXTEND_IMM26_U13 ( .A(offset26_in[15]), .Z(imm26_32[21]) );
  BUF_X32 EXTEND_IMM26_U12 ( .A(offset26_in[16]), .Z(imm26_32[22]) );
  BUF_X32 EXTEND_IMM26_U11 ( .A(offset26_in[17]), .Z(imm26_32[23]) );
  BUF_X32 EXTEND_IMM26_U10 ( .A(offset26_in[18]), .Z(imm26_32[24]) );
  BUF_X32 EXTEND_IMM26_U9 ( .A(offset26_in[19]), .Z(imm26_32[25]) );
  BUF_X32 EXTEND_IMM26_U8 ( .A(offset26_in[20]), .Z(imm26_32[26]) );
  BUF_X32 EXTEND_IMM26_U7 ( .A(offset26_in[21]), .Z(imm26_32[27]) );
  BUF_X32 EXTEND_IMM26_U6 ( .A(offset26_in[22]), .Z(imm26_32[28]) );
  BUF_X32 EXTEND_IMM26_U5 ( .A(offset26_in[23]), .Z(imm26_32[29]) );
  BUF_X32 EXTEND_IMM26_U4 ( .A(offset26_in[24]), .Z(imm26_32[30]) );
  BUF_X32 EXTEND_IMM26_U3 ( .A(offset26_in[25]), .Z(imm26_32[31]) );
  BUF_X4 EXTEND_IMM26_SELECT_EXTEND_U1 ( .A(offset26_in[0]), .Z(imm26_32[0])
         );
  INV_X4 CHOOSE_IMMEDIATE_U3 ( .A(branch_in), .ZN(CHOOSE_IMMEDIATE_n3) );
  INV_X4 CHOOSE_IMMEDIATE_U2 ( .A(CHOOSE_IMMEDIATE_n3), .ZN(
        CHOOSE_IMMEDIATE_n1) );
  INV_X4 CHOOSE_IMMEDIATE_U1 ( .A(CHOOSE_IMMEDIATE_n3), .ZN(
        CHOOSE_IMMEDIATE_n2) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_0__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_0__MUX_n4), .ZN(leapAddr_out[0]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_0__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n1), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_0__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_0__MUX_U1 ( .A1(imm26_32[0]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_0__MUX_n1), .B1(imm16_32[0]), .B2(
        CHOOSE_IMMEDIATE_n1), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_0__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_1__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_1__MUX_n4), .ZN(leapAddr_out[1]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_1__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n1), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_1__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_1__MUX_U1 ( .A1(imm26_32[1]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_1__MUX_n1), .B1(imm16_32[1]), .B2(
        CHOOSE_IMMEDIATE_n1), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_1__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_2__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_2__MUX_n4), .ZN(leapAddr_out[2]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_2__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n1), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_2__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_2__MUX_U1 ( .A1(imm26_32[2]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_2__MUX_n1), .B1(imm16_32[2]), .B2(
        CHOOSE_IMMEDIATE_n1), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_2__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_3__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_3__MUX_n4), .ZN(leapAddr_out[3]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_3__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n1), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_3__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_3__MUX_U1 ( .A1(imm26_32[3]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_3__MUX_n1), .B1(imm16_32[3]), .B2(
        CHOOSE_IMMEDIATE_n1), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_3__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_4__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_4__MUX_n4), .ZN(leapAddr_out[4]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_4__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n1), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_4__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_4__MUX_U1 ( .A1(imm26_32[4]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_4__MUX_n1), .B1(imm16_32[4]), .B2(
        CHOOSE_IMMEDIATE_n1), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_4__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_5__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_5__MUX_n4), .ZN(leapAddr_out[5]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_5__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n1), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_5__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_5__MUX_U1 ( .A1(imm26_32[5]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_5__MUX_n1), .B1(imm16_32[5]), .B2(
        CHOOSE_IMMEDIATE_n1), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_5__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_6__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_6__MUX_n4), .ZN(leapAddr_out[6]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_6__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n1), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_6__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_6__MUX_U1 ( .A1(imm26_32[6]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_6__MUX_n1), .B1(imm16_32[6]), .B2(
        CHOOSE_IMMEDIATE_n1), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_6__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_7__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_7__MUX_n4), .ZN(leapAddr_out[7]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_7__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n1), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_7__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_7__MUX_U1 ( .A1(imm26_32[7]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_7__MUX_n1), .B1(imm16_32[7]), .B2(
        CHOOSE_IMMEDIATE_n1), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_7__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_8__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_8__MUX_n4), .ZN(leapAddr_out[8]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_8__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n1), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_8__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_8__MUX_U1 ( .A1(imm26_32[8]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_8__MUX_n1), .B1(imm16_32[8]), .B2(
        CHOOSE_IMMEDIATE_n1), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_8__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_9__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_9__MUX_n4), .ZN(leapAddr_out[9]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_9__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n1), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_9__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_9__MUX_U1 ( .A1(imm26_32[9]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_9__MUX_n1), .B1(imm16_32[9]), .B2(
        CHOOSE_IMMEDIATE_n1), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_9__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_10__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_10__MUX_n4), .ZN(leapAddr_out[10]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_10__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n1), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_10__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_10__MUX_U1 ( .A1(imm26_32[10]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_10__MUX_n1), .B1(imm16_32[10]), .B2(
        CHOOSE_IMMEDIATE_n1), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_10__MUX_n4)
         );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_11__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_11__MUX_n4), .ZN(leapAddr_out[11]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_11__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n1), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_11__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_11__MUX_U1 ( .A1(imm26_32[11]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_11__MUX_n1), .B1(imm16_32[11]), .B2(
        CHOOSE_IMMEDIATE_n1), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_11__MUX_n4)
         );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_12__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_12__MUX_n4), .ZN(leapAddr_out[12]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_12__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n2), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_12__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_12__MUX_U1 ( .A1(imm26_32[12]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_12__MUX_n1), .B1(imm16_32[12]), .B2(
        CHOOSE_IMMEDIATE_n2), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_12__MUX_n4)
         );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_13__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_13__MUX_n4), .ZN(leapAddr_out[13]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_13__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n2), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_13__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_13__MUX_U1 ( .A1(imm26_32[13]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_13__MUX_n1), .B1(imm16_32[13]), .B2(
        CHOOSE_IMMEDIATE_n2), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_13__MUX_n4)
         );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_14__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_14__MUX_n4), .ZN(leapAddr_out[14]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_14__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n2), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_14__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_14__MUX_U1 ( .A1(imm26_32[14]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_14__MUX_n1), .B1(imm16_32[14]), .B2(
        CHOOSE_IMMEDIATE_n2), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_14__MUX_n4)
         );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_15__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_15__MUX_n4), .ZN(leapAddr_out[15]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_15__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n2), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_15__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_15__MUX_U1 ( .A1(imm26_32[15]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_15__MUX_n1), .B1(imm16_32[15]), .B2(
        CHOOSE_IMMEDIATE_n2), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_15__MUX_n4)
         );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_16__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_16__MUX_n4), .ZN(leapAddr_out[16]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_16__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n2), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_16__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_16__MUX_U1 ( .A1(imm26_32[16]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_16__MUX_n1), .B1(imm16_32[16]), .B2(
        CHOOSE_IMMEDIATE_n2), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_16__MUX_n4)
         );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_17__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_17__MUX_n4), .ZN(leapAddr_out[17]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_17__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n2), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_17__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_17__MUX_U1 ( .A1(imm26_32[17]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_17__MUX_n1), .B1(imm16_32[17]), .B2(
        CHOOSE_IMMEDIATE_n2), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_17__MUX_n4)
         );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_18__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_18__MUX_n4), .ZN(leapAddr_out[18]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_18__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n2), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_18__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_18__MUX_U1 ( .A1(imm26_32[18]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_18__MUX_n1), .B1(imm16_32[18]), .B2(
        CHOOSE_IMMEDIATE_n2), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_18__MUX_n4)
         );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_19__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_19__MUX_n4), .ZN(leapAddr_out[19]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_19__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n2), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_19__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_19__MUX_U1 ( .A1(imm26_32[19]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_19__MUX_n1), .B1(imm16_32[19]), .B2(
        CHOOSE_IMMEDIATE_n2), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_19__MUX_n4)
         );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_20__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_20__MUX_n4), .ZN(leapAddr_out[20]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_20__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n2), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_20__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_20__MUX_U1 ( .A1(imm26_32[20]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_20__MUX_n1), .B1(imm16_32[20]), .B2(
        CHOOSE_IMMEDIATE_n2), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_20__MUX_n4)
         );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_21__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_21__MUX_n4), .ZN(leapAddr_out[21]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_21__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n2), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_21__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_21__MUX_U1 ( .A1(imm26_32[21]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_21__MUX_n1), .B1(imm16_32[21]), .B2(
        CHOOSE_IMMEDIATE_n2), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_21__MUX_n4)
         );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_22__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_22__MUX_n4), .ZN(leapAddr_out[22]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_22__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n2), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_22__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_22__MUX_U1 ( .A1(imm26_32[22]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_22__MUX_n1), .B1(imm16_32[22]), .B2(
        CHOOSE_IMMEDIATE_n2), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_22__MUX_n4)
         );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_23__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_23__MUX_n4), .ZN(leapAddr_out[23]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_23__MUX_U2 ( .A(CHOOSE_IMMEDIATE_n2), 
        .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_23__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_23__MUX_U1 ( .A1(imm26_32[23]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_23__MUX_n1), .B1(imm16_32[23]), .B2(
        CHOOSE_IMMEDIATE_n2), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_23__MUX_n4)
         );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_24__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_24__MUX_n4), .ZN(leapAddr_out[24]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_24__MUX_U2 ( .A(branch_in), .ZN(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_24__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_24__MUX_U1 ( .A1(imm26_32[24]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_24__MUX_n1), .B1(imm16_32[24]), .B2(
        branch_in), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_24__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_25__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_25__MUX_n4), .ZN(leapAddr_out[25]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_25__MUX_U2 ( .A(branch_in), .ZN(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_25__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_25__MUX_U1 ( .A1(imm26_32[25]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_25__MUX_n1), .B1(imm16_32[25]), .B2(
        branch_in), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_25__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_26__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_26__MUX_n4), .ZN(leapAddr_out[26]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_26__MUX_U2 ( .A(branch_in), .ZN(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_26__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_26__MUX_U1 ( .A1(imm26_32[26]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_26__MUX_n1), .B1(imm16_32[26]), .B2(
        branch_in), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_26__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_27__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_27__MUX_n4), .ZN(leapAddr_out[27]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_27__MUX_U2 ( .A(branch_in), .ZN(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_27__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_27__MUX_U1 ( .A1(imm26_32[27]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_27__MUX_n1), .B1(imm16_32[27]), .B2(
        branch_in), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_27__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_28__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_28__MUX_n4), .ZN(leapAddr_out[28]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_28__MUX_U2 ( .A(branch_in), .ZN(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_28__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_28__MUX_U1 ( .A1(imm26_32[28]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_28__MUX_n1), .B1(imm16_32[28]), .B2(
        branch_in), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_28__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_29__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_29__MUX_n4), .ZN(leapAddr_out[29]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_29__MUX_U2 ( .A(branch_in), .ZN(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_29__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_29__MUX_U1 ( .A1(imm26_32[29]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_29__MUX_n1), .B1(imm16_32[29]), .B2(
        branch_in), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_29__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_30__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_30__MUX_n4), .ZN(leapAddr_out[30]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_30__MUX_U2 ( .A(branch_in), .ZN(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_30__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_30__MUX_U1 ( .A1(imm26_32[30]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_30__MUX_n1), .B1(imm16_32[30]), .B2(
        branch_in), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_30__MUX_n4) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_31__MUX_U3 ( .A(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_31__MUX_n4), .ZN(leapAddr_out[31]) );
  INV_X4 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_31__MUX_U2 ( .A(branch_in), .ZN(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_31__MUX_n1) );
  AOI22_X2 CHOOSE_IMMEDIATE_MUX2TO1_32BIT_31__MUX_U1 ( .A1(imm26_32[31]), .A2(
        CHOOSE_IMMEDIATE_MUX2TO1_32BIT_31__MUX_n1), .B1(imm16_32[31]), .B2(
        branch_in), .ZN(CHOOSE_IMMEDIATE_MUX2TO1_32BIT_31__MUX_n4) );
endmodule

